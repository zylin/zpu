-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0bba",
     1 => x"f0040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"d5040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0bbd",
    73 => x"89040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0bbcec",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80fc",
   162 => x"cc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"bcef0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0bbd",
   169 => x"bd040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0bbd",
   177 => x"a5040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80fcdc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053351",
   258 => x"bb893f71",
   259 => x"b00c833d",
   260 => x"0d04fd3d",
   261 => x"0d818cc0",
   262 => x"0852f881",
   263 => x"c08e800b",
   264 => x"80fce808",
   265 => x"55537180",
   266 => x"2e80f738",
   267 => x"7281ff06",
   268 => x"84150c80",
   269 => x"fcbc3370",
   270 => x"81ff0651",
   271 => x"5271802e",
   272 => x"80c23872",
   273 => x"9f2a7310",
   274 => x"0753818c",
   275 => x"c4337081",
   276 => x"ff065152",
   277 => x"71802ed4",
   278 => x"38800b81",
   279 => x"8cc43494",
   280 => x"993f80fc",
   281 => x"b8335473",
   282 => x"80e23880",
   283 => x"fce80873",
   284 => x"81ff0684",
   285 => x"120c80fc",
   286 => x"bc337081",
   287 => x"ff065153",
   288 => x"5471c038",
   289 => x"72812a73",
   290 => x"9f2b0753",
   291 => x"ffbc3972",
   292 => x"812a739f",
   293 => x"2b075380",
   294 => x"fd51b8e0",
   295 => x"3f80fce8",
   296 => x"08547281",
   297 => x"ff068415",
   298 => x"0c80fcbc",
   299 => x"337081ff",
   300 => x"06535471",
   301 => x"802ed838",
   302 => x"729f2a73",
   303 => x"10075380",
   304 => x"fd51b8b8",
   305 => x"3f80fce8",
   306 => x"0854d739",
   307 => x"800bb00c",
   308 => x"853d0d04",
   309 => x"fb3d0d8a",
   310 => x"51b4a03f",
   311 => x"8b823fac",
   312 => x"b2530b0b",
   313 => x"80e69852",
   314 => x"0b0b80e6",
   315 => x"a8518b83",
   316 => x"3facc953",
   317 => x"0b0b80e6",
   318 => x"b0520b0b",
   319 => x"80e6cc51",
   320 => x"8af13f90",
   321 => x"f4530b0b",
   322 => x"80e6d452",
   323 => x"0b0b80e6",
   324 => x"e4518adf",
   325 => x"3fb4da53",
   326 => x"0b0b80e6",
   327 => x"ec520b0b",
   328 => x"80f2e051",
   329 => x"8acd3fb6",
   330 => x"c2530b0b",
   331 => x"80e78452",
   332 => x"0b0b80e6",
   333 => x"fc518abb",
   334 => x"3fb8e353",
   335 => x"0b0b80e7",
   336 => x"90520b0b",
   337 => x"80e7b051",
   338 => x"8aa93fb9",
   339 => x"ce530b0b",
   340 => x"80e7b852",
   341 => x"0b0b80e7",
   342 => x"dc518a97",
   343 => x"3fba8753",
   344 => x"0b0b80e7",
   345 => x"e4520b0b",
   346 => x"80e88051",
   347 => x"8a853fba",
   348 => x"bd530b0b",
   349 => x"80e88852",
   350 => x"0b0b80e8",
   351 => x"ac5189f3",
   352 => x"3fb9a353",
   353 => x"0b0b80e8",
   354 => x"b4520b0b",
   355 => x"80e8cc51",
   356 => x"89e13fb9",
   357 => x"bc530b0b",
   358 => x"80e8d452",
   359 => x"0b0b80e8",
   360 => x"f05189cf",
   361 => x"3fb7b853",
   362 => x"0b0b80e8",
   363 => x"f8520b0b",
   364 => x"80e99051",
   365 => x"89bd3fb8",
   366 => x"8e530b0b",
   367 => x"80e99852",
   368 => x"0b0b80e9",
   369 => x"b45189ab",
   370 => x"3f91cd53",
   371 => x"0b0b80e9",
   372 => x"bc520b0b",
   373 => x"80e9d051",
   374 => x"89993f91",
   375 => x"8d530b0b",
   376 => x"80e9d852",
   377 => x"0b0b80ea",
   378 => x"80518987",
   379 => x"3fb3bb53",
   380 => x"0b0b80ea",
   381 => x"88520b0b",
   382 => x"80ea9c51",
   383 => x"88f53f88",
   384 => x"92530b0b",
   385 => x"80eaa452",
   386 => x"0b0b80ea",
   387 => x"b45188e3",
   388 => x"3fa6eb53",
   389 => x"0b0b80ea",
   390 => x"b8520b0b",
   391 => x"80eacc51",
   392 => x"88d13fa9",
   393 => x"f3530b0b",
   394 => x"80ead052",
   395 => x"0b0b80ea",
   396 => x"f85188bf",
   397 => x"3fb4ae53",
   398 => x"0b0b80eb",
   399 => x"80520b0b",
   400 => x"80eb9051",
   401 => x"88ad3f92",
   402 => x"c7530b0b",
   403 => x"80eb9452",
   404 => x"0b0b80eb",
   405 => x"ac51889b",
   406 => x"3faaad53",
   407 => x"0b0b80eb",
   408 => x"b4520b0b",
   409 => x"80ebc051",
   410 => x"88893fab",
   411 => x"dc530b0b",
   412 => x"80ebc452",
   413 => x"0b0b80eb",
   414 => x"ec5187f7",
   415 => x"3faaad53",
   416 => x"0b0b80eb",
   417 => x"f4520b0b",
   418 => x"80ec9451",
   419 => x"87e53fac",
   420 => x"a2530b0b",
   421 => x"80ec9852",
   422 => x"0b0b80ec",
   423 => x"a85187d3",
   424 => x"3f90c053",
   425 => x"0b0b80f6",
   426 => x"d8520b0b",
   427 => x"80e69051",
   428 => x"87c13f8e",
   429 => x"a53f8898",
   430 => x"3f810b81",
   431 => x"a4b43481",
   432 => x"8cc43370",
   433 => x"81ff0655",
   434 => x"557381ea",
   435 => x"38b58f3f",
   436 => x"b00881d3",
   437 => x"3888873f",
   438 => x"80fce808",
   439 => x"70087084",
   440 => x"2a810651",
   441 => x"55567380",
   442 => x"2e80f238",
   443 => x"f881c08e",
   444 => x"8055818c",
   445 => x"c008802e",
   446 => x"81833874",
   447 => x"81ff0684",
   448 => x"170c80fc",
   449 => x"bc337081",
   450 => x"ff065154",
   451 => x"73802e80",
   452 => x"c138749f",
   453 => x"2a751007",
   454 => x"55818cc4",
   455 => x"337081ff",
   456 => x"06515473",
   457 => x"802ed438",
   458 => x"800b818c",
   459 => x"c4348eca",
   460 => x"3f80fcb8",
   461 => x"335675a5",
   462 => x"3880fce8",
   463 => x"087581ff",
   464 => x"0684120c",
   465 => x"80fcbc33",
   466 => x"7081ff06",
   467 => x"51555673",
   468 => x"c1387481",
   469 => x"2a759f2b",
   470 => x"0755ffbd",
   471 => x"3981a4b4",
   472 => x"335574fe",
   473 => x"da38873d",
   474 => x"0d047481",
   475 => x"2a759f2b",
   476 => x"075580fd",
   477 => x"51b3853f",
   478 => x"80fce808",
   479 => x"567481ff",
   480 => x"0684170c",
   481 => x"80fcbc33",
   482 => x"7081ff06",
   483 => x"57547580",
   484 => x"2ed83874",
   485 => x"9f2a7510",
   486 => x"075580fd",
   487 => x"51b2dd3f",
   488 => x"80fce808",
   489 => x"56d739b3",
   490 => x"c83fb008",
   491 => x"81ff0651",
   492 => x"879a3ffe",
   493 => x"a039800b",
   494 => x"818cc434",
   495 => x"8dbc3fb3",
   496 => x"9d3fb008",
   497 => x"802efe8d",
   498 => x"38dd3980",
   499 => x"3d0d0b0b",
   500 => x"80ecb051",
   501 => x"aebf3f8c",
   502 => x"51aea03f",
   503 => x"0b0b80ec",
   504 => x"b451aeb1",
   505 => x"3f818cc0",
   506 => x"08802e8e",
   507 => x"380b0b80",
   508 => x"eccc51ae",
   509 => x"a03f823d",
   510 => x"0d040b0b",
   511 => x"80ecd851",
   512 => x"ae933f81",
   513 => x"0a51ae8d",
   514 => x"3f0b0b80",
   515 => x"ecec51ae",
   516 => x"843f0b0b",
   517 => x"80ed9451",
   518 => x"adfb3f80",
   519 => x"e451afbf",
   520 => x"3f0b0b80",
   521 => x"eda851ad",
   522 => x"ec3f0b0b",
   523 => x"80edb051",
   524 => x"ade33f0b",
   525 => x"0b80edbc",
   526 => x"51adda3f",
   527 => x"823d0d04",
   528 => x"ff893f8b",
   529 => x"953f800b",
   530 => x"b00c04fe",
   531 => x"3d0d80fc",
   532 => x"ec089811",
   533 => x"0870842a",
   534 => x"70810651",
   535 => x"53535370",
   536 => x"802e8d38",
   537 => x"71ef0698",
   538 => x"140c810b",
   539 => x"818cc434",
   540 => x"843d0d04",
   541 => x"803d0d0b",
   542 => x"0b80edc4",
   543 => x"51ad963f",
   544 => x"8a51acf7",
   545 => x"3f800bb0",
   546 => x"0c823d0d",
   547 => x"04f93d0d",
   548 => x"81518994",
   549 => x"3fb00855",
   550 => x"8251898c",
   551 => x"3f74b008",
   552 => x"075399cc",
   553 => x"57fce297",
   554 => x"f6805872",
   555 => x"802e9038",
   556 => x"74755457",
   557 => x"80548077",
   558 => x"0774b008",
   559 => x"07595776",
   560 => x"5177529b",
   561 => x"fa3f72b0",
   562 => x"0c893d0d",
   563 => x"04fb3d0d",
   564 => x"815187a2",
   565 => x"3fb00856",
   566 => x"81538252",
   567 => x"8051a5a8",
   568 => x"3f80fcc8",
   569 => x"08558975",
   570 => x"0c80fce8",
   571 => x"08841108",
   572 => x"70810a07",
   573 => x"84130c55",
   574 => x"557551af",
   575 => x"d93f80fc",
   576 => x"e8088411",
   577 => x"0870fe0a",
   578 => x"0684130c",
   579 => x"55558153",
   580 => x"82528051",
   581 => x"a4f23f80",
   582 => x"fcc80855",
   583 => x"89750c80",
   584 => x"fce80884",
   585 => x"11087081",
   586 => x"0a078413",
   587 => x"0c555575",
   588 => x"51afa33f",
   589 => x"80fce808",
   590 => x"84110870",
   591 => x"fe0a0684",
   592 => x"130c5555",
   593 => x"ff9239fe",
   594 => x"3d0d8151",
   595 => x"86a83f80",
   596 => x"fce80884",
   597 => x"11087081",
   598 => x"0a078413",
   599 => x"0c5353b0",
   600 => x"0851aef2",
   601 => x"3f80fce8",
   602 => x"08841108",
   603 => x"70fe0a06",
   604 => x"7084140c",
   605 => x"b00c5353",
   606 => x"843d0d04",
   607 => x"fc3d0d80",
   608 => x"fce80870",
   609 => x"08810a06",
   610 => x"818cc00c",
   611 => x"54af913f",
   612 => x"afb53f8a",
   613 => x"c53f938c",
   614 => x"3f80fcec",
   615 => x"08981108",
   616 => x"70880798",
   617 => x"130c5555",
   618 => x"818cc008",
   619 => x"80d53888",
   620 => x"800b81a5",
   621 => x"900cfc93",
   622 => x"3f818cc0",
   623 => x"08802e80",
   624 => x"d3388153",
   625 => x"82528051",
   626 => x"a3be3f80",
   627 => x"fcc80855",
   628 => x"89750c80",
   629 => x"fce80884",
   630 => x"11087081",
   631 => x"0a078413",
   632 => x"0c555580",
   633 => x"51adef3f",
   634 => x"80fce808",
   635 => x"84110870",
   636 => x"fe0a0684",
   637 => x"130c5555",
   638 => x"80fcc808",
   639 => x"5580750c",
   640 => x"b0ab3fbd",
   641 => x"e50b81a5",
   642 => x"900cfbbf",
   643 => x"3f818cc0",
   644 => x"08ffaf38",
   645 => x"80c3930b",
   646 => x"81a5900c",
   647 => x"f5b63f81",
   648 => x"53825280",
   649 => x"51a2e13f",
   650 => x"80fcc808",
   651 => x"5589750c",
   652 => x"80fce808",
   653 => x"84110870",
   654 => x"810a0784",
   655 => x"130c5555",
   656 => x"8051ad92",
   657 => x"3f80fce8",
   658 => x"08841108",
   659 => x"70fe0a06",
   660 => x"84130c55",
   661 => x"5580fcc8",
   662 => x"08558075",
   663 => x"0cafce3f",
   664 => x"800b81a4",
   665 => x"ac34800b",
   666 => x"81a4a834",
   667 => x"800b81a4",
   668 => x"b00c04fc",
   669 => x"3d0d81a4",
   670 => x"a8335372",
   671 => x"a72680c5",
   672 => x"38765272",
   673 => x"10101073",
   674 => x"1005818c",
   675 => x"c80551b4",
   676 => x"b73f7752",
   677 => x"81a4a833",
   678 => x"70902971",
   679 => x"31701010",
   680 => x"818fd805",
   681 => x"535654b4",
   682 => x"9f3f81a4",
   683 => x"a8337010",
   684 => x"1081a2b8",
   685 => x"057a710c",
   686 => x"54810553",
   687 => x"7281a4a8",
   688 => x"34863d0d",
   689 => x"0480eddc",
   690 => x"51a8ca3f",
   691 => x"863d0d04",
   692 => x"803d0d80",
   693 => x"edf851a8",
   694 => x"bc3f823d",
   695 => x"0d04fe3d",
   696 => x"0d81a4b0",
   697 => x"08537285",
   698 => x"38843d0d",
   699 => x"04722db0",
   700 => x"0853800b",
   701 => x"81a4b00c",
   702 => x"b0088c38",
   703 => x"80edf851",
   704 => x"a8933f84",
   705 => x"3d0d0480",
   706 => x"f9a851a8",
   707 => x"883f7283",
   708 => x"ffff26aa",
   709 => x"3881ff73",
   710 => x"27963872",
   711 => x"529051a8",
   712 => x"973f8a51",
   713 => x"a7d53f80",
   714 => x"edf851a7",
   715 => x"e83fd439",
   716 => x"72528851",
   717 => x"a8823f8a",
   718 => x"51a7c03f",
   719 => x"ea397252",
   720 => x"a051a7f4",
   721 => x"3f8a51a7",
   722 => x"b23fdc39",
   723 => x"fa3d0d02",
   724 => x"a3053356",
   725 => x"758d2e80",
   726 => x"f4387588",
   727 => x"32703077",
   728 => x"80ff3270",
   729 => x"30728025",
   730 => x"71802507",
   731 => x"54515658",
   732 => x"55749538",
   733 => x"9f76278c",
   734 => x"3881a4ac",
   735 => x"335580ce",
   736 => x"7527ae38",
   737 => x"883d0d04",
   738 => x"81a4ac33",
   739 => x"5675802e",
   740 => x"f3388851",
   741 => x"a6e53fa0",
   742 => x"51a6e03f",
   743 => x"8851a6db",
   744 => x"3f81a4ac",
   745 => x"33ff0557",
   746 => x"7681a4ac",
   747 => x"34883d0d",
   748 => x"047551a6",
   749 => x"c63f81a4",
   750 => x"ac338111",
   751 => x"55577381",
   752 => x"a4ac3475",
   753 => x"81a3d818",
   754 => x"34883d0d",
   755 => x"048a51a6",
   756 => x"aa3f81a4",
   757 => x"ac338111",
   758 => x"56547481",
   759 => x"a4ac3480",
   760 => x"0b81a3d8",
   761 => x"15348056",
   762 => x"800b81a3",
   763 => x"d8173356",
   764 => x"5474a02e",
   765 => x"83388154",
   766 => x"74802e90",
   767 => x"3873802e",
   768 => x"8b388116",
   769 => x"7081ff06",
   770 => x"5757dd39",
   771 => x"75802ebf",
   772 => x"38800b81",
   773 => x"a4a83355",
   774 => x"55747427",
   775 => x"ab387357",
   776 => x"74101010",
   777 => x"75100576",
   778 => x"5481a3d8",
   779 => x"53818cc8",
   780 => x"0551b2e0",
   781 => x"3fb00880",
   782 => x"2ea63881",
   783 => x"157081ff",
   784 => x"06565476",
   785 => x"7526d938",
   786 => x"80edfc51",
   787 => x"a5c73f80",
   788 => x"edf851a5",
   789 => x"c03f800b",
   790 => x"81a4ac34",
   791 => x"883d0d04",
   792 => x"74101081",
   793 => x"a2b80570",
   794 => x"0881a4b0",
   795 => x"0c56800b",
   796 => x"81a4ac34",
   797 => x"e739f73d",
   798 => x"0d02af05",
   799 => x"3359800b",
   800 => x"81a3d833",
   801 => x"81a3d859",
   802 => x"555673a0",
   803 => x"2e098106",
   804 => x"96388116",
   805 => x"7081ff06",
   806 => x"81a3d811",
   807 => x"70335359",
   808 => x"575473a0",
   809 => x"2eec3880",
   810 => x"58777927",
   811 => x"80ea3880",
   812 => x"77335654",
   813 => x"74742e83",
   814 => x"38815474",
   815 => x"a02e9a38",
   816 => x"7380c538",
   817 => x"74a02e91",
   818 => x"38811870",
   819 => x"81ff0659",
   820 => x"55787826",
   821 => x"da3880c0",
   822 => x"39811670",
   823 => x"81ff0681",
   824 => x"a3d81170",
   825 => x"33575257",
   826 => x"5773a02e",
   827 => x"098106d9",
   828 => x"38811670",
   829 => x"81ff0681",
   830 => x"a3d81170",
   831 => x"33575257",
   832 => x"5773a02e",
   833 => x"d438c239",
   834 => x"81167081",
   835 => x"ff0681a3",
   836 => x"d8115957",
   837 => x"55ff9839",
   838 => x"80538b3d",
   839 => x"fc055276",
   840 => x"51b5b63f",
   841 => x"8b3d0d04",
   842 => x"f73d0d02",
   843 => x"af053359",
   844 => x"800b81a3",
   845 => x"d83381a3",
   846 => x"d8595556",
   847 => x"73a02e09",
   848 => x"81069638",
   849 => x"81167081",
   850 => x"ff0681a3",
   851 => x"d8117033",
   852 => x"53595754",
   853 => x"73a02eec",
   854 => x"38805877",
   855 => x"792780ea",
   856 => x"38807733",
   857 => x"56547474",
   858 => x"2e833881",
   859 => x"5474a02e",
   860 => x"9a387380",
   861 => x"c53874a0",
   862 => x"2e913881",
   863 => x"187081ff",
   864 => x"06595578",
   865 => x"7826da38",
   866 => x"80c03981",
   867 => x"167081ff",
   868 => x"0681a3d8",
   869 => x"11703357",
   870 => x"52575773",
   871 => x"a02e0981",
   872 => x"06d93881",
   873 => x"167081ff",
   874 => x"0681a3d8",
   875 => x"11703357",
   876 => x"52575773",
   877 => x"a02ed438",
   878 => x"c2398116",
   879 => x"7081ff06",
   880 => x"81a3d811",
   881 => x"595755ff",
   882 => x"98399053",
   883 => x"8b3dfc05",
   884 => x"527651b7",
   885 => x"a13f8b3d",
   886 => x"0d04fc3d",
   887 => x"0d8a51a2",
   888 => x"9a3f80ee",
   889 => x"9051a2ad",
   890 => x"3f800b81",
   891 => x"a4a83353",
   892 => x"53727227",
   893 => x"80f53872",
   894 => x"10101073",
   895 => x"1005818c",
   896 => x"c8057052",
   897 => x"54a28e3f",
   898 => x"72842b70",
   899 => x"7431822b",
   900 => x"818fd811",
   901 => x"33515355",
   902 => x"71802eb7",
   903 => x"387351ae",
   904 => x"943fb008",
   905 => x"81ff0652",
   906 => x"71892693",
   907 => x"38a051a1",
   908 => x"ca3f8112",
   909 => x"7081ff06",
   910 => x"53548972",
   911 => x"27ef3880",
   912 => x"eea851a1",
   913 => x"d03f7473",
   914 => x"31822b81",
   915 => x"8fd80551",
   916 => x"a1c33f8a",
   917 => x"51a1a43f",
   918 => x"81137081",
   919 => x"ff0681a4",
   920 => x"a8335454",
   921 => x"55717326",
   922 => x"ff8d388a",
   923 => x"51a18c3f",
   924 => x"81a4a833",
   925 => x"b00c863d",
   926 => x"0d04fe3d",
   927 => x"0d81a588",
   928 => x"22ff0551",
   929 => x"7081a588",
   930 => x"237083ff",
   931 => x"ff065170",
   932 => x"80c43881",
   933 => x"a58c3351",
   934 => x"7081ff2e",
   935 => x"b9387010",
   936 => x"101081a4",
   937 => x"b8055271",
   938 => x"3381a58c",
   939 => x"34fe7234",
   940 => x"81a58c33",
   941 => x"70101010",
   942 => x"81a4b805",
   943 => x"52538211",
   944 => x"2281a588",
   945 => x"23841208",
   946 => x"53722d81",
   947 => x"a5882251",
   948 => x"70802eff",
   949 => x"be38843d",
   950 => x"0d04ff3d",
   951 => x"0d8a5271",
   952 => x"10101081",
   953 => x"a4b00551",
   954 => x"fe7134ff",
   955 => x"127081ff",
   956 => x"06535171",
   957 => x"ea38ff0b",
   958 => x"81a58c34",
   959 => x"833d0d04",
   960 => x"fe3d0d02",
   961 => x"93053302",
   962 => x"84059705",
   963 => x"33545271",
   964 => x"842e80d1",
   965 => x"38718424",
   966 => x"91387181",
   967 => x"2eac3880",
   968 => x"eeac519f",
   969 => x"f03f843d",
   970 => x"0d047180",
   971 => x"d52e0981",
   972 => x"06ed3880",
   973 => x"eeb8519f",
   974 => x"dc3f728c",
   975 => x"26b33872",
   976 => x"101080f3",
   977 => x"ac055271",
   978 => x"080480ee",
   979 => x"c4519fc5",
   980 => x"3ffa1352",
   981 => x"7180db26",
   982 => x"98387110",
   983 => x"1080f3e0",
   984 => x"05527108",
   985 => x"0480eed0",
   986 => x"519faa3f",
   987 => x"728f2e8c",
   988 => x"3880eedc",
   989 => x"519f9e3f",
   990 => x"843d0d04",
   991 => x"80eeec51",
   992 => x"9f933f84",
   993 => x"3d0d0480",
   994 => x"ef84519f",
   995 => x"883f843d",
   996 => x"0d0480ef",
   997 => x"94519efd",
   998 => x"3f843d0d",
   999 => x"0480efac",
  1000 => x"519ef23f",
  1001 => x"843d0d04",
  1002 => x"80efbc51",
  1003 => x"9ee73f84",
  1004 => x"3d0d0480",
  1005 => x"efdc519e",
  1006 => x"dc3f843d",
  1007 => x"0d0480ef",
  1008 => x"f8519ed1",
  1009 => x"3f843d0d",
  1010 => x"0480f094",
  1011 => x"519ec63f",
  1012 => x"843d0d04",
  1013 => x"80f0a851",
  1014 => x"9ebb3f84",
  1015 => x"3d0d0480",
  1016 => x"f0c4519e",
  1017 => x"b03f843d",
  1018 => x"0d0480f0",
  1019 => x"d4519ea5",
  1020 => x"3f843d0d",
  1021 => x"0480f0e4",
  1022 => x"519e9a3f",
  1023 => x"843d0d04",
  1024 => x"80f18451",
  1025 => x"9e8f3f84",
  1026 => x"3d0d0480",
  1027 => x"f198519e",
  1028 => x"843f843d",
  1029 => x"0d0480f1",
  1030 => x"b4519df9",
  1031 => x"3f843d0d",
  1032 => x"0480f1cc",
  1033 => x"519dee3f",
  1034 => x"843d0d04",
  1035 => x"80f1e051",
  1036 => x"9de33f84",
  1037 => x"3d0d0480",
  1038 => x"f1f0519d",
  1039 => x"d83f843d",
  1040 => x"0d0480f2",
  1041 => x"84519dcd",
  1042 => x"3f843d0d",
  1043 => x"0480f294",
  1044 => x"519dc23f",
  1045 => x"843d0d04",
  1046 => x"80f2ac51",
  1047 => x"9db73f84",
  1048 => x"3d0d0480",
  1049 => x"f2c0519d",
  1050 => x"ac3f843d",
  1051 => x"0d0480f2",
  1052 => x"d0519da1",
  1053 => x"3f843d0d",
  1054 => x"04f73d0d",
  1055 => x"02b30533",
  1056 => x"7c7008c0",
  1057 => x"80800659",
  1058 => x"545a8056",
  1059 => x"75832b77",
  1060 => x"07bfe080",
  1061 => x"07707084",
  1062 => x"05520871",
  1063 => x"088c2abf",
  1064 => x"fe800679",
  1065 => x"0771982a",
  1066 => x"728c2a9f",
  1067 => x"ff067385",
  1068 => x"2a708f06",
  1069 => x"759f0656",
  1070 => x"51585d58",
  1071 => x"52555874",
  1072 => x"8d388116",
  1073 => x"568f7627",
  1074 => x"c3388b3d",
  1075 => x"0d0480f2",
  1076 => x"e8519cc1",
  1077 => x"3f75519e",
  1078 => x"863f8452",
  1079 => x"b008519f",
  1080 => x"c73f80f2",
  1081 => x"f4519cad",
  1082 => x"3f745288",
  1083 => x"519cc93f",
  1084 => x"8452b008",
  1085 => x"519fb13f",
  1086 => x"80f2fc51",
  1087 => x"9c973f78",
  1088 => x"5290519c",
  1089 => x"b33f8652",
  1090 => x"b008519f",
  1091 => x"9b3f80f3",
  1092 => x"84519c81",
  1093 => x"3f72519d",
  1094 => x"c63f8452",
  1095 => x"b008519f",
  1096 => x"873f80f3",
  1097 => x"8c519bed",
  1098 => x"3f73519d",
  1099 => x"b23f8452",
  1100 => x"b008519e",
  1101 => x"f33f80f3",
  1102 => x"94519bd9",
  1103 => x"3f7752a0",
  1104 => x"519bf53f",
  1105 => x"8a52b008",
  1106 => x"519edd3f",
  1107 => x"7992388a",
  1108 => x"519ba83f",
  1109 => x"8116568f",
  1110 => x"7627feb0",
  1111 => x"38feeb39",
  1112 => x"7881ff06",
  1113 => x"527451fb",
  1114 => x"973f8a51",
  1115 => x"9b8d3fe4",
  1116 => x"39f83d0d",
  1117 => x"02ab0533",
  1118 => x"59805675",
  1119 => x"852be090",
  1120 => x"11e08012",
  1121 => x"0870982a",
  1122 => x"718c2a9f",
  1123 => x"ff067285",
  1124 => x"2a708f06",
  1125 => x"749f0655",
  1126 => x"51585b53",
  1127 => x"56595574",
  1128 => x"802e81a1",
  1129 => x"3875bf26",
  1130 => x"81a93880",
  1131 => x"f39c519a",
  1132 => x"e43f7551",
  1133 => x"9ca93f86",
  1134 => x"52b00851",
  1135 => x"9dea3f80",
  1136 => x"f2f4519a",
  1137 => x"d03f7452",
  1138 => x"88519aec",
  1139 => x"3f8452b0",
  1140 => x"08519dd4",
  1141 => x"3f80f2fc",
  1142 => x"519aba3f",
  1143 => x"76529051",
  1144 => x"9ad63f86",
  1145 => x"52b00851",
  1146 => x"9dbe3f80",
  1147 => x"f384519a",
  1148 => x"a43f7251",
  1149 => x"9be93f84",
  1150 => x"52b00851",
  1151 => x"9daa3f80",
  1152 => x"f38c519a",
  1153 => x"903f7351",
  1154 => x"9bd53f84",
  1155 => x"52b00851",
  1156 => x"9d963f80",
  1157 => x"f3945199",
  1158 => x"fc3f7708",
  1159 => x"c0808006",
  1160 => x"52a0519a",
  1161 => x"933f8a52",
  1162 => x"b008519c",
  1163 => x"fb3f7881",
  1164 => x"ac388a51",
  1165 => x"99c53f80",
  1166 => x"5374812e",
  1167 => x"81d93876",
  1168 => x"862e81b5",
  1169 => x"38811656",
  1170 => x"80ff7627",
  1171 => x"fead388a",
  1172 => x"3d0d0480",
  1173 => x"f3a45199",
  1174 => x"bc3fc016",
  1175 => x"519b803f",
  1176 => x"8652b008",
  1177 => x"519cc13f",
  1178 => x"80f2f451",
  1179 => x"99a73f74",
  1180 => x"52885199",
  1181 => x"c33f8452",
  1182 => x"b008519c",
  1183 => x"ab3f80f2",
  1184 => x"fc519991",
  1185 => x"3f765290",
  1186 => x"5199ad3f",
  1187 => x"8652b008",
  1188 => x"519c953f",
  1189 => x"80f38451",
  1190 => x"98fb3f72",
  1191 => x"519ac03f",
  1192 => x"8452b008",
  1193 => x"519c813f",
  1194 => x"80f38c51",
  1195 => x"98e73f73",
  1196 => x"519aac3f",
  1197 => x"8452b008",
  1198 => x"519bed3f",
  1199 => x"80f39451",
  1200 => x"98d33f77",
  1201 => x"08c08080",
  1202 => x"0652a051",
  1203 => x"98ea3f8a",
  1204 => x"52b00851",
  1205 => x"9bd23f78",
  1206 => x"802efed6",
  1207 => x"387681ff",
  1208 => x"06527451",
  1209 => x"f89a3f8a",
  1210 => x"5198903f",
  1211 => x"80537481",
  1212 => x"2e098106",
  1213 => x"fec9389f",
  1214 => x"39728106",
  1215 => x"5776802e",
  1216 => x"fec33878",
  1217 => x"527751fa",
  1218 => x"f03f8116",
  1219 => x"5680ff76",
  1220 => x"27fce838",
  1221 => x"feb93974",
  1222 => x"5376862e",
  1223 => x"098106fe",
  1224 => x"a438d639",
  1225 => x"803d0d80",
  1226 => x"fce40851",
  1227 => x"b1710c81",
  1228 => x"800b8412",
  1229 => x"0c823d0d",
  1230 => x"04fe3d0d",
  1231 => x"74028405",
  1232 => x"97053302",
  1233 => x"88059b05",
  1234 => x"3388130c",
  1235 => x"8c120c53",
  1236 => x"8c130870",
  1237 => x"812a8106",
  1238 => x"515271f4",
  1239 => x"388c1308",
  1240 => x"7081ff06",
  1241 => x"b00c5184",
  1242 => x"3d0d04fb",
  1243 => x"3d0d800b",
  1244 => x"80f6d052",
  1245 => x"56979e3f",
  1246 => x"75557410",
  1247 => x"5381d052",
  1248 => x"80fce408",
  1249 => x"51ffb23f",
  1250 => x"b008872a",
  1251 => x"70810651",
  1252 => x"5473802e",
  1253 => x"99388115",
  1254 => x"7081ff06",
  1255 => x"70982b52",
  1256 => x"56547380",
  1257 => x"25d43875",
  1258 => x"b00c873d",
  1259 => x"0d0480f6",
  1260 => x"dc5196e1",
  1261 => x"3f745288",
  1262 => x"5196fd3f",
  1263 => x"80f6e851",
  1264 => x"96d33f81",
  1265 => x"167083ff",
  1266 => x"ff068117",
  1267 => x"7081ff06",
  1268 => x"70982b52",
  1269 => x"58525754",
  1270 => x"738025ff",
  1271 => x"9d38c839",
  1272 => x"f33d0d7f",
  1273 => x"02840580",
  1274 => x"c3053302",
  1275 => x"880580c6",
  1276 => x"052280f6",
  1277 => x"f8545b55",
  1278 => x"58969a3f",
  1279 => x"785197df",
  1280 => x"3f80f784",
  1281 => x"51968e3f",
  1282 => x"73528851",
  1283 => x"96aa3f80",
  1284 => x"ecb05196",
  1285 => x"803f8057",
  1286 => x"76792781",
  1287 => x"91387310",
  1288 => x"8e3d5c5a",
  1289 => x"79538190",
  1290 => x"527751fe",
  1291 => x"8c3f7688",
  1292 => x"2a539052",
  1293 => x"7751fe81",
  1294 => x"3f7681ff",
  1295 => x"06539052",
  1296 => x"7751fdf5",
  1297 => x"3f811a53",
  1298 => x"81905277",
  1299 => x"51fdea3f",
  1300 => x"805380e0",
  1301 => x"527751fd",
  1302 => x"e03fb008",
  1303 => x"872a8106",
  1304 => x"54738a38",
  1305 => x"88180870",
  1306 => x"81ff065d",
  1307 => x"567b81ff",
  1308 => x"0680f9a8",
  1309 => x"5256959d",
  1310 => x"3f755288",
  1311 => x"5195b93f",
  1312 => x"80eed851",
  1313 => x"958f3fe0",
  1314 => x"165480df",
  1315 => x"7427b638",
  1316 => x"76870670",
  1317 => x"1c5755a0",
  1318 => x"76347487",
  1319 => x"2eb93881",
  1320 => x"177083ff",
  1321 => x"ff065855",
  1322 => x"787726fe",
  1323 => x"f73880e0",
  1324 => x"0b8c190c",
  1325 => x"8c180870",
  1326 => x"812a8106",
  1327 => x"585a76f4",
  1328 => x"388f3d0d",
  1329 => x"04768706",
  1330 => x"701c5555",
  1331 => x"75743474",
  1332 => x"872e0981",
  1333 => x"06c9387a",
  1334 => x"5194ba3f",
  1335 => x"8a51949b",
  1336 => x"3f811770",
  1337 => x"83ffff06",
  1338 => x"58557877",
  1339 => x"26feb538",
  1340 => x"ffbc39fb",
  1341 => x"3d0d8151",
  1342 => x"eefc3f82",
  1343 => x"51f0a93f",
  1344 => x"b00881ff",
  1345 => x"06568351",
  1346 => x"eeec3fb0",
  1347 => x"0883ffff",
  1348 => x"0680fce4",
  1349 => x"08565473",
  1350 => x"84388180",
  1351 => x"54735375",
  1352 => x"527451fd",
  1353 => x"bb3f73b0",
  1354 => x"0c873d0d",
  1355 => x"04fb3d0d",
  1356 => x"8151eff4",
  1357 => x"3fb00853",
  1358 => x"8251efec",
  1359 => x"3fb00856",
  1360 => x"b0088338",
  1361 => x"905672fc",
  1362 => x"06557581",
  1363 => x"2e80f138",
  1364 => x"80547376",
  1365 => x"27aa3873",
  1366 => x"83065372",
  1367 => x"802eae38",
  1368 => x"80f9a851",
  1369 => x"93af3f74",
  1370 => x"70840556",
  1371 => x"0852a051",
  1372 => x"93c63fa0",
  1373 => x"5193843f",
  1374 => x"81145475",
  1375 => x"7426d838",
  1376 => x"8a5192f7",
  1377 => x"3f800bb0",
  1378 => x"0c873d0d",
  1379 => x"0480f7a0",
  1380 => x"5193823f",
  1381 => x"7452a051",
  1382 => x"939e3f80",
  1383 => x"f8e85192",
  1384 => x"f43f80f9",
  1385 => x"a85192ed",
  1386 => x"3f747084",
  1387 => x"05560852",
  1388 => x"a0519384",
  1389 => x"3fa05192",
  1390 => x"c23f8114",
  1391 => x"54ffbc39",
  1392 => x"80f9a851",
  1393 => x"92cf3f74",
  1394 => x"0852a051",
  1395 => x"92ea3f8a",
  1396 => x"5192a83f",
  1397 => x"800bb00c",
  1398 => x"873d0d04",
  1399 => x"fc3d0d81",
  1400 => x"51eec53f",
  1401 => x"b0085282",
  1402 => x"51ed8b3f",
  1403 => x"b00881ff",
  1404 => x"06725653",
  1405 => x"83547280",
  1406 => x"2ea13873",
  1407 => x"51eea93f",
  1408 => x"81147081",
  1409 => x"ff06ff15",
  1410 => x"7081ff06",
  1411 => x"b0087970",
  1412 => x"84055b0c",
  1413 => x"56525552",
  1414 => x"72e13872",
  1415 => x"b00c863d",
  1416 => x"0d04803d",
  1417 => x"0d8c5191",
  1418 => x"d23f800b",
  1419 => x"b00c823d",
  1420 => x"0d04803d",
  1421 => x"0d80fcf4",
  1422 => x"0851f8bb",
  1423 => x"9586a171",
  1424 => x"0c810bb0",
  1425 => x"0c823d0d",
  1426 => x"04803d0d",
  1427 => x"8151eca6",
  1428 => x"3fb00881",
  1429 => x"ff0651f6",
  1430 => x"983f800b",
  1431 => x"b00c823d",
  1432 => x"0d04ff3d",
  1433 => x"0d80fcc0",
  1434 => x"08a01108",
  1435 => x"7080ff0a",
  1436 => x"06a0130c",
  1437 => x"5252bbc8",
  1438 => x"80800ba0",
  1439 => x"130c833d",
  1440 => x"0d04ff3d",
  1441 => x"0d028f05",
  1442 => x"3370982b",
  1443 => x"80fcc008",
  1444 => x"52b0120c",
  1445 => x"51833d0d",
  1446 => x"04ff3d0d",
  1447 => x"80fcc008",
  1448 => x"52a41208",
  1449 => x"70892a70",
  1450 => x"81065151",
  1451 => x"5170802e",
  1452 => x"f038b412",
  1453 => x"0870902a",
  1454 => x"b00c5183",
  1455 => x"3d0d04f8",
  1456 => x"3d0d7a7c",
  1457 => x"5755ff9a",
  1458 => x"3f80fce8",
  1459 => x"08841108",
  1460 => x"82808007",
  1461 => x"84120c84",
  1462 => x"1108fdff",
  1463 => x"ff068412",
  1464 => x"0c841108",
  1465 => x"81808007",
  1466 => x"84120c84",
  1467 => x"1108feff",
  1468 => x"ff068412",
  1469 => x"0c53900b",
  1470 => x"893d3494",
  1471 => x"0284059d",
  1472 => x"05348002",
  1473 => x"84059e05",
  1474 => x"3480e102",
  1475 => x"84059f05",
  1476 => x"34883d80",
  1477 => x"fcc00854",
  1478 => x"57a41308",
  1479 => x"70882a81",
  1480 => x"06515271",
  1481 => x"802ef238",
  1482 => x"8751fed6",
  1483 => x"3f800b80",
  1484 => x"f7ab3353",
  1485 => x"53727227",
  1486 => x"99387154",
  1487 => x"76137033",
  1488 => x"5252febe",
  1489 => x"3f811370",
  1490 => x"81ff0654",
  1491 => x"52737326",
  1492 => x"eb38fec5",
  1493 => x"3f800b80",
  1494 => x"f7ab3353",
  1495 => x"53727227",
  1496 => x"93387154",
  1497 => x"feb33f81",
  1498 => x"137081ff",
  1499 => x"06545273",
  1500 => x"7326f138",
  1501 => x"74882a54",
  1502 => x"73893d34",
  1503 => x"74028405",
  1504 => x"9d053474",
  1505 => x"882b7698",
  1506 => x"2a075271",
  1507 => x"0284059e",
  1508 => x"05347490",
  1509 => x"2b76902a",
  1510 => x"07547302",
  1511 => x"84059f05",
  1512 => x"3474982b",
  1513 => x"76882a07",
  1514 => x"53728a3d",
  1515 => x"34750284",
  1516 => x"05a10534",
  1517 => x"80fcc008",
  1518 => x"53a41308",
  1519 => x"70882a81",
  1520 => x"06565274",
  1521 => x"802ef238",
  1522 => x"8251fdb6",
  1523 => x"3f800b80",
  1524 => x"f7a63353",
  1525 => x"53727227",
  1526 => x"99387154",
  1527 => x"76137033",
  1528 => x"5256fd9e",
  1529 => x"3f811370",
  1530 => x"81ff0654",
  1531 => x"55737326",
  1532 => x"eb38fda5",
  1533 => x"3f800b80",
  1534 => x"f7a63353",
  1535 => x"53727227",
  1536 => x"93387154",
  1537 => x"fd933f81",
  1538 => x"137081ff",
  1539 => x"06545273",
  1540 => x"7326f138",
  1541 => x"8a0b893d",
  1542 => x"34ff8c02",
  1543 => x"84059d05",
  1544 => x"3480fcc0",
  1545 => x"0853a413",
  1546 => x"0870882a",
  1547 => x"81065556",
  1548 => x"73802ef2",
  1549 => x"388851fc",
  1550 => x"c93f800b",
  1551 => x"80f7ac33",
  1552 => x"53537272",
  1553 => x"27993871",
  1554 => x"54761370",
  1555 => x"335255fc",
  1556 => x"b13f8113",
  1557 => x"7081ff06",
  1558 => x"54527373",
  1559 => x"26eb38fc",
  1560 => x"b83f800b",
  1561 => x"80f7ac33",
  1562 => x"53537272",
  1563 => x"27933871",
  1564 => x"54fca63f",
  1565 => x"81137081",
  1566 => x"ff065456",
  1567 => x"737326f1",
  1568 => x"388a0b89",
  1569 => x"3d34ff8c",
  1570 => x"0284059d",
  1571 => x"053480fc",
  1572 => x"c00853a4",
  1573 => x"13087088",
  1574 => x"2a810655",
  1575 => x"5573802e",
  1576 => x"f2388951",
  1577 => x"fbdc3f80",
  1578 => x"0b80f7ad",
  1579 => x"33535372",
  1580 => x"72279938",
  1581 => x"71547613",
  1582 => x"70335252",
  1583 => x"fbc43f81",
  1584 => x"137081ff",
  1585 => x"06545673",
  1586 => x"7326eb38",
  1587 => x"fbcb3f80",
  1588 => x"0b80f7ad",
  1589 => x"33535372",
  1590 => x"72279338",
  1591 => x"7154fbb9",
  1592 => x"3f811370",
  1593 => x"81ff0654",
  1594 => x"57737326",
  1595 => x"f13880fc",
  1596 => x"e8088411",
  1597 => x"0880c080",
  1598 => x"0784120c",
  1599 => x"841108ff",
  1600 => x"bfff0684",
  1601 => x"120c5480",
  1602 => x"0bb00c8a",
  1603 => x"3d0d04f8",
  1604 => x"3d0d02ab",
  1605 => x"0533893d",
  1606 => x"80fcc008",
  1607 => x"565856a4",
  1608 => x"14087088",
  1609 => x"2a810651",
  1610 => x"5372802e",
  1611 => x"f2387581",
  1612 => x"800751fa",
  1613 => x"cd3f800b",
  1614 => x"80f7a417",
  1615 => x"33545473",
  1616 => x"73279538",
  1617 => x"72558051",
  1618 => x"fab83f81",
  1619 => x"147081ff",
  1620 => x"06555374",
  1621 => x"7426ef38",
  1622 => x"fabf3f80",
  1623 => x"0b80f7a4",
  1624 => x"17337081",
  1625 => x"ff065557",
  1626 => x"54737327",
  1627 => x"9a387255",
  1628 => x"761453fa",
  1629 => x"a43fb008",
  1630 => x"73348114",
  1631 => x"7081ff06",
  1632 => x"55537474",
  1633 => x"26ea3875",
  1634 => x"81ff0680",
  1635 => x"f9a85255",
  1636 => x"8b833f80",
  1637 => x"54737527",
  1638 => x"99387317",
  1639 => x"70335353",
  1640 => x"88518b94",
  1641 => x"3f811470",
  1642 => x"81ff0655",
  1643 => x"56747426",
  1644 => x"e9388a51",
  1645 => x"8ac53f8a",
  1646 => x"3d0d04fe",
  1647 => x"3d0d80fc",
  1648 => x"e8088411",
  1649 => x"08708180",
  1650 => x"80078413",
  1651 => x"0c548411",
  1652 => x"0870feff",
  1653 => x"ff068413",
  1654 => x"0c5452f9",
  1655 => x"853f80f7",
  1656 => x"b0518ab1",
  1657 => x"3f8751fe",
  1658 => x"a63f80f7",
  1659 => x"c0518aa5",
  1660 => x"3f8251fe",
  1661 => x"9a3f80f7",
  1662 => x"d0518a99",
  1663 => x"3f8551fe",
  1664 => x"8e3f80f7",
  1665 => x"e0518a8d",
  1666 => x"3f8651fe",
  1667 => x"823f80f7",
  1668 => x"f0518a81",
  1669 => x"3f8851fd",
  1670 => x"f63f80f8",
  1671 => x"805189f5",
  1672 => x"3f8951fd",
  1673 => x"ea3f800b",
  1674 => x"b00c843d",
  1675 => x"0d04fe3d",
  1676 => x"0d80fce8",
  1677 => x"08841108",
  1678 => x"820a0784",
  1679 => x"120c7008",
  1680 => x"70902a84",
  1681 => x"130870fd",
  1682 => x"0a068415",
  1683 => x"0c5481ff",
  1684 => x"ff06b00c",
  1685 => x"5353843d",
  1686 => x"0d04ff3d",
  1687 => x"0d80fcc8",
  1688 => x"08700870",
  1689 => x"81ff0651",
  1690 => x"51527189",
  1691 => x"268c3871",
  1692 => x"101080f9",
  1693 => x"d0055271",
  1694 => x"080480f8",
  1695 => x"90518995",
  1696 => x"3f8a5188",
  1697 => x"f63f800b",
  1698 => x"b00c833d",
  1699 => x"0d0480e8",
  1700 => x"ac518981",
  1701 => x"3f8a5188",
  1702 => x"e23f800b",
  1703 => x"b00c833d",
  1704 => x"0d0480f8",
  1705 => x"985188ed",
  1706 => x"3f8a5188",
  1707 => x"ce3f800b",
  1708 => x"b00c833d",
  1709 => x"0d0480f8",
  1710 => x"a05188d9",
  1711 => x"3f8a5188",
  1712 => x"ba3f800b",
  1713 => x"b00c833d",
  1714 => x"0d0480f8",
  1715 => x"ac5188c5",
  1716 => x"3f8a5188",
  1717 => x"a63f800b",
  1718 => x"b00c833d",
  1719 => x"0d0480f8",
  1720 => x"b45188b1",
  1721 => x"3f8a5188",
  1722 => x"923f800b",
  1723 => x"b00c833d",
  1724 => x"0d0480f8",
  1725 => x"bc51889d",
  1726 => x"3f8a5187",
  1727 => x"fe3f800b",
  1728 => x"b00c833d",
  1729 => x"0d0480f8",
  1730 => x"c4518889",
  1731 => x"3f8a5187",
  1732 => x"ea3f800b",
  1733 => x"b00c833d",
  1734 => x"0d0480f8",
  1735 => x"cc5187f5",
  1736 => x"3f8a5187",
  1737 => x"d63f800b",
  1738 => x"b00c833d",
  1739 => x"0d0480f8",
  1740 => x"d45187e1",
  1741 => x"3f8a5187",
  1742 => x"c23f800b",
  1743 => x"b00c833d",
  1744 => x"0d04fe3d",
  1745 => x"0d80fcc8",
  1746 => x"08841108",
  1747 => x"80f8dc53",
  1748 => x"545287c1",
  1749 => x"3f72822a",
  1750 => x"81065189",
  1751 => x"823f80f8",
  1752 => x"ec5187b1",
  1753 => x"3f72812a",
  1754 => x"81065188",
  1755 => x"f23f80f9",
  1756 => x"805187a1",
  1757 => x"3f728106",
  1758 => x"5188e43f",
  1759 => x"8a5186fb",
  1760 => x"3f72b00c",
  1761 => x"843d0d04",
  1762 => x"fe3d0d02",
  1763 => x"93053302",
  1764 => x"84059705",
  1765 => x"3380fcc8",
  1766 => x"08555351",
  1767 => x"80730c76",
  1768 => x"88140c70",
  1769 => x"832b7207",
  1770 => x"8c140c72",
  1771 => x"085170fb",
  1772 => x"3870b00c",
  1773 => x"843d0d04",
  1774 => x"fe3d0d80",
  1775 => x"f9945186",
  1776 => x"d43f80fc",
  1777 => x"c808a011",
  1778 => x"085353a0",
  1779 => x"5186e93f",
  1780 => x"80fcc808",
  1781 => x"a4110853",
  1782 => x"53a05186",
  1783 => x"db3f80f9",
  1784 => x"ac5186b1",
  1785 => x"3f80fcc8",
  1786 => x"08a81108",
  1787 => x"5353a051",
  1788 => x"86c63f80",
  1789 => x"fcc808ac",
  1790 => x"11085353",
  1791 => x"a05186b8",
  1792 => x"3f8a5185",
  1793 => x"f63f800b",
  1794 => x"b00c843d",
  1795 => x"0d04fc3d",
  1796 => x"0d80fcc8",
  1797 => x"089c1108",
  1798 => x"7081ff06",
  1799 => x"80f9c454",
  1800 => x"57535385",
  1801 => x"f03f7451",
  1802 => x"87b53f8a",
  1803 => x"5185cc3f",
  1804 => x"800bff16",
  1805 => x"55537274",
  1806 => x"25a23872",
  1807 => x"101080fc",
  1808 => x"c4080570",
  1809 => x"08525287",
  1810 => x"963f8a51",
  1811 => x"85ad3f81",
  1812 => x"137081ff",
  1813 => x"06545273",
  1814 => x"7324e038",
  1815 => x"74b00c86",
  1816 => x"3d0d04fd",
  1817 => x"3d0d8151",
  1818 => x"e08c3fb0",
  1819 => x"0881ff06",
  1820 => x"528251e1",
  1821 => x"b33fb008",
  1822 => x"81ff0653",
  1823 => x"8351e1a8",
  1824 => x"3f80fcc8",
  1825 => x"08548074",
  1826 => x"0cb00888",
  1827 => x"150c7183",
  1828 => x"2b73078c",
  1829 => x"150c7308",
  1830 => x"5271fb38",
  1831 => x"71b00c85",
  1832 => x"3d0d04ff",
  1833 => x"3d0d8151",
  1834 => x"dfcc3f80",
  1835 => x"fcc808b0",
  1836 => x"0890120c",
  1837 => x"5282720c",
  1838 => x"833d0d04",
  1839 => x"803d0d80",
  1840 => x"fcc80851",
  1841 => x"80710c70",
  1842 => x"b00c823d",
  1843 => x"0d04fd3d",
  1844 => x"0d800b80",
  1845 => x"fcc80854",
  1846 => x"5480730c",
  1847 => x"fecac090",
  1848 => x"860b8814",
  1849 => x"0c73832b",
  1850 => x"82078c14",
  1851 => x"0c720852",
  1852 => x"71fb3881",
  1853 => x"147081ff",
  1854 => x"065551a2",
  1855 => x"7427da38",
  1856 => x"71b00c85",
  1857 => x"3d0d04fd",
  1858 => x"3d0d800b",
  1859 => x"80fcc808",
  1860 => x"54548073",
  1861 => x"0c880a0b",
  1862 => x"88140c73",
  1863 => x"832b8107",
  1864 => x"8c140c72",
  1865 => x"085271fb",
  1866 => x"38811470",
  1867 => x"81ff0655",
  1868 => x"51a27427",
  1869 => x"dd3871b0",
  1870 => x"0c853d0d",
  1871 => x"04fe3d0d",
  1872 => x"8151deb2",
  1873 => x"3f80fcc8",
  1874 => x"08538073",
  1875 => x"0c810b88",
  1876 => x"140cb008",
  1877 => x"832b8ff8",
  1878 => x"06708207",
  1879 => x"8c150c52",
  1880 => x"72085271",
  1881 => x"fb388973",
  1882 => x"0c71b00c",
  1883 => x"843d0d04",
  1884 => x"d88a3f04",
  1885 => x"fb3d0d77",
  1886 => x"79555580",
  1887 => x"56757524",
  1888 => x"ab388074",
  1889 => x"249d3880",
  1890 => x"53735274",
  1891 => x"5180e13f",
  1892 => x"b0085475",
  1893 => x"802e8538",
  1894 => x"b0083054",
  1895 => x"73b00c87",
  1896 => x"3d0d0473",
  1897 => x"30768132",
  1898 => x"5754dc39",
  1899 => x"74305581",
  1900 => x"56738025",
  1901 => x"d238ec39",
  1902 => x"fa3d0d78",
  1903 => x"7a575580",
  1904 => x"57767524",
  1905 => x"a438759f",
  1906 => x"2c548153",
  1907 => x"75743274",
  1908 => x"31527451",
  1909 => x"9b3fb008",
  1910 => x"5476802e",
  1911 => x"8538b008",
  1912 => x"305473b0",
  1913 => x"0c883d0d",
  1914 => x"04743055",
  1915 => x"8157d739",
  1916 => x"fc3d0d76",
  1917 => x"78535481",
  1918 => x"53807473",
  1919 => x"26525572",
  1920 => x"802e9838",
  1921 => x"70802ea9",
  1922 => x"38807224",
  1923 => x"a4387110",
  1924 => x"73107572",
  1925 => x"26535452",
  1926 => x"72ea3873",
  1927 => x"51788338",
  1928 => x"745170b0",
  1929 => x"0c863d0d",
  1930 => x"0472812a",
  1931 => x"72812a53",
  1932 => x"5372802e",
  1933 => x"e6387174",
  1934 => x"26ef3873",
  1935 => x"72317574",
  1936 => x"0774812a",
  1937 => x"74812a55",
  1938 => x"555654e5",
  1939 => x"39101010",
  1940 => x"10101010",
  1941 => x"10101010",
  1942 => x"10101010",
  1943 => x"10101010",
  1944 => x"10101010",
  1945 => x"10101010",
  1946 => x"10101010",
  1947 => x"53510473",
  1948 => x"81ff0673",
  1949 => x"83060981",
  1950 => x"05830510",
  1951 => x"10102b07",
  1952 => x"72fc060c",
  1953 => x"5151043c",
  1954 => x"04727280",
  1955 => x"728106ff",
  1956 => x"05097206",
  1957 => x"05711052",
  1958 => x"720a100a",
  1959 => x"5372ed38",
  1960 => x"51515351",
  1961 => x"04b008b4",
  1962 => x"08b80875",
  1963 => x"75bbb82d",
  1964 => x"5050b008",
  1965 => x"56b80cb4",
  1966 => x"0cb00c51",
  1967 => x"04b008b4",
  1968 => x"08b80875",
  1969 => x"75baf42d",
  1970 => x"5050b008",
  1971 => x"56b80cb4",
  1972 => x"0cb00c51",
  1973 => x"04b008b4",
  1974 => x"08b80890",
  1975 => x"cb2db80c",
  1976 => x"b40cb00c",
  1977 => x"04ff3d0d",
  1978 => x"028f0533",
  1979 => x"80fcf808",
  1980 => x"52710c80",
  1981 => x"0bb00c83",
  1982 => x"3d0d04ff",
  1983 => x"3d0d028f",
  1984 => x"05335181",
  1985 => x"a5900852",
  1986 => x"712db008",
  1987 => x"81ff06b0",
  1988 => x"0c833d0d",
  1989 => x"04fe3d0d",
  1990 => x"74703353",
  1991 => x"5371802e",
  1992 => x"93388113",
  1993 => x"725281a5",
  1994 => x"90085353",
  1995 => x"712d7233",
  1996 => x"5271ef38",
  1997 => x"843d0d04",
  1998 => x"f43d0d7f",
  1999 => x"028405bb",
  2000 => x"05335557",
  2001 => x"880b8c3d",
  2002 => x"5b598953",
  2003 => x"80fa9c52",
  2004 => x"795185e6",
  2005 => x"3f73792e",
  2006 => x"80ff3878",
  2007 => x"5673902e",
  2008 => x"80ec3802",
  2009 => x"a7055876",
  2010 => x"8f065473",
  2011 => x"892680c2",
  2012 => x"387518b0",
  2013 => x"15555573",
  2014 => x"75347684",
  2015 => x"2aff1770",
  2016 => x"81ff0658",
  2017 => x"555775df",
  2018 => x"38781a55",
  2019 => x"75753479",
  2020 => x"70335555",
  2021 => x"73802e93",
  2022 => x"38811574",
  2023 => x"5281a590",
  2024 => x"08575575",
  2025 => x"2d743354",
  2026 => x"73ef3878",
  2027 => x"b00c8e3d",
  2028 => x"0d047518",
  2029 => x"b7155555",
  2030 => x"73753476",
  2031 => x"842aff17",
  2032 => x"7081ff06",
  2033 => x"58555775",
  2034 => x"ff9d38ff",
  2035 => x"bc398470",
  2036 => x"575902a7",
  2037 => x"0558ff8f",
  2038 => x"39827057",
  2039 => x"59f439f1",
  2040 => x"3d0d618d",
  2041 => x"3d705b5c",
  2042 => x"5a807a56",
  2043 => x"57767a24",
  2044 => x"81853878",
  2045 => x"17548a52",
  2046 => x"7451848c",
  2047 => x"3fb008b0",
  2048 => x"05537274",
  2049 => x"34811757",
  2050 => x"8a527451",
  2051 => x"83d53fb0",
  2052 => x"0855b008",
  2053 => x"de38b008",
  2054 => x"779f2a18",
  2055 => x"70812c5a",
  2056 => x"56568078",
  2057 => x"259e3878",
  2058 => x"17ff0555",
  2059 => x"75197033",
  2060 => x"55537433",
  2061 => x"73347375",
  2062 => x"348116ff",
  2063 => x"16565677",
  2064 => x"7624e938",
  2065 => x"76195880",
  2066 => x"7834807a",
  2067 => x"24177081",
  2068 => x"ff067c70",
  2069 => x"33565755",
  2070 => x"5672802e",
  2071 => x"93388115",
  2072 => x"735281a5",
  2073 => x"90085855",
  2074 => x"762d7433",
  2075 => x"5372ef38",
  2076 => x"73b00c91",
  2077 => x"3d0d04ad",
  2078 => x"7b3402ad",
  2079 => x"057a3071",
  2080 => x"19565659",
  2081 => x"8a527451",
  2082 => x"82fe3fb0",
  2083 => x"08b00553",
  2084 => x"72743481",
  2085 => x"17578a52",
  2086 => x"745182c7",
  2087 => x"3fb00855",
  2088 => x"b008fecf",
  2089 => x"38feef39",
  2090 => x"fd3d0d02",
  2091 => x"97053302",
  2092 => x"84059b05",
  2093 => x"33555372",
  2094 => x"74279738",
  2095 => x"a05181a5",
  2096 => x"90085271",
  2097 => x"2d811370",
  2098 => x"81ff0654",
  2099 => x"52737326",
  2100 => x"eb38853d",
  2101 => x"0d04ff3d",
  2102 => x"0d80fcec",
  2103 => x"08741015",
  2104 => x"70822b94",
  2105 => x"130c5252",
  2106 => x"850b9813",
  2107 => x"0c981208",
  2108 => x"70810651",
  2109 => x"5170f638",
  2110 => x"833d0d04",
  2111 => x"fd3d0d80",
  2112 => x"fcec0876",
  2113 => x"80e1d429",
  2114 => x"94120c54",
  2115 => x"850b9815",
  2116 => x"0c981408",
  2117 => x"70810651",
  2118 => x"5372f638",
  2119 => x"853d0d04",
  2120 => x"803d0d80",
  2121 => x"fcec0851",
  2122 => x"870b8412",
  2123 => x"0cff0ba4",
  2124 => x"120ca70b",
  2125 => x"a8120c80",
  2126 => x"e1d40b94",
  2127 => x"120c870b",
  2128 => x"98120c82",
  2129 => x"3d0d0480",
  2130 => x"3d0d80fc",
  2131 => x"f0085180",
  2132 => x"ec0b8c12",
  2133 => x"0c830b88",
  2134 => x"120c823d",
  2135 => x"0d04803d",
  2136 => x"0d80fcf0",
  2137 => x"08841108",
  2138 => x"8106b00c",
  2139 => x"51823d0d",
  2140 => x"04ff3d0d",
  2141 => x"80fcf008",
  2142 => x"52841208",
  2143 => x"70810651",
  2144 => x"5170802e",
  2145 => x"f4387108",
  2146 => x"7081ff06",
  2147 => x"b00c5183",
  2148 => x"3d0d04fe",
  2149 => x"3d0d0293",
  2150 => x"05335372",
  2151 => x"8a2e9c38",
  2152 => x"80fcf008",
  2153 => x"52841208",
  2154 => x"70892a70",
  2155 => x"81065151",
  2156 => x"5170f238",
  2157 => x"72720c84",
  2158 => x"3d0d0480",
  2159 => x"fcf00852",
  2160 => x"84120870",
  2161 => x"892a7081",
  2162 => x"06515151",
  2163 => x"70f2388d",
  2164 => x"720c8412",
  2165 => x"0870892a",
  2166 => x"70810651",
  2167 => x"515170c5",
  2168 => x"38d239bc",
  2169 => x"0802bc0c",
  2170 => x"fd3d0d80",
  2171 => x"53bc088c",
  2172 => x"050852bc",
  2173 => x"08880508",
  2174 => x"51f7f53f",
  2175 => x"b00870b0",
  2176 => x"0c54853d",
  2177 => x"0dbc0c04",
  2178 => x"bc0802bc",
  2179 => x"0cfd3d0d",
  2180 => x"8153bc08",
  2181 => x"8c050852",
  2182 => x"bc088805",
  2183 => x"0851f7d0",
  2184 => x"3fb00870",
  2185 => x"b00c5485",
  2186 => x"3d0dbc0c",
  2187 => x"04803d0d",
  2188 => x"86518496",
  2189 => x"3f8151a1",
  2190 => x"d33ffc3d",
  2191 => x"0d767079",
  2192 => x"7b555555",
  2193 => x"558f7227",
  2194 => x"8c387275",
  2195 => x"07830651",
  2196 => x"70802ea7",
  2197 => x"38ff1252",
  2198 => x"71ff2e98",
  2199 => x"38727081",
  2200 => x"05543374",
  2201 => x"70810556",
  2202 => x"34ff1252",
  2203 => x"71ff2e09",
  2204 => x"8106ea38",
  2205 => x"74b00c86",
  2206 => x"3d0d0474",
  2207 => x"51727084",
  2208 => x"05540871",
  2209 => x"70840553",
  2210 => x"0c727084",
  2211 => x"05540871",
  2212 => x"70840553",
  2213 => x"0c727084",
  2214 => x"05540871",
  2215 => x"70840553",
  2216 => x"0c727084",
  2217 => x"05540871",
  2218 => x"70840553",
  2219 => x"0cf01252",
  2220 => x"718f26c9",
  2221 => x"38837227",
  2222 => x"95387270",
  2223 => x"84055408",
  2224 => x"71708405",
  2225 => x"530cfc12",
  2226 => x"52718326",
  2227 => x"ed387054",
  2228 => x"ff8339fd",
  2229 => x"3d0d7553",
  2230 => x"84d81308",
  2231 => x"802e8a38",
  2232 => x"805372b0",
  2233 => x"0c853d0d",
  2234 => x"04818052",
  2235 => x"72518d9b",
  2236 => x"3fb00884",
  2237 => x"d8140cff",
  2238 => x"53b00880",
  2239 => x"2ee438b0",
  2240 => x"08549f53",
  2241 => x"80747084",
  2242 => x"05560cff",
  2243 => x"13538073",
  2244 => x"24ce3880",
  2245 => x"74708405",
  2246 => x"560cff13",
  2247 => x"53728025",
  2248 => x"e338ffbc",
  2249 => x"39fd3d0d",
  2250 => x"75775553",
  2251 => x"9f74278d",
  2252 => x"3896730c",
  2253 => x"ff5271b0",
  2254 => x"0c853d0d",
  2255 => x"0484d813",
  2256 => x"08527180",
  2257 => x"2e933873",
  2258 => x"10101270",
  2259 => x"0879720c",
  2260 => x"515271b0",
  2261 => x"0c853d0d",
  2262 => x"047251fe",
  2263 => x"f63fff52",
  2264 => x"b008d338",
  2265 => x"84d81308",
  2266 => x"74101011",
  2267 => x"70087a72",
  2268 => x"0c515152",
  2269 => x"dd39f93d",
  2270 => x"0d797b58",
  2271 => x"56769f26",
  2272 => x"80e83884",
  2273 => x"d8160854",
  2274 => x"73802eaa",
  2275 => x"38761010",
  2276 => x"14700855",
  2277 => x"5573802e",
  2278 => x"ba388058",
  2279 => x"73812e8f",
  2280 => x"3873ff2e",
  2281 => x"a3388075",
  2282 => x"0c765173",
  2283 => x"2d805877",
  2284 => x"b00c893d",
  2285 => x"0d047551",
  2286 => x"fe993fff",
  2287 => x"58b008ef",
  2288 => x"3884d816",
  2289 => x"0854c639",
  2290 => x"96760c81",
  2291 => x"0bb00c89",
  2292 => x"3d0d0475",
  2293 => x"5181ed3f",
  2294 => x"7653b008",
  2295 => x"52755181",
  2296 => x"ad3fb008",
  2297 => x"b00c893d",
  2298 => x"0d049676",
  2299 => x"0cff0bb0",
  2300 => x"0c893d0d",
  2301 => x"04fc3d0d",
  2302 => x"76785653",
  2303 => x"ff54749f",
  2304 => x"26b13884",
  2305 => x"d8130852",
  2306 => x"71802eae",
  2307 => x"38741010",
  2308 => x"12700853",
  2309 => x"53815471",
  2310 => x"802e9838",
  2311 => x"825471ff",
  2312 => x"2e913883",
  2313 => x"5471812e",
  2314 => x"8a388073",
  2315 => x"0c745171",
  2316 => x"2d805473",
  2317 => x"b00c863d",
  2318 => x"0d047251",
  2319 => x"fd953fb0",
  2320 => x"08f13884",
  2321 => x"d8130852",
  2322 => x"c439ff3d",
  2323 => x"0d735280",
  2324 => x"fcfc0851",
  2325 => x"fea03f83",
  2326 => x"3d0d04fe",
  2327 => x"3d0d7553",
  2328 => x"745280fc",
  2329 => x"fc0851fd",
  2330 => x"bc3f843d",
  2331 => x"0d04803d",
  2332 => x"0d80fcfc",
  2333 => x"0851fcdb",
  2334 => x"3f823d0d",
  2335 => x"04ff3d0d",
  2336 => x"735280fc",
  2337 => x"fc0851fe",
  2338 => x"ec3f833d",
  2339 => x"0d04fc3d",
  2340 => x"0d800b81",
  2341 => x"a5980c78",
  2342 => x"5277519c",
  2343 => x"aa3fb008",
  2344 => x"54b008ff",
  2345 => x"2e883873",
  2346 => x"b00c863d",
  2347 => x"0d0481a5",
  2348 => x"98085574",
  2349 => x"802ef038",
  2350 => x"7675710c",
  2351 => x"5373b00c",
  2352 => x"863d0d04",
  2353 => x"9bfc3f04",
  2354 => x"fc3d0d76",
  2355 => x"70797073",
  2356 => x"07830654",
  2357 => x"54545570",
  2358 => x"80c33871",
  2359 => x"70087009",
  2360 => x"70f7fbfd",
  2361 => x"ff130670",
  2362 => x"f8848281",
  2363 => x"80065151",
  2364 => x"53535470",
  2365 => x"a6388414",
  2366 => x"72747084",
  2367 => x"05560c70",
  2368 => x"08700970",
  2369 => x"f7fbfdff",
  2370 => x"130670f8",
  2371 => x"84828180",
  2372 => x"06515153",
  2373 => x"53547080",
  2374 => x"2edc3873",
  2375 => x"52717081",
  2376 => x"05533351",
  2377 => x"70737081",
  2378 => x"05553470",
  2379 => x"f03874b0",
  2380 => x"0c863d0d",
  2381 => x"04fd3d0d",
  2382 => x"75707183",
  2383 => x"06535552",
  2384 => x"70b83871",
  2385 => x"70087009",
  2386 => x"f7fbfdff",
  2387 => x"120670f8",
  2388 => x"84828180",
  2389 => x"06515152",
  2390 => x"53709d38",
  2391 => x"84137008",
  2392 => x"7009f7fb",
  2393 => x"fdff1206",
  2394 => x"70f88482",
  2395 => x"81800651",
  2396 => x"51525370",
  2397 => x"802ee538",
  2398 => x"72527133",
  2399 => x"5170802e",
  2400 => x"8a388112",
  2401 => x"70335252",
  2402 => x"70f83871",
  2403 => x"7431b00c",
  2404 => x"853d0d04",
  2405 => x"fa3d0d78",
  2406 => x"7a7c7054",
  2407 => x"55555272",
  2408 => x"802e80d9",
  2409 => x"38717407",
  2410 => x"83065170",
  2411 => x"802e80d4",
  2412 => x"38ff1353",
  2413 => x"72ff2eb1",
  2414 => x"38713374",
  2415 => x"33565174",
  2416 => x"712e0981",
  2417 => x"06a93872",
  2418 => x"802e8187",
  2419 => x"387081ff",
  2420 => x"06517080",
  2421 => x"2e80fc38",
  2422 => x"81128115",
  2423 => x"ff155555",
  2424 => x"5272ff2e",
  2425 => x"098106d1",
  2426 => x"38713374",
  2427 => x"33565170",
  2428 => x"81ff0675",
  2429 => x"81ff0671",
  2430 => x"71315152",
  2431 => x"5270b00c",
  2432 => x"883d0d04",
  2433 => x"71745755",
  2434 => x"83732788",
  2435 => x"38710874",
  2436 => x"082e8838",
  2437 => x"74765552",
  2438 => x"ff9739fc",
  2439 => x"13537280",
  2440 => x"2eb13874",
  2441 => x"087009f7",
  2442 => x"fbfdff12",
  2443 => x"0670f884",
  2444 => x"82818006",
  2445 => x"51515170",
  2446 => x"9a388415",
  2447 => x"84175755",
  2448 => x"837327d0",
  2449 => x"38740876",
  2450 => x"082ed038",
  2451 => x"74765552",
  2452 => x"fedf3980",
  2453 => x"0bb00c88",
  2454 => x"3d0d04f3",
  2455 => x"3d0d6062",
  2456 => x"64725a5a",
  2457 => x"5e5e805c",
  2458 => x"76708105",
  2459 => x"583380fa",
  2460 => x"b1113370",
  2461 => x"832a7081",
  2462 => x"06515555",
  2463 => x"5672e938",
  2464 => x"75ad2e82",
  2465 => x"883875ab",
  2466 => x"2e828438",
  2467 => x"77307079",
  2468 => x"07802579",
  2469 => x"90327030",
  2470 => x"70720780",
  2471 => x"25730753",
  2472 => x"57575153",
  2473 => x"72802e87",
  2474 => x"3875b02e",
  2475 => x"81eb3877",
  2476 => x"8a388858",
  2477 => x"75b02e83",
  2478 => x"388a5881",
  2479 => x"0a5a7b84",
  2480 => x"38fe0a5a",
  2481 => x"77527951",
  2482 => x"f6be3fb0",
  2483 => x"0878537a",
  2484 => x"525bf68f",
  2485 => x"3fb0085a",
  2486 => x"807080fa",
  2487 => x"b1183370",
  2488 => x"822a7081",
  2489 => x"06515656",
  2490 => x"5a557280",
  2491 => x"2e80c138",
  2492 => x"d0165675",
  2493 => x"782580d7",
  2494 => x"38807924",
  2495 => x"757b2607",
  2496 => x"53729338",
  2497 => x"747a2e80",
  2498 => x"eb387a76",
  2499 => x"2580ed38",
  2500 => x"72802e80",
  2501 => x"e738ff77",
  2502 => x"70810559",
  2503 => x"33575980",
  2504 => x"fab11633",
  2505 => x"70822a70",
  2506 => x"81065154",
  2507 => x"5472c138",
  2508 => x"73830653",
  2509 => x"72802e97",
  2510 => x"38738106",
  2511 => x"c9175553",
  2512 => x"728538ff",
  2513 => x"a9165473",
  2514 => x"56777624",
  2515 => x"ffab3880",
  2516 => x"792480f0",
  2517 => x"387b802e",
  2518 => x"84387430",
  2519 => x"557c802e",
  2520 => x"8c38ff17",
  2521 => x"53788338",
  2522 => x"7d53727d",
  2523 => x"0c74b00c",
  2524 => x"8f3d0d04",
  2525 => x"8153757b",
  2526 => x"24ff9538",
  2527 => x"81757929",
  2528 => x"17787081",
  2529 => x"055a3358",
  2530 => x"5659ff93",
  2531 => x"39815c76",
  2532 => x"70810558",
  2533 => x"3356fdf4",
  2534 => x"39807733",
  2535 => x"54547280",
  2536 => x"f82eb238",
  2537 => x"7280d832",
  2538 => x"70307080",
  2539 => x"25760751",
  2540 => x"51537280",
  2541 => x"2efdf838",
  2542 => x"81173382",
  2543 => x"18585690",
  2544 => x"58fdf839",
  2545 => x"810a557b",
  2546 => x"8438fe0a",
  2547 => x"557f53a2",
  2548 => x"730cff89",
  2549 => x"398154cc",
  2550 => x"39fd3d0d",
  2551 => x"77547653",
  2552 => x"755280fc",
  2553 => x"fc0851fc",
  2554 => x"f23f853d",
  2555 => x"0d04f33d",
  2556 => x"0d606264",
  2557 => x"725a5a5d",
  2558 => x"5d805e76",
  2559 => x"70810558",
  2560 => x"3380fab1",
  2561 => x"11337083",
  2562 => x"2a708106",
  2563 => x"51555556",
  2564 => x"72e93875",
  2565 => x"ad2e81ff",
  2566 => x"3875ab2e",
  2567 => x"81fb3877",
  2568 => x"30707907",
  2569 => x"80257990",
  2570 => x"32703070",
  2571 => x"72078025",
  2572 => x"73075357",
  2573 => x"57515372",
  2574 => x"802e8738",
  2575 => x"75b02e81",
  2576 => x"e238778a",
  2577 => x"38885875",
  2578 => x"b02e8338",
  2579 => x"8a587752",
  2580 => x"ff51f38f",
  2581 => x"3fb00878",
  2582 => x"535aff51",
  2583 => x"f3aa3fb0",
  2584 => x"085b8070",
  2585 => x"5a5580fa",
  2586 => x"b1163370",
  2587 => x"822a7081",
  2588 => x"06515454",
  2589 => x"72802e80",
  2590 => x"c138d016",
  2591 => x"56757825",
  2592 => x"80d73880",
  2593 => x"7924757b",
  2594 => x"26075372",
  2595 => x"9338747a",
  2596 => x"2e80eb38",
  2597 => x"7a762580",
  2598 => x"ed387280",
  2599 => x"2e80e738",
  2600 => x"ff777081",
  2601 => x"05593357",
  2602 => x"5980fab1",
  2603 => x"16337082",
  2604 => x"2a708106",
  2605 => x"51545472",
  2606 => x"c1387383",
  2607 => x"06537280",
  2608 => x"2e973873",
  2609 => x"8106c917",
  2610 => x"55537285",
  2611 => x"38ffa916",
  2612 => x"54735677",
  2613 => x"7624ffab",
  2614 => x"38807924",
  2615 => x"8189387d",
  2616 => x"802e8438",
  2617 => x"7430557b",
  2618 => x"802e8c38",
  2619 => x"ff175378",
  2620 => x"83387c53",
  2621 => x"727c0c74",
  2622 => x"b00c8f3d",
  2623 => x"0d048153",
  2624 => x"757b24ff",
  2625 => x"95388175",
  2626 => x"79291778",
  2627 => x"7081055a",
  2628 => x"33585659",
  2629 => x"ff933981",
  2630 => x"5e767081",
  2631 => x"05583356",
  2632 => x"fdfd3980",
  2633 => x"77335454",
  2634 => x"7280f82e",
  2635 => x"80c33872",
  2636 => x"80d83270",
  2637 => x"30708025",
  2638 => x"76075151",
  2639 => x"5372802e",
  2640 => x"fe803881",
  2641 => x"17338218",
  2642 => x"58569070",
  2643 => x"5358ff51",
  2644 => x"f1913fb0",
  2645 => x"0878535a",
  2646 => x"ff51f1ac",
  2647 => x"3fb0085b",
  2648 => x"80705a55",
  2649 => x"fe8039ff",
  2650 => x"605455a2",
  2651 => x"730cfef7",
  2652 => x"398154ff",
  2653 => x"ba39fd3d",
  2654 => x"0d775476",
  2655 => x"53755280",
  2656 => x"fcfc0851",
  2657 => x"fce83f85",
  2658 => x"3d0d04f3",
  2659 => x"3d0d7f61",
  2660 => x"8b1170f8",
  2661 => x"065c5555",
  2662 => x"5e729626",
  2663 => x"83389059",
  2664 => x"80792474",
  2665 => x"7a260753",
  2666 => x"80547274",
  2667 => x"2e098106",
  2668 => x"80cb387d",
  2669 => x"518bca3f",
  2670 => x"7883f726",
  2671 => x"80c63878",
  2672 => x"832a7010",
  2673 => x"10108184",
  2674 => x"b8058c11",
  2675 => x"0859595a",
  2676 => x"76782e83",
  2677 => x"b0388417",
  2678 => x"08fc0656",
  2679 => x"8c170888",
  2680 => x"1808718c",
  2681 => x"120c8812",
  2682 => x"0c587517",
  2683 => x"84110881",
  2684 => x"0784120c",
  2685 => x"537d518b",
  2686 => x"893f8817",
  2687 => x"5473b00c",
  2688 => x"8f3d0d04",
  2689 => x"78892a79",
  2690 => x"832a5b53",
  2691 => x"72802ebf",
  2692 => x"3878862a",
  2693 => x"b8055a84",
  2694 => x"7327b438",
  2695 => x"80db135a",
  2696 => x"947327ab",
  2697 => x"38788c2a",
  2698 => x"80ee055a",
  2699 => x"80d47327",
  2700 => x"9e38788f",
  2701 => x"2a80f705",
  2702 => x"5a82d473",
  2703 => x"27913878",
  2704 => x"922a80fc",
  2705 => x"055a8ad4",
  2706 => x"73278438",
  2707 => x"80fe5a79",
  2708 => x"10101081",
  2709 => x"84b8058c",
  2710 => x"11085855",
  2711 => x"76752ea3",
  2712 => x"38841708",
  2713 => x"fc06707a",
  2714 => x"31555673",
  2715 => x"8f2488d5",
  2716 => x"38738025",
  2717 => x"fee6388c",
  2718 => x"17085776",
  2719 => x"752e0981",
  2720 => x"06df3881",
  2721 => x"1a5a8184",
  2722 => x"c8085776",
  2723 => x"8184c02e",
  2724 => x"82c03884",
  2725 => x"1708fc06",
  2726 => x"707a3155",
  2727 => x"56738f24",
  2728 => x"81f93881",
  2729 => x"84c00b81",
  2730 => x"84cc0c81",
  2731 => x"84c00b81",
  2732 => x"84c80c73",
  2733 => x"8025feb2",
  2734 => x"3883ff76",
  2735 => x"2783df38",
  2736 => x"75892a76",
  2737 => x"832a5553",
  2738 => x"72802ebf",
  2739 => x"3875862a",
  2740 => x"b8055484",
  2741 => x"7327b438",
  2742 => x"80db1354",
  2743 => x"947327ab",
  2744 => x"38758c2a",
  2745 => x"80ee0554",
  2746 => x"80d47327",
  2747 => x"9e38758f",
  2748 => x"2a80f705",
  2749 => x"5482d473",
  2750 => x"27913875",
  2751 => x"922a80fc",
  2752 => x"05548ad4",
  2753 => x"73278438",
  2754 => x"80fe5473",
  2755 => x"10101081",
  2756 => x"84b80588",
  2757 => x"11085658",
  2758 => x"74782e86",
  2759 => x"cf388415",
  2760 => x"08fc0653",
  2761 => x"7573278d",
  2762 => x"38881508",
  2763 => x"5574782e",
  2764 => x"098106ea",
  2765 => x"388c1508",
  2766 => x"8184b80b",
  2767 => x"84050871",
  2768 => x"8c1a0c76",
  2769 => x"881a0c78",
  2770 => x"88130c78",
  2771 => x"8c180c5d",
  2772 => x"58795380",
  2773 => x"7a2483e6",
  2774 => x"3872822c",
  2775 => x"81712b5c",
  2776 => x"537a7c26",
  2777 => x"8198387b",
  2778 => x"7b065372",
  2779 => x"82f13879",
  2780 => x"fc068405",
  2781 => x"5a7a1070",
  2782 => x"7d06545b",
  2783 => x"7282e038",
  2784 => x"841a5af1",
  2785 => x"3988178c",
  2786 => x"11085858",
  2787 => x"76782e09",
  2788 => x"8106fcc2",
  2789 => x"38821a5a",
  2790 => x"fdec3978",
  2791 => x"17798107",
  2792 => x"84190c70",
  2793 => x"8184cc0c",
  2794 => x"708184c8",
  2795 => x"0c8184c0",
  2796 => x"0b8c120c",
  2797 => x"8c110888",
  2798 => x"120c7481",
  2799 => x"0784120c",
  2800 => x"74117571",
  2801 => x"0c51537d",
  2802 => x"5187b73f",
  2803 => x"881754fc",
  2804 => x"ac398184",
  2805 => x"b80b8405",
  2806 => x"087a545c",
  2807 => x"798025fe",
  2808 => x"f83882da",
  2809 => x"397a097c",
  2810 => x"06708184",
  2811 => x"b80b8405",
  2812 => x"0c5c7a10",
  2813 => x"5b7a7c26",
  2814 => x"85387a85",
  2815 => x"b8388184",
  2816 => x"b80b8805",
  2817 => x"08708412",
  2818 => x"08fc0670",
  2819 => x"7c317c72",
  2820 => x"268f7225",
  2821 => x"0757575c",
  2822 => x"5d557280",
  2823 => x"2e80db38",
  2824 => x"797a1681",
  2825 => x"84b0081b",
  2826 => x"90115a55",
  2827 => x"575b8184",
  2828 => x"ac08ff2e",
  2829 => x"8838a08f",
  2830 => x"13e08006",
  2831 => x"5776527d",
  2832 => x"5186c03f",
  2833 => x"b00854b0",
  2834 => x"08ff2e90",
  2835 => x"38b00876",
  2836 => x"27829938",
  2837 => x"748184b8",
  2838 => x"2e829138",
  2839 => x"8184b80b",
  2840 => x"88050855",
  2841 => x"841508fc",
  2842 => x"06707a31",
  2843 => x"7a72268f",
  2844 => x"72250752",
  2845 => x"55537283",
  2846 => x"e6387479",
  2847 => x"81078417",
  2848 => x"0c791670",
  2849 => x"8184b80b",
  2850 => x"88050c75",
  2851 => x"81078412",
  2852 => x"0c547e52",
  2853 => x"5785eb3f",
  2854 => x"881754fa",
  2855 => x"e0397583",
  2856 => x"2a705454",
  2857 => x"80742481",
  2858 => x"9b387282",
  2859 => x"2c81712b",
  2860 => x"8184bc08",
  2861 => x"07708184",
  2862 => x"b80b8405",
  2863 => x"0c751010",
  2864 => x"108184b8",
  2865 => x"05881108",
  2866 => x"585a5d53",
  2867 => x"778c180c",
  2868 => x"7488180c",
  2869 => x"7688190c",
  2870 => x"768c160c",
  2871 => x"fcf33979",
  2872 => x"7a101010",
  2873 => x"8184b805",
  2874 => x"7057595d",
  2875 => x"8c150857",
  2876 => x"76752ea3",
  2877 => x"38841708",
  2878 => x"fc06707a",
  2879 => x"31555673",
  2880 => x"8f2483ca",
  2881 => x"38738025",
  2882 => x"8481388c",
  2883 => x"17085776",
  2884 => x"752e0981",
  2885 => x"06df3888",
  2886 => x"15811b70",
  2887 => x"8306555b",
  2888 => x"5572c938",
  2889 => x"7c830653",
  2890 => x"72802efd",
  2891 => x"b838ff1d",
  2892 => x"f819595d",
  2893 => x"88180878",
  2894 => x"2eea38fd",
  2895 => x"b539831a",
  2896 => x"53fc9639",
  2897 => x"83147082",
  2898 => x"2c81712b",
  2899 => x"8184bc08",
  2900 => x"07708184",
  2901 => x"b80b8405",
  2902 => x"0c761010",
  2903 => x"108184b8",
  2904 => x"05881108",
  2905 => x"595b5e51",
  2906 => x"53fee139",
  2907 => x"8183fc08",
  2908 => x"1758b008",
  2909 => x"762e818d",
  2910 => x"388184ac",
  2911 => x"08ff2e83",
  2912 => x"ec387376",
  2913 => x"31188183",
  2914 => x"fc0c7387",
  2915 => x"06705753",
  2916 => x"72802e88",
  2917 => x"38887331",
  2918 => x"70155556",
  2919 => x"76149fff",
  2920 => x"06a08071",
  2921 => x"31177054",
  2922 => x"7f535753",
  2923 => x"83d53fb0",
  2924 => x"0853b008",
  2925 => x"ff2e81a0",
  2926 => x"388183fc",
  2927 => x"08167081",
  2928 => x"83fc0c74",
  2929 => x"758184b8",
  2930 => x"0b88050c",
  2931 => x"74763118",
  2932 => x"70810751",
  2933 => x"5556587b",
  2934 => x"8184b82e",
  2935 => x"839c3879",
  2936 => x"8f2682cb",
  2937 => x"38810b84",
  2938 => x"150c8415",
  2939 => x"08fc0670",
  2940 => x"7a317a72",
  2941 => x"268f7225",
  2942 => x"07525553",
  2943 => x"72802efc",
  2944 => x"f93880db",
  2945 => x"39b0089f",
  2946 => x"ff065372",
  2947 => x"feeb3877",
  2948 => x"8183fc0c",
  2949 => x"8184b80b",
  2950 => x"8805087b",
  2951 => x"18810784",
  2952 => x"120c5581",
  2953 => x"84a80878",
  2954 => x"27863877",
  2955 => x"8184a80c",
  2956 => x"8184a408",
  2957 => x"7827fcac",
  2958 => x"38778184",
  2959 => x"a40c8415",
  2960 => x"08fc0670",
  2961 => x"7a317a72",
  2962 => x"268f7225",
  2963 => x"07525553",
  2964 => x"72802efc",
  2965 => x"a5388839",
  2966 => x"80745456",
  2967 => x"fedb397d",
  2968 => x"51829f3f",
  2969 => x"800bb00c",
  2970 => x"8f3d0d04",
  2971 => x"73538074",
  2972 => x"24a93872",
  2973 => x"822c8171",
  2974 => x"2b8184bc",
  2975 => x"08077081",
  2976 => x"84b80b84",
  2977 => x"050c5d53",
  2978 => x"778c180c",
  2979 => x"7488180c",
  2980 => x"7688190c",
  2981 => x"768c160c",
  2982 => x"f9b73983",
  2983 => x"1470822c",
  2984 => x"81712b81",
  2985 => x"84bc0807",
  2986 => x"708184b8",
  2987 => x"0b84050c",
  2988 => x"5e5153d4",
  2989 => x"397b7b06",
  2990 => x"5372fca3",
  2991 => x"38841a7b",
  2992 => x"105c5af1",
  2993 => x"39ff1a81",
  2994 => x"11515af7",
  2995 => x"b9397817",
  2996 => x"79810784",
  2997 => x"190c8c18",
  2998 => x"08881908",
  2999 => x"718c120c",
  3000 => x"88120c59",
  3001 => x"708184cc",
  3002 => x"0c708184",
  3003 => x"c80c8184",
  3004 => x"c00b8c12",
  3005 => x"0c8c1108",
  3006 => x"88120c74",
  3007 => x"81078412",
  3008 => x"0c741175",
  3009 => x"710c5153",
  3010 => x"f9bd3975",
  3011 => x"17841108",
  3012 => x"81078412",
  3013 => x"0c538c17",
  3014 => x"08881808",
  3015 => x"718c120c",
  3016 => x"88120c58",
  3017 => x"7d5180da",
  3018 => x"3f881754",
  3019 => x"f5cf3972",
  3020 => x"84150cf4",
  3021 => x"1af80670",
  3022 => x"841e0881",
  3023 => x"0607841e",
  3024 => x"0c701d54",
  3025 => x"5b850b84",
  3026 => x"140c850b",
  3027 => x"88140c8f",
  3028 => x"7b27fdcf",
  3029 => x"38881c52",
  3030 => x"7d518290",
  3031 => x"3f8184b8",
  3032 => x"0b880508",
  3033 => x"8183fc08",
  3034 => x"5955fdb7",
  3035 => x"39778183",
  3036 => x"fc0c7381",
  3037 => x"84ac0cfc",
  3038 => x"91397284",
  3039 => x"150cfda3",
  3040 => x"390404fd",
  3041 => x"3d0d800b",
  3042 => x"81a5980c",
  3043 => x"765186cb",
  3044 => x"3fb00853",
  3045 => x"b008ff2e",
  3046 => x"883872b0",
  3047 => x"0c853d0d",
  3048 => x"0481a598",
  3049 => x"08547380",
  3050 => x"2ef03875",
  3051 => x"74710c52",
  3052 => x"72b00c85",
  3053 => x"3d0d04fb",
  3054 => x"3d0d7770",
  3055 => x"5256c23f",
  3056 => x"8184b80b",
  3057 => x"88050884",
  3058 => x"1108fc06",
  3059 => x"707b319f",
  3060 => x"ef05e080",
  3061 => x"06e08005",
  3062 => x"565653a0",
  3063 => x"80742494",
  3064 => x"38805275",
  3065 => x"51ff9c3f",
  3066 => x"8184c008",
  3067 => x"155372b0",
  3068 => x"082e8f38",
  3069 => x"7551ff8a",
  3070 => x"3f805372",
  3071 => x"b00c873d",
  3072 => x"0d047330",
  3073 => x"527551fe",
  3074 => x"fa3fb008",
  3075 => x"ff2ea838",
  3076 => x"8184b80b",
  3077 => x"88050875",
  3078 => x"75318107",
  3079 => x"84120c53",
  3080 => x"8183fc08",
  3081 => x"74318183",
  3082 => x"fc0c7551",
  3083 => x"fed43f81",
  3084 => x"0bb00c87",
  3085 => x"3d0d0480",
  3086 => x"527551fe",
  3087 => x"c63f8184",
  3088 => x"b80b8805",
  3089 => x"08b00871",
  3090 => x"3156538f",
  3091 => x"7525ffa4",
  3092 => x"38b00881",
  3093 => x"84ac0831",
  3094 => x"8183fc0c",
  3095 => x"74810784",
  3096 => x"140c7551",
  3097 => x"fe9c3f80",
  3098 => x"53ff9039",
  3099 => x"f63d0d7c",
  3100 => x"7e545b72",
  3101 => x"802e8283",
  3102 => x"387a51fe",
  3103 => x"843ff813",
  3104 => x"84110870",
  3105 => x"fe067013",
  3106 => x"841108fc",
  3107 => x"065d5859",
  3108 => x"54588184",
  3109 => x"c008752e",
  3110 => x"82de3878",
  3111 => x"84160c80",
  3112 => x"73810654",
  3113 => x"5a727a2e",
  3114 => x"81d53878",
  3115 => x"15841108",
  3116 => x"81065153",
  3117 => x"72a03878",
  3118 => x"17577981",
  3119 => x"e6388815",
  3120 => x"08537281",
  3121 => x"84c02e82",
  3122 => x"f9388c15",
  3123 => x"08708c15",
  3124 => x"0c738812",
  3125 => x"0c567681",
  3126 => x"0784190c",
  3127 => x"76187771",
  3128 => x"0c537981",
  3129 => x"913883ff",
  3130 => x"772781c8",
  3131 => x"3876892a",
  3132 => x"77832a56",
  3133 => x"5372802e",
  3134 => x"bf387686",
  3135 => x"2ab80555",
  3136 => x"847327b4",
  3137 => x"3880db13",
  3138 => x"55947327",
  3139 => x"ab38768c",
  3140 => x"2a80ee05",
  3141 => x"5580d473",
  3142 => x"279e3876",
  3143 => x"8f2a80f7",
  3144 => x"055582d4",
  3145 => x"73279138",
  3146 => x"76922a80",
  3147 => x"fc05558a",
  3148 => x"d4732784",
  3149 => x"3880fe55",
  3150 => x"74101010",
  3151 => x"8184b805",
  3152 => x"88110855",
  3153 => x"5673762e",
  3154 => x"82b33884",
  3155 => x"1408fc06",
  3156 => x"53767327",
  3157 => x"8d388814",
  3158 => x"08547376",
  3159 => x"2e098106",
  3160 => x"ea388c14",
  3161 => x"08708c1a",
  3162 => x"0c74881a",
  3163 => x"0c788812",
  3164 => x"0c56778c",
  3165 => x"150c7a51",
  3166 => x"fc883f8c",
  3167 => x"3d0d0477",
  3168 => x"08787131",
  3169 => x"59770588",
  3170 => x"19085457",
  3171 => x"728184c0",
  3172 => x"2e80e038",
  3173 => x"8c180870",
  3174 => x"8c150c73",
  3175 => x"88120c56",
  3176 => x"fe893988",
  3177 => x"15088c16",
  3178 => x"08708c13",
  3179 => x"0c578817",
  3180 => x"0cfea339",
  3181 => x"76832a70",
  3182 => x"54558075",
  3183 => x"24819838",
  3184 => x"72822c81",
  3185 => x"712b8184",
  3186 => x"bc080781",
  3187 => x"84b80b84",
  3188 => x"050c5374",
  3189 => x"10101081",
  3190 => x"84b80588",
  3191 => x"11085556",
  3192 => x"758c190c",
  3193 => x"7388190c",
  3194 => x"7788170c",
  3195 => x"778c150c",
  3196 => x"ff843981",
  3197 => x"5afdb439",
  3198 => x"78177381",
  3199 => x"06545772",
  3200 => x"98387708",
  3201 => x"78713159",
  3202 => x"77058c19",
  3203 => x"08881a08",
  3204 => x"718c120c",
  3205 => x"88120c57",
  3206 => x"57768107",
  3207 => x"84190c77",
  3208 => x"8184b80b",
  3209 => x"88050c81",
  3210 => x"84b40877",
  3211 => x"26fec738",
  3212 => x"8184b008",
  3213 => x"527a51fa",
  3214 => x"fe3f7a51",
  3215 => x"fac43ffe",
  3216 => x"ba398178",
  3217 => x"8c150c78",
  3218 => x"88150c73",
  3219 => x"8c1a0c73",
  3220 => x"881a0c5a",
  3221 => x"fd803983",
  3222 => x"1570822c",
  3223 => x"81712b81",
  3224 => x"84bc0807",
  3225 => x"8184b80b",
  3226 => x"84050c51",
  3227 => x"53741010",
  3228 => x"108184b8",
  3229 => x"05881108",
  3230 => x"5556fee4",
  3231 => x"39745380",
  3232 => x"7524a738",
  3233 => x"72822c81",
  3234 => x"712b8184",
  3235 => x"bc080781",
  3236 => x"84b80b84",
  3237 => x"050c5375",
  3238 => x"8c190c73",
  3239 => x"88190c77",
  3240 => x"88170c77",
  3241 => x"8c150cfd",
  3242 => x"cd398315",
  3243 => x"70822c81",
  3244 => x"712b8184",
  3245 => x"bc080781",
  3246 => x"84b80b84",
  3247 => x"050c5153",
  3248 => x"d639810b",
  3249 => x"b00c0480",
  3250 => x"3d0d7281",
  3251 => x"2e893880",
  3252 => x"0bb00c82",
  3253 => x"3d0d0473",
  3254 => x"51b23ffe",
  3255 => x"3d0d81a5",
  3256 => x"94085170",
  3257 => x"8a3881a5",
  3258 => x"9c7081a5",
  3259 => x"940c5170",
  3260 => x"75125252",
  3261 => x"ff537087",
  3262 => x"fb808026",
  3263 => x"88387081",
  3264 => x"a5940c71",
  3265 => x"5372b00c",
  3266 => x"843d0d04",
  3267 => x"00ff3900",
  3268 => x"68656c70",
  3269 => x"00000000",
  3270 => x"73797374",
  3271 => x"656d2072",
  3272 => x"65736574",
  3273 => x"00000000",
  3274 => x"72657365",
  3275 => x"74000000",
  3276 => x"73686f77",
  3277 => x"20737973",
  3278 => x"74656d20",
  3279 => x"696e666f",
  3280 => x"203c7665",
  3281 => x"72626f73",
  3282 => x"653e0000",
  3283 => x"73797369",
  3284 => x"6e666f00",
  3285 => x"7265706f",
  3286 => x"72742076",
  3287 => x"65727369",
  3288 => x"6f6e0000",
  3289 => x"76657273",
  3290 => x"696f6e00",
  3291 => x"72656e61",
  3292 => x"20636f6e",
  3293 => x"74726f6c",
  3294 => x"6c657220",
  3295 => x"73746174",
  3296 => x"75730000",
  3297 => x"72656e61",
  3298 => x"20737461",
  3299 => x"74757300",
  3300 => x"3c636861",
  3301 => x"6e6e656c",
  3302 => x"3e203c68",
  3303 => x"6967683e",
  3304 => x"203c6c6f",
  3305 => x"775f636f",
  3306 => x"6e666967",
  3307 => x"3e000000",
  3308 => x"636f6e66",
  3309 => x"69670000",
  3310 => x"646f2063",
  3311 => x"6f6d706c",
  3312 => x"65746520",
  3313 => x"64656d6f",
  3314 => x"20636f6e",
  3315 => x"66696720",
  3316 => x"666f7220",
  3317 => x"52454e41",
  3318 => x"00000000",
  3319 => x"64656d6f",
  3320 => x"00000000",
  3321 => x"73657420",
  3322 => x"52454e41",
  3323 => x"20746f20",
  3324 => x"706f7765",
  3325 => x"7220646f",
  3326 => x"776e206d",
  3327 => x"6f646500",
  3328 => x"706f6666",
  3329 => x"00000000",
  3330 => x"73657420",
  3331 => x"72656e61",
  3332 => x"20636861",
  3333 => x"6e6e656c",
  3334 => x"20302074",
  3335 => x"6f20666f",
  3336 => x"6c6c6f77",
  3337 => x"6572206d",
  3338 => x"6f646500",
  3339 => x"666f6c6c",
  3340 => x"6f770000",
  3341 => x"3c74696d",
  3342 => x"653e2061",
  3343 => x"63746976",
  3344 => x"61746520",
  3345 => x"52454e41",
  3346 => x"00000000",
  3347 => x"61637175",
  3348 => x"69726500",
  3349 => x"73657420",
  3350 => x"52454e41",
  3351 => x"20636f6e",
  3352 => x"74726f6c",
  3353 => x"6c657220",
  3354 => x"746f2049",
  3355 => x"444c4500",
  3356 => x"73746f70",
  3357 => x"00000000",
  3358 => x"7072696e",
  3359 => x"74207472",
  3360 => x"69676765",
  3361 => x"72206368",
  3362 => x"61696e73",
  3363 => x"00000000",
  3364 => x"63686169",
  3365 => x"6e730000",
  3366 => x"7072696e",
  3367 => x"74207361",
  3368 => x"6d706c65",
  3369 => x"64205245",
  3370 => x"4e412074",
  3371 => x"6f6b656e",
  3372 => x"73000000",
  3373 => x"746f6b65",
  3374 => x"6e000000",
  3375 => x"74726f75",
  3376 => x"626c6573",
  3377 => x"65617263",
  3378 => x"68205245",
  3379 => x"4e410000",
  3380 => x"74726f75",
  3381 => x"626c6500",
  3382 => x"696e6974",
  3383 => x"616c697a",
  3384 => x"65204444",
  3385 => x"53206368",
  3386 => x"6970203c",
  3387 => x"66726571",
  3388 => x"2074756e",
  3389 => x"696e6720",
  3390 => x"776f7264",
  3391 => x"3e000000",
  3392 => x"64647369",
  3393 => x"6e697400",
  3394 => x"72656164",
  3395 => x"20646473",
  3396 => x"20726567",
  3397 => x"69737465",
  3398 => x"72730000",
  3399 => x"64647369",
  3400 => x"6e666f00",
  3401 => x"72756e6e",
  3402 => x"696e6720",
  3403 => x"6c696768",
  3404 => x"74000000",
  3405 => x"72756e00",
  3406 => x"63686563",
  3407 => x"6b204932",
  3408 => x"43206164",
  3409 => x"64726573",
  3410 => x"73000000",
  3411 => x"69326300",
  3412 => x"72656164",
  3413 => x"20454550",
  3414 => x"524f4d20",
  3415 => x"3c627573",
  3416 => x"3e203c69",
  3417 => x"32635f61",
  3418 => x"6464723e",
  3419 => x"203c6c65",
  3420 => x"6e677468",
  3421 => x"3e000000",
  3422 => x"65657072",
  3423 => x"6f6d0000",
  3424 => x"72656164",
  3425 => x"20616463",
  3426 => x"2076616c",
  3427 => x"75650000",
  3428 => x"61646300",
  3429 => x"67656e65",
  3430 => x"72617465",
  3431 => x"20746573",
  3432 => x"7420696d",
  3433 => x"70756c73",
  3434 => x"65000000",
  3435 => x"74657374",
  3436 => x"67656e00",
  3437 => x"616c6961",
  3438 => x"7320666f",
  3439 => x"72207800",
  3440 => x"6d656d00",
  3441 => x"77726974",
  3442 => x"6520776f",
  3443 => x"7264203c",
  3444 => x"61646472",
  3445 => x"3e203c6c",
  3446 => x"656e6774",
  3447 => x"683e203c",
  3448 => x"76616c75",
  3449 => x"65287329",
  3450 => x"3e000000",
  3451 => x"776d656d",
  3452 => x"00000000",
  3453 => x"6558616d",
  3454 => x"696e6520",
  3455 => x"6d656d6f",
  3456 => x"7279203c",
  3457 => x"61646472",
  3458 => x"3e203c6c",
  3459 => x"656e6774",
  3460 => x"683e0000",
  3461 => x"78000000",
  3462 => x"636c6561",
  3463 => x"72207363",
  3464 => x"7265656e",
  3465 => x"00000000",
  3466 => x"636c6561",
  3467 => x"72000000",
  3468 => x"0a0a0000",
  3469 => x"72656e61",
  3470 => x"3320636f",
  3471 => x"6e74726f",
  3472 => x"6c6c6572",
  3473 => x"20626f61",
  3474 => x"72640000",
  3475 => x"20286f6e",
  3476 => x"2073696d",
  3477 => x"290a0000",
  3478 => x"0a485720",
  3479 => x"73796e74",
  3480 => x"68657369",
  3481 => x"7a65643a",
  3482 => x"20000000",
  3483 => x"0a535720",
  3484 => x"636f6d70",
  3485 => x"696c6564",
  3486 => x"2020203a",
  3487 => x"204a616e",
  3488 => x"20203220",
  3489 => x"32303132",
  3490 => x"20203134",
  3491 => x"3a32313a",
  3492 => x"30320000",
  3493 => x"0a737973",
  3494 => x"74656d20",
  3495 => x"636c6f63",
  3496 => x"6b20203a",
  3497 => x"20000000",
  3498 => x"204d487a",
  3499 => x"0a000000",
  3500 => x"44454255",
  3501 => x"47204d4f",
  3502 => x"44450000",
  3503 => x"204f4e0a",
  3504 => x"00000000",
  3505 => x"56312e30",
  3506 => x"2d31322e",
  3507 => x"32303131",
  3508 => x"5f524f45",
  3509 => x"5f5a5055",
  3510 => x"00000000",
  3511 => x"4552524f",
  3512 => x"523a2074",
  3513 => x"6f6f206d",
  3514 => x"75636820",
  3515 => x"636f6d6d",
  3516 => x"616e6473",
  3517 => x"2e0a0000",
  3518 => x"3e200000",
  3519 => x"636f6d6d",
  3520 => x"616e6420",
  3521 => x"6e6f7420",
  3522 => x"666f756e",
  3523 => x"642e0a00",
  3524 => x"73757070",
  3525 => x"6f727465",
  3526 => x"6420636f",
  3527 => x"6d6d616e",
  3528 => x"64733a0a",
  3529 => x"0a000000",
  3530 => x"202d2000",
  3531 => x"76656e64",
  3532 => x"6f723f20",
  3533 => x"20000000",
  3534 => x"485a4452",
  3535 => x"20202020",
  3536 => x"20000000",
  3537 => x"67616973",
  3538 => x"6c657220",
  3539 => x"20000000",
  3540 => x"45534120",
  3541 => x"20202020",
  3542 => x"20000000",
  3543 => x"756e6b6e",
  3544 => x"6f776e20",
  3545 => x"64657669",
  3546 => x"63650000",
  3547 => x"4c656f6e",
  3548 => x"32204d65",
  3549 => x"6d6f7279",
  3550 => x"20436f6e",
  3551 => x"74726f6c",
  3552 => x"6c657200",
  3553 => x"56474120",
  3554 => x"636f6e74",
  3555 => x"726f6c6c",
  3556 => x"65720000",
  3557 => x"53504920",
  3558 => x"4d656d6f",
  3559 => x"72792043",
  3560 => x"6f6e7472",
  3561 => x"6f6c6c65",
  3562 => x"72000000",
  3563 => x"53504920",
  3564 => x"436f6e74",
  3565 => x"726f6c6c",
  3566 => x"65720000",
  3567 => x"414d4241",
  3568 => x"20577261",
  3569 => x"70706572",
  3570 => x"20666f72",
  3571 => x"204f4320",
  3572 => x"4932432d",
  3573 => x"6d617374",
  3574 => x"65720000",
  3575 => x"47522031",
  3576 => x"302f3130",
  3577 => x"30204d62",
  3578 => x"69742045",
  3579 => x"74686572",
  3580 => x"6e657420",
  3581 => x"4d414300",
  3582 => x"47656e65",
  3583 => x"72616c20",
  3584 => x"50757270",
  3585 => x"6f736520",
  3586 => x"492f4f20",
  3587 => x"706f7274",
  3588 => x"00000000",
  3589 => x"4d6f6475",
  3590 => x"6c617220",
  3591 => x"54696d65",
  3592 => x"7220556e",
  3593 => x"69740000",
  3594 => x"4475616c",
  3595 => x"2d706f72",
  3596 => x"74204148",
  3597 => x"42205352",
  3598 => x"414d206d",
  3599 => x"6f64756c",
  3600 => x"65000000",
  3601 => x"47656e65",
  3602 => x"72696320",
  3603 => x"55415254",
  3604 => x"00000000",
  3605 => x"4148422f",
  3606 => x"41504220",
  3607 => x"42726964",
  3608 => x"67650000",
  3609 => x"64696666",
  3610 => x"6572656e",
  3611 => x"7469616c",
  3612 => x"20637572",
  3613 => x"72656e74",
  3614 => x"206d6f6e",
  3615 => x"69746f72",
  3616 => x"00000000",
  3617 => x"64656275",
  3618 => x"67207472",
  3619 => x"61636572",
  3620 => x"206d656d",
  3621 => x"6f727900",
  3622 => x"4541444f",
  3623 => x"47533130",
  3624 => x"32206469",
  3625 => x"73706c61",
  3626 => x"79206472",
  3627 => x"69766572",
  3628 => x"00000000",
  3629 => x"64656275",
  3630 => x"67206275",
  3631 => x"66666572",
  3632 => x"20636f6e",
  3633 => x"74726f6c",
  3634 => x"00000000",
  3635 => x"52454e41",
  3636 => x"3320636f",
  3637 => x"6e74726f",
  3638 => x"6c6c6572",
  3639 => x"00000000",
  3640 => x"53465020",
  3641 => x"636f6e74",
  3642 => x"726f6c6c",
  3643 => x"65720000",
  3644 => x"5a505520",
  3645 => x"4d656d6f",
  3646 => x"72792077",
  3647 => x"72617070",
  3648 => x"65720000",
  3649 => x"5a505520",
  3650 => x"41484220",
  3651 => x"57726170",
  3652 => x"70657200",
  3653 => x"6265616d",
  3654 => x"20706f73",
  3655 => x"6974696f",
  3656 => x"6e206d6f",
  3657 => x"6e69746f",
  3658 => x"72000000",
  3659 => x"74726967",
  3660 => x"67657220",
  3661 => x"67656e65",
  3662 => x"7261746f",
  3663 => x"72000000",
  3664 => x"64656275",
  3665 => x"6720636f",
  3666 => x"6e736f6c",
  3667 => x"65000000",
  3668 => x"44434d20",
  3669 => x"70686173",
  3670 => x"65207368",
  3671 => x"69667420",
  3672 => x"636f6e74",
  3673 => x"726f6c00",
  3674 => x"20206170",
  3675 => x"62736c76",
  3676 => x"00000000",
  3677 => x"76656e64",
  3678 => x"20307800",
  3679 => x"64657620",
  3680 => x"30780000",
  3681 => x"76657220",
  3682 => x"00000000",
  3683 => x"69727120",
  3684 => x"00000000",
  3685 => x"61646472",
  3686 => x"20307800",
  3687 => x"6168626d",
  3688 => x"73740000",
  3689 => x"61686273",
  3690 => x"6c760000",
  3691 => x"00000f71",
  3692 => x"00001042",
  3693 => x"00001037",
  3694 => x"0000106e",
  3695 => x"00001063",
  3696 => x"00001058",
  3697 => x"0000104d",
  3698 => x"00001016",
  3699 => x"0000100b",
  3700 => x"00001000",
  3701 => x"00000ff5",
  3702 => x"0000102c",
  3703 => x"00001021",
  3704 => x"00000fea",
  3705 => x"00000f71",
  3706 => x"00000f71",
  3707 => x"00000f71",
  3708 => x"00000f71",
  3709 => x"00000f71",
  3710 => x"00000fdf",
  3711 => x"00000f71",
  3712 => x"00000f71",
  3713 => x"00000fd4",
  3714 => x"00000f71",
  3715 => x"00000fc9",
  3716 => x"00000f71",
  3717 => x"00000f71",
  3718 => x"00000f71",
  3719 => x"00000f71",
  3720 => x"00000f71",
  3721 => x"00000f71",
  3722 => x"00000f71",
  3723 => x"00000f71",
  3724 => x"00000fbe",
  3725 => x"00000f71",
  3726 => x"00000f71",
  3727 => x"00000fb3",
  3728 => x"00000f71",
  3729 => x"00000f71",
  3730 => x"00000f71",
  3731 => x"00000f71",
  3732 => x"00000f71",
  3733 => x"00000f71",
  3734 => x"00000f71",
  3735 => x"00000f71",
  3736 => x"00000f71",
  3737 => x"00000f71",
  3738 => x"00000fa8",
  3739 => x"00000f71",
  3740 => x"00000f71",
  3741 => x"00000f71",
  3742 => x"00000f71",
  3743 => x"00000f9d",
  3744 => x"00000f71",
  3745 => x"00000f71",
  3746 => x"00000f71",
  3747 => x"00000f71",
  3748 => x"00000f71",
  3749 => x"00000f71",
  3750 => x"00000f71",
  3751 => x"00000f71",
  3752 => x"00000f71",
  3753 => x"00000f71",
  3754 => x"00000f71",
  3755 => x"00000f71",
  3756 => x"00000f71",
  3757 => x"00000f71",
  3758 => x"00000f71",
  3759 => x"00000f71",
  3760 => x"00000f71",
  3761 => x"00000f71",
  3762 => x"00000f71",
  3763 => x"00000f71",
  3764 => x"00000f71",
  3765 => x"00000f71",
  3766 => x"00000f71",
  3767 => x"00000f92",
  3768 => x"00000f71",
  3769 => x"00000f71",
  3770 => x"00000f71",
  3771 => x"00000f71",
  3772 => x"00000f71",
  3773 => x"00000f71",
  3774 => x"00000f71",
  3775 => x"00000f71",
  3776 => x"00000f71",
  3777 => x"00000f71",
  3778 => x"00000f71",
  3779 => x"00000f71",
  3780 => x"00000f71",
  3781 => x"00000f71",
  3782 => x"00000f71",
  3783 => x"00000f71",
  3784 => x"00000f71",
  3785 => x"00000f71",
  3786 => x"00000f71",
  3787 => x"00000f71",
  3788 => x"00000f71",
  3789 => x"00000f71",
  3790 => x"00000f71",
  3791 => x"00000f71",
  3792 => x"00000f71",
  3793 => x"00000f71",
  3794 => x"00000f71",
  3795 => x"00000f87",
  3796 => x"69326320",
  3797 => x"464d430a",
  3798 => x"00000000",
  3799 => x"61646472",
  3800 => x"6573733a",
  3801 => x"20307800",
  3802 => x"2020202d",
  3803 => x"2d3e2020",
  3804 => x"2041434b",
  3805 => x"0a000000",
  3806 => x"72656164",
  3807 => x"20646174",
  3808 => x"61202800",
  3809 => x"20627974",
  3810 => x"65732920",
  3811 => x"66726f6d",
  3812 => x"20493243",
  3813 => x"2d616464",
  3814 => x"72657373",
  3815 => x"20307800",
  3816 => x"0a307800",
  3817 => x"02020606",
  3818 => x"06040304",
  3819 => x"02020102",
  3820 => x"636f6e74",
  3821 => x"726f6c20",
  3822 => x"2020203a",
  3823 => x"20000000",
  3824 => x"66726571",
  3825 => x"75656e63",
  3826 => x"7920203a",
  3827 => x"20000000",
  3828 => x"75706461",
  3829 => x"74652063",
  3830 => x"6c6b203a",
  3831 => x"20000000",
  3832 => x"72616d70",
  3833 => x"20726174",
  3834 => x"6520203a",
  3835 => x"20000000",
  3836 => x"49206d75",
  3837 => x"6c742072",
  3838 => x"6567203a",
  3839 => x"20000000",
  3840 => x"51206d75",
  3841 => x"6c742072",
  3842 => x"6567203a",
  3843 => x"20000000",
  3844 => x"554e4b4e",
  3845 => x"4f574e00",
  3846 => x"69646c65",
  3847 => x"00000000",
  3848 => x"636f6e66",
  3849 => x"69677572",
  3850 => x"65000000",
  3851 => x"64657465",
  3852 => x"63740000",
  3853 => x"61717569",
  3854 => x"72650000",
  3855 => x"616e616c",
  3856 => x"797a6500",
  3857 => x"64657369",
  3858 => x"72650000",
  3859 => x"72656164",
  3860 => x"6f757400",
  3861 => x"72656164",
  3862 => x"6c616700",
  3863 => x"66617374",
  3864 => x"20747269",
  3865 => x"67676572",
  3866 => x"203a2000",
  3867 => x"0a736c6f",
  3868 => x"77207472",
  3869 => x"69676765",
  3870 => x"72203a20",
  3871 => x"00000000",
  3872 => x"0a6f7665",
  3873 => x"72666c6f",
  3874 => x"77202020",
  3875 => x"20203a20",
  3876 => x"00000000",
  3877 => x"66617374",
  3878 => x"20747269",
  3879 => x"67676572",
  3880 => x"20636861",
  3881 => x"696e3a20",
  3882 => x"30780000",
  3883 => x"0a736c6f",
  3884 => x"77207472",
  3885 => x"69676765",
  3886 => x"72206368",
  3887 => x"61696e3a",
  3888 => x"20307800",
  3889 => x"746f6b65",
  3890 => x"6e733a20",
  3891 => x"00000000",
  3892 => x"00001aa2",
  3893 => x"00001ab6",
  3894 => x"00001a7a",
  3895 => x"00001aca",
  3896 => x"00001ade",
  3897 => x"00001af2",
  3898 => x"00001b06",
  3899 => x"00001b1a",
  3900 => x"00001b2e",
  3901 => x"00001a8e",
  3902 => x"30622020",
  3903 => x"20202020",
  3904 => x"20202020",
  3905 => x"20202020",
  3906 => x"20202020",
  3907 => x"20202020",
  3908 => x"20202020",
  3909 => x"20202020",
  3910 => x"20200000",
  3911 => x"20202020",
  3912 => x"20202020",
  3913 => x"00000000",
  3914 => x"79657300",
  3915 => x"6e6f0000",
  3916 => x"00202020",
  3917 => x"20202020",
  3918 => x"20202828",
  3919 => x"28282820",
  3920 => x"20202020",
  3921 => x"20202020",
  3922 => x"20202020",
  3923 => x"20202020",
  3924 => x"20881010",
  3925 => x"10101010",
  3926 => x"10101010",
  3927 => x"10101010",
  3928 => x"10040404",
  3929 => x"04040404",
  3930 => x"04040410",
  3931 => x"10101010",
  3932 => x"10104141",
  3933 => x"41414141",
  3934 => x"01010101",
  3935 => x"01010101",
  3936 => x"01010101",
  3937 => x"01010101",
  3938 => x"01010101",
  3939 => x"10101010",
  3940 => x"10104242",
  3941 => x"42424242",
  3942 => x"02020202",
  3943 => x"02020202",
  3944 => x"02020202",
  3945 => x"02020202",
  3946 => x"02020202",
  3947 => x"10101010",
  3948 => x"20000000",
  3949 => x"00000000",
  3950 => x"00000000",
  3951 => x"00000000",
  3952 => x"00000000",
  3953 => x"00000000",
  3954 => x"00000000",
  3955 => x"00000000",
  3956 => x"00000000",
  3957 => x"00000000",
  3958 => x"00000000",
  3959 => x"00000000",
  3960 => x"00000000",
  3961 => x"00000000",
  3962 => x"00000000",
  3963 => x"00000000",
  3964 => x"00000000",
  3965 => x"00000000",
  3966 => x"00000000",
  3967 => x"00000000",
  3968 => x"00000000",
  3969 => x"00000000",
  3970 => x"00000000",
  3971 => x"00000000",
  3972 => x"00000000",
  3973 => x"00000000",
  3974 => x"00000000",
  3975 => x"00000000",
  3976 => x"00000000",
  3977 => x"00000000",
  3978 => x"00000000",
  3979 => x"00000000",
  3980 => x"00000000",
  3981 => x"43000000",
  3982 => x"00000000",
  3983 => x"00000000",
  3984 => x"80000b00",
  3985 => x"10000000",
  3986 => x"80000d00",
  3987 => x"00ffffff",
  3988 => x"ff00ffff",
  3989 => x"ffff00ff",
  3990 => x"ffffff00",
  3991 => x"00000000",
  3992 => x"00000000",
  3993 => x"80000a00",
  3994 => x"80000400",
  3995 => x"80000200",
  3996 => x"80000100",
  3997 => x"80000004",
  3998 => x"80000000",
  3999 => x"00003e80",
  4000 => x"00000000",
  4001 => x"000040e8",
  4002 => x"00004144",
  4003 => x"000041a0",
  4004 => x"00000000",
  4005 => x"00000000",
  4006 => x"00000000",
  4007 => x"00000000",
  4008 => x"00000000",
  4009 => x"00000000",
  4010 => x"00000000",
  4011 => x"00000000",
  4012 => x"00000000",
  4013 => x"00003e34",
  4014 => x"00000000",
  4015 => x"00000000",
  4016 => x"00000000",
  4017 => x"00000000",
  4018 => x"00000000",
  4019 => x"00000000",
  4020 => x"00000000",
  4021 => x"00000000",
  4022 => x"00000000",
  4023 => x"00000000",
  4024 => x"00000000",
  4025 => x"00000000",
  4026 => x"00000000",
  4027 => x"00000000",
  4028 => x"00000000",
  4029 => x"00000000",
  4030 => x"00000000",
  4031 => x"00000000",
  4032 => x"00000000",
  4033 => x"00000000",
  4034 => x"00000000",
  4035 => x"00000000",
  4036 => x"00000000",
  4037 => x"00000000",
  4038 => x"00000000",
  4039 => x"00000000",
  4040 => x"00000000",
  4041 => x"00000000",
  4042 => x"00000001",
  4043 => x"330eabcd",
  4044 => x"1234e66d",
  4045 => x"deec0005",
  4046 => x"000b0000",
  4047 => x"00000000",
  4048 => x"00000000",
  4049 => x"00000000",
  4050 => x"00000000",
  4051 => x"00000000",
  4052 => x"00000000",
  4053 => x"00000000",
  4054 => x"00000000",
  4055 => x"00000000",
  4056 => x"00000000",
  4057 => x"00000000",
  4058 => x"00000000",
  4059 => x"00000000",
  4060 => x"00000000",
  4061 => x"00000000",
  4062 => x"00000000",
  4063 => x"00000000",
  4064 => x"00000000",
  4065 => x"00000000",
  4066 => x"00000000",
  4067 => x"00000000",
  4068 => x"00000000",
  4069 => x"00000000",
  4070 => x"00000000",
  4071 => x"00000000",
  4072 => x"00000000",
  4073 => x"00000000",
  4074 => x"00000000",
  4075 => x"00000000",
  4076 => x"00000000",
  4077 => x"00000000",
  4078 => x"00000000",
  4079 => x"00000000",
  4080 => x"00000000",
  4081 => x"00000000",
  4082 => x"00000000",
  4083 => x"00000000",
  4084 => x"00000000",
  4085 => x"00000000",
  4086 => x"00000000",
  4087 => x"00000000",
  4088 => x"00000000",
  4089 => x"00000000",
  4090 => x"00000000",
  4091 => x"00000000",
  4092 => x"00000000",
  4093 => x"00000000",
  4094 => x"00000000",
  4095 => x"00000000",
  4096 => x"00000000",
  4097 => x"00000000",
  4098 => x"00000000",
  4099 => x"00000000",
  4100 => x"00000000",
  4101 => x"00000000",
  4102 => x"00000000",
  4103 => x"00000000",
  4104 => x"00000000",
  4105 => x"00000000",
  4106 => x"00000000",
  4107 => x"00000000",
  4108 => x"00000000",
  4109 => x"00000000",
  4110 => x"00000000",
  4111 => x"00000000",
  4112 => x"00000000",
  4113 => x"00000000",
  4114 => x"00000000",
  4115 => x"00000000",
  4116 => x"00000000",
  4117 => x"00000000",
  4118 => x"00000000",
  4119 => x"00000000",
  4120 => x"00000000",
  4121 => x"00000000",
  4122 => x"00000000",
  4123 => x"00000000",
  4124 => x"00000000",
  4125 => x"00000000",
  4126 => x"00000000",
  4127 => x"00000000",
  4128 => x"00000000",
  4129 => x"00000000",
  4130 => x"00000000",
  4131 => x"00000000",
  4132 => x"00000000",
  4133 => x"00000000",
  4134 => x"00000000",
  4135 => x"00000000",
  4136 => x"00000000",
  4137 => x"00000000",
  4138 => x"00000000",
  4139 => x"00000000",
  4140 => x"00000000",
  4141 => x"00000000",
  4142 => x"00000000",
  4143 => x"00000000",
  4144 => x"00000000",
  4145 => x"00000000",
  4146 => x"00000000",
  4147 => x"00000000",
  4148 => x"00000000",
  4149 => x"00000000",
  4150 => x"00000000",
  4151 => x"00000000",
  4152 => x"00000000",
  4153 => x"00000000",
  4154 => x"00000000",
  4155 => x"00000000",
  4156 => x"00000000",
  4157 => x"00000000",
  4158 => x"00000000",
  4159 => x"00000000",
  4160 => x"00000000",
  4161 => x"00000000",
  4162 => x"00000000",
  4163 => x"00000000",
  4164 => x"00000000",
  4165 => x"00000000",
  4166 => x"00000000",
  4167 => x"00000000",
  4168 => x"00000000",
  4169 => x"00000000",
  4170 => x"00000000",
  4171 => x"00000000",
  4172 => x"00000000",
  4173 => x"00000000",
  4174 => x"00000000",
  4175 => x"00000000",
  4176 => x"00000000",
  4177 => x"00000000",
  4178 => x"00000000",
  4179 => x"00000000",
  4180 => x"00000000",
  4181 => x"00000000",
  4182 => x"00000000",
  4183 => x"00000000",
  4184 => x"00000000",
  4185 => x"00000000",
  4186 => x"00000000",
  4187 => x"00000000",
  4188 => x"00000000",
  4189 => x"00000000",
  4190 => x"00000000",
  4191 => x"00000000",
  4192 => x"00000000",
  4193 => x"00000000",
  4194 => x"00000000",
  4195 => x"00000000",
  4196 => x"00000000",
  4197 => x"00000000",
  4198 => x"00000000",
  4199 => x"00000000",
  4200 => x"00000000",
  4201 => x"00000000",
  4202 => x"00000000",
  4203 => x"00000000",
  4204 => x"00000000",
  4205 => x"00000000",
  4206 => x"00000000",
  4207 => x"00000000",
  4208 => x"00000000",
  4209 => x"00000000",
  4210 => x"00000000",
  4211 => x"00000000",
  4212 => x"00000000",
  4213 => x"00000000",
  4214 => x"00000000",
  4215 => x"00000000",
  4216 => x"00000000",
  4217 => x"00000000",
  4218 => x"00000000",
  4219 => x"00000000",
  4220 => x"00000000",
  4221 => x"00000000",
  4222 => x"00000000",
  4223 => x"00000000",
  4224 => x"00000000",
  4225 => x"00000000",
  4226 => x"00000000",
  4227 => x"00000000",
  4228 => x"00000000",
  4229 => x"00000000",
  4230 => x"00000000",
  4231 => x"00000000",
  4232 => x"00000000",
  4233 => x"00000000",
  4234 => x"00000000",
  4235 => x"ffffffff",
  4236 => x"00000000",
  4237 => x"00020000",
  4238 => x"00000000",
  4239 => x"00000000",
  4240 => x"00004238",
  4241 => x"00004238",
  4242 => x"00004240",
  4243 => x"00004240",
  4244 => x"00004248",
  4245 => x"00004248",
  4246 => x"00004250",
  4247 => x"00004250",
  4248 => x"00004258",
  4249 => x"00004258",
  4250 => x"00004260",
  4251 => x"00004260",
  4252 => x"00004268",
  4253 => x"00004268",
  4254 => x"00004270",
  4255 => x"00004270",
  4256 => x"00004278",
  4257 => x"00004278",
  4258 => x"00004280",
  4259 => x"00004280",
  4260 => x"00004288",
  4261 => x"00004288",
  4262 => x"00004290",
  4263 => x"00004290",
  4264 => x"00004298",
  4265 => x"00004298",
  4266 => x"000042a0",
  4267 => x"000042a0",
  4268 => x"000042a8",
  4269 => x"000042a8",
  4270 => x"000042b0",
  4271 => x"000042b0",
  4272 => x"000042b8",
  4273 => x"000042b8",
  4274 => x"000042c0",
  4275 => x"000042c0",
  4276 => x"000042c8",
  4277 => x"000042c8",
  4278 => x"000042d0",
  4279 => x"000042d0",
  4280 => x"000042d8",
  4281 => x"000042d8",
  4282 => x"000042e0",
  4283 => x"000042e0",
  4284 => x"000042e8",
  4285 => x"000042e8",
  4286 => x"000042f0",
  4287 => x"000042f0",
  4288 => x"000042f8",
  4289 => x"000042f8",
  4290 => x"00004300",
  4291 => x"00004300",
  4292 => x"00004308",
  4293 => x"00004308",
  4294 => x"00004310",
  4295 => x"00004310",
  4296 => x"00004318",
  4297 => x"00004318",
  4298 => x"00004320",
  4299 => x"00004320",
  4300 => x"00004328",
  4301 => x"00004328",
  4302 => x"00004330",
  4303 => x"00004330",
  4304 => x"00004338",
  4305 => x"00004338",
  4306 => x"00004340",
  4307 => x"00004340",
  4308 => x"00004348",
  4309 => x"00004348",
  4310 => x"00004350",
  4311 => x"00004350",
  4312 => x"00004358",
  4313 => x"00004358",
  4314 => x"00004360",
  4315 => x"00004360",
  4316 => x"00004368",
  4317 => x"00004368",
  4318 => x"00004370",
  4319 => x"00004370",
  4320 => x"00004378",
  4321 => x"00004378",
  4322 => x"00004380",
  4323 => x"00004380",
  4324 => x"00004388",
  4325 => x"00004388",
  4326 => x"00004390",
  4327 => x"00004390",
  4328 => x"00004398",
  4329 => x"00004398",
  4330 => x"000043a0",
  4331 => x"000043a0",
  4332 => x"000043a8",
  4333 => x"000043a8",
  4334 => x"000043b0",
  4335 => x"000043b0",
  4336 => x"000043b8",
  4337 => x"000043b8",
  4338 => x"000043c0",
  4339 => x"000043c0",
  4340 => x"000043c8",
  4341 => x"000043c8",
  4342 => x"000043d0",
  4343 => x"000043d0",
  4344 => x"000043d8",
  4345 => x"000043d8",
  4346 => x"000043e0",
  4347 => x"000043e0",
  4348 => x"000043e8",
  4349 => x"000043e8",
  4350 => x"000043f0",
  4351 => x"000043f0",
  4352 => x"000043f8",
  4353 => x"000043f8",
  4354 => x"00004400",
  4355 => x"00004400",
  4356 => x"00004408",
  4357 => x"00004408",
  4358 => x"00004410",
  4359 => x"00004410",
  4360 => x"00004418",
  4361 => x"00004418",
  4362 => x"00004420",
  4363 => x"00004420",
  4364 => x"00004428",
  4365 => x"00004428",
  4366 => x"00004430",
  4367 => x"00004430",
  4368 => x"00004438",
  4369 => x"00004438",
  4370 => x"00004440",
  4371 => x"00004440",
  4372 => x"00004448",
  4373 => x"00004448",
  4374 => x"00004450",
  4375 => x"00004450",
  4376 => x"00004458",
  4377 => x"00004458",
  4378 => x"00004460",
  4379 => x"00004460",
  4380 => x"00004468",
  4381 => x"00004468",
  4382 => x"00004470",
  4383 => x"00004470",
  4384 => x"00004478",
  4385 => x"00004478",
  4386 => x"00004480",
  4387 => x"00004480",
  4388 => x"00004488",
  4389 => x"00004488",
  4390 => x"00004490",
  4391 => x"00004490",
  4392 => x"00004498",
  4393 => x"00004498",
  4394 => x"000044a0",
  4395 => x"000044a0",
  4396 => x"000044a8",
  4397 => x"000044a8",
  4398 => x"000044b0",
  4399 => x"000044b0",
  4400 => x"000044b8",
  4401 => x"000044b8",
  4402 => x"000044c0",
  4403 => x"000044c0",
  4404 => x"000044c8",
  4405 => x"000044c8",
  4406 => x"000044d0",
  4407 => x"000044d0",
  4408 => x"000044d8",
  4409 => x"000044d8",
  4410 => x"000044e0",
  4411 => x"000044e0",
  4412 => x"000044e8",
  4413 => x"000044e8",
  4414 => x"000044f0",
  4415 => x"000044f0",
  4416 => x"000044f8",
  4417 => x"000044f8",
  4418 => x"00004500",
  4419 => x"00004500",
  4420 => x"00004508",
  4421 => x"00004508",
  4422 => x"00004510",
  4423 => x"00004510",
  4424 => x"00004518",
  4425 => x"00004518",
  4426 => x"00004520",
  4427 => x"00004520",
  4428 => x"00004528",
  4429 => x"00004528",
  4430 => x"00004530",
  4431 => x"00004530",
  4432 => x"00004538",
  4433 => x"00004538",
  4434 => x"00004540",
  4435 => x"00004540",
  4436 => x"00004548",
  4437 => x"00004548",
  4438 => x"00004550",
  4439 => x"00004550",
  4440 => x"00004558",
  4441 => x"00004558",
  4442 => x"00004560",
  4443 => x"00004560",
  4444 => x"00004568",
  4445 => x"00004568",
  4446 => x"00004570",
  4447 => x"00004570",
  4448 => x"00004578",
  4449 => x"00004578",
  4450 => x"00004580",
  4451 => x"00004580",
  4452 => x"00004588",
  4453 => x"00004588",
  4454 => x"00004590",
  4455 => x"00004590",
  4456 => x"00004598",
  4457 => x"00004598",
  4458 => x"000045a0",
  4459 => x"000045a0",
  4460 => x"000045a8",
  4461 => x"000045a8",
  4462 => x"000045b0",
  4463 => x"000045b0",
  4464 => x"000045b8",
  4465 => x"000045b8",
  4466 => x"000045c0",
  4467 => x"000045c0",
  4468 => x"000045c8",
  4469 => x"000045c8",
  4470 => x"000045d0",
  4471 => x"000045d0",
  4472 => x"000045d8",
  4473 => x"000045d8",
  4474 => x"000045e0",
  4475 => x"000045e0",
  4476 => x"000045e8",
  4477 => x"000045e8",
  4478 => x"000045f0",
  4479 => x"000045f0",
  4480 => x"000045f8",
  4481 => x"000045f8",
  4482 => x"00004600",
  4483 => x"00004600",
  4484 => x"00004608",
  4485 => x"00004608",
  4486 => x"00004610",
  4487 => x"00004610",
  4488 => x"00004618",
  4489 => x"00004618",
  4490 => x"00004620",
  4491 => x"00004620",
  4492 => x"00004628",
  4493 => x"00004628",
  4494 => x"00004630",
  4495 => x"00004630",
	--others => x"00dead00" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
