-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0ba7980c",
     3 => x"3a0b0b0b",
     4 => x"a4e10400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0ba5a12d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba7",
   162 => x"84738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8a",
   171 => x"ba2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8b",
   179 => x"ec2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0ba7940c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f9e",
   257 => x"c13f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104a7",
   280 => x"9408802e",
   281 => x"a138a798",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"b7800c82",
   286 => x"a0800bb7",
   287 => x"840c8290",
   288 => x"800bb788",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0bb7",
   292 => x"800cf880",
   293 => x"8082800b",
   294 => x"b7840cf8",
   295 => x"80808480",
   296 => x"0bb7880c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0bb780",
   300 => x"0c80c0a8",
   301 => x"80940bb7",
   302 => x"840c0b0b",
   303 => x"0ba6f00b",
   304 => x"b7880c04",
   305 => x"ff3d0db7",
   306 => x"8c335170",
   307 => x"a338a7a0",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"a7a00c70",
   312 => x"2da7a008",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0bb78c34",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0bb6",
   319 => x"fc08802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0bb6fc",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"ff3d0d8a",
   330 => x"5271f880",
   331 => x"8090800c",
   332 => x"f8808090",
   333 => x"84085183",
   334 => x"fd3f8c08",
   335 => x"028c0cf9",
   336 => x"3d0d800b",
   337 => x"8c08fc05",
   338 => x"0c8c0888",
   339 => x"05088025",
   340 => x"ab388c08",
   341 => x"88050830",
   342 => x"8c088805",
   343 => x"0c800b8c",
   344 => x"08f4050c",
   345 => x"8c08fc05",
   346 => x"08883881",
   347 => x"0b8c08f4",
   348 => x"050c8c08",
   349 => x"f405088c",
   350 => x"08fc050c",
   351 => x"8c088c05",
   352 => x"088025ab",
   353 => x"388c088c",
   354 => x"0508308c",
   355 => x"088c050c",
   356 => x"800b8c08",
   357 => x"f0050c8c",
   358 => x"08fc0508",
   359 => x"8838810b",
   360 => x"8c08f005",
   361 => x"0c8c08f0",
   362 => x"05088c08",
   363 => x"fc050c80",
   364 => x"538c088c",
   365 => x"0508528c",
   366 => x"08880508",
   367 => x"5181a73f",
   368 => x"8008708c",
   369 => x"08f8050c",
   370 => x"548c08fc",
   371 => x"0508802e",
   372 => x"8c388c08",
   373 => x"f8050830",
   374 => x"8c08f805",
   375 => x"0c8c08f8",
   376 => x"05087080",
   377 => x"0c54893d",
   378 => x"0d8c0c04",
   379 => x"8c08028c",
   380 => x"0cfb3d0d",
   381 => x"800b8c08",
   382 => x"fc050c8c",
   383 => x"08880508",
   384 => x"80259338",
   385 => x"8c088805",
   386 => x"08308c08",
   387 => x"88050c81",
   388 => x"0b8c08fc",
   389 => x"050c8c08",
   390 => x"8c050880",
   391 => x"258c388c",
   392 => x"088c0508",
   393 => x"308c088c",
   394 => x"050c8153",
   395 => x"8c088c05",
   396 => x"08528c08",
   397 => x"88050851",
   398 => x"ad3f8008",
   399 => x"708c08f8",
   400 => x"050c548c",
   401 => x"08fc0508",
   402 => x"802e8c38",
   403 => x"8c08f805",
   404 => x"08308c08",
   405 => x"f8050c8c",
   406 => x"08f80508",
   407 => x"70800c54",
   408 => x"873d0d8c",
   409 => x"0c048c08",
   410 => x"028c0cfd",
   411 => x"3d0d810b",
   412 => x"8c08fc05",
   413 => x"0c800b8c",
   414 => x"08f8050c",
   415 => x"8c088c05",
   416 => x"088c0888",
   417 => x"050827ac",
   418 => x"388c08fc",
   419 => x"0508802e",
   420 => x"a338800b",
   421 => x"8c088c05",
   422 => x"08249938",
   423 => x"8c088c05",
   424 => x"08108c08",
   425 => x"8c050c8c",
   426 => x"08fc0508",
   427 => x"108c08fc",
   428 => x"050cc939",
   429 => x"8c08fc05",
   430 => x"08802e80",
   431 => x"c9388c08",
   432 => x"8c05088c",
   433 => x"08880508",
   434 => x"26a1388c",
   435 => x"08880508",
   436 => x"8c088c05",
   437 => x"08318c08",
   438 => x"88050c8c",
   439 => x"08f80508",
   440 => x"8c08fc05",
   441 => x"08078c08",
   442 => x"f8050c8c",
   443 => x"08fc0508",
   444 => x"812a8c08",
   445 => x"fc050c8c",
   446 => x"088c0508",
   447 => x"812a8c08",
   448 => x"8c050cff",
   449 => x"af398c08",
   450 => x"90050880",
   451 => x"2e8f388c",
   452 => x"08880508",
   453 => x"708c08f4",
   454 => x"050c518d",
   455 => x"398c08f8",
   456 => x"0508708c",
   457 => x"08f4050c",
   458 => x"518c08f4",
   459 => x"0508800c",
   460 => x"853d0d8c",
   461 => x"0c04803d",
   462 => x"0d865182",
   463 => x"fd3f8151",
   464 => x"96dc3ffd",
   465 => x"3d0d7553",
   466 => x"84d81308",
   467 => x"802e8a38",
   468 => x"80537280",
   469 => x"0c853d0d",
   470 => x"04818052",
   471 => x"725183d2",
   472 => x"3f800884",
   473 => x"d8140cff",
   474 => x"53800880",
   475 => x"2ee43880",
   476 => x"08549f53",
   477 => x"80747084",
   478 => x"05560cff",
   479 => x"13538073",
   480 => x"24ce3880",
   481 => x"74708405",
   482 => x"560cff13",
   483 => x"53728025",
   484 => x"e338ffbc",
   485 => x"39fd3d0d",
   486 => x"75775553",
   487 => x"9f74278d",
   488 => x"3896730c",
   489 => x"ff527180",
   490 => x"0c853d0d",
   491 => x"0484d813",
   492 => x"08527180",
   493 => x"2e933873",
   494 => x"10101270",
   495 => x"0879720c",
   496 => x"51527180",
   497 => x"0c853d0d",
   498 => x"047251fe",
   499 => x"f63fff52",
   500 => x"8008d338",
   501 => x"84d81308",
   502 => x"74101011",
   503 => x"70087a72",
   504 => x"0c515152",
   505 => x"dd39f93d",
   506 => x"0d797b58",
   507 => x"56769f26",
   508 => x"80e83884",
   509 => x"d8160854",
   510 => x"73802eaa",
   511 => x"38761010",
   512 => x"14700855",
   513 => x"5573802e",
   514 => x"ba388058",
   515 => x"73812e8f",
   516 => x"3873ff2e",
   517 => x"a3388075",
   518 => x"0c765173",
   519 => x"2d805877",
   520 => x"800c893d",
   521 => x"0d047551",
   522 => x"fe993fff",
   523 => x"588008ef",
   524 => x"3884d816",
   525 => x"0854c639",
   526 => x"96760c81",
   527 => x"0b800c89",
   528 => x"3d0d0475",
   529 => x"5181e73f",
   530 => x"76538008",
   531 => x"52755181",
   532 => x"a93f8008",
   533 => x"800c893d",
   534 => x"0d049676",
   535 => x"0cff0b80",
   536 => x"0c893d0d",
   537 => x"04fc3d0d",
   538 => x"76785653",
   539 => x"ff54749f",
   540 => x"26b13884",
   541 => x"d8130852",
   542 => x"71802eae",
   543 => x"38741010",
   544 => x"12700853",
   545 => x"53815471",
   546 => x"802e9838",
   547 => x"825471ff",
   548 => x"2e913883",
   549 => x"5471812e",
   550 => x"8a388073",
   551 => x"0c745171",
   552 => x"2d805473",
   553 => x"800c863d",
   554 => x"0d047251",
   555 => x"fd953f80",
   556 => x"08f13884",
   557 => x"d8130852",
   558 => x"c439ff3d",
   559 => x"0d7352a7",
   560 => x"a40851fe",
   561 => x"a13f833d",
   562 => x"0d04fe3d",
   563 => x"0d755374",
   564 => x"52a7a408",
   565 => x"51fdbe3f",
   566 => x"843d0d04",
   567 => x"803d0da7",
   568 => x"a40851fc",
   569 => x"de3f823d",
   570 => x"0d04ff3d",
   571 => x"0d7352a7",
   572 => x"a40851fe",
   573 => x"f03f833d",
   574 => x"0d04fc3d",
   575 => x"0d800bb7",
   576 => x"980c7852",
   577 => x"77519297",
   578 => x"3f800854",
   579 => x"8008ff2e",
   580 => x"88387380",
   581 => x"0c863d0d",
   582 => x"04b79808",
   583 => x"5574802e",
   584 => x"f1387675",
   585 => x"710c5373",
   586 => x"800c863d",
   587 => x"0d0491ea",
   588 => x"3f04f33d",
   589 => x"0d7f618b",
   590 => x"1170f806",
   591 => x"5c55555e",
   592 => x"72962683",
   593 => x"38905980",
   594 => x"7924747a",
   595 => x"26075380",
   596 => x"5472742e",
   597 => x"09810680",
   598 => x"ca387d51",
   599 => x"8b963f78",
   600 => x"83f72680",
   601 => x"c5387883",
   602 => x"2a701010",
   603 => x"10aee005",
   604 => x"8c110859",
   605 => x"595a7678",
   606 => x"2e83a738",
   607 => x"841708fc",
   608 => x"06568c17",
   609 => x"08881808",
   610 => x"718c120c",
   611 => x"88120c58",
   612 => x"75178411",
   613 => x"08810784",
   614 => x"120c537d",
   615 => x"518ad63f",
   616 => x"88175473",
   617 => x"800c8f3d",
   618 => x"0d047889",
   619 => x"2a79832a",
   620 => x"5b537280",
   621 => x"2ebf3878",
   622 => x"862ab805",
   623 => x"5a847327",
   624 => x"b43880db",
   625 => x"135a9473",
   626 => x"27ab3878",
   627 => x"8c2a80ee",
   628 => x"055a80d4",
   629 => x"73279e38",
   630 => x"788f2a80",
   631 => x"f7055a82",
   632 => x"d4732791",
   633 => x"3878922a",
   634 => x"80fc055a",
   635 => x"8ad47327",
   636 => x"843880fe",
   637 => x"5a791010",
   638 => x"10aee005",
   639 => x"8c110858",
   640 => x"5576752e",
   641 => x"a3388417",
   642 => x"08fc0670",
   643 => x"7a315556",
   644 => x"738f2488",
   645 => x"aa387380",
   646 => x"25fee738",
   647 => x"8c170857",
   648 => x"76752e09",
   649 => x"8106df38",
   650 => x"811a5aae",
   651 => x"f0085776",
   652 => x"aee82e82",
   653 => x"b7388417",
   654 => x"08fc0670",
   655 => x"7a315556",
   656 => x"738f2481",
   657 => x"f338aee8",
   658 => x"0baef40c",
   659 => x"aee80bae",
   660 => x"f00c7380",
   661 => x"25feb938",
   662 => x"83ff7627",
   663 => x"83d23875",
   664 => x"892a7683",
   665 => x"2a555372",
   666 => x"802ebf38",
   667 => x"75862ab8",
   668 => x"05548473",
   669 => x"27b43880",
   670 => x"db135494",
   671 => x"7327ab38",
   672 => x"758c2a80",
   673 => x"ee055480",
   674 => x"d473279e",
   675 => x"38758f2a",
   676 => x"80f70554",
   677 => x"82d47327",
   678 => x"91387592",
   679 => x"2a80fc05",
   680 => x"548ad473",
   681 => x"27843880",
   682 => x"fe547310",
   683 => x"1010aee0",
   684 => x"05881108",
   685 => x"56587478",
   686 => x"2e86af38",
   687 => x"841508fc",
   688 => x"06537573",
   689 => x"278d3888",
   690 => x"15085574",
   691 => x"782e0981",
   692 => x"06ea388c",
   693 => x"1508aee0",
   694 => x"0b840508",
   695 => x"718c1a0c",
   696 => x"76881a0c",
   697 => x"7888130c",
   698 => x"788c180c",
   699 => x"5d587953",
   700 => x"807a2483",
   701 => x"d7387282",
   702 => x"2c81712b",
   703 => x"5c537a7c",
   704 => x"26819338",
   705 => x"7b7b0653",
   706 => x"7282e338",
   707 => x"79fc0684",
   708 => x"055a7a10",
   709 => x"707d0654",
   710 => x"5b7282d2",
   711 => x"38841a5a",
   712 => x"f1398817",
   713 => x"8c110858",
   714 => x"5876782e",
   715 => x"098106fc",
   716 => x"cb38821a",
   717 => x"5afdf439",
   718 => x"78177981",
   719 => x"0784190c",
   720 => x"70aef40c",
   721 => x"70aef00c",
   722 => x"aee80b8c",
   723 => x"120c8c11",
   724 => x"0888120c",
   725 => x"74810784",
   726 => x"120c7411",
   727 => x"75710c51",
   728 => x"537d5187",
   729 => x"903f8817",
   730 => x"54fcb839",
   731 => x"aee00b84",
   732 => x"05087a54",
   733 => x"5c798025",
   734 => x"fefc3882",
   735 => x"cf397a09",
   736 => x"7c0670ae",
   737 => x"e00b8405",
   738 => x"0c5c7a10",
   739 => x"5b7a7c26",
   740 => x"85387a85",
   741 => x"9a38aee0",
   742 => x"0b880508",
   743 => x"70841208",
   744 => x"fc06707c",
   745 => x"317c7226",
   746 => x"8f722507",
   747 => x"57575c5d",
   748 => x"5572802e",
   749 => x"80d73879",
   750 => x"7a16aed8",
   751 => x"081b9011",
   752 => x"5a55575b",
   753 => x"aed408ff",
   754 => x"2e8838a0",
   755 => x"8f13e080",
   756 => x"06577652",
   757 => x"7d51869e",
   758 => x"3f800854",
   759 => x"8008ff2e",
   760 => x"8f388008",
   761 => x"7627828f",
   762 => x"3874aee0",
   763 => x"2e828838",
   764 => x"aee00b88",
   765 => x"05085584",
   766 => x"1508fc06",
   767 => x"707a317a",
   768 => x"72268f72",
   769 => x"25075255",
   770 => x"537283d1",
   771 => x"38747981",
   772 => x"0784170c",
   773 => x"791670ae",
   774 => x"e00b8805",
   775 => x"0c758107",
   776 => x"84120c54",
   777 => x"7e525785",
   778 => x"cc3f8817",
   779 => x"54faf439",
   780 => x"75832a70",
   781 => x"54548074",
   782 => x"24819738",
   783 => x"72822c81",
   784 => x"712baee4",
   785 => x"080770ae",
   786 => x"e00b8405",
   787 => x"0c751010",
   788 => x"10aee005",
   789 => x"88110858",
   790 => x"5a5d5377",
   791 => x"8c180c74",
   792 => x"88180c76",
   793 => x"88190c76",
   794 => x"8c160cfd",
   795 => x"8139797a",
   796 => x"101010ae",
   797 => x"e0057057",
   798 => x"595d8c15",
   799 => x"08577675",
   800 => x"2ea33884",
   801 => x"1708fc06",
   802 => x"707a3155",
   803 => x"56738f24",
   804 => x"83b63873",
   805 => x"802583ea",
   806 => x"388c1708",
   807 => x"5776752e",
   808 => x"098106df",
   809 => x"38881581",
   810 => x"1b708306",
   811 => x"555b5572",
   812 => x"c9387c83",
   813 => x"06537280",
   814 => x"2efdc338",
   815 => x"ff1df819",
   816 => x"595d8818",
   817 => x"08782eea",
   818 => x"38fdbf39",
   819 => x"831a53fc",
   820 => x"a5398314",
   821 => x"70822c81",
   822 => x"712baee4",
   823 => x"080770ae",
   824 => x"e00b8405",
   825 => x"0c761010",
   826 => x"10aee005",
   827 => x"88110859",
   828 => x"5b5e5153",
   829 => x"fee539ae",
   830 => x"a4081758",
   831 => x"8008762e",
   832 => x"818738ae",
   833 => x"d408ff2e",
   834 => x"83d83873",
   835 => x"763118ae",
   836 => x"a40c7387",
   837 => x"06705753",
   838 => x"72802e88",
   839 => x"38887331",
   840 => x"70155556",
   841 => x"76149fff",
   842 => x"06a08071",
   843 => x"31177054",
   844 => x"7f535753",
   845 => x"83c03f80",
   846 => x"08538008",
   847 => x"ff2e8196",
   848 => x"38aea408",
   849 => x"1670aea4",
   850 => x"0c7475ae",
   851 => x"e00b8805",
   852 => x"0c747631",
   853 => x"18708107",
   854 => x"51555658",
   855 => x"7baee02e",
   856 => x"838b3879",
   857 => x"8f2682be",
   858 => x"38810b84",
   859 => x"150c8415",
   860 => x"08fc0670",
   861 => x"7a317a72",
   862 => x"268f7225",
   863 => x"07525553",
   864 => x"72802efd",
   865 => x"883880d5",
   866 => x"3980089f",
   867 => x"ff065372",
   868 => x"fef13877",
   869 => x"aea40cae",
   870 => x"e00b8805",
   871 => x"087b1881",
   872 => x"0784120c",
   873 => x"55aed008",
   874 => x"78278538",
   875 => x"77aed00c",
   876 => x"aecc0878",
   877 => x"27fcc038",
   878 => x"77aecc0c",
   879 => x"841508fc",
   880 => x"06707a31",
   881 => x"7a72268f",
   882 => x"72250752",
   883 => x"55537280",
   884 => x"2efcba38",
   885 => x"88398074",
   886 => x"5456fee5",
   887 => x"397d5182",
   888 => x"943f800b",
   889 => x"800c8f3d",
   890 => x"0d047353",
   891 => x"807424a7",
   892 => x"3872822c",
   893 => x"81712bae",
   894 => x"e4080770",
   895 => x"aee00b84",
   896 => x"050c5d53",
   897 => x"778c180c",
   898 => x"7488180c",
   899 => x"7688190c",
   900 => x"768c160c",
   901 => x"f9d83983",
   902 => x"1470822c",
   903 => x"81712bae",
   904 => x"e4080770",
   905 => x"aee00b84",
   906 => x"050c5e51",
   907 => x"53d6397b",
   908 => x"7b065372",
   909 => x"fcb83884",
   910 => x"1a7b105c",
   911 => x"5af139ff",
   912 => x"1a811151",
   913 => x"5af7e439",
   914 => x"78177981",
   915 => x"0784190c",
   916 => x"8c180888",
   917 => x"1908718c",
   918 => x"120c8812",
   919 => x"0c5970ae",
   920 => x"f40c70ae",
   921 => x"f00caee8",
   922 => x"0b8c120c",
   923 => x"8c110888",
   924 => x"120c7481",
   925 => x"0784120c",
   926 => x"74117571",
   927 => x"0c5153f9",
   928 => x"e0397517",
   929 => x"84110881",
   930 => x"0784120c",
   931 => x"538c1708",
   932 => x"88180871",
   933 => x"8c120c88",
   934 => x"120c587d",
   935 => x"5180d63f",
   936 => x"881754f5",
   937 => x"fe397284",
   938 => x"150cf41a",
   939 => x"f8067084",
   940 => x"1e088106",
   941 => x"07841e0c",
   942 => x"701d545b",
   943 => x"850b8414",
   944 => x"0c850b88",
   945 => x"140c8f7b",
   946 => x"27fdda38",
   947 => x"881c527d",
   948 => x"5182823f",
   949 => x"aee00b88",
   950 => x"0508aea4",
   951 => x"085955fd",
   952 => x"c43977ae",
   953 => x"a40c73ae",
   954 => x"d40cfca6",
   955 => x"39728415",
   956 => x"0cfdb239",
   957 => x"0404fd3d",
   958 => x"0d800bb7",
   959 => x"980c7651",
   960 => x"86b23f80",
   961 => x"08538008",
   962 => x"ff2e8838",
   963 => x"72800c85",
   964 => x"3d0d04b7",
   965 => x"98085473",
   966 => x"802ef138",
   967 => x"7574710c",
   968 => x"5272800c",
   969 => x"853d0d04",
   970 => x"fb3d0d77",
   971 => x"705256c4",
   972 => x"3faee00b",
   973 => x"88050884",
   974 => x"1108fc06",
   975 => x"707b319f",
   976 => x"ef05e080",
   977 => x"06e08005",
   978 => x"565653a0",
   979 => x"80742493",
   980 => x"38805275",
   981 => x"51ff9f3f",
   982 => x"aee80815",
   983 => x"53728008",
   984 => x"2e8f3875",
   985 => x"51ff8e3f",
   986 => x"80537280",
   987 => x"0c873d0d",
   988 => x"04733052",
   989 => x"7551fefe",
   990 => x"3f8008ff",
   991 => x"2ea538ae",
   992 => x"e00b8805",
   993 => x"08757531",
   994 => x"81078412",
   995 => x"0c53aea4",
   996 => x"087431ae",
   997 => x"a40c7551",
   998 => x"fedb3f81",
   999 => x"0b800c87",
  1000 => x"3d0d0480",
  1001 => x"527551fe",
  1002 => x"cd3faee0",
  1003 => x"0b880508",
  1004 => x"80087131",
  1005 => x"56538f75",
  1006 => x"25ffa838",
  1007 => x"8008aed4",
  1008 => x"0831aea4",
  1009 => x"0c748107",
  1010 => x"84140c75",
  1011 => x"51fea63f",
  1012 => x"8053ff96",
  1013 => x"39f63d0d",
  1014 => x"7c7e545b",
  1015 => x"72802e82",
  1016 => x"80387a51",
  1017 => x"fe8e3ff8",
  1018 => x"13841108",
  1019 => x"70fe0670",
  1020 => x"13841108",
  1021 => x"fc065d58",
  1022 => x"595458ae",
  1023 => x"e808752e",
  1024 => x"82d83878",
  1025 => x"84160c80",
  1026 => x"73810654",
  1027 => x"5a727a2e",
  1028 => x"81d33878",
  1029 => x"15841108",
  1030 => x"81065153",
  1031 => x"729f3878",
  1032 => x"17577981",
  1033 => x"e3388815",
  1034 => x"085372ae",
  1035 => x"e82e82f1",
  1036 => x"388c1508",
  1037 => x"708c150c",
  1038 => x"7388120c",
  1039 => x"56768107",
  1040 => x"84190c76",
  1041 => x"1877710c",
  1042 => x"53798190",
  1043 => x"3883ff77",
  1044 => x"2781c638",
  1045 => x"76892a77",
  1046 => x"832a5653",
  1047 => x"72802ebf",
  1048 => x"3876862a",
  1049 => x"b8055584",
  1050 => x"7327b438",
  1051 => x"80db1355",
  1052 => x"947327ab",
  1053 => x"38768c2a",
  1054 => x"80ee0555",
  1055 => x"80d47327",
  1056 => x"9e38768f",
  1057 => x"2a80f705",
  1058 => x"5582d473",
  1059 => x"27913876",
  1060 => x"922a80fc",
  1061 => x"05558ad4",
  1062 => x"73278438",
  1063 => x"80fe5574",
  1064 => x"101010ae",
  1065 => x"e0058811",
  1066 => x"08555673",
  1067 => x"762e82a9",
  1068 => x"38841408",
  1069 => x"fc065376",
  1070 => x"73278d38",
  1071 => x"88140854",
  1072 => x"73762e09",
  1073 => x"8106ea38",
  1074 => x"8c140870",
  1075 => x"8c1a0c74",
  1076 => x"881a0c78",
  1077 => x"88120c56",
  1078 => x"778c150c",
  1079 => x"7a51fc95",
  1080 => x"3f8c3d0d",
  1081 => x"04770878",
  1082 => x"71315977",
  1083 => x"05881908",
  1084 => x"545772ae",
  1085 => x"e82e80dd",
  1086 => x"388c1808",
  1087 => x"708c150c",
  1088 => x"7388120c",
  1089 => x"56fe8c39",
  1090 => x"8815088c",
  1091 => x"1608708c",
  1092 => x"130c5788",
  1093 => x"170cfea5",
  1094 => x"3976832a",
  1095 => x"70545580",
  1096 => x"75248192",
  1097 => x"3872822c",
  1098 => x"81712bae",
  1099 => x"e40807ae",
  1100 => x"e00b8405",
  1101 => x"0c537410",
  1102 => x"1010aee0",
  1103 => x"05881108",
  1104 => x"5556758c",
  1105 => x"190c7388",
  1106 => x"190c7788",
  1107 => x"170c778c",
  1108 => x"150cff88",
  1109 => x"39815afd",
  1110 => x"ba397817",
  1111 => x"73810654",
  1112 => x"57729838",
  1113 => x"77087871",
  1114 => x"31597705",
  1115 => x"8c190888",
  1116 => x"1a08718c",
  1117 => x"120c8812",
  1118 => x"0c575776",
  1119 => x"81078419",
  1120 => x"0c77aee0",
  1121 => x"0b88050c",
  1122 => x"aedc0877",
  1123 => x"26fecd38",
  1124 => x"aed80852",
  1125 => x"7a51fb90",
  1126 => x"3f7a51fa",
  1127 => x"d83ffec1",
  1128 => x"3981788c",
  1129 => x"150c7888",
  1130 => x"150c738c",
  1131 => x"1a0c7388",
  1132 => x"1a0c5afd",
  1133 => x"88398315",
  1134 => x"70822c81",
  1135 => x"712baee4",
  1136 => x"0807aee0",
  1137 => x"0b84050c",
  1138 => x"51537410",
  1139 => x"1010aee0",
  1140 => x"05881108",
  1141 => x"5556feea",
  1142 => x"39745380",
  1143 => x"7524a538",
  1144 => x"72822c81",
  1145 => x"712baee4",
  1146 => x"0807aee0",
  1147 => x"0b84050c",
  1148 => x"53758c19",
  1149 => x"0c738819",
  1150 => x"0c778817",
  1151 => x"0c778c15",
  1152 => x"0cfdd939",
  1153 => x"83157082",
  1154 => x"2c81712b",
  1155 => x"aee40807",
  1156 => x"aee00b84",
  1157 => x"050c5153",
  1158 => x"d839810b",
  1159 => x"800c0480",
  1160 => x"3d0d7281",
  1161 => x"2e893880",
  1162 => x"0b800c82",
  1163 => x"3d0d0473",
  1164 => x"5180eb3f",
  1165 => x"fe3d0db7",
  1166 => x"90085170",
  1167 => x"8838b79c",
  1168 => x"70b7900c",
  1169 => x"51707512",
  1170 => x"5252ff53",
  1171 => x"7087fb80",
  1172 => x"80268738",
  1173 => x"70b7900c",
  1174 => x"71537280",
  1175 => x"0c843d0d",
  1176 => x"04fd3d0d",
  1177 => x"800ba798",
  1178 => x"08545472",
  1179 => x"812e9838",
  1180 => x"73b7940c",
  1181 => x"e3e93fe3",
  1182 => x"873fb6e8",
  1183 => x"528151e5",
  1184 => x"a33f8008",
  1185 => x"519e3f72",
  1186 => x"b7940ce3",
  1187 => x"d23fe2f0",
  1188 => x"3fb6e852",
  1189 => x"8151e58c",
  1190 => x"3f800851",
  1191 => x"873f00ff",
  1192 => x"3900ff39",
  1193 => x"f73d0d7b",
  1194 => x"a7a40882",
  1195 => x"c811085a",
  1196 => x"545a7780",
  1197 => x"2e80d938",
  1198 => x"81881884",
  1199 => x"1908ff05",
  1200 => x"81712b59",
  1201 => x"55598074",
  1202 => x"2480e938",
  1203 => x"807424b5",
  1204 => x"3873822b",
  1205 => x"78118805",
  1206 => x"56568180",
  1207 => x"19087706",
  1208 => x"5372802e",
  1209 => x"b5387816",
  1210 => x"70085353",
  1211 => x"79517408",
  1212 => x"53722dff",
  1213 => x"14fc17fc",
  1214 => x"1779812c",
  1215 => x"5a575754",
  1216 => x"738025d6",
  1217 => x"38770858",
  1218 => x"77ffad38",
  1219 => x"a7a40853",
  1220 => x"bc1308a5",
  1221 => x"387951ff",
  1222 => x"853f7408",
  1223 => x"53722dff",
  1224 => x"14fc17fc",
  1225 => x"1779812c",
  1226 => x"5a575754",
  1227 => x"738025ff",
  1228 => x"a938d239",
  1229 => x"8057ff94",
  1230 => x"397251bc",
  1231 => x"13085372",
  1232 => x"2d7951fe",
  1233 => x"d93fff3d",
  1234 => x"0db6f00b",
  1235 => x"fc057008",
  1236 => x"525270ff",
  1237 => x"2e913870",
  1238 => x"2dfc1270",
  1239 => x"08525270",
  1240 => x"ff2e0981",
  1241 => x"06f13883",
  1242 => x"3d0d0404",
  1243 => x"e2d63f04",
  1244 => x"00000040",
  1245 => x"43000000",
  1246 => x"64756d6d",
  1247 => x"792e6578",
  1248 => x"65000000",
  1249 => x"00ffffff",
  1250 => x"ff00ffff",
  1251 => x"ffff00ff",
  1252 => x"ffffff00",
  1253 => x"00000000",
  1254 => x"00000000",
  1255 => x"00000000",
  1256 => x"00001b78",
  1257 => x"000013a8",
  1258 => x"00000000",
  1259 => x"00001610",
  1260 => x"0000166c",
  1261 => x"000016c8",
  1262 => x"00000000",
  1263 => x"00000000",
  1264 => x"00000000",
  1265 => x"00000000",
  1266 => x"00000000",
  1267 => x"00000000",
  1268 => x"00000000",
  1269 => x"00000000",
  1270 => x"00000000",
  1271 => x"00001374",
  1272 => x"00000000",
  1273 => x"00000000",
  1274 => x"00000000",
  1275 => x"00000000",
  1276 => x"00000000",
  1277 => x"00000000",
  1278 => x"00000000",
  1279 => x"00000000",
  1280 => x"00000000",
  1281 => x"00000000",
  1282 => x"00000000",
  1283 => x"00000000",
  1284 => x"00000000",
  1285 => x"00000000",
  1286 => x"00000000",
  1287 => x"00000000",
  1288 => x"00000000",
  1289 => x"00000000",
  1290 => x"00000000",
  1291 => x"00000000",
  1292 => x"00000000",
  1293 => x"00000000",
  1294 => x"00000000",
  1295 => x"00000000",
  1296 => x"00000000",
  1297 => x"00000000",
  1298 => x"00000000",
  1299 => x"00000000",
  1300 => x"00000001",
  1301 => x"330eabcd",
  1302 => x"1234e66d",
  1303 => x"deec0005",
  1304 => x"000b0000",
  1305 => x"00000000",
  1306 => x"00000000",
  1307 => x"00000000",
  1308 => x"00000000",
  1309 => x"00000000",
  1310 => x"00000000",
  1311 => x"00000000",
  1312 => x"00000000",
  1313 => x"00000000",
  1314 => x"00000000",
  1315 => x"00000000",
  1316 => x"00000000",
  1317 => x"00000000",
  1318 => x"00000000",
  1319 => x"00000000",
  1320 => x"00000000",
  1321 => x"00000000",
  1322 => x"00000000",
  1323 => x"00000000",
  1324 => x"00000000",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00000000",
  1329 => x"00000000",
  1330 => x"00000000",
  1331 => x"00000000",
  1332 => x"00000000",
  1333 => x"00000000",
  1334 => x"00000000",
  1335 => x"00000000",
  1336 => x"00000000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"00000000",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"00000000",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000000",
  1404 => x"00000000",
  1405 => x"00000000",
  1406 => x"00000000",
  1407 => x"00000000",
  1408 => x"00000000",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00000000",
  1414 => x"00000000",
  1415 => x"00000000",
  1416 => x"00000000",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"00000000",
  1420 => x"00000000",
  1421 => x"00000000",
  1422 => x"00000000",
  1423 => x"00000000",
  1424 => x"00000000",
  1425 => x"00000000",
  1426 => x"00000000",
  1427 => x"00000000",
  1428 => x"00000000",
  1429 => x"00000000",
  1430 => x"00000000",
  1431 => x"00000000",
  1432 => x"00000000",
  1433 => x"00000000",
  1434 => x"00000000",
  1435 => x"00000000",
  1436 => x"00000000",
  1437 => x"00000000",
  1438 => x"00000000",
  1439 => x"00000000",
  1440 => x"00000000",
  1441 => x"00000000",
  1442 => x"00000000",
  1443 => x"00000000",
  1444 => x"00000000",
  1445 => x"00000000",
  1446 => x"00000000",
  1447 => x"00000000",
  1448 => x"00000000",
  1449 => x"00000000",
  1450 => x"00000000",
  1451 => x"00000000",
  1452 => x"00000000",
  1453 => x"00000000",
  1454 => x"00000000",
  1455 => x"00000000",
  1456 => x"00000000",
  1457 => x"00000000",
  1458 => x"00000000",
  1459 => x"00000000",
  1460 => x"00000000",
  1461 => x"00000000",
  1462 => x"00000000",
  1463 => x"00000000",
  1464 => x"00000000",
  1465 => x"00000000",
  1466 => x"00000000",
  1467 => x"00000000",
  1468 => x"00000000",
  1469 => x"00000000",
  1470 => x"00000000",
  1471 => x"00000000",
  1472 => x"00000000",
  1473 => x"00000000",
  1474 => x"00000000",
  1475 => x"00000000",
  1476 => x"00000000",
  1477 => x"00000000",
  1478 => x"00000000",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000000",
  1483 => x"00000000",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"00000000",
  1492 => x"00000000",
  1493 => x"ffffffff",
  1494 => x"00000000",
  1495 => x"00020000",
  1496 => x"00000000",
  1497 => x"00000000",
  1498 => x"00001760",
  1499 => x"00001760",
  1500 => x"00001768",
  1501 => x"00001768",
  1502 => x"00001770",
  1503 => x"00001770",
  1504 => x"00001778",
  1505 => x"00001778",
  1506 => x"00001780",
  1507 => x"00001780",
  1508 => x"00001788",
  1509 => x"00001788",
  1510 => x"00001790",
  1511 => x"00001790",
  1512 => x"00001798",
  1513 => x"00001798",
  1514 => x"000017a0",
  1515 => x"000017a0",
  1516 => x"000017a8",
  1517 => x"000017a8",
  1518 => x"000017b0",
  1519 => x"000017b0",
  1520 => x"000017b8",
  1521 => x"000017b8",
  1522 => x"000017c0",
  1523 => x"000017c0",
  1524 => x"000017c8",
  1525 => x"000017c8",
  1526 => x"000017d0",
  1527 => x"000017d0",
  1528 => x"000017d8",
  1529 => x"000017d8",
  1530 => x"000017e0",
  1531 => x"000017e0",
  1532 => x"000017e8",
  1533 => x"000017e8",
  1534 => x"000017f0",
  1535 => x"000017f0",
  1536 => x"000017f8",
  1537 => x"000017f8",
  1538 => x"00001800",
  1539 => x"00001800",
  1540 => x"00001808",
  1541 => x"00001808",
  1542 => x"00001810",
  1543 => x"00001810",
  1544 => x"00001818",
  1545 => x"00001818",
  1546 => x"00001820",
  1547 => x"00001820",
  1548 => x"00001828",
  1549 => x"00001828",
  1550 => x"00001830",
  1551 => x"00001830",
  1552 => x"00001838",
  1553 => x"00001838",
  1554 => x"00001840",
  1555 => x"00001840",
  1556 => x"00001848",
  1557 => x"00001848",
  1558 => x"00001850",
  1559 => x"00001850",
  1560 => x"00001858",
  1561 => x"00001858",
  1562 => x"00001860",
  1563 => x"00001860",
  1564 => x"00001868",
  1565 => x"00001868",
  1566 => x"00001870",
  1567 => x"00001870",
  1568 => x"00001878",
  1569 => x"00001878",
  1570 => x"00001880",
  1571 => x"00001880",
  1572 => x"00001888",
  1573 => x"00001888",
  1574 => x"00001890",
  1575 => x"00001890",
  1576 => x"00001898",
  1577 => x"00001898",
  1578 => x"000018a0",
  1579 => x"000018a0",
  1580 => x"000018a8",
  1581 => x"000018a8",
  1582 => x"000018b0",
  1583 => x"000018b0",
  1584 => x"000018b8",
  1585 => x"000018b8",
  1586 => x"000018c0",
  1587 => x"000018c0",
  1588 => x"000018c8",
  1589 => x"000018c8",
  1590 => x"000018d0",
  1591 => x"000018d0",
  1592 => x"000018d8",
  1593 => x"000018d8",
  1594 => x"000018e0",
  1595 => x"000018e0",
  1596 => x"000018e8",
  1597 => x"000018e8",
  1598 => x"000018f0",
  1599 => x"000018f0",
  1600 => x"000018f8",
  1601 => x"000018f8",
  1602 => x"00001900",
  1603 => x"00001900",
  1604 => x"00001908",
  1605 => x"00001908",
  1606 => x"00001910",
  1607 => x"00001910",
  1608 => x"00001918",
  1609 => x"00001918",
  1610 => x"00001920",
  1611 => x"00001920",
  1612 => x"00001928",
  1613 => x"00001928",
  1614 => x"00001930",
  1615 => x"00001930",
  1616 => x"00001938",
  1617 => x"00001938",
  1618 => x"00001940",
  1619 => x"00001940",
  1620 => x"00001948",
  1621 => x"00001948",
  1622 => x"00001950",
  1623 => x"00001950",
  1624 => x"00001958",
  1625 => x"00001958",
  1626 => x"00001960",
  1627 => x"00001960",
  1628 => x"00001968",
  1629 => x"00001968",
  1630 => x"00001970",
  1631 => x"00001970",
  1632 => x"00001978",
  1633 => x"00001978",
  1634 => x"00001980",
  1635 => x"00001980",
  1636 => x"00001988",
  1637 => x"00001988",
  1638 => x"00001990",
  1639 => x"00001990",
  1640 => x"00001998",
  1641 => x"00001998",
  1642 => x"000019a0",
  1643 => x"000019a0",
  1644 => x"000019a8",
  1645 => x"000019a8",
  1646 => x"000019b0",
  1647 => x"000019b0",
  1648 => x"000019b8",
  1649 => x"000019b8",
  1650 => x"000019c0",
  1651 => x"000019c0",
  1652 => x"000019c8",
  1653 => x"000019c8",
  1654 => x"000019d0",
  1655 => x"000019d0",
  1656 => x"000019d8",
  1657 => x"000019d8",
  1658 => x"000019e0",
  1659 => x"000019e0",
  1660 => x"000019e8",
  1661 => x"000019e8",
  1662 => x"000019f0",
  1663 => x"000019f0",
  1664 => x"000019f8",
  1665 => x"000019f8",
  1666 => x"00001a00",
  1667 => x"00001a00",
  1668 => x"00001a08",
  1669 => x"00001a08",
  1670 => x"00001a10",
  1671 => x"00001a10",
  1672 => x"00001a18",
  1673 => x"00001a18",
  1674 => x"00001a20",
  1675 => x"00001a20",
  1676 => x"00001a28",
  1677 => x"00001a28",
  1678 => x"00001a30",
  1679 => x"00001a30",
  1680 => x"00001a38",
  1681 => x"00001a38",
  1682 => x"00001a40",
  1683 => x"00001a40",
  1684 => x"00001a48",
  1685 => x"00001a48",
  1686 => x"00001a50",
  1687 => x"00001a50",
  1688 => x"00001a58",
  1689 => x"00001a58",
  1690 => x"00001a60",
  1691 => x"00001a60",
  1692 => x"00001a68",
  1693 => x"00001a68",
  1694 => x"00001a70",
  1695 => x"00001a70",
  1696 => x"00001a78",
  1697 => x"00001a78",
  1698 => x"00001a80",
  1699 => x"00001a80",
  1700 => x"00001a88",
  1701 => x"00001a88",
  1702 => x"00001a90",
  1703 => x"00001a90",
  1704 => x"00001a98",
  1705 => x"00001a98",
  1706 => x"00001aa0",
  1707 => x"00001aa0",
  1708 => x"00001aa8",
  1709 => x"00001aa8",
  1710 => x"00001ab0",
  1711 => x"00001ab0",
  1712 => x"00001ab8",
  1713 => x"00001ab8",
  1714 => x"00001ac0",
  1715 => x"00001ac0",
  1716 => x"00001ac8",
  1717 => x"00001ac8",
  1718 => x"00001ad0",
  1719 => x"00001ad0",
  1720 => x"00001ad8",
  1721 => x"00001ad8",
  1722 => x"00001ae0",
  1723 => x"00001ae0",
  1724 => x"00001ae8",
  1725 => x"00001ae8",
  1726 => x"00001af0",
  1727 => x"00001af0",
  1728 => x"00001af8",
  1729 => x"00001af8",
  1730 => x"00001b00",
  1731 => x"00001b00",
  1732 => x"00001b08",
  1733 => x"00001b08",
  1734 => x"00001b10",
  1735 => x"00001b10",
  1736 => x"00001b18",
  1737 => x"00001b18",
  1738 => x"00001b20",
  1739 => x"00001b20",
  1740 => x"00001b28",
  1741 => x"00001b28",
  1742 => x"00001b30",
  1743 => x"00001b30",
  1744 => x"00001b38",
  1745 => x"00001b38",
  1746 => x"00001b40",
  1747 => x"00001b40",
  1748 => x"00001b48",
  1749 => x"00001b48",
  1750 => x"00001b50",
  1751 => x"00001b50",
  1752 => x"00001b58",
  1753 => x"00001b58",
  1754 => x"00001378",
  1755 => x"ffffffff",
  1756 => x"00000000",
  1757 => x"ffffffff",
  1758 => x"00000000",
  1759 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
