# ====================================================================
#
#      phi_opencores_ethmac_drivers.cdl
#
#      Ethernet drivers - support for Opencores ethermac controller
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Gaisler Research, (Konrad Eisele<eiselekd@web.de>)
# Contributors:	  Zylin AS, (Edgar Grimberg<edgar.grimberg@zylin.com>)
# Date:           2005-01-20
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ZPU_OPENCORES_PHI {

    display       "PHI opencores ethernet driver"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_ZYLIN_ZPU_PHI
    
    requires      CYGPKG_DEVS_ETH_OPENCORES_ETHERMAC
    description   "Ethernet driver for ethermac in on a Zylin Phi Board."

    include_dir   cyg/io
    compile       -library=libextras.a if_opencores.c

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_OPENCORES_ETHERMAC_INL <cyg/io/devs_eth_zpu_opencores_phi.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_OPENCORES_ETHERMAC_CFG <pkgconf/devs_eth_zpu_opencores_phi.h>"
        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }
    
    # Arguably this should do in the generic package
    # but then there is a logic loop so you can never enable it.

    cdl_interface CYGINT_DEVS_ETH_OPENCORES_ETHERMAC_REQUIRED {
        display   "opencores ethermac driver required"
    }

    cdl_component CYGPKG_DEVS_ETH_ZPU_OPENCORES_PHI_ETH0 {
        display       "Ethernet port 0 driver"
        flavor        bool
        default_value 1

        implements    CYGHWR_NET_DRIVERS
        implements    CYGHWR_NET_DRIVER_ETH0
        implements    CYGINT_DEVS_ETH_OPENCORES_ETHERMAC_REQUIRED
    
        cdl_option CYGPKG_DEVS_ETH_ZPU_OPENCORES_PHI_ETH0_NAME {
            display       "Device name for the ethernet driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                          This option sets the name of the ethernet device for the
                          ethernet port."
       }
    
        cdl_option CYGPKG_DEVS_ETH_ZPU_OPENCORES_PHI_ETH0_ESA {
            display       "The ethernet station address (MAC)"
            flavor        data
            default_value {"{0x00, 0x00, 0x5E, 0x21, 0x00, 0x01}"}
            description   "A static ethernet station address. 
                          Caution: Booting two systems with the same MAC on the same
                          network, will cause severe conflicts."
       }
    }

    cdl_component CYGPKG_DEVS_ETH_ZPU_OPENCORES_PHI_OPTIONS {
        display "Opencores ethermac driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_ZPU_OPENCORES_PHI_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the opencores ethermac driver package.
                These flags are used in addition
                to the set of global flags."
        }
    }

}

# EOF phi_opencores_ethmac_drivers.cdl
