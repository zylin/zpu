-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0b91800c",
     3 => x"3a0b0b0b",
     4 => x"8ec60400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b8f862d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b90",
   162 => x"ec738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8a",
   171 => x"ca2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8b",
   179 => x"fc2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0b90fc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f88",
   257 => x"a63f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"53510490",
   280 => x"fc08802e",
   281 => x"a1389180",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"98a40c82",
   286 => x"a0800b98",
   287 => x"a80c8290",
   288 => x"800b98ac",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0b98",
   292 => x"a40cf880",
   293 => x"8082800b",
   294 => x"98a80cf8",
   295 => x"80808480",
   296 => x"0b98ac0c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0b98a4",
   300 => x"0c80c0a8",
   301 => x"80940b98",
   302 => x"a80c0b0b",
   303 => x"0b90d80b",
   304 => x"98ac0c04",
   305 => x"ff3d0d98",
   306 => x"b0335170",
   307 => x"a3389188",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"91880c70",
   312 => x"2d918808",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0b98b034",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0b98",
   319 => x"a008802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0b98a0",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"ff3d0d8c",
   330 => x"80838052",
   331 => x"71f88080",
   332 => x"90840c71",
   333 => x"9f2a7210",
   334 => x"0770f880",
   335 => x"8090840c",
   336 => x"709f2a71",
   337 => x"10075152",
   338 => x"e3398c08",
   339 => x"028c0cf9",
   340 => x"3d0d800b",
   341 => x"8c08fc05",
   342 => x"0c8c0888",
   343 => x"05088025",
   344 => x"ab388c08",
   345 => x"88050830",
   346 => x"8c088805",
   347 => x"0c800b8c",
   348 => x"08f4050c",
   349 => x"8c08fc05",
   350 => x"08883881",
   351 => x"0b8c08f4",
   352 => x"050c8c08",
   353 => x"f405088c",
   354 => x"08fc050c",
   355 => x"8c088c05",
   356 => x"088025ab",
   357 => x"388c088c",
   358 => x"0508308c",
   359 => x"088c050c",
   360 => x"800b8c08",
   361 => x"f0050c8c",
   362 => x"08fc0508",
   363 => x"8838810b",
   364 => x"8c08f005",
   365 => x"0c8c08f0",
   366 => x"05088c08",
   367 => x"fc050c80",
   368 => x"538c088c",
   369 => x"0508528c",
   370 => x"08880508",
   371 => x"5181a73f",
   372 => x"8008708c",
   373 => x"08f8050c",
   374 => x"548c08fc",
   375 => x"0508802e",
   376 => x"8c388c08",
   377 => x"f8050830",
   378 => x"8c08f805",
   379 => x"0c8c08f8",
   380 => x"05087080",
   381 => x"0c54893d",
   382 => x"0d8c0c04",
   383 => x"8c08028c",
   384 => x"0cfb3d0d",
   385 => x"800b8c08",
   386 => x"fc050c8c",
   387 => x"08880508",
   388 => x"80259338",
   389 => x"8c088805",
   390 => x"08308c08",
   391 => x"88050c81",
   392 => x"0b8c08fc",
   393 => x"050c8c08",
   394 => x"8c050880",
   395 => x"258c388c",
   396 => x"088c0508",
   397 => x"308c088c",
   398 => x"050c8153",
   399 => x"8c088c05",
   400 => x"08528c08",
   401 => x"88050851",
   402 => x"ad3f8008",
   403 => x"708c08f8",
   404 => x"050c548c",
   405 => x"08fc0508",
   406 => x"802e8c38",
   407 => x"8c08f805",
   408 => x"08308c08",
   409 => x"f8050c8c",
   410 => x"08f80508",
   411 => x"70800c54",
   412 => x"873d0d8c",
   413 => x"0c048c08",
   414 => x"028c0cfd",
   415 => x"3d0d810b",
   416 => x"8c08fc05",
   417 => x"0c800b8c",
   418 => x"08f8050c",
   419 => x"8c088c05",
   420 => x"088c0888",
   421 => x"050827ac",
   422 => x"388c08fc",
   423 => x"0508802e",
   424 => x"a338800b",
   425 => x"8c088c05",
   426 => x"08249938",
   427 => x"8c088c05",
   428 => x"08108c08",
   429 => x"8c050c8c",
   430 => x"08fc0508",
   431 => x"108c08fc",
   432 => x"050cc939",
   433 => x"8c08fc05",
   434 => x"08802e80",
   435 => x"c9388c08",
   436 => x"8c05088c",
   437 => x"08880508",
   438 => x"26a1388c",
   439 => x"08880508",
   440 => x"8c088c05",
   441 => x"08318c08",
   442 => x"88050c8c",
   443 => x"08f80508",
   444 => x"8c08fc05",
   445 => x"08078c08",
   446 => x"f8050c8c",
   447 => x"08fc0508",
   448 => x"812a8c08",
   449 => x"fc050c8c",
   450 => x"088c0508",
   451 => x"812a8c08",
   452 => x"8c050cff",
   453 => x"af398c08",
   454 => x"90050880",
   455 => x"2e8f388c",
   456 => x"08880508",
   457 => x"708c08f4",
   458 => x"050c518d",
   459 => x"398c08f8",
   460 => x"0508708c",
   461 => x"08f4050c",
   462 => x"518c08f4",
   463 => x"0508800c",
   464 => x"853d0d8c",
   465 => x"0c04fd3d",
   466 => x"0d800b91",
   467 => x"80085454",
   468 => x"72812e98",
   469 => x"387398b4",
   470 => x"0cfa843f",
   471 => x"f9a23f91",
   472 => x"8c528151",
   473 => x"fbbe3f80",
   474 => x"08519e3f",
   475 => x"7298b40c",
   476 => x"f9ed3ff9",
   477 => x"8b3f918c",
   478 => x"528151fb",
   479 => x"a73f8008",
   480 => x"51873f00",
   481 => x"ff3900ff",
   482 => x"39f73d0d",
   483 => x"7b919008",
   484 => x"82c81108",
   485 => x"5a545a77",
   486 => x"802e80d9",
   487 => x"38818818",
   488 => x"841908ff",
   489 => x"0581712b",
   490 => x"59555980",
   491 => x"742480e9",
   492 => x"38807424",
   493 => x"b5387382",
   494 => x"2b781188",
   495 => x"05565681",
   496 => x"80190877",
   497 => x"06537280",
   498 => x"2eb53878",
   499 => x"16700853",
   500 => x"53795174",
   501 => x"0853722d",
   502 => x"ff14fc17",
   503 => x"fc177981",
   504 => x"2c5a5757",
   505 => x"54738025",
   506 => x"d6387708",
   507 => x"5877ffad",
   508 => x"38919008",
   509 => x"53bc1308",
   510 => x"a5387951",
   511 => x"ff853f74",
   512 => x"0853722d",
   513 => x"ff14fc17",
   514 => x"fc177981",
   515 => x"2c5a5757",
   516 => x"54738025",
   517 => x"ffa938d2",
   518 => x"398057ff",
   519 => x"94397251",
   520 => x"bc130853",
   521 => x"722d7951",
   522 => x"fed93fff",
   523 => x"3d0d9894",
   524 => x"0bfc0570",
   525 => x"08525270",
   526 => x"ff2e9138",
   527 => x"702dfc12",
   528 => x"70085252",
   529 => x"70ff2e09",
   530 => x"8106f138",
   531 => x"833d0d04",
   532 => x"04f8f13f",
   533 => x"04000000",
   534 => x"00000040",
   535 => x"64756d6d",
   536 => x"792e6578",
   537 => x"65000000",
   538 => x"43000000",
   539 => x"00ffffff",
   540 => x"ff00ffff",
   541 => x"ffff00ff",
   542 => x"ffffff00",
   543 => x"00000000",
   544 => x"00000000",
   545 => x"00000000",
   546 => x"00000c1c",
   547 => x"0000085c",
   548 => x"00000894",
   549 => x"00000000",
   550 => x"00000afc",
   551 => x"00000b58",
   552 => x"00000bb4",
   553 => x"00000000",
   554 => x"00000000",
   555 => x"00000000",
   556 => x"00000000",
   557 => x"00000000",
   558 => x"00000000",
   559 => x"00000000",
   560 => x"00000000",
   561 => x"00000000",
   562 => x"00000868",
   563 => x"00000000",
   564 => x"00000000",
   565 => x"00000000",
   566 => x"00000000",
   567 => x"00000000",
   568 => x"00000000",
   569 => x"00000000",
   570 => x"00000000",
   571 => x"00000000",
   572 => x"00000000",
   573 => x"00000000",
   574 => x"00000000",
   575 => x"00000000",
   576 => x"00000000",
   577 => x"00000000",
   578 => x"00000000",
   579 => x"00000000",
   580 => x"00000000",
   581 => x"00000000",
   582 => x"00000000",
   583 => x"00000000",
   584 => x"00000000",
   585 => x"00000000",
   586 => x"00000000",
   587 => x"00000000",
   588 => x"00000000",
   589 => x"00000000",
   590 => x"00000000",
   591 => x"00000001",
   592 => x"330eabcd",
   593 => x"1234e66d",
   594 => x"deec0005",
   595 => x"000b0000",
   596 => x"00000000",
   597 => x"00000000",
   598 => x"00000000",
   599 => x"00000000",
   600 => x"00000000",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000000",
   605 => x"00000000",
   606 => x"00000000",
   607 => x"00000000",
   608 => x"00000000",
   609 => x"00000000",
   610 => x"00000000",
   611 => x"00000000",
   612 => x"00000000",
   613 => x"00000000",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000000",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000000",
   653 => x"00000000",
   654 => x"00000000",
   655 => x"00000000",
   656 => x"00000000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"ffffffff",
   773 => x"00000000",
   774 => x"ffffffff",
   775 => x"00000000",
   776 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
