-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0bb38c0c",
     3 => x"3a0b0b0b",
     4 => x"a6be0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0ba6fe2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bb2",
   162 => x"f8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0ba1",
   171 => x"a92d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0ba2",
   179 => x"db2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bb3880c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33fa0",
   257 => x"9e3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104b3",
   280 => x"8808802e",
   281 => x"a138b38c",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"bac80c82",
   286 => x"a0800bba",
   287 => x"cc0c8290",
   288 => x"800bbad0",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0bba",
   292 => x"c80cf880",
   293 => x"8082800b",
   294 => x"bacc0cf8",
   295 => x"80808480",
   296 => x"0bbad00c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0bbac8",
   300 => x"0c80c0a8",
   301 => x"80940bba",
   302 => x"cc0c0b0b",
   303 => x"0ba8d00b",
   304 => x"bad00c04",
   305 => x"ff3d0dba",
   306 => x"d4335170",
   307 => x"a338b394",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"b3940c70",
   312 => x"2db39408",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0bbad434",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0bba",
   319 => x"c408802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0bbac4",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"f83d0d7a",
   330 => x"7c595380",
   331 => x"73565776",
   332 => x"732480dc",
   333 => x"38771754",
   334 => x"8a527451",
   335 => x"96c63f80",
   336 => x"08b00553",
   337 => x"72743481",
   338 => x"17578a52",
   339 => x"7451968f",
   340 => x"3f800855",
   341 => x"8008de38",
   342 => x"8008779f",
   343 => x"2a187081",
   344 => x"2c5b5656",
   345 => x"8079259e",
   346 => x"387717ff",
   347 => x"05557518",
   348 => x"70335553",
   349 => x"74337334",
   350 => x"73753481",
   351 => x"16ff1656",
   352 => x"56787624",
   353 => x"e9387618",
   354 => x"56807634",
   355 => x"8a3d0d04",
   356 => x"ad787081",
   357 => x"055a3472",
   358 => x"30781855",
   359 => x"558a5274",
   360 => x"5195e13f",
   361 => x"8008b005",
   362 => x"53727434",
   363 => x"8117578a",
   364 => x"52745195",
   365 => x"aa3f8008",
   366 => x"558008fe",
   367 => x"f838ff98",
   368 => x"39f93d0d",
   369 => x"79707133",
   370 => x"7081ff06",
   371 => x"54555555",
   372 => x"70802eb0",
   373 => x"38b3ac08",
   374 => x"527281ff",
   375 => x"06811555",
   376 => x"53728a2e",
   377 => x"80f13884",
   378 => x"12087082",
   379 => x"2a810652",
   380 => x"5770802e",
   381 => x"f2387272",
   382 => x"0c733370",
   383 => x"81ff0659",
   384 => x"5377d638",
   385 => x"74753352",
   386 => x"5670802e",
   387 => x"80c53870",
   388 => x"b3a40859",
   389 => x"538116ba",
   390 => x"dc337081",
   391 => x"ff067010",
   392 => x"1011bae0",
   393 => x"337081ff",
   394 => x"06729029",
   395 => x"1170882b",
   396 => x"7a077f0c",
   397 => x"53595954",
   398 => x"54585672",
   399 => x"8a2ebd38",
   400 => x"7380cf2e",
   401 => x"b7388115",
   402 => x"5372bae0",
   403 => x"34753353",
   404 => x"72c33889",
   405 => x"3d0d0484",
   406 => x"12087082",
   407 => x"2a810657",
   408 => x"5875802e",
   409 => x"f2388d72",
   410 => x"0c841208",
   411 => x"70822a81",
   412 => x"06525770",
   413 => x"802efeef",
   414 => x"38fefb39",
   415 => x"71a32697",
   416 => x"38811752",
   417 => x"71badc34",
   418 => x"800bbae0",
   419 => x"34753353",
   420 => x"72ff8238",
   421 => x"ffbd3980",
   422 => x"0bbadc34",
   423 => x"800bbae0",
   424 => x"34eb39e9",
   425 => x"3d0db3a4",
   426 => x"0855800b",
   427 => x"84160cfe",
   428 => x"800a0b88",
   429 => x"160c800b",
   430 => x"badc3480",
   431 => x"0bbae034",
   432 => x"943d7053",
   433 => x"b3980884",
   434 => x"11085355",
   435 => x"5cfcd53f",
   436 => x"abd80bab",
   437 => x"d833555a",
   438 => x"73802e80",
   439 => x"c738b3a4",
   440 => x"0874575b",
   441 => x"811abadc",
   442 => x"337081ff",
   443 => x"06701010",
   444 => x"11bae033",
   445 => x"7081ff06",
   446 => x"72902911",
   447 => x"70882b7d",
   448 => x"07620c44",
   449 => x"5c5c4257",
   450 => x"5a5a758a",
   451 => x"2e87a538",
   452 => x"7680cf2e",
   453 => x"879e3881",
   454 => x"185776ba",
   455 => x"e0347933",
   456 => x"5675c138",
   457 => x"7b7c3355",
   458 => x"5a73802e",
   459 => x"80c738b3",
   460 => x"a4087457",
   461 => x"5b811aba",
   462 => x"dc337081",
   463 => x"ff067010",
   464 => x"1011bae0",
   465 => x"337081ff",
   466 => x"06729029",
   467 => x"1170882b",
   468 => x"7d07620c",
   469 => x"465c5c57",
   470 => x"575a5a75",
   471 => x"8a2e86ef",
   472 => x"387680cf",
   473 => x"2e86e838",
   474 => x"81185978",
   475 => x"bae03479",
   476 => x"335675c1",
   477 => x"38abe80b",
   478 => x"abe83355",
   479 => x"5a73802e",
   480 => x"80c738b3",
   481 => x"a4087457",
   482 => x"5b811aba",
   483 => x"dc337081",
   484 => x"ff067010",
   485 => x"1011bae0",
   486 => x"337081ff",
   487 => x"06729029",
   488 => x"1170882b",
   489 => x"7d07620c",
   490 => x"445c5c42",
   491 => x"575a5a75",
   492 => x"8a2e85e4",
   493 => x"387680cf",
   494 => x"2e85dd38",
   495 => x"81185675",
   496 => x"bae03479",
   497 => x"335675c1",
   498 => x"38890a5c",
   499 => x"8070933d",
   500 => x"028c0580",
   501 => x"c1054142",
   502 => x"5e5f7cbf",
   503 => x"065a7982",
   504 => x"aa38abd0",
   505 => x"0babd033",
   506 => x"555a7380",
   507 => x"2e80c738",
   508 => x"b3a40874",
   509 => x"575b811a",
   510 => x"badc3370",
   511 => x"81ff0670",
   512 => x"101011ba",
   513 => x"e0337081",
   514 => x"ff067290",
   515 => x"29117088",
   516 => x"2b7d0762",
   517 => x"0c535c5c",
   518 => x"57575a5a",
   519 => x"758a2e82",
   520 => x"f8387680",
   521 => x"cf2e82f1",
   522 => x"38811859",
   523 => x"78bae034",
   524 => x"79335675",
   525 => x"c1387b56",
   526 => x"8b53a8d4",
   527 => x"527f5194",
   528 => x"e43f8857",
   529 => x"758f0654",
   530 => x"73892682",
   531 => x"b038761e",
   532 => x"b0155555",
   533 => x"73753475",
   534 => x"842aff18",
   535 => x"7081ff06",
   536 => x"595c5676",
   537 => x"df387f60",
   538 => x"33555a73",
   539 => x"802e80c7",
   540 => x"38b3a408",
   541 => x"74575b81",
   542 => x"1abadc33",
   543 => x"7081ff06",
   544 => x"70101011",
   545 => x"bae03370",
   546 => x"81ff0672",
   547 => x"90291170",
   548 => x"882b7d07",
   549 => x"620c535c",
   550 => x"5c57575a",
   551 => x"5a758a2e",
   552 => x"84ed3876",
   553 => x"80cf2e84",
   554 => x"e6388118",
   555 => x"5574bae0",
   556 => x"34793356",
   557 => x"75c138ab",
   558 => x"ec0babec",
   559 => x"33555a73",
   560 => x"802e80c7",
   561 => x"38b3a408",
   562 => x"74575b81",
   563 => x"1abadc33",
   564 => x"7081ff06",
   565 => x"70101011",
   566 => x"bae03370",
   567 => x"81ff0672",
   568 => x"90291170",
   569 => x"882b7d07",
   570 => x"620c535c",
   571 => x"5c57575a",
   572 => x"5a758a2e",
   573 => x"84b43876",
   574 => x"80cf2e84",
   575 => x"ad388118",
   576 => x"5776bae0",
   577 => x"34793356",
   578 => x"75c1387b",
   579 => x"7c082e81",
   580 => x"a438abf0",
   581 => x"0babf033",
   582 => x"555a7380",
   583 => x"2e80c738",
   584 => x"b3a40874",
   585 => x"575b811a",
   586 => x"badc3370",
   587 => x"81ff0670",
   588 => x"101011ba",
   589 => x"e0337081",
   590 => x"ff067290",
   591 => x"29117088",
   592 => x"2b7d0762",
   593 => x"0c535c5c",
   594 => x"57575a5a",
   595 => x"758a2e82",
   596 => x"93387680",
   597 => x"cf2e828c",
   598 => x"38811856",
   599 => x"75bae034",
   600 => x"79335675",
   601 => x"c138811f",
   602 => x"5f821c81",
   603 => x"1e5e5c8f",
   604 => x"ff7d27fc",
   605 => x"e5387e80",
   606 => x"0c993d0d",
   607 => x"04761eb7",
   608 => x"15555573",
   609 => x"75347584",
   610 => x"2aff1870",
   611 => x"81ff0659",
   612 => x"5c5676fd",
   613 => x"af38fdce",
   614 => x"3974a326",
   615 => x"81ed3881",
   616 => x"195776ba",
   617 => x"dc34800b",
   618 => x"bae03479",
   619 => x"335675fc",
   620 => x"c538fd82",
   621 => x"39841c5a",
   622 => x"797a082e",
   623 => x"098106fe",
   624 => x"d138abf4",
   625 => x"0babf433",
   626 => x"555a7380",
   627 => x"2eff9a38",
   628 => x"b3a40874",
   629 => x"811cbadc",
   630 => x"337081ff",
   631 => x"06701010",
   632 => x"11bae033",
   633 => x"7081ff06",
   634 => x"72902911",
   635 => x"70882b78",
   636 => x"07790c53",
   637 => x"5e5e5959",
   638 => x"5c5c575b",
   639 => x"758a2e80",
   640 => x"c7387680",
   641 => x"cf2e80c0",
   642 => x"38811859",
   643 => x"78bae034",
   644 => x"79335675",
   645 => x"802efed1",
   646 => x"38811aba",
   647 => x"dc337081",
   648 => x"ff067010",
   649 => x"1011bae0",
   650 => x"337081ff",
   651 => x"06729029",
   652 => x"1170882b",
   653 => x"7d07620c",
   654 => x"535c5c57",
   655 => x"575a5a75",
   656 => x"8a2e0981",
   657 => x"06ffbb38",
   658 => x"74a32682",
   659 => x"90388119",
   660 => x"5877badc",
   661 => x"34800bba",
   662 => x"e0347933",
   663 => x"5675ffb9",
   664 => x"38fe8639",
   665 => x"74a32697",
   666 => x"38811955",
   667 => x"74badc34",
   668 => x"800bbae0",
   669 => x"34793356",
   670 => x"75fdab38",
   671 => x"fde83980",
   672 => x"0bbadc34",
   673 => x"800bbae0",
   674 => x"34eb3980",
   675 => x"0bbadc34",
   676 => x"800bbae0",
   677 => x"34fe9439",
   678 => x"74a32680",
   679 => x"e5388119",
   680 => x"5574badc",
   681 => x"34800bba",
   682 => x"e0347933",
   683 => x"5675f9d9",
   684 => x"38fa9639",
   685 => x"74a326be",
   686 => x"38811956",
   687 => x"75badc34",
   688 => x"800bbae0",
   689 => x"34793356",
   690 => x"75f89938",
   691 => x"f8d63974",
   692 => x"a3269738",
   693 => x"81195877",
   694 => x"badc3480",
   695 => x"0bbae034",
   696 => x"79335675",
   697 => x"f8cf38f9",
   698 => x"8c39800b",
   699 => x"badc3480",
   700 => x"0bbae034",
   701 => x"eb39800b",
   702 => x"badc3480",
   703 => x"0bbae034",
   704 => x"c439800b",
   705 => x"badc3480",
   706 => x"0bbae034",
   707 => x"ff9c3974",
   708 => x"a326be38",
   709 => x"81195877",
   710 => x"badc3480",
   711 => x"0bbae034",
   712 => x"79335675",
   713 => x"fad138fb",
   714 => x"8e3974a3",
   715 => x"26973881",
   716 => x"195675ba",
   717 => x"dc34800b",
   718 => x"bae03479",
   719 => x"335675fb",
   720 => x"8a38fbc7",
   721 => x"39800bba",
   722 => x"dc34800b",
   723 => x"bae034eb",
   724 => x"39800bba",
   725 => x"dc34800b",
   726 => x"bae034c4",
   727 => x"39800bba",
   728 => x"dc34800b",
   729 => x"bae034fd",
   730 => x"f139ec3d",
   731 => x"0db18451",
   732 => x"f4cf3fb1",
   733 => x"a051f4c9",
   734 => x"3f913d70",
   735 => x"53b39808",
   736 => x"84110853",
   737 => x"555cf39c",
   738 => x"3f7b51f4",
   739 => x"b43fabec",
   740 => x"51f4ae3f",
   741 => x"f68d3f80",
   742 => x"088f3d5a",
   743 => x"568b53a8",
   744 => x"d4527851",
   745 => x"8dff3f88",
   746 => x"028405b5",
   747 => x"05595775",
   748 => x"8f065473",
   749 => x"892684c9",
   750 => x"387618b0",
   751 => x"15555573",
   752 => x"75347584",
   753 => x"2aff1870",
   754 => x"81ff0659",
   755 => x"565676df",
   756 => x"38787933",
   757 => x"55577380",
   758 => x"2ea83873",
   759 => x"b3ac0856",
   760 => x"56811757",
   761 => x"758a2e84",
   762 => x"b4388415",
   763 => x"0870822a",
   764 => x"81065e58",
   765 => x"7c802ef2",
   766 => x"3875750c",
   767 => x"76335675",
   768 => x"e0387879",
   769 => x"33555a73",
   770 => x"802e80c7",
   771 => x"3873b3a4",
   772 => x"085c5681",
   773 => x"1abadc33",
   774 => x"7081ff06",
   775 => x"70101011",
   776 => x"bae03370",
   777 => x"81ff0672",
   778 => x"90291170",
   779 => x"882b7d07",
   780 => x"620c5a5c",
   781 => x"5c40575a",
   782 => x"5a758a2e",
   783 => x"84843876",
   784 => x"80cf2e83",
   785 => x"fd388118",
   786 => x"5776bae0",
   787 => x"34793356",
   788 => x"75c138b3",
   789 => x"98088411",
   790 => x"085a56fe",
   791 => x"817925a8",
   792 => x"38b3a808",
   793 => x"55800b84",
   794 => x"170cb0ea",
   795 => x"0b94160c",
   796 => x"850b9816",
   797 => x"0c981508",
   798 => x"81065a79",
   799 => x"f8388416",
   800 => x"085877fe",
   801 => x"8124de38",
   802 => x"83ffff5a",
   803 => x"fe810b84",
   804 => x"1708565b",
   805 => x"7481fe24",
   806 => x"80c63880",
   807 => x"0b88170c",
   808 => x"f4813f80",
   809 => x"0883ffff",
   810 => x"0655747a",
   811 => x"278b3874",
   812 => x"b3980884",
   813 => x"11085d55",
   814 => x"5aabd051",
   815 => x"f2833f7b",
   816 => x"527451f0",
   817 => x"df3f7b51",
   818 => x"f1f73f74",
   819 => x"802e8399",
   820 => x"38b39808",
   821 => x"84110856",
   822 => x"5681fe75",
   823 => x"25ffbc38",
   824 => x"8416085d",
   825 => x"84160857",
   826 => x"7681fe24",
   827 => x"80c43880",
   828 => x"0b88170c",
   829 => x"f3ad3f80",
   830 => x"0883ffff",
   831 => x"0655747a",
   832 => x"278b3874",
   833 => x"b3980884",
   834 => x"11085d57",
   835 => x"5aabd051",
   836 => x"f1af3f7b",
   837 => x"527451f0",
   838 => x"8b3f7b51",
   839 => x"f1a33f74",
   840 => x"82d238b3",
   841 => x"98088411",
   842 => x"08585681",
   843 => x"fe7725ff",
   844 => x"be388416",
   845 => x"08598079",
   846 => x"7c315957",
   847 => x"767825ae",
   848 => x"38b3a808",
   849 => x"55800b84",
   850 => x"170cb0ea",
   851 => x"0b94160c",
   852 => x"850b9816",
   853 => x"0c981508",
   854 => x"70810651",
   855 => x"5473f638",
   856 => x"81177083",
   857 => x"ffff0658",
   858 => x"54777724",
   859 => x"d838b1ac",
   860 => x"51f0ce3f",
   861 => x"7b527c51",
   862 => x"efaa3f7b",
   863 => x"51f0c23f",
   864 => x"b1bc51f0",
   865 => x"bc3f7b52",
   866 => x"7851ef98",
   867 => x"3f7b51f0",
   868 => x"b03fb1cc",
   869 => x"51f0aa3f",
   870 => x"7b52787d",
   871 => x"31705258",
   872 => x"ef823f7b",
   873 => x"51f09a3f",
   874 => x"b1dc51f0",
   875 => x"943f7b52",
   876 => x"779f2a18",
   877 => x"70812c52",
   878 => x"59eee93f",
   879 => x"7b51f081",
   880 => x"3fb1ec51",
   881 => x"effb3f7b",
   882 => x"527951ee",
   883 => x"d73f7b51",
   884 => x"efef3fb1",
   885 => x"fc51efe9",
   886 => x"3f7b527a",
   887 => x"51eec53f",
   888 => x"7b51efdd",
   889 => x"3fb28c51",
   890 => x"efd73f7b",
   891 => x"52b39808",
   892 => x"84110852",
   893 => x"5deead3f",
   894 => x"7b51efc5",
   895 => x"3f963d0d",
   896 => x"047618b7",
   897 => x"15555573",
   898 => x"75347584",
   899 => x"2aff1870",
   900 => x"81ff0659",
   901 => x"565676fb",
   902 => x"9638fbb5",
   903 => x"39841508",
   904 => x"70822a81",
   905 => x"06595b77",
   906 => x"802ef238",
   907 => x"8d750c84",
   908 => x"15087082",
   909 => x"2a81065e",
   910 => x"587c802e",
   911 => x"fbac38fb",
   912 => x"b83974a3",
   913 => x"26973881",
   914 => x"195675ba",
   915 => x"dc34800b",
   916 => x"bae03479",
   917 => x"335675fb",
   918 => x"ba38fbf7",
   919 => x"39800bba",
   920 => x"dc34800b",
   921 => x"bae034eb",
   922 => x"39b39808",
   923 => x"8411085e",
   924 => x"56fcf139",
   925 => x"b3980856",
   926 => x"fdb839f7",
   927 => x"3d0db3a0",
   928 => x"08700881",
   929 => x"0a06bad8",
   930 => x"0c55890a",
   931 => x"53f0800a",
   932 => x"5472730c",
   933 => x"8413ff15",
   934 => x"55537380",
   935 => x"25f338b3",
   936 => x"a8085487",
   937 => x"0b84150c",
   938 => x"b3a40853",
   939 => x"800b8414",
   940 => x"0cfe800a",
   941 => x"0b88140c",
   942 => x"800bbadc",
   943 => x"34800bba",
   944 => x"e034b3ac",
   945 => x"0854b60b",
   946 => x"8c150c83",
   947 => x"0b88150c",
   948 => x"81ff0b88",
   949 => x"160cb39c",
   950 => x"0854ff0b",
   951 => x"84150cfc",
   952 => x"94800b88",
   953 => x"150c82d0",
   954 => x"affdfb0b",
   955 => x"8c150c80",
   956 => x"c0740c73",
   957 => x"0870862a",
   958 => x"81065155",
   959 => x"74f53890",
   960 => x"14087083",
   961 => x"2a810651",
   962 => x"5372f438",
   963 => x"81fc8081",
   964 => x"0b90150c",
   965 => x"90140870",
   966 => x"832a8106",
   967 => x"515372f4",
   968 => x"3880fdc0",
   969 => x"810b9015",
   970 => x"0caba051",
   971 => x"ed933f72",
   972 => x"b3a40856",
   973 => x"5473882b",
   974 => x"750c8114",
   975 => x"54979074",
   976 => x"26f33880",
   977 => x"0bbadc34",
   978 => x"800bbae0",
   979 => x"34b29c51",
   980 => x"ecef3fba",
   981 => x"d808802e",
   982 => x"81ff38b2",
   983 => x"a451ece1",
   984 => x"3fb2b451",
   985 => x"ecdb3ff8",
   986 => x"813f800b",
   987 => x"b3a80855",
   988 => x"55bfa9bc",
   989 => x"0b94150c",
   990 => x"850b9815",
   991 => x"0c981408",
   992 => x"70810651",
   993 => x"5372f638",
   994 => x"bfa9bc0b",
   995 => x"94150c85",
   996 => x"0b98150c",
   997 => x"98140870",
   998 => x"81065153",
   999 => x"72f638bf",
  1000 => x"a9bc0b94",
  1001 => x"150c850b",
  1002 => x"98150c98",
  1003 => x"14087081",
  1004 => x"06515372",
  1005 => x"f638bfa9",
  1006 => x"bc0b9415",
  1007 => x"0c850b98",
  1008 => x"150c9814",
  1009 => x"08708106",
  1010 => x"515372f6",
  1011 => x"38bfa9bc",
  1012 => x"0b94150c",
  1013 => x"850b9815",
  1014 => x"0c981408",
  1015 => x"70810651",
  1016 => x"5372f638",
  1017 => x"bfa9bc0b",
  1018 => x"94150c85",
  1019 => x"0b98150c",
  1020 => x"98140870",
  1021 => x"81065153",
  1022 => x"72f63881",
  1023 => x"15558a75",
  1024 => x"26feee38",
  1025 => x"72b3a408",
  1026 => x"56547388",
  1027 => x"2b750c81",
  1028 => x"14549790",
  1029 => x"7426f338",
  1030 => x"800bbadc",
  1031 => x"34800bba",
  1032 => x"e034ecff",
  1033 => x"3fb3a008",
  1034 => x"70087087",
  1035 => x"2a810651",
  1036 => x"56547480",
  1037 => x"2e8a38b3",
  1038 => x"98085380",
  1039 => x"0b84140c",
  1040 => x"73087084",
  1041 => x"2a810655",
  1042 => x"5373802e",
  1043 => x"d538b398",
  1044 => x"0854800b",
  1045 => x"88150cca",
  1046 => x"39b2d851",
  1047 => x"fe80398c",
  1048 => x"08028c0c",
  1049 => x"fd3d0d80",
  1050 => x"538c088c",
  1051 => x"0508528c",
  1052 => x"08880508",
  1053 => x"5182de3f",
  1054 => x"80087080",
  1055 => x"0c54853d",
  1056 => x"0d8c0c04",
  1057 => x"8c08028c",
  1058 => x"0cfd3d0d",
  1059 => x"81538c08",
  1060 => x"8c050852",
  1061 => x"8c088805",
  1062 => x"085182b9",
  1063 => x"3f800870",
  1064 => x"800c5485",
  1065 => x"3d0d8c0c",
  1066 => x"048c0802",
  1067 => x"8c0cf93d",
  1068 => x"0d800b8c",
  1069 => x"08fc050c",
  1070 => x"8c088805",
  1071 => x"088025ab",
  1072 => x"388c0888",
  1073 => x"0508308c",
  1074 => x"0888050c",
  1075 => x"800b8c08",
  1076 => x"f4050c8c",
  1077 => x"08fc0508",
  1078 => x"8838810b",
  1079 => x"8c08f405",
  1080 => x"0c8c08f4",
  1081 => x"05088c08",
  1082 => x"fc050c8c",
  1083 => x"088c0508",
  1084 => x"8025ab38",
  1085 => x"8c088c05",
  1086 => x"08308c08",
  1087 => x"8c050c80",
  1088 => x"0b8c08f0",
  1089 => x"050c8c08",
  1090 => x"fc050888",
  1091 => x"38810b8c",
  1092 => x"08f0050c",
  1093 => x"8c08f005",
  1094 => x"088c08fc",
  1095 => x"050c8053",
  1096 => x"8c088c05",
  1097 => x"08528c08",
  1098 => x"88050851",
  1099 => x"81a73f80",
  1100 => x"08708c08",
  1101 => x"f8050c54",
  1102 => x"8c08fc05",
  1103 => x"08802e8c",
  1104 => x"388c08f8",
  1105 => x"0508308c",
  1106 => x"08f8050c",
  1107 => x"8c08f805",
  1108 => x"0870800c",
  1109 => x"54893d0d",
  1110 => x"8c0c048c",
  1111 => x"08028c0c",
  1112 => x"fb3d0d80",
  1113 => x"0b8c08fc",
  1114 => x"050c8c08",
  1115 => x"88050880",
  1116 => x"2593388c",
  1117 => x"08880508",
  1118 => x"308c0888",
  1119 => x"050c810b",
  1120 => x"8c08fc05",
  1121 => x"0c8c088c",
  1122 => x"05088025",
  1123 => x"8c388c08",
  1124 => x"8c050830",
  1125 => x"8c088c05",
  1126 => x"0c81538c",
  1127 => x"088c0508",
  1128 => x"528c0888",
  1129 => x"050851ad",
  1130 => x"3f800870",
  1131 => x"8c08f805",
  1132 => x"0c548c08",
  1133 => x"fc050880",
  1134 => x"2e8c388c",
  1135 => x"08f80508",
  1136 => x"308c08f8",
  1137 => x"050c8c08",
  1138 => x"f8050870",
  1139 => x"800c5487",
  1140 => x"3d0d8c0c",
  1141 => x"048c0802",
  1142 => x"8c0cfd3d",
  1143 => x"0d810b8c",
  1144 => x"08fc050c",
  1145 => x"800b8c08",
  1146 => x"f8050c8c",
  1147 => x"088c0508",
  1148 => x"8c088805",
  1149 => x"0827ac38",
  1150 => x"8c08fc05",
  1151 => x"08802ea3",
  1152 => x"38800b8c",
  1153 => x"088c0508",
  1154 => x"2499388c",
  1155 => x"088c0508",
  1156 => x"108c088c",
  1157 => x"050c8c08",
  1158 => x"fc050810",
  1159 => x"8c08fc05",
  1160 => x"0cc9398c",
  1161 => x"08fc0508",
  1162 => x"802e80c9",
  1163 => x"388c088c",
  1164 => x"05088c08",
  1165 => x"88050826",
  1166 => x"a1388c08",
  1167 => x"8805088c",
  1168 => x"088c0508",
  1169 => x"318c0888",
  1170 => x"050c8c08",
  1171 => x"f805088c",
  1172 => x"08fc0508",
  1173 => x"078c08f8",
  1174 => x"050c8c08",
  1175 => x"fc050881",
  1176 => x"2a8c08fc",
  1177 => x"050c8c08",
  1178 => x"8c050881",
  1179 => x"2a8c088c",
  1180 => x"050cffaf",
  1181 => x"398c0890",
  1182 => x"0508802e",
  1183 => x"8f388c08",
  1184 => x"88050870",
  1185 => x"8c08f405",
  1186 => x"0c518d39",
  1187 => x"8c08f805",
  1188 => x"08708c08",
  1189 => x"f4050c51",
  1190 => x"8c08f405",
  1191 => x"08800c85",
  1192 => x"3d0d8c0c",
  1193 => x"04fc3d0d",
  1194 => x"7670797b",
  1195 => x"55555555",
  1196 => x"8f72278c",
  1197 => x"38727507",
  1198 => x"83065170",
  1199 => x"802ea738",
  1200 => x"ff125271",
  1201 => x"ff2e9838",
  1202 => x"72708105",
  1203 => x"54337470",
  1204 => x"81055634",
  1205 => x"ff125271",
  1206 => x"ff2e0981",
  1207 => x"06ea3874",
  1208 => x"800c863d",
  1209 => x"0d047451",
  1210 => x"72708405",
  1211 => x"54087170",
  1212 => x"8405530c",
  1213 => x"72708405",
  1214 => x"54087170",
  1215 => x"8405530c",
  1216 => x"72708405",
  1217 => x"54087170",
  1218 => x"8405530c",
  1219 => x"72708405",
  1220 => x"54087170",
  1221 => x"8405530c",
  1222 => x"f0125271",
  1223 => x"8f26c938",
  1224 => x"83722795",
  1225 => x"38727084",
  1226 => x"05540871",
  1227 => x"70840553",
  1228 => x"0cfc1252",
  1229 => x"718326ed",
  1230 => x"387054ff",
  1231 => x"8339fd3d",
  1232 => x"0d800bb3",
  1233 => x"8c085454",
  1234 => x"72812e98",
  1235 => x"3873bae4",
  1236 => x"0ce28c3f",
  1237 => x"e1aa3fb3",
  1238 => x"b0528151",
  1239 => x"f69d3f80",
  1240 => x"08519e3f",
  1241 => x"72bae40c",
  1242 => x"e1f53fe1",
  1243 => x"933fb3b0",
  1244 => x"528151f6",
  1245 => x"863f8008",
  1246 => x"51873f00",
  1247 => x"ff3900ff",
  1248 => x"39f73d0d",
  1249 => x"7bb3b408",
  1250 => x"82c81108",
  1251 => x"5a545a77",
  1252 => x"802e80d9",
  1253 => x"38818818",
  1254 => x"841908ff",
  1255 => x"0581712b",
  1256 => x"59555980",
  1257 => x"742480e9",
  1258 => x"38807424",
  1259 => x"b5387382",
  1260 => x"2b781188",
  1261 => x"05565681",
  1262 => x"80190877",
  1263 => x"06537280",
  1264 => x"2eb53878",
  1265 => x"16700853",
  1266 => x"53795174",
  1267 => x"0853722d",
  1268 => x"ff14fc17",
  1269 => x"fc177981",
  1270 => x"2c5a5757",
  1271 => x"54738025",
  1272 => x"d6387708",
  1273 => x"5877ffad",
  1274 => x"38b3b408",
  1275 => x"53bc1308",
  1276 => x"a5387951",
  1277 => x"ff853f74",
  1278 => x"0853722d",
  1279 => x"ff14fc17",
  1280 => x"fc177981",
  1281 => x"2c5a5757",
  1282 => x"54738025",
  1283 => x"ffa938d2",
  1284 => x"398057ff",
  1285 => x"94397251",
  1286 => x"bc130853",
  1287 => x"722d7951",
  1288 => x"fed93fff",
  1289 => x"3d0dbab8",
  1290 => x"0bfc0570",
  1291 => x"08525270",
  1292 => x"ff2e9138",
  1293 => x"702dfc12",
  1294 => x"70085252",
  1295 => x"70ff2e09",
  1296 => x"8106f138",
  1297 => x"833d0d04",
  1298 => x"04e0f93f",
  1299 => x"04000000",
  1300 => x"00000040",
  1301 => x"30782020",
  1302 => x"20202020",
  1303 => x"20200000",
  1304 => x"0a677265",
  1305 => x"74682072",
  1306 => x"65676973",
  1307 => x"74657273",
  1308 => x"3a000000",
  1309 => x"0a636f6e",
  1310 => x"74726f6c",
  1311 => x"3a202020",
  1312 => x"20202000",
  1313 => x"0a737461",
  1314 => x"7475733a",
  1315 => x"20202020",
  1316 => x"20202000",
  1317 => x"0a6d6163",
  1318 => x"5f6d7362",
  1319 => x"3a202020",
  1320 => x"20202000",
  1321 => x"0a6d6163",
  1322 => x"5f6c7362",
  1323 => x"3a202020",
  1324 => x"20202000",
  1325 => x"0a6d6469",
  1326 => x"6f5f636f",
  1327 => x"6e74726f",
  1328 => x"6c3a2000",
  1329 => x"0a74785f",
  1330 => x"706f696e",
  1331 => x"7465723a",
  1332 => x"20202000",
  1333 => x"0a72785f",
  1334 => x"706f696e",
  1335 => x"7465723a",
  1336 => x"20202000",
  1337 => x"0a656463",
  1338 => x"6c5f6970",
  1339 => x"3a202020",
  1340 => x"20202000",
  1341 => x"0a686173",
  1342 => x"685f6d73",
  1343 => x"623a2020",
  1344 => x"20202000",
  1345 => x"0a686173",
  1346 => x"685f6c73",
  1347 => x"623a2020",
  1348 => x"20202000",
  1349 => x"0a6d6469",
  1350 => x"6f207068",
  1351 => x"79207265",
  1352 => x"67697374",
  1353 => x"65727300",
  1354 => x"0a206d64",
  1355 => x"696f2070",
  1356 => x"68793a20",
  1357 => x"00000000",
  1358 => x"0a202072",
  1359 => x"65673a20",
  1360 => x"00000000",
  1361 => x"2d3e2000",
  1362 => x"0a677265",
  1363 => x"74682d3e",
  1364 => x"636f6e74",
  1365 => x"726f6c20",
  1366 => x"3a000000",
  1367 => x"0a677265",
  1368 => x"74682d3e",
  1369 => x"73746174",
  1370 => x"75732020",
  1371 => x"3a000000",
  1372 => x"0a646573",
  1373 => x"63722d3e",
  1374 => x"636f6e74",
  1375 => x"726f6c20",
  1376 => x"3a000000",
  1377 => x"77726974",
  1378 => x"65206164",
  1379 => x"64726573",
  1380 => x"733a2000",
  1381 => x"20206c65",
  1382 => x"6e677468",
  1383 => x"3a200000",
  1384 => x"0a0a0000",
  1385 => x"72656164",
  1386 => x"20206164",
  1387 => x"64726573",
  1388 => x"733a2000",
  1389 => x"20206578",
  1390 => x"70656374",
  1391 => x"3a200000",
  1392 => x"2020676f",
  1393 => x"743a2000",
  1394 => x"20657272",
  1395 => x"6f720000",
  1396 => x"0a000000",
  1397 => x"206f6b00",
  1398 => x"70686173",
  1399 => x"65207368",
  1400 => x"69667420",
  1401 => x"3a200000",
  1402 => x"20202020",
  1403 => x"20000000",
  1404 => x"21000000",
  1405 => x"2e000000",
  1406 => x"44445220",
  1407 => x"6d656d6f",
  1408 => x"72792069",
  1409 => x"6e666f00",
  1410 => x"0a617574",
  1411 => x"6f20745f",
  1412 => x"52455245",
  1413 => x"5348203a",
  1414 => x"00000000",
  1415 => x"0a636c6f",
  1416 => x"636b2065",
  1417 => x"6e61626c",
  1418 => x"6520203a",
  1419 => x"00000000",
  1420 => x"0a696e69",
  1421 => x"74616c69",
  1422 => x"7a652020",
  1423 => x"2020203a",
  1424 => x"00000000",
  1425 => x"0a636f6c",
  1426 => x"756d6e20",
  1427 => x"73697a65",
  1428 => x"2020203a",
  1429 => x"00000000",
  1430 => x"0a62616e",
  1431 => x"6b73697a",
  1432 => x"65202020",
  1433 => x"2020203a",
  1434 => x"00000000",
  1435 => x"4d627974",
  1436 => x"65000000",
  1437 => x"0a745f52",
  1438 => x"43442020",
  1439 => x"20202020",
  1440 => x"2020203a",
  1441 => x"00000000",
  1442 => x"0a745f52",
  1443 => x"46432020",
  1444 => x"20202020",
  1445 => x"2020203a",
  1446 => x"00000000",
  1447 => x"0a745f52",
  1448 => x"50202020",
  1449 => x"20202020",
  1450 => x"2020203a",
  1451 => x"00000000",
  1452 => x"0a726566",
  1453 => x"72657368",
  1454 => x"20656e2e",
  1455 => x"2020203a",
  1456 => x"00000000",
  1457 => x"0a444452",
  1458 => x"20667265",
  1459 => x"7175656e",
  1460 => x"6379203a",
  1461 => x"00000000",
  1462 => x"0a444452",
  1463 => x"20646174",
  1464 => x"61207769",
  1465 => x"6474683a",
  1466 => x"00000000",
  1467 => x"0a6d6f62",
  1468 => x"696c6520",
  1469 => x"73757070",
  1470 => x"6f72743a",
  1471 => x"00000000",
  1472 => x"0a73656c",
  1473 => x"66207265",
  1474 => x"66726573",
  1475 => x"6820203a",
  1476 => x"00000000",
  1477 => x"756e6b6e",
  1478 => x"6f776e00",
  1479 => x"20617272",
  1480 => x"61790000",
  1481 => x"0a74656d",
  1482 => x"702d636f",
  1483 => x"6d702072",
  1484 => x"6566723a",
  1485 => x"00000000",
  1486 => x"c2b04300",
  1487 => x"0a647269",
  1488 => x"76652073",
  1489 => x"7472656e",
  1490 => x"6774683a",
  1491 => x"00000000",
  1492 => x"0a706f77",
  1493 => x"65722073",
  1494 => x"6176696e",
  1495 => x"6720203a",
  1496 => x"00000000",
  1497 => x"0a745f58",
  1498 => x"50202020",
  1499 => x"20202020",
  1500 => x"2020203a",
  1501 => x"00000000",
  1502 => x"0a745f58",
  1503 => x"53522020",
  1504 => x"20202020",
  1505 => x"2020203a",
  1506 => x"00000000",
  1507 => x"0a745f43",
  1508 => x"4b452020",
  1509 => x"20202020",
  1510 => x"2020203a",
  1511 => x"00000000",
  1512 => x"0a434153",
  1513 => x"206c6174",
  1514 => x"656e6379",
  1515 => x"2020203a",
  1516 => x"00000000",
  1517 => x"0a6d6f62",
  1518 => x"696c6520",
  1519 => x"656e6162",
  1520 => x"6c65643a",
  1521 => x"00000000",
  1522 => x"0a737461",
  1523 => x"74757320",
  1524 => x"72656164",
  1525 => x"2020203a",
  1526 => x"00000000",
  1527 => x"332f3400",
  1528 => x"38350000",
  1529 => x"68616c66",
  1530 => x"00000000",
  1531 => x"34303639",
  1532 => x"00000000",
  1533 => x"20353132",
  1534 => x"00000000",
  1535 => x"66756c6c",
  1536 => x"00000000",
  1537 => x"37300000",
  1538 => x"34350000",
  1539 => x"31303234",
  1540 => x"00000000",
  1541 => x"31350000",
  1542 => x"312f3400",
  1543 => x"32303438",
  1544 => x"00000000",
  1545 => x"312f3800",
  1546 => x"312f3200",
  1547 => x"312f3100",
  1548 => x"64656570",
  1549 => x"20706f77",
  1550 => x"65722064",
  1551 => x"6f776e00",
  1552 => x"636c6f63",
  1553 => x"6b207374",
  1554 => x"6f700000",
  1555 => x"73656c66",
  1556 => x"20726566",
  1557 => x"72657368",
  1558 => x"00000000",
  1559 => x"706f7765",
  1560 => x"7220646f",
  1561 => x"776e0000",
  1562 => x"6e6f6e65",
  1563 => x"00000000",
  1564 => x"61646472",
  1565 => x"6573733a",
  1566 => x"20000000",
  1567 => x"20646174",
  1568 => x"613a2000",
  1569 => x"0a0a4443",
  1570 => x"4d207068",
  1571 => x"61736520",
  1572 => x"73686966",
  1573 => x"74207465",
  1574 => x"7374696e",
  1575 => x"67000000",
  1576 => x"0a696e69",
  1577 => x"7469616c",
  1578 => x"3a200000",
  1579 => x"0a6c6f77",
  1580 => x"3a202020",
  1581 => x"20202020",
  1582 => x"20200000",
  1583 => x"0a686967",
  1584 => x"683a2020",
  1585 => x"20202020",
  1586 => x"20200000",
  1587 => x"0a646966",
  1588 => x"663a2020",
  1589 => x"20202020",
  1590 => x"20200000",
  1591 => x"0a646966",
  1592 => x"662f323a",
  1593 => x"20202020",
  1594 => x"20200000",
  1595 => x"0a6d696e",
  1596 => x"5f657272",
  1597 => x"3a202020",
  1598 => x"20200000",
  1599 => x"0a6d696e",
  1600 => x"5f657272",
  1601 => x"5f706f73",
  1602 => x"3a200000",
  1603 => x"0a66696e",
  1604 => x"616c3a20",
  1605 => x"20202020",
  1606 => x"20200000",
  1607 => x"74657374",
  1608 => x"2e632000",
  1609 => x"286f6e20",
  1610 => x"73696d75",
  1611 => x"6c61746f",
  1612 => x"72290a00",
  1613 => x"636f6d70",
  1614 => x"696c6564",
  1615 => x"3a204175",
  1616 => x"67203237",
  1617 => x"20323031",
  1618 => x"30202031",
  1619 => x"333a3536",
  1620 => x"3a33320a",
  1621 => x"00000000",
  1622 => x"286f6e20",
  1623 => x"68617264",
  1624 => x"77617265",
  1625 => x"290a0000",
  1626 => x"64756d6d",
  1627 => x"792e6578",
  1628 => x"65000000",
  1629 => x"43000000",
  1630 => x"00ffffff",
  1631 => x"ff00ffff",
  1632 => x"ffff00ff",
  1633 => x"ffffff00",
  1634 => x"00000000",
  1635 => x"00000000",
  1636 => x"00000000",
  1637 => x"00001d40",
  1638 => x"80000e00",
  1639 => x"80000c00",
  1640 => x"80000800",
  1641 => x"80000600",
  1642 => x"80000200",
  1643 => x"80000100",
  1644 => x"00001968",
  1645 => x"000019b8",
  1646 => x"00000000",
  1647 => x"00001c20",
  1648 => x"00001c7c",
  1649 => x"00001cd8",
  1650 => x"00000000",
  1651 => x"00000000",
  1652 => x"00000000",
  1653 => x"00000000",
  1654 => x"00000000",
  1655 => x"00000000",
  1656 => x"00000000",
  1657 => x"00000000",
  1658 => x"00000000",
  1659 => x"00001974",
  1660 => x"00000000",
  1661 => x"00000000",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00000000",
  1666 => x"00000000",
  1667 => x"00000000",
  1668 => x"00000000",
  1669 => x"00000000",
  1670 => x"00000000",
  1671 => x"00000000",
  1672 => x"00000000",
  1673 => x"00000000",
  1674 => x"00000000",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00000000",
  1678 => x"00000000",
  1679 => x"00000000",
  1680 => x"00000000",
  1681 => x"00000000",
  1682 => x"00000000",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000001",
  1689 => x"330eabcd",
  1690 => x"1234e66d",
  1691 => x"deec0005",
  1692 => x"000b0000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"00000000",
  1717 => x"00000000",
  1718 => x"00000000",
  1719 => x"00000000",
  1720 => x"00000000",
  1721 => x"00000000",
  1722 => x"00000000",
  1723 => x"00000000",
  1724 => x"00000000",
  1725 => x"00000000",
  1726 => x"00000000",
  1727 => x"00000000",
  1728 => x"00000000",
  1729 => x"00000000",
  1730 => x"00000000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"00000000",
  1737 => x"00000000",
  1738 => x"00000000",
  1739 => x"00000000",
  1740 => x"00000000",
  1741 => x"00000000",
  1742 => x"00000000",
  1743 => x"00000000",
  1744 => x"00000000",
  1745 => x"00000000",
  1746 => x"00000000",
  1747 => x"00000000",
  1748 => x"00000000",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000000",
  1785 => x"00000000",
  1786 => x"00000000",
  1787 => x"00000000",
  1788 => x"00000000",
  1789 => x"00000000",
  1790 => x"00000000",
  1791 => x"00000000",
  1792 => x"00000000",
  1793 => x"00000000",
  1794 => x"00000000",
  1795 => x"00000000",
  1796 => x"00000000",
  1797 => x"00000000",
  1798 => x"00000000",
  1799 => x"00000000",
  1800 => x"00000000",
  1801 => x"00000000",
  1802 => x"00000000",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"00000000",
  1807 => x"00000000",
  1808 => x"00000000",
  1809 => x"00000000",
  1810 => x"00000000",
  1811 => x"00000000",
  1812 => x"00000000",
  1813 => x"00000000",
  1814 => x"00000000",
  1815 => x"00000000",
  1816 => x"00000000",
  1817 => x"00000000",
  1818 => x"00000000",
  1819 => x"00000000",
  1820 => x"00000000",
  1821 => x"00000000",
  1822 => x"00000000",
  1823 => x"00000000",
  1824 => x"00000000",
  1825 => x"00000000",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00000000",
  1829 => x"00000000",
  1830 => x"00000000",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000000",
  1834 => x"00000000",
  1835 => x"00000000",
  1836 => x"00000000",
  1837 => x"00000000",
  1838 => x"00000000",
  1839 => x"00000000",
  1840 => x"00000000",
  1841 => x"00000000",
  1842 => x"00000000",
  1843 => x"00000000",
  1844 => x"00000000",
  1845 => x"00000000",
  1846 => x"00000000",
  1847 => x"00000000",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00000000",
  1853 => x"00000000",
  1854 => x"00000000",
  1855 => x"00000000",
  1856 => x"00000000",
  1857 => x"00000000",
  1858 => x"00000000",
  1859 => x"00000000",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"00000000",
  1868 => x"00000000",
  1869 => x"ffffffff",
  1870 => x"00000000",
  1871 => x"ffffffff",
  1872 => x"00000000",
  1873 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
