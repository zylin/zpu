-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0bbd9c0c",
     3 => x"3a0b0b0b",
     4 => x"aed50400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0baf992d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bbd",
   162 => x"88738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b92",
   171 => x"c02d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b93",
   179 => x"f22d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bbd980c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81fb3fa8",
   257 => x"b93f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104bd",
   280 => x"9808802e",
   281 => x"a338bd9c",
   282 => x"08822ebd",
   283 => x"38838080",
   284 => x"0b0b0b80",
   285 => x"cda00c82",
   286 => x"a0800b80",
   287 => x"cda40c82",
   288 => x"90800b80",
   289 => x"cda80c04",
   290 => x"f8808080",
   291 => x"a40b0b0b",
   292 => x"80cda00c",
   293 => x"f8808082",
   294 => x"800b80cd",
   295 => x"a40cf880",
   296 => x"8084800b",
   297 => x"80cda80c",
   298 => x"0480c0a8",
   299 => x"808c0b0b",
   300 => x"0b80cda0",
   301 => x"0c80c0a8",
   302 => x"80940b80",
   303 => x"cda40c0b",
   304 => x"0b0bb0ec",
   305 => x"0b80cda8",
   306 => x"0c04ff3d",
   307 => x"0d80cdac",
   308 => x"335170a4",
   309 => x"38bda408",
   310 => x"70085252",
   311 => x"70802e92",
   312 => x"388412bd",
   313 => x"a40c702d",
   314 => x"bda40870",
   315 => x"08525270",
   316 => x"f038810b",
   317 => x"80cdac34",
   318 => x"833d0d04",
   319 => x"04803d0d",
   320 => x"0b0b80cd",
   321 => x"9c08802e",
   322 => x"8e380b0b",
   323 => x"0b0b800b",
   324 => x"802e0981",
   325 => x"06853882",
   326 => x"3d0d040b",
   327 => x"0b80cd9c",
   328 => x"510b0b0b",
   329 => x"f5da3f82",
   330 => x"3d0d0404",
   331 => x"ff3d0d02",
   332 => x"8f053370",
   333 => x"5252868f",
   334 => x"3f715187",
   335 => x"813f7180",
   336 => x"0c833d0d",
   337 => x"04ff3d0d",
   338 => x"028f0533",
   339 => x"bdac0871",
   340 => x"710c5380",
   341 => x"0c833d0d",
   342 => x"04f63d0d",
   343 => x"bdb40870",
   344 => x"08810a06",
   345 => x"80cdb00c",
   346 => x"5485ac3f",
   347 => x"85c43f8a",
   348 => x"c55380cd",
   349 => x"b0088438",
   350 => x"8aac5372",
   351 => x"80cdb40c",
   352 => x"86993fbd",
   353 => x"a80854fa",
   354 => x"c98e868c",
   355 => x"740c7308",
   356 => x"70842a81",
   357 => x"06545672",
   358 => x"f538bdb0",
   359 => x"08738412",
   360 => x"0c549480",
   361 => x"0b88150c",
   362 => x"82d0affd",
   363 => x"fb0b8c15",
   364 => x"0c80c074",
   365 => x"0c730870",
   366 => x"862a8106",
   367 => x"545672f5",
   368 => x"38901408",
   369 => x"70832a81",
   370 => x"06545672",
   371 => x"f43881fc",
   372 => x"80810b90",
   373 => x"150c9014",
   374 => x"0870832a",
   375 => x"81065456",
   376 => x"72f43883",
   377 => x"f0820b90",
   378 => x"150c9014",
   379 => x"0870832a",
   380 => x"81065456",
   381 => x"72f43890",
   382 => x"14087096",
   383 => x"2a810654",
   384 => x"5672d338",
   385 => x"90140870",
   386 => x"832a8106",
   387 => x"545672f4",
   388 => x"3880fdc0",
   389 => x"810b9015",
   390 => x"0cbc8051",
   391 => x"828d3f80",
   392 => x"cdb00880",
   393 => x"2e81f038",
   394 => x"bc885181",
   395 => x"fe3fbc94",
   396 => x"5181f83f",
   397 => x"b3b05181",
   398 => x"f23f8054",
   399 => x"800bfa80",
   400 => x"8080840c",
   401 => x"bbea0b85",
   402 => x"0a0cbdb0",
   403 => x"0853850a",
   404 => x"0b94140c",
   405 => x"91730c85",
   406 => x"0a08708b",
   407 => x"2a810656",
   408 => x"5374f438",
   409 => x"b2d85181",
   410 => x"c23fbdb0",
   411 => x"08700853",
   412 => x"53a05181",
   413 => x"d93fb2ec",
   414 => x"5181b03f",
   415 => x"bdb00884",
   416 => x"11085356",
   417 => x"a05181c6",
   418 => x"3fb38051",
   419 => x"819d3f85",
   420 => x"0a0852a0",
   421 => x"5181b73f",
   422 => x"81147081",
   423 => x"ff065555",
   424 => x"937427ff",
   425 => x"9738f881",
   426 => x"c08e8054",
   427 => x"a00bbdb4",
   428 => x"08565680",
   429 => x"cdb00880",
   430 => x"2eab3873",
   431 => x"81ff0684",
   432 => x"160c739f",
   433 => x"2a741007",
   434 => x"5475802e",
   435 => x"9538ff16",
   436 => x"7481ff06",
   437 => x"84170c74",
   438 => x"9f2a7510",
   439 => x"07555675",
   440 => x"ed3888d8",
   441 => x"3f7381ff",
   442 => x"0684160c",
   443 => x"739f2a74",
   444 => x"10075480",
   445 => x"fd5181fd",
   446 => x"3fbdb408",
   447 => x"7481ff06",
   448 => x"84120c55",
   449 => x"739f2a74",
   450 => x"10075480",
   451 => x"fd5181e5",
   452 => x"3fbdb408",
   453 => x"55cf39bc",
   454 => x"b851903f",
   455 => x"bc94518b",
   456 => x"3fb3b051",
   457 => x"863f8054",
   458 => x"fe9239fe",
   459 => x"3d0d7470",
   460 => x"33535371",
   461 => x"802e9338",
   462 => x"81137252",
   463 => x"80cdb408",
   464 => x"5353712d",
   465 => x"72335271",
   466 => x"ef38843d",
   467 => x"0d04f43d",
   468 => x"0d7f0284",
   469 => x"05bb0533",
   470 => x"5557a00b",
   471 => x"8c3d5b59",
   472 => x"8b53bcec",
   473 => x"52795187",
   474 => x"e03f7388",
   475 => x"2e818038",
   476 => x"78567390",
   477 => x"2e80ed38",
   478 => x"02a90558",
   479 => x"768f0654",
   480 => x"73892680",
   481 => x"c3387518",
   482 => x"b0155555",
   483 => x"73753476",
   484 => x"842aff17",
   485 => x"7081ff06",
   486 => x"58555775",
   487 => x"df388e3d",
   488 => x"7905f605",
   489 => x"57757734",
   490 => x"79703355",
   491 => x"5573802e",
   492 => x"93388115",
   493 => x"745280cd",
   494 => x"b4085755",
   495 => x"752d7433",
   496 => x"5473ef38",
   497 => x"8e3d0d04",
   498 => x"7518b715",
   499 => x"55557375",
   500 => x"3476842a",
   501 => x"ff177081",
   502 => x"ff065855",
   503 => x"5775ff9c",
   504 => x"38ffbb39",
   505 => x"84705759",
   506 => x"02a90558",
   507 => x"ff8e3982",
   508 => x"705759f4",
   509 => x"39fd3d0d",
   510 => x"bdbc0876",
   511 => x"b0ea2994",
   512 => x"120c5485",
   513 => x"0b98150c",
   514 => x"98140870",
   515 => x"81065153",
   516 => x"72f63885",
   517 => x"3d0d0480",
   518 => x"3d0dbdbc",
   519 => x"0851870b",
   520 => x"84120cb0",
   521 => x"ea0ba412",
   522 => x"0c870ba8",
   523 => x"120c823d",
   524 => x"0d04803d",
   525 => x"0dbdc008",
   526 => x"51b60b8c",
   527 => x"120c830b",
   528 => x"88120c82",
   529 => x"3d0d04fe",
   530 => x"3d0d0293",
   531 => x"05335372",
   532 => x"8a2e9d38",
   533 => x"bdc00852",
   534 => x"84120870",
   535 => x"822a7081",
   536 => x"06515151",
   537 => x"70802ef0",
   538 => x"3872720c",
   539 => x"843d0d04",
   540 => x"bdc00852",
   541 => x"84120870",
   542 => x"822a7081",
   543 => x"06515151",
   544 => x"70802ef0",
   545 => x"388d720c",
   546 => x"84120870",
   547 => x"822a7081",
   548 => x"06515151",
   549 => x"70802ec0",
   550 => x"38cf3980",
   551 => x"3d0dbdb8",
   552 => x"0851800b",
   553 => x"84120cfe",
   554 => x"800a0b88",
   555 => x"120c800b",
   556 => x"80cdb834",
   557 => x"800b80cd",
   558 => x"bc34823d",
   559 => x"0d04fa3d",
   560 => x"0d02a305",
   561 => x"33bdb808",
   562 => x"80cdb833",
   563 => x"7081ff06",
   564 => x"70101011",
   565 => x"80cdbc33",
   566 => x"7081ff06",
   567 => x"72902911",
   568 => x"70882b78",
   569 => x"07770c53",
   570 => x"5b5b5555",
   571 => x"59545473",
   572 => x"8a2e9838",
   573 => x"7480cf2e",
   574 => x"9238738c",
   575 => x"2ea43881",
   576 => x"16537280",
   577 => x"cdbc3488",
   578 => x"3d0d0471",
   579 => x"a326a338",
   580 => x"81175271",
   581 => x"80cdb834",
   582 => x"800b80cd",
   583 => x"bc34883d",
   584 => x"0d048052",
   585 => x"71882b73",
   586 => x"0c811252",
   587 => x"97907226",
   588 => x"f338800b",
   589 => x"80cdb834",
   590 => x"800b80cd",
   591 => x"bc34df39",
   592 => x"8c08028c",
   593 => x"0cf93d0d",
   594 => x"800b8c08",
   595 => x"fc050c8c",
   596 => x"08880508",
   597 => x"8025ab38",
   598 => x"8c088805",
   599 => x"08308c08",
   600 => x"88050c80",
   601 => x"0b8c08f4",
   602 => x"050c8c08",
   603 => x"fc050888",
   604 => x"38810b8c",
   605 => x"08f4050c",
   606 => x"8c08f405",
   607 => x"088c08fc",
   608 => x"050c8c08",
   609 => x"8c050880",
   610 => x"25ab388c",
   611 => x"088c0508",
   612 => x"308c088c",
   613 => x"050c800b",
   614 => x"8c08f005",
   615 => x"0c8c08fc",
   616 => x"05088838",
   617 => x"810b8c08",
   618 => x"f0050c8c",
   619 => x"08f00508",
   620 => x"8c08fc05",
   621 => x"0c80538c",
   622 => x"088c0508",
   623 => x"528c0888",
   624 => x"05085181",
   625 => x"a73f8008",
   626 => x"708c08f8",
   627 => x"050c548c",
   628 => x"08fc0508",
   629 => x"802e8c38",
   630 => x"8c08f805",
   631 => x"08308c08",
   632 => x"f8050c8c",
   633 => x"08f80508",
   634 => x"70800c54",
   635 => x"893d0d8c",
   636 => x"0c048c08",
   637 => x"028c0cfb",
   638 => x"3d0d800b",
   639 => x"8c08fc05",
   640 => x"0c8c0888",
   641 => x"05088025",
   642 => x"93388c08",
   643 => x"88050830",
   644 => x"8c088805",
   645 => x"0c810b8c",
   646 => x"08fc050c",
   647 => x"8c088c05",
   648 => x"0880258c",
   649 => x"388c088c",
   650 => x"0508308c",
   651 => x"088c050c",
   652 => x"81538c08",
   653 => x"8c050852",
   654 => x"8c088805",
   655 => x"0851ad3f",
   656 => x"8008708c",
   657 => x"08f8050c",
   658 => x"548c08fc",
   659 => x"0508802e",
   660 => x"8c388c08",
   661 => x"f8050830",
   662 => x"8c08f805",
   663 => x"0c8c08f8",
   664 => x"05087080",
   665 => x"0c54873d",
   666 => x"0d8c0c04",
   667 => x"8c08028c",
   668 => x"0cfd3d0d",
   669 => x"810b8c08",
   670 => x"fc050c80",
   671 => x"0b8c08f8",
   672 => x"050c8c08",
   673 => x"8c05088c",
   674 => x"08880508",
   675 => x"27ac388c",
   676 => x"08fc0508",
   677 => x"802ea338",
   678 => x"800b8c08",
   679 => x"8c050824",
   680 => x"99388c08",
   681 => x"8c050810",
   682 => x"8c088c05",
   683 => x"0c8c08fc",
   684 => x"0508108c",
   685 => x"08fc050c",
   686 => x"c9398c08",
   687 => x"fc050880",
   688 => x"2e80c938",
   689 => x"8c088c05",
   690 => x"088c0888",
   691 => x"050826a1",
   692 => x"388c0888",
   693 => x"05088c08",
   694 => x"8c050831",
   695 => x"8c088805",
   696 => x"0c8c08f8",
   697 => x"05088c08",
   698 => x"fc050807",
   699 => x"8c08f805",
   700 => x"0c8c08fc",
   701 => x"0508812a",
   702 => x"8c08fc05",
   703 => x"0c8c088c",
   704 => x"0508812a",
   705 => x"8c088c05",
   706 => x"0cffaf39",
   707 => x"8c089005",
   708 => x"08802e8f",
   709 => x"388c0888",
   710 => x"0508708c",
   711 => x"08f4050c",
   712 => x"518d398c",
   713 => x"08f80508",
   714 => x"708c08f4",
   715 => x"050c518c",
   716 => x"08f40508",
   717 => x"800c853d",
   718 => x"0d8c0c04",
   719 => x"803d0d86",
   720 => x"5184963f",
   721 => x"815198ce",
   722 => x"3ffc3d0d",
   723 => x"7670797b",
   724 => x"55555555",
   725 => x"8f72278c",
   726 => x"38727507",
   727 => x"83065170",
   728 => x"802ea738",
   729 => x"ff125271",
   730 => x"ff2e9838",
   731 => x"72708105",
   732 => x"54337470",
   733 => x"81055634",
   734 => x"ff125271",
   735 => x"ff2e0981",
   736 => x"06ea3874",
   737 => x"800c863d",
   738 => x"0d047451",
   739 => x"72708405",
   740 => x"54087170",
   741 => x"8405530c",
   742 => x"72708405",
   743 => x"54087170",
   744 => x"8405530c",
   745 => x"72708405",
   746 => x"54087170",
   747 => x"8405530c",
   748 => x"72708405",
   749 => x"54087170",
   750 => x"8405530c",
   751 => x"f0125271",
   752 => x"8f26c938",
   753 => x"83722795",
   754 => x"38727084",
   755 => x"05540871",
   756 => x"70840553",
   757 => x"0cfc1252",
   758 => x"718326ed",
   759 => x"387054ff",
   760 => x"8339fd3d",
   761 => x"0d755384",
   762 => x"d8130880",
   763 => x"2e8a3880",
   764 => x"5372800c",
   765 => x"853d0d04",
   766 => x"81805272",
   767 => x"5183d43f",
   768 => x"800884d8",
   769 => x"140cff53",
   770 => x"8008802e",
   771 => x"e4388008",
   772 => x"549f5380",
   773 => x"74708405",
   774 => x"560cff13",
   775 => x"53807324",
   776 => x"ce388074",
   777 => x"70840556",
   778 => x"0cff1353",
   779 => x"728025e3",
   780 => x"38ffbc39",
   781 => x"fd3d0d75",
   782 => x"7755539f",
   783 => x"74278d38",
   784 => x"96730cff",
   785 => x"5271800c",
   786 => x"853d0d04",
   787 => x"84d81308",
   788 => x"5271802e",
   789 => x"93387310",
   790 => x"10127008",
   791 => x"79720c51",
   792 => x"5271800c",
   793 => x"853d0d04",
   794 => x"7251fef6",
   795 => x"3fff5280",
   796 => x"08d33884",
   797 => x"d8130874",
   798 => x"10101170",
   799 => x"087a720c",
   800 => x"515152dd",
   801 => x"39f93d0d",
   802 => x"797b5856",
   803 => x"769f2680",
   804 => x"e83884d8",
   805 => x"16085473",
   806 => x"802eaa38",
   807 => x"76101014",
   808 => x"70085555",
   809 => x"73802eba",
   810 => x"38805873",
   811 => x"812e8f38",
   812 => x"73ff2ea3",
   813 => x"3880750c",
   814 => x"7651732d",
   815 => x"80587780",
   816 => x"0c893d0d",
   817 => x"047551fe",
   818 => x"993fff58",
   819 => x"8008ef38",
   820 => x"84d81608",
   821 => x"54c63996",
   822 => x"760c810b",
   823 => x"800c893d",
   824 => x"0d047551",
   825 => x"81e93f76",
   826 => x"53800852",
   827 => x"755181a9",
   828 => x"3f800880",
   829 => x"0c893d0d",
   830 => x"0496760c",
   831 => x"ff0b800c",
   832 => x"893d0d04",
   833 => x"fc3d0d76",
   834 => x"785653ff",
   835 => x"54749f26",
   836 => x"b13884d8",
   837 => x"13085271",
   838 => x"802eae38",
   839 => x"74101012",
   840 => x"70085353",
   841 => x"81547180",
   842 => x"2e983882",
   843 => x"5471ff2e",
   844 => x"91388354",
   845 => x"71812e8a",
   846 => x"3880730c",
   847 => x"7451712d",
   848 => x"80547380",
   849 => x"0c863d0d",
   850 => x"047251fd",
   851 => x"953f8008",
   852 => x"f13884d8",
   853 => x"130852c4",
   854 => x"39ff3d0d",
   855 => x"7352bdc4",
   856 => x"0851fea1",
   857 => x"3f833d0d",
   858 => x"04fe3d0d",
   859 => x"75537452",
   860 => x"bdc40851",
   861 => x"fdbe3f84",
   862 => x"3d0d0480",
   863 => x"3d0dbdc4",
   864 => x"0851fcde",
   865 => x"3f823d0d",
   866 => x"04ff3d0d",
   867 => x"7352bdc4",
   868 => x"0851fef0",
   869 => x"3f833d0d",
   870 => x"04fc3d0d",
   871 => x"800b80cd",
   872 => x"c80c7852",
   873 => x"775192e7",
   874 => x"3f800854",
   875 => x"8008ff2e",
   876 => x"88387380",
   877 => x"0c863d0d",
   878 => x"0480cdc8",
   879 => x"08557480",
   880 => x"2ef03876",
   881 => x"75710c53",
   882 => x"73800c86",
   883 => x"3d0d0492",
   884 => x"b93f04f3",
   885 => x"3d0d7f61",
   886 => x"8b1170f8",
   887 => x"065c5555",
   888 => x"5e729626",
   889 => x"83389059",
   890 => x"80792474",
   891 => x"7a260753",
   892 => x"80547274",
   893 => x"2e098106",
   894 => x"80cb387d",
   895 => x"518bca3f",
   896 => x"7883f726",
   897 => x"80c63878",
   898 => x"832a7010",
   899 => x"101080c5",
   900 => x"80058c11",
   901 => x"0859595a",
   902 => x"76782e83",
   903 => x"b0388417",
   904 => x"08fc0656",
   905 => x"8c170888",
   906 => x"1808718c",
   907 => x"120c8812",
   908 => x"0c587517",
   909 => x"84110881",
   910 => x"0784120c",
   911 => x"537d518b",
   912 => x"893f8817",
   913 => x"5473800c",
   914 => x"8f3d0d04",
   915 => x"78892a79",
   916 => x"832a5b53",
   917 => x"72802ebf",
   918 => x"3878862a",
   919 => x"b8055a84",
   920 => x"7327b438",
   921 => x"80db135a",
   922 => x"947327ab",
   923 => x"38788c2a",
   924 => x"80ee055a",
   925 => x"80d47327",
   926 => x"9e38788f",
   927 => x"2a80f705",
   928 => x"5a82d473",
   929 => x"27913878",
   930 => x"922a80fc",
   931 => x"055a8ad4",
   932 => x"73278438",
   933 => x"80fe5a79",
   934 => x"10101080",
   935 => x"c580058c",
   936 => x"11085855",
   937 => x"76752ea3",
   938 => x"38841708",
   939 => x"fc06707a",
   940 => x"31555673",
   941 => x"8f2488d5",
   942 => x"38738025",
   943 => x"fee6388c",
   944 => x"17085776",
   945 => x"752e0981",
   946 => x"06df3881",
   947 => x"1a5a80c5",
   948 => x"90085776",
   949 => x"80c5882e",
   950 => x"82c03884",
   951 => x"1708fc06",
   952 => x"707a3155",
   953 => x"56738f24",
   954 => x"81f93880",
   955 => x"c5880b80",
   956 => x"c5940c80",
   957 => x"c5880b80",
   958 => x"c5900c73",
   959 => x"8025feb2",
   960 => x"3883ff76",
   961 => x"2783df38",
   962 => x"75892a76",
   963 => x"832a5553",
   964 => x"72802ebf",
   965 => x"3875862a",
   966 => x"b8055484",
   967 => x"7327b438",
   968 => x"80db1354",
   969 => x"947327ab",
   970 => x"38758c2a",
   971 => x"80ee0554",
   972 => x"80d47327",
   973 => x"9e38758f",
   974 => x"2a80f705",
   975 => x"5482d473",
   976 => x"27913875",
   977 => x"922a80fc",
   978 => x"05548ad4",
   979 => x"73278438",
   980 => x"80fe5473",
   981 => x"10101080",
   982 => x"c5800588",
   983 => x"11085658",
   984 => x"74782e86",
   985 => x"cf388415",
   986 => x"08fc0653",
   987 => x"7573278d",
   988 => x"38881508",
   989 => x"5574782e",
   990 => x"098106ea",
   991 => x"388c1508",
   992 => x"80c5800b",
   993 => x"84050871",
   994 => x"8c1a0c76",
   995 => x"881a0c78",
   996 => x"88130c78",
   997 => x"8c180c5d",
   998 => x"58795380",
   999 => x"7a2483e6",
  1000 => x"3872822c",
  1001 => x"81712b5c",
  1002 => x"537a7c26",
  1003 => x"8198387b",
  1004 => x"7b065372",
  1005 => x"82f13879",
  1006 => x"fc068405",
  1007 => x"5a7a1070",
  1008 => x"7d06545b",
  1009 => x"7282e038",
  1010 => x"841a5af1",
  1011 => x"3988178c",
  1012 => x"11085858",
  1013 => x"76782e09",
  1014 => x"8106fcc2",
  1015 => x"38821a5a",
  1016 => x"fdec3978",
  1017 => x"17798107",
  1018 => x"84190c70",
  1019 => x"80c5940c",
  1020 => x"7080c590",
  1021 => x"0c80c588",
  1022 => x"0b8c120c",
  1023 => x"8c110888",
  1024 => x"120c7481",
  1025 => x"0784120c",
  1026 => x"74117571",
  1027 => x"0c51537d",
  1028 => x"5187b73f",
  1029 => x"881754fc",
  1030 => x"ac3980c5",
  1031 => x"800b8405",
  1032 => x"087a545c",
  1033 => x"798025fe",
  1034 => x"f83882da",
  1035 => x"397a097c",
  1036 => x"067080c5",
  1037 => x"800b8405",
  1038 => x"0c5c7a10",
  1039 => x"5b7a7c26",
  1040 => x"85387a85",
  1041 => x"b83880c5",
  1042 => x"800b8805",
  1043 => x"08708412",
  1044 => x"08fc0670",
  1045 => x"7c317c72",
  1046 => x"268f7225",
  1047 => x"0757575c",
  1048 => x"5d557280",
  1049 => x"2e80db38",
  1050 => x"797a1680",
  1051 => x"c4f8081b",
  1052 => x"90115a55",
  1053 => x"575b80c4",
  1054 => x"f408ff2e",
  1055 => x"8838a08f",
  1056 => x"13e08006",
  1057 => x"5776527d",
  1058 => x"5186c03f",
  1059 => x"80085480",
  1060 => x"08ff2e90",
  1061 => x"38800876",
  1062 => x"27829938",
  1063 => x"7480c580",
  1064 => x"2e829138",
  1065 => x"80c5800b",
  1066 => x"88050855",
  1067 => x"841508fc",
  1068 => x"06707a31",
  1069 => x"7a72268f",
  1070 => x"72250752",
  1071 => x"55537283",
  1072 => x"e6387479",
  1073 => x"81078417",
  1074 => x"0c791670",
  1075 => x"80c5800b",
  1076 => x"88050c75",
  1077 => x"81078412",
  1078 => x"0c547e52",
  1079 => x"5785eb3f",
  1080 => x"881754fa",
  1081 => x"e0397583",
  1082 => x"2a705454",
  1083 => x"80742481",
  1084 => x"9b387282",
  1085 => x"2c81712b",
  1086 => x"80c58408",
  1087 => x"077080c5",
  1088 => x"800b8405",
  1089 => x"0c751010",
  1090 => x"1080c580",
  1091 => x"05881108",
  1092 => x"585a5d53",
  1093 => x"778c180c",
  1094 => x"7488180c",
  1095 => x"7688190c",
  1096 => x"768c160c",
  1097 => x"fcf33979",
  1098 => x"7a101010",
  1099 => x"80c58005",
  1100 => x"7057595d",
  1101 => x"8c150857",
  1102 => x"76752ea3",
  1103 => x"38841708",
  1104 => x"fc06707a",
  1105 => x"31555673",
  1106 => x"8f2483ca",
  1107 => x"38738025",
  1108 => x"8481388c",
  1109 => x"17085776",
  1110 => x"752e0981",
  1111 => x"06df3888",
  1112 => x"15811b70",
  1113 => x"8306555b",
  1114 => x"5572c938",
  1115 => x"7c830653",
  1116 => x"72802efd",
  1117 => x"b838ff1d",
  1118 => x"f819595d",
  1119 => x"88180878",
  1120 => x"2eea38fd",
  1121 => x"b539831a",
  1122 => x"53fc9639",
  1123 => x"83147082",
  1124 => x"2c81712b",
  1125 => x"80c58408",
  1126 => x"077080c5",
  1127 => x"800b8405",
  1128 => x"0c761010",
  1129 => x"1080c580",
  1130 => x"05881108",
  1131 => x"595b5e51",
  1132 => x"53fee139",
  1133 => x"80c4c408",
  1134 => x"17588008",
  1135 => x"762e818d",
  1136 => x"3880c4f4",
  1137 => x"08ff2e83",
  1138 => x"ec387376",
  1139 => x"311880c4",
  1140 => x"c40c7387",
  1141 => x"06705753",
  1142 => x"72802e88",
  1143 => x"38887331",
  1144 => x"70155556",
  1145 => x"76149fff",
  1146 => x"06a08071",
  1147 => x"31177054",
  1148 => x"7f535753",
  1149 => x"83d53f80",
  1150 => x"08538008",
  1151 => x"ff2e81a0",
  1152 => x"3880c4c4",
  1153 => x"08167080",
  1154 => x"c4c40c74",
  1155 => x"7580c580",
  1156 => x"0b88050c",
  1157 => x"74763118",
  1158 => x"70810751",
  1159 => x"5556587b",
  1160 => x"80c5802e",
  1161 => x"839c3879",
  1162 => x"8f2682cb",
  1163 => x"38810b84",
  1164 => x"150c8415",
  1165 => x"08fc0670",
  1166 => x"7a317a72",
  1167 => x"268f7225",
  1168 => x"07525553",
  1169 => x"72802efc",
  1170 => x"f93880db",
  1171 => x"3980089f",
  1172 => x"ff065372",
  1173 => x"feeb3877",
  1174 => x"80c4c40c",
  1175 => x"80c5800b",
  1176 => x"8805087b",
  1177 => x"18810784",
  1178 => x"120c5580",
  1179 => x"c4f00878",
  1180 => x"27863877",
  1181 => x"80c4f00c",
  1182 => x"80c4ec08",
  1183 => x"7827fcac",
  1184 => x"387780c4",
  1185 => x"ec0c8415",
  1186 => x"08fc0670",
  1187 => x"7a317a72",
  1188 => x"268f7225",
  1189 => x"07525553",
  1190 => x"72802efc",
  1191 => x"a5388839",
  1192 => x"80745456",
  1193 => x"fedb397d",
  1194 => x"51829f3f",
  1195 => x"800b800c",
  1196 => x"8f3d0d04",
  1197 => x"73538074",
  1198 => x"24a93872",
  1199 => x"822c8171",
  1200 => x"2b80c584",
  1201 => x"08077080",
  1202 => x"c5800b84",
  1203 => x"050c5d53",
  1204 => x"778c180c",
  1205 => x"7488180c",
  1206 => x"7688190c",
  1207 => x"768c160c",
  1208 => x"f9b73983",
  1209 => x"1470822c",
  1210 => x"81712b80",
  1211 => x"c5840807",
  1212 => x"7080c580",
  1213 => x"0b84050c",
  1214 => x"5e5153d4",
  1215 => x"397b7b06",
  1216 => x"5372fca3",
  1217 => x"38841a7b",
  1218 => x"105c5af1",
  1219 => x"39ff1a81",
  1220 => x"11515af7",
  1221 => x"b9397817",
  1222 => x"79810784",
  1223 => x"190c8c18",
  1224 => x"08881908",
  1225 => x"718c120c",
  1226 => x"88120c59",
  1227 => x"7080c594",
  1228 => x"0c7080c5",
  1229 => x"900c80c5",
  1230 => x"880b8c12",
  1231 => x"0c8c1108",
  1232 => x"88120c74",
  1233 => x"81078412",
  1234 => x"0c741175",
  1235 => x"710c5153",
  1236 => x"f9bd3975",
  1237 => x"17841108",
  1238 => x"81078412",
  1239 => x"0c538c17",
  1240 => x"08881808",
  1241 => x"718c120c",
  1242 => x"88120c58",
  1243 => x"7d5180da",
  1244 => x"3f881754",
  1245 => x"f5cf3972",
  1246 => x"84150cf4",
  1247 => x"1af80670",
  1248 => x"841e0881",
  1249 => x"0607841e",
  1250 => x"0c701d54",
  1251 => x"5b850b84",
  1252 => x"140c850b",
  1253 => x"88140c8f",
  1254 => x"7b27fdcf",
  1255 => x"38881c52",
  1256 => x"7d518290",
  1257 => x"3f80c580",
  1258 => x"0b880508",
  1259 => x"80c4c408",
  1260 => x"5955fdb7",
  1261 => x"397780c4",
  1262 => x"c40c7380",
  1263 => x"c4f40cfc",
  1264 => x"91397284",
  1265 => x"150cfda3",
  1266 => x"390404fd",
  1267 => x"3d0d800b",
  1268 => x"80cdc80c",
  1269 => x"765186cc",
  1270 => x"3f800853",
  1271 => x"8008ff2e",
  1272 => x"88387280",
  1273 => x"0c853d0d",
  1274 => x"0480cdc8",
  1275 => x"08547380",
  1276 => x"2ef03875",
  1277 => x"74710c52",
  1278 => x"72800c85",
  1279 => x"3d0d04fb",
  1280 => x"3d0d7770",
  1281 => x"5256c23f",
  1282 => x"80c5800b",
  1283 => x"88050884",
  1284 => x"1108fc06",
  1285 => x"707b319f",
  1286 => x"ef05e080",
  1287 => x"06e08005",
  1288 => x"565653a0",
  1289 => x"80742494",
  1290 => x"38805275",
  1291 => x"51ff9c3f",
  1292 => x"80c58808",
  1293 => x"15537280",
  1294 => x"082e8f38",
  1295 => x"7551ff8a",
  1296 => x"3f805372",
  1297 => x"800c873d",
  1298 => x"0d047330",
  1299 => x"527551fe",
  1300 => x"fa3f8008",
  1301 => x"ff2ea838",
  1302 => x"80c5800b",
  1303 => x"88050875",
  1304 => x"75318107",
  1305 => x"84120c53",
  1306 => x"80c4c408",
  1307 => x"743180c4",
  1308 => x"c40c7551",
  1309 => x"fed43f81",
  1310 => x"0b800c87",
  1311 => x"3d0d0480",
  1312 => x"527551fe",
  1313 => x"c63f80c5",
  1314 => x"800b8805",
  1315 => x"08800871",
  1316 => x"3156538f",
  1317 => x"7525ffa4",
  1318 => x"38800880",
  1319 => x"c4f40831",
  1320 => x"80c4c40c",
  1321 => x"74810784",
  1322 => x"140c7551",
  1323 => x"fe9c3f80",
  1324 => x"53ff9039",
  1325 => x"f63d0d7c",
  1326 => x"7e545b72",
  1327 => x"802e8283",
  1328 => x"387a51fe",
  1329 => x"843ff813",
  1330 => x"84110870",
  1331 => x"fe067013",
  1332 => x"841108fc",
  1333 => x"065d5859",
  1334 => x"545880c5",
  1335 => x"8808752e",
  1336 => x"82de3878",
  1337 => x"84160c80",
  1338 => x"73810654",
  1339 => x"5a727a2e",
  1340 => x"81d53878",
  1341 => x"15841108",
  1342 => x"81065153",
  1343 => x"72a03878",
  1344 => x"17577981",
  1345 => x"e6388815",
  1346 => x"08537280",
  1347 => x"c5882e82",
  1348 => x"f9388c15",
  1349 => x"08708c15",
  1350 => x"0c738812",
  1351 => x"0c567681",
  1352 => x"0784190c",
  1353 => x"76187771",
  1354 => x"0c537981",
  1355 => x"913883ff",
  1356 => x"772781c8",
  1357 => x"3876892a",
  1358 => x"77832a56",
  1359 => x"5372802e",
  1360 => x"bf387686",
  1361 => x"2ab80555",
  1362 => x"847327b4",
  1363 => x"3880db13",
  1364 => x"55947327",
  1365 => x"ab38768c",
  1366 => x"2a80ee05",
  1367 => x"5580d473",
  1368 => x"279e3876",
  1369 => x"8f2a80f7",
  1370 => x"055582d4",
  1371 => x"73279138",
  1372 => x"76922a80",
  1373 => x"fc05558a",
  1374 => x"d4732784",
  1375 => x"3880fe55",
  1376 => x"74101010",
  1377 => x"80c58005",
  1378 => x"88110855",
  1379 => x"5673762e",
  1380 => x"82b33884",
  1381 => x"1408fc06",
  1382 => x"53767327",
  1383 => x"8d388814",
  1384 => x"08547376",
  1385 => x"2e098106",
  1386 => x"ea388c14",
  1387 => x"08708c1a",
  1388 => x"0c74881a",
  1389 => x"0c788812",
  1390 => x"0c56778c",
  1391 => x"150c7a51",
  1392 => x"fc883f8c",
  1393 => x"3d0d0477",
  1394 => x"08787131",
  1395 => x"59770588",
  1396 => x"19085457",
  1397 => x"7280c588",
  1398 => x"2e80e038",
  1399 => x"8c180870",
  1400 => x"8c150c73",
  1401 => x"88120c56",
  1402 => x"fe893988",
  1403 => x"15088c16",
  1404 => x"08708c13",
  1405 => x"0c578817",
  1406 => x"0cfea339",
  1407 => x"76832a70",
  1408 => x"54558075",
  1409 => x"24819838",
  1410 => x"72822c81",
  1411 => x"712b80c5",
  1412 => x"84080780",
  1413 => x"c5800b84",
  1414 => x"050c5374",
  1415 => x"10101080",
  1416 => x"c5800588",
  1417 => x"11085556",
  1418 => x"758c190c",
  1419 => x"7388190c",
  1420 => x"7788170c",
  1421 => x"778c150c",
  1422 => x"ff843981",
  1423 => x"5afdb439",
  1424 => x"78177381",
  1425 => x"06545772",
  1426 => x"98387708",
  1427 => x"78713159",
  1428 => x"77058c19",
  1429 => x"08881a08",
  1430 => x"718c120c",
  1431 => x"88120c57",
  1432 => x"57768107",
  1433 => x"84190c77",
  1434 => x"80c5800b",
  1435 => x"88050c80",
  1436 => x"c4fc0877",
  1437 => x"26fec738",
  1438 => x"80c4f808",
  1439 => x"527a51fa",
  1440 => x"fe3f7a51",
  1441 => x"fac43ffe",
  1442 => x"ba398178",
  1443 => x"8c150c78",
  1444 => x"88150c73",
  1445 => x"8c1a0c73",
  1446 => x"881a0c5a",
  1447 => x"fd803983",
  1448 => x"1570822c",
  1449 => x"81712b80",
  1450 => x"c5840807",
  1451 => x"80c5800b",
  1452 => x"84050c51",
  1453 => x"53741010",
  1454 => x"1080c580",
  1455 => x"05881108",
  1456 => x"5556fee4",
  1457 => x"39745380",
  1458 => x"7524a738",
  1459 => x"72822c81",
  1460 => x"712b80c5",
  1461 => x"84080780",
  1462 => x"c5800b84",
  1463 => x"050c5375",
  1464 => x"8c190c73",
  1465 => x"88190c77",
  1466 => x"88170c77",
  1467 => x"8c150cfd",
  1468 => x"cd398315",
  1469 => x"70822c81",
  1470 => x"712b80c5",
  1471 => x"84080780",
  1472 => x"c5800b84",
  1473 => x"050c5153",
  1474 => x"d639810b",
  1475 => x"800c0480",
  1476 => x"3d0d7281",
  1477 => x"2e893880",
  1478 => x"0b800c82",
  1479 => x"3d0d0473",
  1480 => x"5180f33f",
  1481 => x"fe3d0d80",
  1482 => x"cdc00851",
  1483 => x"708a3880",
  1484 => x"cdcc7080",
  1485 => x"cdc00c51",
  1486 => x"70751252",
  1487 => x"52ff5370",
  1488 => x"87fb8080",
  1489 => x"26883870",
  1490 => x"80cdc00c",
  1491 => x"71537280",
  1492 => x"0c843d0d",
  1493 => x"04fd3d0d",
  1494 => x"800bbd9c",
  1495 => x"08545472",
  1496 => x"812e9a38",
  1497 => x"7380cdc4",
  1498 => x"0cd9f43f",
  1499 => x"d9923f80",
  1500 => x"cd885281",
  1501 => x"51dbe23f",
  1502 => x"800851a0",
  1503 => x"3f7280cd",
  1504 => x"c40cd9db",
  1505 => x"3fd8f93f",
  1506 => x"80cd8852",
  1507 => x"8151dbc9",
  1508 => x"3f800851",
  1509 => x"873f00ff",
  1510 => x"3900ff39",
  1511 => x"f73d0d7b",
  1512 => x"bdc40882",
  1513 => x"c811085a",
  1514 => x"545a7780",
  1515 => x"2e80d938",
  1516 => x"81881884",
  1517 => x"1908ff05",
  1518 => x"81712b59",
  1519 => x"55598074",
  1520 => x"2480e938",
  1521 => x"807424b5",
  1522 => x"3873822b",
  1523 => x"78118805",
  1524 => x"56568180",
  1525 => x"19087706",
  1526 => x"5372802e",
  1527 => x"b5387816",
  1528 => x"70085353",
  1529 => x"79517408",
  1530 => x"53722dff",
  1531 => x"14fc17fc",
  1532 => x"1779812c",
  1533 => x"5a575754",
  1534 => x"738025d6",
  1535 => x"38770858",
  1536 => x"77ffad38",
  1537 => x"bdc40853",
  1538 => x"bc1308a5",
  1539 => x"387951ff",
  1540 => x"853f7408",
  1541 => x"53722dff",
  1542 => x"14fc17fc",
  1543 => x"1779812c",
  1544 => x"5a575754",
  1545 => x"738025ff",
  1546 => x"a938d239",
  1547 => x"8057ff94",
  1548 => x"397251bc",
  1549 => x"13085372",
  1550 => x"2d7951fe",
  1551 => x"d93fff3d",
  1552 => x"0d80cd90",
  1553 => x"0bfc0570",
  1554 => x"08525270",
  1555 => x"ff2e9138",
  1556 => x"702dfc12",
  1557 => x"70085252",
  1558 => x"70ff2e09",
  1559 => x"8106f138",
  1560 => x"833d0d04",
  1561 => x"04d8e33f",
  1562 => x"04000000",
  1563 => x"00000040",
  1564 => x"0a677265",
  1565 => x"74682072",
  1566 => x"65676973",
  1567 => x"74657273",
  1568 => x"3a000000",
  1569 => x"0a636f6e",
  1570 => x"74726f6c",
  1571 => x"3a202020",
  1572 => x"20202000",
  1573 => x"0a737461",
  1574 => x"7475733a",
  1575 => x"20202020",
  1576 => x"20202000",
  1577 => x"0a6d6163",
  1578 => x"5f6d7362",
  1579 => x"3a202020",
  1580 => x"20202000",
  1581 => x"0a6d6163",
  1582 => x"5f6c7362",
  1583 => x"3a202020",
  1584 => x"20202000",
  1585 => x"0a6d6469",
  1586 => x"6f5f636f",
  1587 => x"6e74726f",
  1588 => x"6c3a2000",
  1589 => x"0a74785f",
  1590 => x"706f696e",
  1591 => x"7465723a",
  1592 => x"20202000",
  1593 => x"0a72785f",
  1594 => x"706f696e",
  1595 => x"7465723a",
  1596 => x"20202000",
  1597 => x"0a656463",
  1598 => x"6c5f6970",
  1599 => x"3a202020",
  1600 => x"20202000",
  1601 => x"0a686173",
  1602 => x"685f6d73",
  1603 => x"623a2020",
  1604 => x"20202000",
  1605 => x"0a686173",
  1606 => x"685f6c73",
  1607 => x"623a2020",
  1608 => x"20202000",
  1609 => x"0a6d6469",
  1610 => x"6f207068",
  1611 => x"79207265",
  1612 => x"67697374",
  1613 => x"65727300",
  1614 => x"0a206d64",
  1615 => x"696f2070",
  1616 => x"68793a20",
  1617 => x"00000000",
  1618 => x"0a202072",
  1619 => x"65673a20",
  1620 => x"00000000",
  1621 => x"2d3e2000",
  1622 => x"0a677265",
  1623 => x"74682d3e",
  1624 => x"636f6e74",
  1625 => x"726f6c20",
  1626 => x"3a000000",
  1627 => x"0a677265",
  1628 => x"74682d3e",
  1629 => x"73746174",
  1630 => x"75732020",
  1631 => x"3a000000",
  1632 => x"0a646573",
  1633 => x"63722d3e",
  1634 => x"636f6e74",
  1635 => x"726f6c20",
  1636 => x"3a000000",
  1637 => x"77726974",
  1638 => x"65206164",
  1639 => x"64726573",
  1640 => x"733a2000",
  1641 => x"20206c65",
  1642 => x"6e677468",
  1643 => x"3a200000",
  1644 => x"0a0a0000",
  1645 => x"72656164",
  1646 => x"20206164",
  1647 => x"64726573",
  1648 => x"733a2000",
  1649 => x"20206578",
  1650 => x"70656374",
  1651 => x"3a200000",
  1652 => x"2020676f",
  1653 => x"743a2000",
  1654 => x"20657272",
  1655 => x"6f720000",
  1656 => x"206f6b00",
  1657 => x"70686173",
  1658 => x"65207368",
  1659 => x"69667420",
  1660 => x"202d2020",
  1661 => x"76616c75",
  1662 => x"653a2000",
  1663 => x"20207374",
  1664 => x"61747573",
  1665 => x"3a200000",
  1666 => x"20202020",
  1667 => x"20000000",
  1668 => x"6f6b2020",
  1669 => x"00000000",
  1670 => x"4641494c",
  1671 => x"00000000",
  1672 => x"44445220",
  1673 => x"6d656d6f",
  1674 => x"72792069",
  1675 => x"6e666f00",
  1676 => x"0a0a6175",
  1677 => x"746f2074",
  1678 => x"5f524552",
  1679 => x"45534820",
  1680 => x"3a000000",
  1681 => x"0a636c6f",
  1682 => x"636b2065",
  1683 => x"6e61626c",
  1684 => x"6520203a",
  1685 => x"00000000",
  1686 => x"0a696e69",
  1687 => x"74616c69",
  1688 => x"7a652020",
  1689 => x"2020203a",
  1690 => x"00000000",
  1691 => x"0a636f6c",
  1692 => x"756d6e20",
  1693 => x"73697a65",
  1694 => x"2020203a",
  1695 => x"00000000",
  1696 => x"0a62616e",
  1697 => x"6b73697a",
  1698 => x"65202020",
  1699 => x"2020203a",
  1700 => x"00000000",
  1701 => x"4d627974",
  1702 => x"65000000",
  1703 => x"0a745f52",
  1704 => x"43442020",
  1705 => x"20202020",
  1706 => x"2020203a",
  1707 => x"00000000",
  1708 => x"0a745f52",
  1709 => x"46432020",
  1710 => x"20202020",
  1711 => x"2020203a",
  1712 => x"00000000",
  1713 => x"0a745f52",
  1714 => x"50202020",
  1715 => x"20202020",
  1716 => x"2020203a",
  1717 => x"00000000",
  1718 => x"0a726566",
  1719 => x"72657368",
  1720 => x"20656e2e",
  1721 => x"2020203a",
  1722 => x"00000000",
  1723 => x"0a0a4444",
  1724 => x"52206672",
  1725 => x"65717565",
  1726 => x"6e637920",
  1727 => x"3a000000",
  1728 => x"0a444452",
  1729 => x"20646174",
  1730 => x"61207769",
  1731 => x"6474683a",
  1732 => x"00000000",
  1733 => x"0a6d6f62",
  1734 => x"696c6520",
  1735 => x"73757070",
  1736 => x"6f72743a",
  1737 => x"00000000",
  1738 => x"0a0a7374",
  1739 => x"61747573",
  1740 => x"20726561",
  1741 => x"64202020",
  1742 => x"3a000000",
  1743 => x"0a0a7365",
  1744 => x"6c662072",
  1745 => x"65667265",
  1746 => x"73682020",
  1747 => x"3a000000",
  1748 => x"20353132",
  1749 => x"00000000",
  1750 => x"34303639",
  1751 => x"00000000",
  1752 => x"312f3800",
  1753 => x"20617272",
  1754 => x"61790000",
  1755 => x"0a74656d",
  1756 => x"702d636f",
  1757 => x"6d702072",
  1758 => x"6566723a",
  1759 => x"00000000",
  1760 => x"c2b04300",
  1761 => x"0a647269",
  1762 => x"76652073",
  1763 => x"7472656e",
  1764 => x"6774683a",
  1765 => x"00000000",
  1766 => x"0a706f77",
  1767 => x"65722073",
  1768 => x"6176696e",
  1769 => x"6720203a",
  1770 => x"00000000",
  1771 => x"756e6b6e",
  1772 => x"6f776e00",
  1773 => x"0a745f58",
  1774 => x"50202020",
  1775 => x"20202020",
  1776 => x"2020203a",
  1777 => x"00000000",
  1778 => x"0a745f58",
  1779 => x"53522020",
  1780 => x"20202020",
  1781 => x"2020203a",
  1782 => x"00000000",
  1783 => x"0a745f43",
  1784 => x"4b452020",
  1785 => x"20202020",
  1786 => x"2020203a",
  1787 => x"00000000",
  1788 => x"0a434153",
  1789 => x"206c6174",
  1790 => x"656e6379",
  1791 => x"2020203a",
  1792 => x"00000000",
  1793 => x"0a6d6f62",
  1794 => x"696c6520",
  1795 => x"656e6162",
  1796 => x"6c65643a",
  1797 => x"00000000",
  1798 => x"0a0a7068",
  1799 => x"7920636f",
  1800 => x"6e666967",
  1801 => x"20302020",
  1802 => x"3a000000",
  1803 => x"0a0a7068",
  1804 => x"7920636f",
  1805 => x"6e666967",
  1806 => x"20312020",
  1807 => x"3a000000",
  1808 => x"31303234",
  1809 => x"00000000",
  1810 => x"32303438",
  1811 => x"00000000",
  1812 => x"66756c6c",
  1813 => x"00000000",
  1814 => x"37300000",
  1815 => x"64656570",
  1816 => x"20706f77",
  1817 => x"65722064",
  1818 => x"6f776e00",
  1819 => x"636c6f63",
  1820 => x"6b207374",
  1821 => x"6f700000",
  1822 => x"73656c66",
  1823 => x"20726566",
  1824 => x"72657368",
  1825 => x"00000000",
  1826 => x"706f7765",
  1827 => x"7220646f",
  1828 => x"776e0000",
  1829 => x"6e6f6e65",
  1830 => x"00000000",
  1831 => x"312f3200",
  1832 => x"312f3400",
  1833 => x"312f3100",
  1834 => x"332f3400",
  1835 => x"38350000",
  1836 => x"34350000",
  1837 => x"68616c66",
  1838 => x"00000000",
  1839 => x"31350000",
  1840 => x"61646472",
  1841 => x"6573733a",
  1842 => x"20000000",
  1843 => x"20646174",
  1844 => x"613a2000",
  1845 => x"0a0a4443",
  1846 => x"4d207068",
  1847 => x"61736520",
  1848 => x"73686966",
  1849 => x"74207465",
  1850 => x"7374696e",
  1851 => x"67000000",
  1852 => x"0a696e69",
  1853 => x"7469616c",
  1854 => x"3a200000",
  1855 => x"09000000",
  1856 => x"20202020",
  1857 => x"00000000",
  1858 => x"6c6f7720",
  1859 => x"666f756e",
  1860 => x"64000000",
  1861 => x"68696768",
  1862 => x"20666f75",
  1863 => x"6e640000",
  1864 => x"0a6c6f77",
  1865 => x"3a202020",
  1866 => x"20202020",
  1867 => x"20200000",
  1868 => x"0a686967",
  1869 => x"683a2020",
  1870 => x"20202020",
  1871 => x"20200000",
  1872 => x"0a646966",
  1873 => x"663a2020",
  1874 => x"20202020",
  1875 => x"20200000",
  1876 => x"0a6d696e",
  1877 => x"5f657272",
  1878 => x"3a202020",
  1879 => x"20200000",
  1880 => x"0a6d696e",
  1881 => x"5f657272",
  1882 => x"5f706f73",
  1883 => x"3a200000",
  1884 => x"676f206d",
  1885 => x"696e5f65",
  1886 => x"72726f72",
  1887 => x"00000000",
  1888 => x"0a66696e",
  1889 => x"616c3a20",
  1890 => x"20202020",
  1891 => x"20200000",
  1892 => x"6c6f7720",
  1893 => x"4e4f5420",
  1894 => x"666f756e",
  1895 => x"64000000",
  1896 => x"68696768",
  1897 => x"204e4f54",
  1898 => x"20666f75",
  1899 => x"6e640000",
  1900 => x"676f207a",
  1901 => x"65726f00",
  1902 => x"64617461",
  1903 => x"2076616c",
  1904 => x"69640000",
  1905 => x"6c6f7720",
  1906 => x"20666f75",
  1907 => x"6e640000",
  1908 => x"0a646966",
  1909 => x"662f323a",
  1910 => x"20202020",
  1911 => x"20200000",
  1912 => x"6c6f7720",
  1913 => x"204e4f54",
  1914 => x"20666f75",
  1915 => x"6e640000",
  1916 => x"64617461",
  1917 => x"204e4f54",
  1918 => x"2076616c",
  1919 => x"69640000",
  1920 => x"74657374",
  1921 => x"2e632000",
  1922 => x"286f6e20",
  1923 => x"73696d29",
  1924 => x"0a000000",
  1925 => x"636f6d70",
  1926 => x"696c6564",
  1927 => x"3a204e6f",
  1928 => x"76203138",
  1929 => x"20323031",
  1930 => x"30202031",
  1931 => x"373a3433",
  1932 => x"3a30380a",
  1933 => x"00000000",
  1934 => x"286f6e20",
  1935 => x"68617264",
  1936 => x"77617265",
  1937 => x"290a0000",
  1938 => x"30622020",
  1939 => x"20202020",
  1940 => x"20202020",
  1941 => x"20202020",
  1942 => x"20202020",
  1943 => x"20202020",
  1944 => x"20202020",
  1945 => x"20202020",
  1946 => x"20200000",
  1947 => x"30782020",
  1948 => x"20202020",
  1949 => x"20200000",
  1950 => x"43000000",
  1951 => x"64756d6d",
  1952 => x"792e6578",
  1953 => x"65000000",
  1954 => x"00ffffff",
  1955 => x"ff00ffff",
  1956 => x"ffff00ff",
  1957 => x"ffffff00",
  1958 => x"00000000",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00002698",
  1962 => x"fff00000",
  1963 => x"80000d00",
  1964 => x"80000c00",
  1965 => x"80000800",
  1966 => x"80000600",
  1967 => x"80000200",
  1968 => x"80000100",
  1969 => x"00001ec8",
  1970 => x"00000000",
  1971 => x"00002130",
  1972 => x"0000218c",
  1973 => x"000021e8",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00001e78",
  1984 => x"00000000",
  1985 => x"00000000",
  1986 => x"00000000",
  1987 => x"00000000",
  1988 => x"00000000",
  1989 => x"00000000",
  1990 => x"00000000",
  1991 => x"00000000",
  1992 => x"00000000",
  1993 => x"00000000",
  1994 => x"00000000",
  1995 => x"00000000",
  1996 => x"00000000",
  1997 => x"00000000",
  1998 => x"00000000",
  1999 => x"00000000",
  2000 => x"00000000",
  2001 => x"00000000",
  2002 => x"00000000",
  2003 => x"00000000",
  2004 => x"00000000",
  2005 => x"00000000",
  2006 => x"00000000",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00000000",
  2010 => x"00000000",
  2011 => x"00000000",
  2012 => x"00000001",
  2013 => x"330eabcd",
  2014 => x"1234e66d",
  2015 => x"deec0005",
  2016 => x"000b0000",
  2017 => x"00000000",
  2018 => x"00000000",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00000000",
  2026 => x"00000000",
  2027 => x"00000000",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000000",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"00000000",
  2049 => x"00000000",
  2050 => x"00000000",
  2051 => x"00000000",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"ffffffff",
  2206 => x"00000000",
  2207 => x"00020000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00002280",
  2211 => x"00002280",
  2212 => x"00002288",
  2213 => x"00002288",
  2214 => x"00002290",
  2215 => x"00002290",
  2216 => x"00002298",
  2217 => x"00002298",
  2218 => x"000022a0",
  2219 => x"000022a0",
  2220 => x"000022a8",
  2221 => x"000022a8",
  2222 => x"000022b0",
  2223 => x"000022b0",
  2224 => x"000022b8",
  2225 => x"000022b8",
  2226 => x"000022c0",
  2227 => x"000022c0",
  2228 => x"000022c8",
  2229 => x"000022c8",
  2230 => x"000022d0",
  2231 => x"000022d0",
  2232 => x"000022d8",
  2233 => x"000022d8",
  2234 => x"000022e0",
  2235 => x"000022e0",
  2236 => x"000022e8",
  2237 => x"000022e8",
  2238 => x"000022f0",
  2239 => x"000022f0",
  2240 => x"000022f8",
  2241 => x"000022f8",
  2242 => x"00002300",
  2243 => x"00002300",
  2244 => x"00002308",
  2245 => x"00002308",
  2246 => x"00002310",
  2247 => x"00002310",
  2248 => x"00002318",
  2249 => x"00002318",
  2250 => x"00002320",
  2251 => x"00002320",
  2252 => x"00002328",
  2253 => x"00002328",
  2254 => x"00002330",
  2255 => x"00002330",
  2256 => x"00002338",
  2257 => x"00002338",
  2258 => x"00002340",
  2259 => x"00002340",
  2260 => x"00002348",
  2261 => x"00002348",
  2262 => x"00002350",
  2263 => x"00002350",
  2264 => x"00002358",
  2265 => x"00002358",
  2266 => x"00002360",
  2267 => x"00002360",
  2268 => x"00002368",
  2269 => x"00002368",
  2270 => x"00002370",
  2271 => x"00002370",
  2272 => x"00002378",
  2273 => x"00002378",
  2274 => x"00002380",
  2275 => x"00002380",
  2276 => x"00002388",
  2277 => x"00002388",
  2278 => x"00002390",
  2279 => x"00002390",
  2280 => x"00002398",
  2281 => x"00002398",
  2282 => x"000023a0",
  2283 => x"000023a0",
  2284 => x"000023a8",
  2285 => x"000023a8",
  2286 => x"000023b0",
  2287 => x"000023b0",
  2288 => x"000023b8",
  2289 => x"000023b8",
  2290 => x"000023c0",
  2291 => x"000023c0",
  2292 => x"000023c8",
  2293 => x"000023c8",
  2294 => x"000023d0",
  2295 => x"000023d0",
  2296 => x"000023d8",
  2297 => x"000023d8",
  2298 => x"000023e0",
  2299 => x"000023e0",
  2300 => x"000023e8",
  2301 => x"000023e8",
  2302 => x"000023f0",
  2303 => x"000023f0",
  2304 => x"000023f8",
  2305 => x"000023f8",
  2306 => x"00002400",
  2307 => x"00002400",
  2308 => x"00002408",
  2309 => x"00002408",
  2310 => x"00002410",
  2311 => x"00002410",
  2312 => x"00002418",
  2313 => x"00002418",
  2314 => x"00002420",
  2315 => x"00002420",
  2316 => x"00002428",
  2317 => x"00002428",
  2318 => x"00002430",
  2319 => x"00002430",
  2320 => x"00002438",
  2321 => x"00002438",
  2322 => x"00002440",
  2323 => x"00002440",
  2324 => x"00002448",
  2325 => x"00002448",
  2326 => x"00002450",
  2327 => x"00002450",
  2328 => x"00002458",
  2329 => x"00002458",
  2330 => x"00002460",
  2331 => x"00002460",
  2332 => x"00002468",
  2333 => x"00002468",
  2334 => x"00002470",
  2335 => x"00002470",
  2336 => x"00002478",
  2337 => x"00002478",
  2338 => x"00002480",
  2339 => x"00002480",
  2340 => x"00002488",
  2341 => x"00002488",
  2342 => x"00002490",
  2343 => x"00002490",
  2344 => x"00002498",
  2345 => x"00002498",
  2346 => x"000024a0",
  2347 => x"000024a0",
  2348 => x"000024a8",
  2349 => x"000024a8",
  2350 => x"000024b0",
  2351 => x"000024b0",
  2352 => x"000024b8",
  2353 => x"000024b8",
  2354 => x"000024c0",
  2355 => x"000024c0",
  2356 => x"000024c8",
  2357 => x"000024c8",
  2358 => x"000024d0",
  2359 => x"000024d0",
  2360 => x"000024d8",
  2361 => x"000024d8",
  2362 => x"000024e0",
  2363 => x"000024e0",
  2364 => x"000024e8",
  2365 => x"000024e8",
  2366 => x"000024f0",
  2367 => x"000024f0",
  2368 => x"000024f8",
  2369 => x"000024f8",
  2370 => x"00002500",
  2371 => x"00002500",
  2372 => x"00002508",
  2373 => x"00002508",
  2374 => x"00002510",
  2375 => x"00002510",
  2376 => x"00002518",
  2377 => x"00002518",
  2378 => x"00002520",
  2379 => x"00002520",
  2380 => x"00002528",
  2381 => x"00002528",
  2382 => x"00002530",
  2383 => x"00002530",
  2384 => x"00002538",
  2385 => x"00002538",
  2386 => x"00002540",
  2387 => x"00002540",
  2388 => x"00002548",
  2389 => x"00002548",
  2390 => x"00002550",
  2391 => x"00002550",
  2392 => x"00002558",
  2393 => x"00002558",
  2394 => x"00002560",
  2395 => x"00002560",
  2396 => x"00002568",
  2397 => x"00002568",
  2398 => x"00002570",
  2399 => x"00002570",
  2400 => x"00002578",
  2401 => x"00002578",
  2402 => x"00002580",
  2403 => x"00002580",
  2404 => x"00002588",
  2405 => x"00002588",
  2406 => x"00002590",
  2407 => x"00002590",
  2408 => x"00002598",
  2409 => x"00002598",
  2410 => x"000025a0",
  2411 => x"000025a0",
  2412 => x"000025a8",
  2413 => x"000025a8",
  2414 => x"000025b0",
  2415 => x"000025b0",
  2416 => x"000025b8",
  2417 => x"000025b8",
  2418 => x"000025c0",
  2419 => x"000025c0",
  2420 => x"000025c8",
  2421 => x"000025c8",
  2422 => x"000025d0",
  2423 => x"000025d0",
  2424 => x"000025d8",
  2425 => x"000025d8",
  2426 => x"000025e0",
  2427 => x"000025e0",
  2428 => x"000025e8",
  2429 => x"000025e8",
  2430 => x"000025f0",
  2431 => x"000025f0",
  2432 => x"000025f8",
  2433 => x"000025f8",
  2434 => x"00002600",
  2435 => x"00002600",
  2436 => x"00002608",
  2437 => x"00002608",
  2438 => x"00002610",
  2439 => x"00002610",
  2440 => x"00002618",
  2441 => x"00002618",
  2442 => x"00002620",
  2443 => x"00002620",
  2444 => x"00002628",
  2445 => x"00002628",
  2446 => x"00002630",
  2447 => x"00002630",
  2448 => x"00002638",
  2449 => x"00002638",
  2450 => x"00002640",
  2451 => x"00002640",
  2452 => x"00002648",
  2453 => x"00002648",
  2454 => x"00002650",
  2455 => x"00002650",
  2456 => x"00002658",
  2457 => x"00002658",
  2458 => x"00002660",
  2459 => x"00002660",
  2460 => x"00002668",
  2461 => x"00002668",
  2462 => x"00002670",
  2463 => x"00002670",
  2464 => x"00002678",
  2465 => x"00002678",
  2466 => x"00001e7c",
  2467 => x"ffffffff",
  2468 => x"00000000",
  2469 => x"ffffffff",
  2470 => x"00000000",
  2471 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
