-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b8191",
     1 => x"ff040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b8194",
     9 => x"e7040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b8194",
    73 => x"99040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b8193fc",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b81f5",
   162 => x"e4738306",
   163 => x"10100508",
   164 => x"060b0b81",
   165 => x"93ff0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b8194",
   169 => x"ce040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b8194",
   177 => x"b5040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"81f5f40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053370",
   258 => x"52528191",
   259 => x"e43f7151",
   260 => x"8192d23f",
   261 => x"71b00c83",
   262 => x"3d0d04ff",
   263 => x"3d0d028f",
   264 => x"05337052",
   265 => x"528191c9",
   266 => x"3f715181",
   267 => x"92b73f71",
   268 => x"5180cac3",
   269 => x"3f71b00c",
   270 => x"833d0d04",
   271 => x"ff3d0d81",
   272 => x"f5cc08b8",
   273 => x"11085351",
   274 => x"800bb812",
   275 => x"0c71b00c",
   276 => x"833d0d04",
   277 => x"fa3d0d8a",
   278 => x"51818cb1",
   279 => x"3f96bc3f",
   280 => x"80e0eb53",
   281 => x"81c48c52",
   282 => x"81c4a051",
   283 => x"96c03f80",
   284 => x"f4af5381",
   285 => x"c4a45281",
   286 => x"c4b85196",
   287 => x"b13f80f4",
   288 => x"855381c4",
   289 => x"bc5281c4",
   290 => x"e45196a2",
   291 => x"3f80fcf0",
   292 => x"5381c4ec",
   293 => x"5281c4fc",
   294 => x"5196933f",
   295 => x"80fd8753",
   296 => x"81c58452",
   297 => x"81c5a051",
   298 => x"96843f80",
   299 => x"f6e15381",
   300 => x"c5a85281",
   301 => x"c5c05195",
   302 => x"f53f8180",
   303 => x"e85381c5",
   304 => x"c85281c5",
   305 => x"ec5195e6",
   306 => x"3f90b453",
   307 => x"81c5f452",
   308 => x"81c69051",
   309 => x"95d83f91",
   310 => x"cf5381c6",
   311 => x"945281c6",
   312 => x"b85195ca",
   313 => x"3f8fd253",
   314 => x"81c6c052",
   315 => x"81c6e451",
   316 => x"95bc3f81",
   317 => x"8fda5381",
   318 => x"c6ec5281",
   319 => x"c7945195",
   320 => x"ad3f8191",
   321 => x"875381c7",
   322 => x"9c5281c7",
   323 => x"bc51959e",
   324 => x"3f88bc53",
   325 => x"81c7c452",
   326 => x"81c7e451",
   327 => x"95903f80",
   328 => x"f78c5381",
   329 => x"c7ec5281",
   330 => x"c8805195",
   331 => x"813f80fd",
   332 => x"a25381c8",
   333 => x"885281c7",
   334 => x"b45194f2",
   335 => x"3f8180b4",
   336 => x"5381c8a4",
   337 => x"5281c8b8",
   338 => x"5194e33f",
   339 => x"80feb253",
   340 => x"81c8c052",
   341 => x"81c8e051",
   342 => x"94d43f80",
   343 => x"ff945381",
   344 => x"c8e85281",
   345 => x"c9885194",
   346 => x"c53f818f",
   347 => x"b25381c9",
   348 => x"905281c9",
   349 => x"ac5194b6",
   350 => x"3f818694",
   351 => x"5381c9b4",
   352 => x"5281c9c8",
   353 => x"5194a73f",
   354 => x"81828153",
   355 => x"81c9d052",
   356 => x"81c9f451",
   357 => x"94983f96",
   358 => x"8c5381c9",
   359 => x"fc5281ca",
   360 => x"8c51948a",
   361 => x"3f93bc53",
   362 => x"81ca9052",
   363 => x"81caac51",
   364 => x"93fc3f8f",
   365 => x"b65381ca",
   366 => x"b45281ca",
   367 => x"cc5193ee",
   368 => x"3f93c453",
   369 => x"81cad452",
   370 => x"81cae851",
   371 => x"93e03f80",
   372 => x"d3975381",
   373 => x"caf05281",
   374 => x"cb845193",
   375 => x"d13f80d7",
   376 => x"965381cb",
   377 => x"885281cb",
   378 => x"b05193c2",
   379 => x"3f80fabc",
   380 => x"5381cbb8",
   381 => x"5281cbd8",
   382 => x"5193b33f",
   383 => x"80f9e053",
   384 => x"81cbe052",
   385 => x"81cbf451",
   386 => x"93a43f80",
   387 => x"d9835381",
   388 => x"cbfc5281",
   389 => x"cc945193",
   390 => x"953fbbc5",
   391 => x"5381cc9c",
   392 => x"5281ccb4",
   393 => x"5193873f",
   394 => x"80d9e753",
   395 => x"81ccbc52",
   396 => x"81cce451",
   397 => x"92f83f80",
   398 => x"fae65381",
   399 => x"ccec5281",
   400 => x"ccf85192",
   401 => x"e93f80fc",
   402 => x"975381cc",
   403 => x"fc5281cd",
   404 => x"a45192da",
   405 => x"3f80fae6",
   406 => x"5381cdac",
   407 => x"5281f0d8",
   408 => x"5192cb3f",
   409 => x"80fce053",
   410 => x"81cdcc52",
   411 => x"81cddc51",
   412 => x"92bc3f80",
   413 => x"fadb5381",
   414 => x"defc5281",
   415 => x"c3fc5192",
   416 => x"ad3fa6ad",
   417 => x"5381defc",
   418 => x"5281c484",
   419 => x"51929f3f",
   420 => x"999b3f92",
   421 => x"f93f810b",
   422 => x"829dd834",
   423 => x"8285e833",
   424 => x"7081ff06",
   425 => x"555573b2",
   426 => x"38818bed",
   427 => x"3fb00890",
   428 => x"3892ea3f",
   429 => x"829dd833",
   430 => x"5675e138",
   431 => x"883d0d04",
   432 => x"818be93f",
   433 => x"b00881ff",
   434 => x"065193c8",
   435 => x"3f92ce3f",
   436 => x"829dd833",
   437 => x"5675c538",
   438 => x"e339800b",
   439 => x"8285e834",
   440 => x"99f43f81",
   441 => x"f68c0870",
   442 => x"0870872a",
   443 => x"81065257",
   444 => x"5473802e",
   445 => x"8f387680",
   446 => x"2e819738",
   447 => x"ff177081",
   448 => x"ff065854",
   449 => x"75862a81",
   450 => x"06557480",
   451 => x"2e8f3876",
   452 => x"802e8190",
   453 => x"38ff1770",
   454 => x"81ff0658",
   455 => x"5575852a",
   456 => x"81065473",
   457 => x"802e9638",
   458 => x"76ba3881",
   459 => x"960b81f5",
   460 => x"cc08b811",
   461 => x"08575557",
   462 => x"800bb815",
   463 => x"0c75842a",
   464 => x"81065675",
   465 => x"802efee1",
   466 => x"3876802e",
   467 => x"a138ff17",
   468 => x"7081ff06",
   469 => x"5855818a",
   470 => x"c03fb008",
   471 => x"802efed1",
   472 => x"38fedd39",
   473 => x"ff177081",
   474 => x"ff065855",
   475 => x"d0398196",
   476 => x"0b81f68c",
   477 => x"08841108",
   478 => x"840a0784",
   479 => x"120c5657",
   480 => x"80e4da3f",
   481 => x"818a923f",
   482 => x"b008802e",
   483 => x"fea338fe",
   484 => x"af398196",
   485 => x"76822a83",
   486 => x"06535780",
   487 => x"5180fadb",
   488 => x"3ffee139",
   489 => x"81965780",
   490 => x"5181829f",
   491 => x"3f815181",
   492 => x"82993ffe",
   493 => x"e839fe3d",
   494 => x"0d815194",
   495 => x"8a3fb008",
   496 => x"81ff0681",
   497 => x"f5c00871",
   498 => x"88120c53",
   499 => x"b00c843d",
   500 => x"0d04fc3d",
   501 => x"0d815193",
   502 => x"ee3fb008",
   503 => x"81ff0654",
   504 => x"825193e3",
   505 => x"3fb00881",
   506 => x"ff0681f6",
   507 => x"8c088411",
   508 => x"0870fe8f",
   509 => x"0a067798",
   510 => x"2b075154",
   511 => x"56537280",
   512 => x"2e863871",
   513 => x"810a0752",
   514 => x"7184160c",
   515 => x"71b00c86",
   516 => x"3d0d04ff",
   517 => x"3d0d81f6",
   518 => x"8c087008",
   519 => x"709e2a70",
   520 => x"81065152",
   521 => x"53518152",
   522 => x"70833870",
   523 => x"5271b00c",
   524 => x"833d0d04",
   525 => x"fc3d0d81",
   526 => x"51938c3f",
   527 => x"b00881ff",
   528 => x"0681cde4",
   529 => x"52558184",
   530 => x"de3f81f6",
   531 => x"8c087008",
   532 => x"709e2a70",
   533 => x"81065154",
   534 => x"54548153",
   535 => x"71833871",
   536 => x"5372802e",
   537 => x"80cb3881",
   538 => x"cdf45181",
   539 => x"84b93f81",
   540 => x"cde45181",
   541 => x"84b13f74",
   542 => x"802eac38",
   543 => x"81cdfc51",
   544 => x"8184a43f",
   545 => x"81f68c08",
   546 => x"84110870",
   547 => x"fd0a0655",
   548 => x"53547480",
   549 => x"2e863871",
   550 => x"820a0753",
   551 => x"7284150c",
   552 => x"71b00c86",
   553 => x"3d0d0481",
   554 => x"ce885181",
   555 => x"83f93fcc",
   556 => x"3981ce88",
   557 => x"518183ef",
   558 => x"3f81cdf4",
   559 => x"518183e7",
   560 => x"3f81cde4",
   561 => x"518183df",
   562 => x"3f74ffb0",
   563 => x"38d939fd",
   564 => x"3d0d8151",
   565 => x"91f13fb0",
   566 => x"0881ff06",
   567 => x"81ce9052",
   568 => x"548183c3",
   569 => x"3f73a638",
   570 => x"81c6e451",
   571 => x"8183b83f",
   572 => x"81f68c08",
   573 => x"84110870",
   574 => x"fb0a0684",
   575 => x"130c5353",
   576 => x"8a518183",
   577 => x"883f73b0",
   578 => x"0c853d0d",
   579 => x"0481cea4",
   580 => x"51818393",
   581 => x"3f81f68c",
   582 => x"08841108",
   583 => x"70840a07",
   584 => x"84130c53",
   585 => x"538a5181",
   586 => x"82e33f73",
   587 => x"b00c853d",
   588 => x"0d04f73d",
   589 => x"0d853d54",
   590 => x"965381ce",
   591 => x"b0527351",
   592 => x"8189fc3f",
   593 => x"ad8b3f81",
   594 => x"5190fc3f",
   595 => x"80528051",
   596 => x"aaeb3f73",
   597 => x"53805281",
   598 => x"d68451bf",
   599 => x"aa3f8052",
   600 => x"8151aad9",
   601 => x"3f735382",
   602 => x"5281d684",
   603 => x"51bf983f",
   604 => x"80528251",
   605 => x"aac73f73",
   606 => x"53815281",
   607 => x"d68451bf",
   608 => x"863f8052",
   609 => x"8451aab5",
   610 => x"3f735384",
   611 => x"5281d684",
   612 => x"51bef43f",
   613 => x"80528551",
   614 => x"aaa33f73",
   615 => x"53905281",
   616 => x"d68451be",
   617 => x"e23f8052",
   618 => x"8651aa91",
   619 => x"3f735383",
   620 => x"5281d684",
   621 => x"51bed03f",
   622 => x"8b3d0d04",
   623 => x"fef43f80",
   624 => x"0bb00c04",
   625 => x"fc3d0dab",
   626 => x"973f81be",
   627 => x"94548055",
   628 => x"84527451",
   629 => x"a9e73f80",
   630 => x"53737081",
   631 => x"05553351",
   632 => x"aae13f81",
   633 => x"137081ff",
   634 => x"06515380",
   635 => x"dc7327e9",
   636 => x"38811570",
   637 => x"81ff0656",
   638 => x"53877527",
   639 => x"d338800b",
   640 => x"b00c863d",
   641 => x"0d04fd3d",
   642 => x"0d81f5dc",
   643 => x"337081ff",
   644 => x"06545472",
   645 => x"bf26ab38",
   646 => x"81f5dc33",
   647 => x"7081ff06",
   648 => x"81f5c008",
   649 => x"5288120c",
   650 => x"5480e452",
   651 => x"94865194",
   652 => x"853f81f5",
   653 => x"dc338105",
   654 => x"537281f5",
   655 => x"dc34853d",
   656 => x"0d0480e4",
   657 => x"5294db51",
   658 => x"93ec3f81",
   659 => x"f5dc3381",
   660 => x"05537281",
   661 => x"f5dc3485",
   662 => x"3d0d04fd",
   663 => x"3d0d81f5",
   664 => x"dc337081",
   665 => x"ff065454",
   666 => x"72bf2680",
   667 => x"c83881f5",
   668 => x"dc337081",
   669 => x"ff0681f5",
   670 => x"c0085688",
   671 => x"160c5381",
   672 => x"f5dc3370",
   673 => x"81ff0655",
   674 => x"5373bf2e",
   675 => x"80d03880",
   676 => x"e45294db",
   677 => x"51939f3f",
   678 => x"81f5dc33",
   679 => x"81055372",
   680 => x"81f5dc34",
   681 => x"81f5dc33",
   682 => x"80ff0653",
   683 => x"7281f5dc",
   684 => x"34853d0d",
   685 => x"0481f5dc",
   686 => x"337081ff",
   687 => x"0680ff71",
   688 => x"3181f5c0",
   689 => x"08528812",
   690 => x"0c555381",
   691 => x"f5dc3370",
   692 => x"81ff0655",
   693 => x"5373bf2e",
   694 => x"098106ff",
   695 => x"b23880ce",
   696 => x"905294db",
   697 => x"5192cf3f",
   698 => x"81f5dc33",
   699 => x"81055372",
   700 => x"81f5dc34",
   701 => x"81f5dc33",
   702 => x"80ff0653",
   703 => x"7281f5dc",
   704 => x"34853d0d",
   705 => x"04810b81",
   706 => x"f5c43404",
   707 => x"fd3d0d82",
   708 => x"85e40852",
   709 => x"f881c08e",
   710 => x"800b81f6",
   711 => x"8c085553",
   712 => x"71802e80",
   713 => x"f8387281",
   714 => x"ff068415",
   715 => x"0c81f5dc",
   716 => x"337081ff",
   717 => x"06515271",
   718 => x"802e80c2",
   719 => x"38729f2a",
   720 => x"73100753",
   721 => x"8285e833",
   722 => x"7081ff06",
   723 => x"51527180",
   724 => x"2ed43880",
   725 => x"0b8285e8",
   726 => x"3490fb3f",
   727 => x"81f5c433",
   728 => x"547380e4",
   729 => x"3881f68c",
   730 => x"087381ff",
   731 => x"0684120c",
   732 => x"81f5dc33",
   733 => x"7081ff06",
   734 => x"51535471",
   735 => x"c0387281",
   736 => x"2a739f2b",
   737 => x"0753ffbc",
   738 => x"3972812a",
   739 => x"739f2b07",
   740 => x"5380fd51",
   741 => x"8181a33f",
   742 => x"81f68c08",
   743 => x"547281ff",
   744 => x"0684150c",
   745 => x"81f5dc33",
   746 => x"7081ff06",
   747 => x"53547180",
   748 => x"2ed73872",
   749 => x"9f2a7310",
   750 => x"075380fd",
   751 => x"518180fa",
   752 => x"3f81f68c",
   753 => x"0854d639",
   754 => x"800bb00c",
   755 => x"853d0d04",
   756 => x"fe3d0d81",
   757 => x"f6900898",
   758 => x"11087084",
   759 => x"2a708106",
   760 => x"51535353",
   761 => x"70802e8d",
   762 => x"3871ef06",
   763 => x"98140c81",
   764 => x"0b8285e8",
   765 => x"34843d0d",
   766 => x"04fb3d0d",
   767 => x"81f68c08",
   768 => x"7008810a",
   769 => x"068285e4",
   770 => x"0c548180",
   771 => x"d03f8180",
   772 => x"f23f91df",
   773 => x"3f81f690",
   774 => x"08981108",
   775 => x"88079812",
   776 => x"0c548285",
   777 => x"e4085372",
   778 => x"802e85a9",
   779 => x"388194f7",
   780 => x"0b829ebc",
   781 => x"0c81cec8",
   782 => x"5180fceb",
   783 => x"3f8c5180",
   784 => x"fccb3f81",
   785 => x"ceb05180",
   786 => x"fcdd3f82",
   787 => x"85e40880",
   788 => x"2e81ee38",
   789 => x"81cecc51",
   790 => x"80fccc3f",
   791 => x"8285e408",
   792 => x"5473802e",
   793 => x"82f33881",
   794 => x"f5e00854",
   795 => x"81740c81",
   796 => x"f68c0884",
   797 => x"11087056",
   798 => x"57558053",
   799 => x"73fe8f0a",
   800 => x"0673982b",
   801 => x"07708417",
   802 => x"0c811470",
   803 => x"81ff0651",
   804 => x"54548f73",
   805 => x"27e63875",
   806 => x"84160c81",
   807 => x"f5cc0853",
   808 => x"800bb814",
   809 => x"0c81f5fc",
   810 => x"087008fe",
   811 => x"8006710c",
   812 => x"54a0808d",
   813 => x"0a085180",
   814 => x"fdb73f8a",
   815 => x"5180fbcd",
   816 => x"3f825296",
   817 => x"85518eee",
   818 => x"3ff881c0",
   819 => x"8e800b81",
   820 => x"f68c0856",
   821 => x"548285e4",
   822 => x"08802e81",
   823 => x"d1387381",
   824 => x"ff068416",
   825 => x"0c81f5dc",
   826 => x"337081ff",
   827 => x"06545672",
   828 => x"802e80c2",
   829 => x"38739f2a",
   830 => x"74100754",
   831 => x"8285e833",
   832 => x"7081ff06",
   833 => x"57537580",
   834 => x"2ed43880",
   835 => x"0b8285e8",
   836 => x"348dc33f",
   837 => x"81f5c433",
   838 => x"557484fb",
   839 => x"3881f68c",
   840 => x"087481ff",
   841 => x"0684120c",
   842 => x"81f5dc33",
   843 => x"7081ff06",
   844 => x"55575572",
   845 => x"c0387381",
   846 => x"2a749f2b",
   847 => x"0754ffbc",
   848 => x"3981ced8",
   849 => x"5180fadf",
   850 => x"3f810a51",
   851 => x"80fad83f",
   852 => x"81ceec51",
   853 => x"80fad03f",
   854 => x"81cf9451",
   855 => x"80fac83f",
   856 => x"b45180fc",
   857 => x"8c3f81cf",
   858 => x"a85180fa",
   859 => x"ba3f81cf",
   860 => x"b05180fa",
   861 => x"b23f81cf",
   862 => x"bc5180fa",
   863 => x"aa3f81cf",
   864 => x"c45180fa",
   865 => x"a23f81cf",
   866 => x"e05180fa",
   867 => x"9a3f8285",
   868 => x"e4085473",
   869 => x"fdd13880",
   870 => x"c0397381",
   871 => x"2a749f2b",
   872 => x"075480fd",
   873 => x"5180fd92",
   874 => x"3f81f68c",
   875 => x"08557381",
   876 => x"ff068416",
   877 => x"0c81f5dc",
   878 => x"337081ff",
   879 => x"06565674",
   880 => x"802ed738",
   881 => x"739f2a74",
   882 => x"10075480",
   883 => x"fd5180fc",
   884 => x"e93f81f6",
   885 => x"8c0855d6",
   886 => x"39889b0b",
   887 => x"829ebc0c",
   888 => x"81cfe851",
   889 => x"80f9c03f",
   890 => x"810a5180",
   891 => x"f9b93f81",
   892 => x"d0805180",
   893 => x"f9b13f81",
   894 => x"f5cc0874",
   895 => x"b4120c74",
   896 => x"b8120c55",
   897 => x"81d09851",
   898 => x"80f99c3f",
   899 => x"735180dd",
   900 => x"823fb008",
   901 => x"982b5372",
   902 => x"82c83881",
   903 => x"d0a45180",
   904 => x"f9853f81",
   905 => x"f68c0870",
   906 => x"08709e2a",
   907 => x"81065557",
   908 => x"54815572",
   909 => x"802e81ba",
   910 => x"387481ff",
   911 => x"06841508",
   912 => x"70fd0a06",
   913 => x"58565372",
   914 => x"802e8638",
   915 => x"74820a07",
   916 => x"56758415",
   917 => x"0c730870",
   918 => x"9e2a8106",
   919 => x"54558154",
   920 => x"72833872",
   921 => x"5473802e",
   922 => x"818d3881",
   923 => x"d0b05180",
   924 => x"f8b53f81",
   925 => x"5180f4d3",
   926 => x"3f81f68c",
   927 => x"08841108",
   928 => x"840a0784",
   929 => x"120c5581",
   930 => x"d0bc5180",
   931 => x"f8993f81",
   932 => x"f5cc0854",
   933 => x"800bb815",
   934 => x"0c81f5e0",
   935 => x"08568176",
   936 => x"0c88800b",
   937 => x"829ebc0c",
   938 => x"a7885293",
   939 => x"c4518b86",
   940 => x"3f87e852",
   941 => x"9486518a",
   942 => x"fd3feb98",
   943 => x"3f81f5e0",
   944 => x"08548174",
   945 => x"0c81f68c",
   946 => x"08841108",
   947 => x"70565755",
   948 => x"8053fba8",
   949 => x"3980fce9",
   950 => x"3f9dea3f",
   951 => x"a1f33f72",
   952 => x"5281d684",
   953 => x"51a3cc3f",
   954 => x"88800b82",
   955 => x"9ebc0cfa",
   956 => x"c4397255",
   957 => x"fec33981",
   958 => x"d0c85180",
   959 => x"f7a93f81",
   960 => x"f5cc08b8",
   961 => x"1108810a",
   962 => x"07b8120c",
   963 => x"5481d0b0",
   964 => x"5180f793",
   965 => x"3f815180",
   966 => x"f3b13f81",
   967 => x"f68c0884",
   968 => x"1108840a",
   969 => x"0784120c",
   970 => x"5581d0bc",
   971 => x"5180f6f7",
   972 => x"3f81f5cc",
   973 => x"0854800b",
   974 => x"b8150c81",
   975 => x"f5e00856",
   976 => x"81760c88",
   977 => x"800b829e",
   978 => x"bc0ca788",
   979 => x"5293c451",
   980 => x"89e43f87",
   981 => x"e8529486",
   982 => x"5189db3f",
   983 => x"e9f63ffe",
   984 => x"dc3981d0",
   985 => x"c85180f6",
   986 => x"be3f81f5",
   987 => x"cc08b811",
   988 => x"08810a07",
   989 => x"b8120c56",
   990 => x"81d0a451",
   991 => x"80f6a83f",
   992 => x"81f68c08",
   993 => x"7008709e",
   994 => x"2a810655",
   995 => x"57548155",
   996 => x"72fda638",
   997 => x"fedc3980",
   998 => x"fd983f80",
   999 => x"0b829dd0",
  1000 => x"34800b82",
  1001 => x"9dcc3480",
  1002 => x"0b829dd4",
  1003 => x"0c04fc3d",
  1004 => x"0d829dcc",
  1005 => x"335372a7",
  1006 => x"2680c738",
  1007 => x"76527210",
  1008 => x"10107310",
  1009 => x"058285ec",
  1010 => x"05518182",
  1011 => x"803f7752",
  1012 => x"829dcc33",
  1013 => x"70902971",
  1014 => x"31701010",
  1015 => x"8288fc05",
  1016 => x"53565481",
  1017 => x"81e73f82",
  1018 => x"9dcc3370",
  1019 => x"1010829b",
  1020 => x"dc057a71",
  1021 => x"0c548105",
  1022 => x"5372829d",
  1023 => x"cc34863d",
  1024 => x"0d0481d0",
  1025 => x"d45180f5",
  1026 => x"9e3f863d",
  1027 => x"0d04803d",
  1028 => x"0d81d0f0",
  1029 => x"5180f58f",
  1030 => x"3f823d0d",
  1031 => x"04fe3d0d",
  1032 => x"829dd408",
  1033 => x"53728538",
  1034 => x"843d0d04",
  1035 => x"722db008",
  1036 => x"53800b82",
  1037 => x"9dd40cb0",
  1038 => x"088d3881",
  1039 => x"d0f05180",
  1040 => x"f4e53f84",
  1041 => x"3d0d0481",
  1042 => x"d5ac5180",
  1043 => x"f4d93f72",
  1044 => x"83ffff26",
  1045 => x"af3881ff",
  1046 => x"73279938",
  1047 => x"72529051",
  1048 => x"80f4e73f",
  1049 => x"8a5180f4",
  1050 => x"a43f81d0",
  1051 => x"f05180f4",
  1052 => x"b63fd039",
  1053 => x"72528851",
  1054 => x"80f4cf3f",
  1055 => x"8a5180f4",
  1056 => x"8c3fe739",
  1057 => x"7252a051",
  1058 => x"80f4bf3f",
  1059 => x"8a5180f3",
  1060 => x"fc3fd739",
  1061 => x"fa3d0d02",
  1062 => x"a3053356",
  1063 => x"758d2e80",
  1064 => x"f8387588",
  1065 => x"32703077",
  1066 => x"80ff3270",
  1067 => x"30728025",
  1068 => x"71802507",
  1069 => x"54515658",
  1070 => x"55749538",
  1071 => x"9f76278c",
  1072 => x"38829dd0",
  1073 => x"335580ce",
  1074 => x"7527b138",
  1075 => x"883d0d04",
  1076 => x"829dd033",
  1077 => x"5675802e",
  1078 => x"f3388851",
  1079 => x"80f3ae3f",
  1080 => x"a05180f3",
  1081 => x"a83f8851",
  1082 => x"80f3a23f",
  1083 => x"829dd033",
  1084 => x"ff055776",
  1085 => x"829dd034",
  1086 => x"883d0d04",
  1087 => x"755180f3",
  1088 => x"8c3f829d",
  1089 => x"d0338111",
  1090 => x"55577382",
  1091 => x"9dd03475",
  1092 => x"829cfc18",
  1093 => x"34883d0d",
  1094 => x"048a5180",
  1095 => x"f2ef3f82",
  1096 => x"9dd03381",
  1097 => x"11565474",
  1098 => x"829dd034",
  1099 => x"800b829c",
  1100 => x"fc153480",
  1101 => x"56800b82",
  1102 => x"9cfc1733",
  1103 => x"565474a0",
  1104 => x"2e833881",
  1105 => x"5474802e",
  1106 => x"90387380",
  1107 => x"2e8b3881",
  1108 => x"167081ff",
  1109 => x"065757dd",
  1110 => x"3975802e",
  1111 => x"80c13880",
  1112 => x"0b829dcc",
  1113 => x"33555574",
  1114 => x"7427ac38",
  1115 => x"73577410",
  1116 => x"10107510",
  1117 => x"05765482",
  1118 => x"9cfc5382",
  1119 => x"85ec0551",
  1120 => x"8180963f",
  1121 => x"b008802e",
  1122 => x"a8388115",
  1123 => x"7081ff06",
  1124 => x"56547675",
  1125 => x"26d83881",
  1126 => x"d0f45180",
  1127 => x"f2893f81",
  1128 => x"d0f05180",
  1129 => x"f2813f80",
  1130 => x"0b829dd0",
  1131 => x"34883d0d",
  1132 => x"04741010",
  1133 => x"829bdc05",
  1134 => x"7008829d",
  1135 => x"d40c5680",
  1136 => x"0b829dd0",
  1137 => x"34e739f7",
  1138 => x"3d0d02af",
  1139 => x"05335980",
  1140 => x"0b829cfc",
  1141 => x"33829cfc",
  1142 => x"59555673",
  1143 => x"a02e0981",
  1144 => x"06963881",
  1145 => x"167081ff",
  1146 => x"06829cfc",
  1147 => x"11703353",
  1148 => x"59575473",
  1149 => x"a02eec38",
  1150 => x"80587779",
  1151 => x"2780ea38",
  1152 => x"80773356",
  1153 => x"5474742e",
  1154 => x"83388154",
  1155 => x"74a02e9a",
  1156 => x"387380c5",
  1157 => x"3874a02e",
  1158 => x"91388118",
  1159 => x"7081ff06",
  1160 => x"59557878",
  1161 => x"26da3880",
  1162 => x"c0398116",
  1163 => x"7081ff06",
  1164 => x"829cfc11",
  1165 => x"70335752",
  1166 => x"575773a0",
  1167 => x"2e098106",
  1168 => x"d9388116",
  1169 => x"7081ff06",
  1170 => x"829cfc11",
  1171 => x"70335752",
  1172 => x"575773a0",
  1173 => x"2ed438c2",
  1174 => x"39811670",
  1175 => x"81ff0682",
  1176 => x"9cfc1159",
  1177 => x"5755ff98",
  1178 => x"3980538b",
  1179 => x"3dfc0552",
  1180 => x"76518182",
  1181 => x"e93f8b3d",
  1182 => x"0d04f73d",
  1183 => x"0d02af05",
  1184 => x"3359800b",
  1185 => x"829cfc33",
  1186 => x"829cfc59",
  1187 => x"555673a0",
  1188 => x"2e098106",
  1189 => x"96388116",
  1190 => x"7081ff06",
  1191 => x"829cfc11",
  1192 => x"70335359",
  1193 => x"575473a0",
  1194 => x"2eec3880",
  1195 => x"58777927",
  1196 => x"80ea3880",
  1197 => x"77335654",
  1198 => x"74742e83",
  1199 => x"38815474",
  1200 => x"a02e9a38",
  1201 => x"7380c538",
  1202 => x"74a02e91",
  1203 => x"38811870",
  1204 => x"81ff0659",
  1205 => x"55787826",
  1206 => x"da3880c0",
  1207 => x"39811670",
  1208 => x"81ff0682",
  1209 => x"9cfc1170",
  1210 => x"33575257",
  1211 => x"5773a02e",
  1212 => x"098106d9",
  1213 => x"38811670",
  1214 => x"81ff0682",
  1215 => x"9cfc1170",
  1216 => x"33575257",
  1217 => x"5773a02e",
  1218 => x"d438c239",
  1219 => x"81167081",
  1220 => x"ff06829c",
  1221 => x"fc115957",
  1222 => x"55ff9839",
  1223 => x"90538b3d",
  1224 => x"fc055276",
  1225 => x"518184d3",
  1226 => x"3f8b3d0d",
  1227 => x"04fc3d0d",
  1228 => x"8a5180ee",
  1229 => x"d83f81d1",
  1230 => x"885180ee",
  1231 => x"ea3f800b",
  1232 => x"829dcc33",
  1233 => x"53537272",
  1234 => x"2780fb38",
  1235 => x"72101010",
  1236 => x"73100582",
  1237 => x"85ec0570",
  1238 => x"525480ee",
  1239 => x"ca3f7284",
  1240 => x"2b707431",
  1241 => x"822b8288",
  1242 => x"fc113351",
  1243 => x"53557180",
  1244 => x"2ebb3873",
  1245 => x"5180fbc2",
  1246 => x"3fb00881",
  1247 => x"ff065271",
  1248 => x"89269438",
  1249 => x"a05180ee",
  1250 => x"843f8112",
  1251 => x"7081ff06",
  1252 => x"53548972",
  1253 => x"27ee3881",
  1254 => x"d1a05180",
  1255 => x"ee893f74",
  1256 => x"7331822b",
  1257 => x"8288fc05",
  1258 => x"5180edfb",
  1259 => x"3f8a5180",
  1260 => x"eddb3f81",
  1261 => x"137081ff",
  1262 => x"06829dcc",
  1263 => x"33545455",
  1264 => x"717326ff",
  1265 => x"87388a51",
  1266 => x"80edc23f",
  1267 => x"829dcc33",
  1268 => x"b00c863d",
  1269 => x"0d04fe3d",
  1270 => x"0d829eac",
  1271 => x"22ff0551",
  1272 => x"70829eac",
  1273 => x"237083ff",
  1274 => x"ff065170",
  1275 => x"80c43882",
  1276 => x"9eb03351",
  1277 => x"7081ff2e",
  1278 => x"b9387010",
  1279 => x"1010829d",
  1280 => x"dc055271",
  1281 => x"33829eb0",
  1282 => x"34fe7234",
  1283 => x"829eb033",
  1284 => x"70101010",
  1285 => x"829ddc05",
  1286 => x"52538211",
  1287 => x"22829eac",
  1288 => x"23841208",
  1289 => x"53722d82",
  1290 => x"9eac2251",
  1291 => x"70802eff",
  1292 => x"be38843d",
  1293 => x"0d04f93d",
  1294 => x"0d02aa05",
  1295 => x"22568055",
  1296 => x"74101010",
  1297 => x"829ddc05",
  1298 => x"70335252",
  1299 => x"7081fe2e",
  1300 => x"99388115",
  1301 => x"7081ff06",
  1302 => x"5652748a",
  1303 => x"2e098106",
  1304 => x"df38810b",
  1305 => x"b00c893d",
  1306 => x"0d04829e",
  1307 => x"b0337081",
  1308 => x"ff06829e",
  1309 => x"ac225354",
  1310 => x"587281ff",
  1311 => x"2eb03872",
  1312 => x"832b5470",
  1313 => x"762780de",
  1314 => x"38757131",
  1315 => x"7083ffff",
  1316 => x"0674829d",
  1317 => x"dc173370",
  1318 => x"832b829d",
  1319 => x"de112256",
  1320 => x"58565257",
  1321 => x"577281ff",
  1322 => x"2e098106",
  1323 => x"d6387272",
  1324 => x"34758213",
  1325 => x"23798413",
  1326 => x"0c7781ff",
  1327 => x"06547373",
  1328 => x"2e963876",
  1329 => x"10101082",
  1330 => x"9ddc0553",
  1331 => x"74733480",
  1332 => x"5170b00c",
  1333 => x"893d0d04",
  1334 => x"74829eb0",
  1335 => x"3475829e",
  1336 => x"ac238051",
  1337 => x"ec397076",
  1338 => x"31517082",
  1339 => x"9dde1523",
  1340 => x"ffbc39ff",
  1341 => x"3d0d8a52",
  1342 => x"71101010",
  1343 => x"829dd405",
  1344 => x"51fe7134",
  1345 => x"ff127081",
  1346 => x"ff065351",
  1347 => x"71ea38ff",
  1348 => x"0b829eb0",
  1349 => x"34833d0d",
  1350 => x"04f53d0d",
  1351 => x"7d598a54",
  1352 => x"81028405",
  1353 => x"ba052257",
  1354 => x"5c80e453",
  1355 => x"805280ee",
  1356 => x"e83fb008",
  1357 => x"722e0981",
  1358 => x"06833881",
  1359 => x"5272802e",
  1360 => x"b3387180",
  1361 => x"2e923880",
  1362 => x"e45180ed",
  1363 => x"ed3fff13",
  1364 => x"7081ff06",
  1365 => x"5452d539",
  1366 => x"72802e98",
  1367 => x"3880eecc",
  1368 => x"3fb00881",
  1369 => x"ff065271",
  1370 => x"952e82a7",
  1371 => x"387180c3",
  1372 => x"2e81f838",
  1373 => x"ff147081",
  1374 => x"ff065553",
  1375 => x"73ffaa38",
  1376 => x"75802e81",
  1377 => x"d6388a7c",
  1378 => x"095c5a81",
  1379 => x"5180eebe",
  1380 => x"3f7b5180",
  1381 => x"eeb83f7a",
  1382 => x"5180eeb2",
  1383 => x"3f807055",
  1384 => x"57818055",
  1385 => x"ff157081",
  1386 => x"ff065652",
  1387 => x"9a537580",
  1388 => x"2e913878",
  1389 => x"7081055a",
  1390 => x"33ff1770",
  1391 => x"83ffff06",
  1392 => x"58535372",
  1393 => x"5180ee86",
  1394 => x"3f77802e",
  1395 => x"81b13872",
  1396 => x"882b7432",
  1397 => x"53875472",
  1398 => x"902b5280",
  1399 => x"72248190",
  1400 => x"38721083",
  1401 => x"fffe0653",
  1402 => x"ff145473",
  1403 => x"8025e838",
  1404 => x"7283ffff",
  1405 => x"065474ff",
  1406 => x"ab387780",
  1407 => x"2e818b38",
  1408 => x"73882a51",
  1409 => x"80edc73f",
  1410 => x"7381ff06",
  1411 => x"5180edbe",
  1412 => x"3f80ed85",
  1413 => x"3fb008f9",
  1414 => x"3880ed90",
  1415 => x"3fb00881",
  1416 => x"ff065271",
  1417 => x"862e80f0",
  1418 => x"3871982e",
  1419 => x"80f538ff",
  1420 => x"1a7081ff",
  1421 => x"065b5479",
  1422 => x"fed138fe",
  1423 => x"5271b00c",
  1424 => x"8d3d0d04",
  1425 => x"80ecd23f",
  1426 => x"b008f938",
  1427 => x"80ecdd3f",
  1428 => x"b00881ff",
  1429 => x"06527186",
  1430 => x"2ee33884",
  1431 => x"5180ecee",
  1432 => x"3f80ecb5",
  1433 => x"3fb008dc",
  1434 => x"38e23981",
  1435 => x"58fe9139",
  1436 => x"7210a0a1",
  1437 => x"327083ff",
  1438 => x"ff065452",
  1439 => x"feea3972",
  1440 => x"177081ff",
  1441 => x"065852fe",
  1442 => x"ed397651",
  1443 => x"80ecbf3f",
  1444 => x"feff3980",
  1445 => x"58fde939",
  1446 => x"811c7081",
  1447 => x"ff065d55",
  1448 => x"fdde39ff",
  1449 => x"0bb00c8d",
  1450 => x"3d0d04f6",
  1451 => x"3d0d7c7e",
  1452 => x"5b5980c3",
  1453 => x"578a5581",
  1454 => x"5b805880",
  1455 => x"e4538054",
  1456 => x"777a2482",
  1457 => x"b4387651",
  1458 => x"80ec833f",
  1459 => x"805280eb",
  1460 => x"c83fb008",
  1461 => x"722e0981",
  1462 => x"06833881",
  1463 => x"5272802e",
  1464 => x"81ed3871",
  1465 => x"802e9238",
  1466 => x"80e45180",
  1467 => x"eacc3fff",
  1468 => x"137081ff",
  1469 => x"065452d4",
  1470 => x"3972802e",
  1471 => x"81d13880",
  1472 => x"ebaa3fb0",
  1473 => x"0881ff06",
  1474 => x"5271842e",
  1475 => x"82883871",
  1476 => x"842481cf",
  1477 => x"3871812e",
  1478 => x"09810681",
  1479 => x"b2388657",
  1480 => x"80eb893f",
  1481 => x"b00881ff",
  1482 => x"06537a73",
  1483 => x"2e833895",
  1484 => x"5780eaf8",
  1485 => x"3fb00809",
  1486 => x"7081ff06",
  1487 => x"57527a76",
  1488 => x"2e833895",
  1489 => x"57805380",
  1490 => x"eae23f78",
  1491 => x"1356b008",
  1492 => x"76348113",
  1493 => x"7081ff06",
  1494 => x"70982b58",
  1495 => x"54527580",
  1496 => x"25e53880",
  1497 => x"56781670",
  1498 => x"3370882b",
  1499 => x"76325253",
  1500 => x"53875472",
  1501 => x"902b5280",
  1502 => x"7224818b",
  1503 => x"38721083",
  1504 => x"fffe0653",
  1505 => x"ff145473",
  1506 => x"8025e838",
  1507 => x"7283ffff",
  1508 => x"06811770",
  1509 => x"81ff0670",
  1510 => x"982b5658",
  1511 => x"53547280",
  1512 => x"25c33880",
  1513 => x"ea863fb0",
  1514 => x"0881ff06",
  1515 => x"74882a57",
  1516 => x"5372762e",
  1517 => x"83389557",
  1518 => x"80e9f13f",
  1519 => x"b00881ff",
  1520 => x"067481ff",
  1521 => x"06535675",
  1522 => x"722e80d7",
  1523 => x"389557ff",
  1524 => x"157081ff",
  1525 => x"06565274",
  1526 => x"fde138fe",
  1527 => x"0bb00c8c",
  1528 => x"3d0d0471",
  1529 => x"982e0981",
  1530 => x"06e53886",
  1531 => x"5180e9de",
  1532 => x"3fff0bb0",
  1533 => x"0c8c3d0d",
  1534 => x"04985180",
  1535 => x"e9d03ffd",
  1536 => x"0bb00c8c",
  1537 => x"3d0d0472",
  1538 => x"10a0a132",
  1539 => x"7083ffff",
  1540 => x"065452fe",
  1541 => x"ef398651",
  1542 => x"80e9b33f",
  1543 => x"77b00c8c",
  1544 => x"3d0d0476",
  1545 => x"862e0981",
  1546 => x"06ffa438",
  1547 => x"77848080",
  1548 => x"2982800a",
  1549 => x"0570902c",
  1550 => x"81801b81",
  1551 => x"1e7081ff",
  1552 => x"065f575b",
  1553 => x"595374fc",
  1554 => x"f238ff8f",
  1555 => x"39fe3d0d",
  1556 => x"02930533",
  1557 => x"02840597",
  1558 => x"05335452",
  1559 => x"71842e80",
  1560 => x"ed387184",
  1561 => x"24923871",
  1562 => x"812eaf38",
  1563 => x"81d1a451",
  1564 => x"80e4b43f",
  1565 => x"843d0d04",
  1566 => x"7180d52e",
  1567 => x"098106ec",
  1568 => x"3881d1b0",
  1569 => x"5180e49f",
  1570 => x"3f728a26",
  1571 => x"80cd3872",
  1572 => x"101081d5",
  1573 => x"d8055271",
  1574 => x"080481d1",
  1575 => x"bc5180e4",
  1576 => x"863f729a",
  1577 => x"2e829c38",
  1578 => x"729a2480",
  1579 => x"c638728c",
  1580 => x"2e829c38",
  1581 => x"728c2481",
  1582 => x"ef387286",
  1583 => x"2e098106",
  1584 => x"9a3881d1",
  1585 => x"c85180e3",
  1586 => x"de3f843d",
  1587 => x"0d0481d1",
  1588 => x"d85180e3",
  1589 => x"d23f728f",
  1590 => x"2e8d3881",
  1591 => x"d1e45180",
  1592 => x"e3c53f84",
  1593 => x"3d0d0481",
  1594 => x"d1f45180",
  1595 => x"e3b93f84",
  1596 => x"3d0d0472",
  1597 => x"a82e81e3",
  1598 => x"3872a824",
  1599 => x"818d3872",
  1600 => x"9d2e0981",
  1601 => x"06d53881",
  1602 => x"d28c5180",
  1603 => x"e3993f84",
  1604 => x"3d0d0481",
  1605 => x"d2a85180",
  1606 => x"e38d3f84",
  1607 => x"3d0d0481",
  1608 => x"d2c85180",
  1609 => x"e3813f84",
  1610 => x"3d0d0481",
  1611 => x"d2dc5180",
  1612 => x"e2f53f84",
  1613 => x"3d0d0481",
  1614 => x"d2f85180",
  1615 => x"e2e93f84",
  1616 => x"3d0d0481",
  1617 => x"ceb05180",
  1618 => x"e2dd3f84",
  1619 => x"3d0d0481",
  1620 => x"d3905180",
  1621 => x"e2d13f84",
  1622 => x"3d0d0481",
  1623 => x"d3a45180",
  1624 => x"e2c53f84",
  1625 => x"3d0d0481",
  1626 => x"d3b45180",
  1627 => x"e2b93f84",
  1628 => x"3d0d0481",
  1629 => x"d3cc5180",
  1630 => x"e2ad3f84",
  1631 => x"3d0d0481",
  1632 => x"d3e05180",
  1633 => x"e2a13f84",
  1634 => x"3d0d0472",
  1635 => x"80c52e80",
  1636 => x"d6387280",
  1637 => x"e12e0981",
  1638 => x"06fec038",
  1639 => x"81d3f051",
  1640 => x"80e2843f",
  1641 => x"843d0d04",
  1642 => x"728f2e80",
  1643 => x"c6387291",
  1644 => x"2e098106",
  1645 => x"fea53881",
  1646 => x"d4805180",
  1647 => x"e1e93f84",
  1648 => x"3d0d0481",
  1649 => x"d4945180",
  1650 => x"e1dd3f84",
  1651 => x"3d0d0481",
  1652 => x"d4b05180",
  1653 => x"e1d13f84",
  1654 => x"3d0d0481",
  1655 => x"d4c05180",
  1656 => x"e1c53f84",
  1657 => x"3d0d0481",
  1658 => x"d4e05180",
  1659 => x"e1b93f84",
  1660 => x"3d0d0481",
  1661 => x"d4f85180",
  1662 => x"e1ad3f84",
  1663 => x"3d0d04f7",
  1664 => x"3d0d02b3",
  1665 => x"05337c70",
  1666 => x"08c08080",
  1667 => x"0659545a",
  1668 => x"80567583",
  1669 => x"2b7707bf",
  1670 => x"e0800770",
  1671 => x"70840552",
  1672 => x"0871088c",
  1673 => x"2abffe80",
  1674 => x"06790771",
  1675 => x"982a728c",
  1676 => x"2a9fff06",
  1677 => x"73852a70",
  1678 => x"8f06759f",
  1679 => x"06565158",
  1680 => x"5d585255",
  1681 => x"58748d38",
  1682 => x"8116568f",
  1683 => x"7627c338",
  1684 => x"8b3d0d04",
  1685 => x"81d59451",
  1686 => x"80e0cc3f",
  1687 => x"755180e2",
  1688 => x"903f8452",
  1689 => x"b00851a5",
  1690 => x"cb3f81d5",
  1691 => x"a05180e0",
  1692 => x"b63f7452",
  1693 => x"885180e0",
  1694 => x"d13f8452",
  1695 => x"b00851a5",
  1696 => x"b33f81d5",
  1697 => x"a85180e0",
  1698 => x"9e3f7852",
  1699 => x"905180e0",
  1700 => x"b93f8652",
  1701 => x"b00851a5",
  1702 => x"9b3f81d5",
  1703 => x"b05180e0",
  1704 => x"863f7251",
  1705 => x"80e1ca3f",
  1706 => x"8452b008",
  1707 => x"51a5853f",
  1708 => x"81d5b851",
  1709 => x"80dff03f",
  1710 => x"735180e1",
  1711 => x"b43f8452",
  1712 => x"b00851a4",
  1713 => x"ef3f81d5",
  1714 => x"c05180df",
  1715 => x"da3f7752",
  1716 => x"a05180df",
  1717 => x"f53f8a52",
  1718 => x"b00851a4",
  1719 => x"d73f7993",
  1720 => x"388a5180",
  1721 => x"dfa73f81",
  1722 => x"16568f76",
  1723 => x"27fea338",
  1724 => x"fede3978",
  1725 => x"81ff0652",
  1726 => x"7451fad1",
  1727 => x"3f8a5180",
  1728 => x"df8b3fe3",
  1729 => x"39f83d0d",
  1730 => x"02ab0533",
  1731 => x"59805675",
  1732 => x"852be090",
  1733 => x"11e08012",
  1734 => x"0870982a",
  1735 => x"718c2a9f",
  1736 => x"ff067285",
  1737 => x"2a708f06",
  1738 => x"749f0655",
  1739 => x"51585b53",
  1740 => x"56595574",
  1741 => x"802e81ae",
  1742 => x"3875bf26",
  1743 => x"81b63881",
  1744 => x"d5c85180",
  1745 => x"dee13f75",
  1746 => x"5180e0a5",
  1747 => x"3f8652b0",
  1748 => x"0851a3e0",
  1749 => x"3f81d5a0",
  1750 => x"5180decb",
  1751 => x"3f745288",
  1752 => x"5180dee6",
  1753 => x"3f8452b0",
  1754 => x"0851a3c8",
  1755 => x"3f81d5a8",
  1756 => x"5180deb3",
  1757 => x"3f765290",
  1758 => x"5180dece",
  1759 => x"3f8652b0",
  1760 => x"0851a3b0",
  1761 => x"3f81d5b0",
  1762 => x"5180de9b",
  1763 => x"3f725180",
  1764 => x"dfdf3f84",
  1765 => x"52b00851",
  1766 => x"a39a3f81",
  1767 => x"d5b85180",
  1768 => x"de853f73",
  1769 => x"5180dfc9",
  1770 => x"3f8452b0",
  1771 => x"0851a384",
  1772 => x"3f81d5c0",
  1773 => x"5180ddef",
  1774 => x"3f7708c0",
  1775 => x"80800652",
  1776 => x"a05180de",
  1777 => x"853f8a52",
  1778 => x"b00851a2",
  1779 => x"e73f7881",
  1780 => x"b9388a51",
  1781 => x"80ddb63f",
  1782 => x"80537481",
  1783 => x"2e81e638",
  1784 => x"76862e81",
  1785 => x"c2388116",
  1786 => x"5680ff76",
  1787 => x"27fea038",
  1788 => x"8a3d0d04",
  1789 => x"81d5d051",
  1790 => x"80ddac3f",
  1791 => x"c0165180",
  1792 => x"deef3f86",
  1793 => x"52b00851",
  1794 => x"a2aa3f81",
  1795 => x"d5a05180",
  1796 => x"dd953f74",
  1797 => x"52885180",
  1798 => x"ddb03f84",
  1799 => x"52b00851",
  1800 => x"a2923f81",
  1801 => x"d5a85180",
  1802 => x"dcfd3f76",
  1803 => x"52905180",
  1804 => x"dd983f86",
  1805 => x"52b00851",
  1806 => x"a1fa3f81",
  1807 => x"d5b05180",
  1808 => x"dce53f72",
  1809 => x"5180dea9",
  1810 => x"3f8452b0",
  1811 => x"0851a1e4",
  1812 => x"3f81d5b8",
  1813 => x"5180dccf",
  1814 => x"3f735180",
  1815 => x"de933f84",
  1816 => x"52b00851",
  1817 => x"a1ce3f81",
  1818 => x"d5c05180",
  1819 => x"dcb93f77",
  1820 => x"08c08080",
  1821 => x"0652a051",
  1822 => x"80dccf3f",
  1823 => x"8a52b008",
  1824 => x"51a1b13f",
  1825 => x"78802efe",
  1826 => x"c9387681",
  1827 => x"ff065274",
  1828 => x"51f7ba3f",
  1829 => x"8a5180db",
  1830 => x"f43f8053",
  1831 => x"74812e09",
  1832 => x"8106febc",
  1833 => x"389f3972",
  1834 => x"81065776",
  1835 => x"802efeb6",
  1836 => x"38785277",
  1837 => x"51fac83f",
  1838 => x"81165680",
  1839 => x"ff7627fc",
  1840 => x"ce38feac",
  1841 => x"39745376",
  1842 => x"862e0981",
  1843 => x"06fe9738",
  1844 => x"d639803d",
  1845 => x"0d81f684",
  1846 => x"08519971",
  1847 => x"0c81800b",
  1848 => x"84120c81",
  1849 => x"f6800851",
  1850 => x"99710c81",
  1851 => x"800b8412",
  1852 => x"0c823d0d",
  1853 => x"04fe3d0d",
  1854 => x"74028405",
  1855 => x"97053302",
  1856 => x"88059b05",
  1857 => x"3388130c",
  1858 => x"8c120c53",
  1859 => x"8c130870",
  1860 => x"812a8106",
  1861 => x"515271f4",
  1862 => x"388c1308",
  1863 => x"7081ff06",
  1864 => x"b00c5184",
  1865 => x"3d0d0480",
  1866 => x"3d0d728c",
  1867 => x"11087087",
  1868 => x"2a813281",
  1869 => x"06b00c51",
  1870 => x"51823d0d",
  1871 => x"04fd3d0d",
  1872 => x"02970533",
  1873 => x"5481ec53",
  1874 => x"81905281",
  1875 => x"f6840851",
  1876 => x"ffa33f73",
  1877 => x"53905281",
  1878 => x"f6840851",
  1879 => x"ff973f81",
  1880 => x"ed538190",
  1881 => x"5281f684",
  1882 => x"0851ff89",
  1883 => x"3f805380",
  1884 => x"e05281f6",
  1885 => x"840851fe",
  1886 => x"fc3f81f6",
  1887 => x"84088811",
  1888 => x"08b00c54",
  1889 => x"853d0d04",
  1890 => x"fc3d0d02",
  1891 => x"9b053302",
  1892 => x"84059f05",
  1893 => x"33565481",
  1894 => x"ec538190",
  1895 => x"5281f684",
  1896 => x"0851fed1",
  1897 => x"3f735390",
  1898 => x"5281f684",
  1899 => x"0851fec5",
  1900 => x"3f745380",
  1901 => x"d05281f6",
  1902 => x"840851fe",
  1903 => x"b83f73b0",
  1904 => x"0c863d0d",
  1905 => x"04fe3d0d",
  1906 => x"fe883f81",
  1907 => x"ec538190",
  1908 => x"5281f684",
  1909 => x"0851fe9d",
  1910 => x"3f9d5390",
  1911 => x"5281f684",
  1912 => x"0851fe91",
  1913 => x"3f80c553",
  1914 => x"80d05281",
  1915 => x"f6840851",
  1916 => x"fe833f81",
  1917 => x"ec538190",
  1918 => x"5281f684",
  1919 => x"0851fdf5",
  1920 => x"3fa15390",
  1921 => x"5281f684",
  1922 => x"0851fde9",
  1923 => x"3f895380",
  1924 => x"d05281f6",
  1925 => x"840851fd",
  1926 => x"dc3f81ec",
  1927 => x"53819052",
  1928 => x"81f68408",
  1929 => x"51fdce3f",
  1930 => x"b3539052",
  1931 => x"81f68408",
  1932 => x"51fdc23f",
  1933 => x"885380d0",
  1934 => x"5281f684",
  1935 => x"0851fdb5",
  1936 => x"3f81ec53",
  1937 => x"81905281",
  1938 => x"f6840851",
  1939 => x"fda73fb4",
  1940 => x"53905281",
  1941 => x"f6840851",
  1942 => x"fd9b3f96",
  1943 => x"5380d052",
  1944 => x"81f68408",
  1945 => x"51fd8e3f",
  1946 => x"81ec5381",
  1947 => x"905281f6",
  1948 => x"840851fd",
  1949 => x"803fb653",
  1950 => x"905281f6",
  1951 => x"840851fc",
  1952 => x"f43f80e0",
  1953 => x"5380d052",
  1954 => x"81f68408",
  1955 => x"51fce63f",
  1956 => x"81ec5381",
  1957 => x"905281f6",
  1958 => x"840851fc",
  1959 => x"d83f80c9",
  1960 => x"53905281",
  1961 => x"f6840851",
  1962 => x"fccb3f81",
  1963 => x"c05380d0",
  1964 => x"5281f684",
  1965 => x"0851fcbd",
  1966 => x"3f843d0d",
  1967 => x"04fd3d0d",
  1968 => x"02970533",
  1969 => x"0284059b",
  1970 => x"05337181",
  1971 => x"b00781bf",
  1972 => x"06535454",
  1973 => x"f8808098",
  1974 => x"8071710c",
  1975 => x"73842a90",
  1976 => x"07710c73",
  1977 => x"8f06710c",
  1978 => x"527281f5",
  1979 => x"d0347381",
  1980 => x"f5d43485",
  1981 => x"3d0d04fd",
  1982 => x"3d0d0297",
  1983 => x"053381f5",
  1984 => x"d4335473",
  1985 => x"05870602",
  1986 => x"84059a05",
  1987 => x"2281f5d0",
  1988 => x"33547305",
  1989 => x"7081ff06",
  1990 => x"7281b007",
  1991 => x"54515454",
  1992 => x"f8808098",
  1993 => x"8071710c",
  1994 => x"73842a90",
  1995 => x"07710c73",
  1996 => x"8f06710c",
  1997 => x"527281f5",
  1998 => x"d0347381",
  1999 => x"f5d43485",
  2000 => x"3d0d04ff",
  2001 => x"3d0d028f",
  2002 => x"0533f880",
  2003 => x"8098840c",
  2004 => x"81f5d033",
  2005 => x"81055170",
  2006 => x"81f5d034",
  2007 => x"833d0d04",
  2008 => x"ff3d0d80",
  2009 => x"527181b0",
  2010 => x"0781bf06",
  2011 => x"f8808098",
  2012 => x"800c900b",
  2013 => x"f8808098",
  2014 => x"800c800b",
  2015 => x"f8808098",
  2016 => x"800c8051",
  2017 => x"800bf880",
  2018 => x"8098840c",
  2019 => x"81117081",
  2020 => x"ff065151",
  2021 => x"80e57127",
  2022 => x"eb388112",
  2023 => x"7081ff06",
  2024 => x"53518772",
  2025 => x"27ffbe38",
  2026 => x"81b00bf8",
  2027 => x"80809880",
  2028 => x"0c900bf8",
  2029 => x"80809880",
  2030 => x"0c800bf8",
  2031 => x"80809880",
  2032 => x"0c800b81",
  2033 => x"f5d03480",
  2034 => x"0b81f5d4",
  2035 => x"34833d0d",
  2036 => x"04ff3d0d",
  2037 => x"80c00bf8",
  2038 => x"80809880",
  2039 => x"0c81a10b",
  2040 => x"f8808098",
  2041 => x"800c81c0",
  2042 => x"0bf88080",
  2043 => x"98800c81",
  2044 => x"a40bf880",
  2045 => x"8098800c",
  2046 => x"81a60bf8",
  2047 => x"80809880",
  2048 => x"0c81a20b",
  2049 => x"f8808098",
  2050 => x"800caf0b",
  2051 => x"f8808098",
  2052 => x"800ca50b",
  2053 => x"f8808098",
  2054 => x"800c8181",
  2055 => x"0bf88080",
  2056 => x"98800c9d",
  2057 => x"0bf88080",
  2058 => x"98800c81",
  2059 => x"fa0bf880",
  2060 => x"8098800c",
  2061 => x"800bf880",
  2062 => x"8098800c",
  2063 => x"80527181",
  2064 => x"b00781bf",
  2065 => x"06f88080",
  2066 => x"98800c90",
  2067 => x"0bf88080",
  2068 => x"98800c80",
  2069 => x"0bf88080",
  2070 => x"98800c80",
  2071 => x"51800bf8",
  2072 => x"80809884",
  2073 => x"0c811170",
  2074 => x"81ff0651",
  2075 => x"5180e571",
  2076 => x"27eb3881",
  2077 => x"127081ff",
  2078 => x"06535187",
  2079 => x"7227ffbe",
  2080 => x"3881b00b",
  2081 => x"f8808098",
  2082 => x"800c900b",
  2083 => x"f8808098",
  2084 => x"800c800b",
  2085 => x"f8808098",
  2086 => x"800c800b",
  2087 => x"81f5d034",
  2088 => x"800b81f5",
  2089 => x"d43481af",
  2090 => x"0bf88080",
  2091 => x"98800c83",
  2092 => x"3d0d0480",
  2093 => x"3d0d028f",
  2094 => x"05337382",
  2095 => x"9eb40c51",
  2096 => x"70829eb8",
  2097 => x"34823d0d",
  2098 => x"04ee3d0d",
  2099 => x"64028405",
  2100 => x"80d70533",
  2101 => x"02880580",
  2102 => x"db053359",
  2103 => x"57598076",
  2104 => x"81067781",
  2105 => x"2a810678",
  2106 => x"832b8180",
  2107 => x"0679822a",
  2108 => x"8106575e",
  2109 => x"415f5d81",
  2110 => x"ff42727d",
  2111 => x"2e098106",
  2112 => x"83387c42",
  2113 => x"768a2e83",
  2114 => x"b9388819",
  2115 => x"08557480",
  2116 => x"2e83a438",
  2117 => x"8519335a",
  2118 => x"ff53767a",
  2119 => x"268e3884",
  2120 => x"19335473",
  2121 => x"77268538",
  2122 => x"76743153",
  2123 => x"74137033",
  2124 => x"54587281",
  2125 => x"ff06831a",
  2126 => x"3370982b",
  2127 => x"81ff0a11",
  2128 => x"9b2a8105",
  2129 => x"5b454240",
  2130 => x"81537483",
  2131 => x"38745372",
  2132 => x"81ff0643",
  2133 => x"807a81ff",
  2134 => x"06545cff",
  2135 => x"54767326",
  2136 => x"8b388419",
  2137 => x"33537673",
  2138 => x"2783f438",
  2139 => x"737481ff",
  2140 => x"06555380",
  2141 => x"5a797324",
  2142 => x"ab38747a",
  2143 => x"2e098106",
  2144 => x"82e13860",
  2145 => x"982b81ff",
  2146 => x"0a119b2a",
  2147 => x"821b3371",
  2148 => x"71291170",
  2149 => x"81ff0678",
  2150 => x"71298c1f",
  2151 => x"08055245",
  2152 => x"5d575d53",
  2153 => x"7f630570",
  2154 => x"81ff0670",
  2155 => x"612b7081",
  2156 => x"ff067b62",
  2157 => x"2b7081ff",
  2158 => x"067b832a",
  2159 => x"81065f53",
  2160 => x"58525e42",
  2161 => x"5578802e",
  2162 => x"8f3881f5",
  2163 => x"d0336105",
  2164 => x"567580e6",
  2165 => x"2483c538",
  2166 => x"7f782961",
  2167 => x"3041577c",
  2168 => x"7e2c982b",
  2169 => x"70982c55",
  2170 => x"55737725",
  2171 => x"818238ff",
  2172 => x"1c7d8106",
  2173 => x"5a537c73",
  2174 => x"2e83c438",
  2175 => x"7e86a638",
  2176 => x"6184eb38",
  2177 => x"7d802e82",
  2178 => x"a4387914",
  2179 => x"70337058",
  2180 => x"54558055",
  2181 => x"78752e85",
  2182 => x"3872842a",
  2183 => x"5675832a",
  2184 => x"70810651",
  2185 => x"5372802e",
  2186 => x"843881c0",
  2187 => x"5575822a",
  2188 => x"70810651",
  2189 => x"5372802e",
  2190 => x"853874b0",
  2191 => x"07557581",
  2192 => x"2a708106",
  2193 => x"51537280",
  2194 => x"2e853874",
  2195 => x"8c075575",
  2196 => x"81065372",
  2197 => x"802e8538",
  2198 => x"74830755",
  2199 => x"7451f9e3",
  2200 => x"3f771498",
  2201 => x"2b70982c",
  2202 => x"55567674",
  2203 => x"24ff9b38",
  2204 => x"62802e95",
  2205 => x"3861ff1d",
  2206 => x"54547c73",
  2207 => x"2e81fb38",
  2208 => x"7351f9bf",
  2209 => x"3f7e81ea",
  2210 => x"387f5281",
  2211 => x"51f8e83f",
  2212 => x"811d7081",
  2213 => x"ff065e54",
  2214 => x"7b7d26fe",
  2215 => x"c2386052",
  2216 => x"7b307098",
  2217 => x"2b70982c",
  2218 => x"53585bf8",
  2219 => x"ca3f6053",
  2220 => x"72b00c94",
  2221 => x"3d0d0482",
  2222 => x"1933851a",
  2223 => x"335b53fc",
  2224 => x"f13981f5",
  2225 => x"d4335372",
  2226 => x"8726819a",
  2227 => x"38811356",
  2228 => x"80527581",
  2229 => x"ff0651f7",
  2230 => x"e43f8053",
  2231 => x"72b00c94",
  2232 => x"3d0d0473",
  2233 => x"802eaf38",
  2234 => x"ff147081",
  2235 => x"ff06555a",
  2236 => x"7381ff2e",
  2237 => x"a1387470",
  2238 => x"81055633",
  2239 => x"7c057083",
  2240 => x"ffff06ff",
  2241 => x"167081ff",
  2242 => x"06575c5d",
  2243 => x"537381ff",
  2244 => x"2e098106",
  2245 => x"e1386098",
  2246 => x"2b81ff0a",
  2247 => x"119b2a70",
  2248 => x"7e291e8c",
  2249 => x"1c08055c",
  2250 => x"4255fcf8",
  2251 => x"39791470",
  2252 => x"335259f8",
  2253 => x"8e3f7714",
  2254 => x"982b7098",
  2255 => x"2c555673",
  2256 => x"7725feac",
  2257 => x"38791470",
  2258 => x"335259f7",
  2259 => x"f63f7714",
  2260 => x"982b7098",
  2261 => x"2c555676",
  2262 => x"7424d238",
  2263 => x"fe923976",
  2264 => x"733154fc",
  2265 => x"87398052",
  2266 => x"8051f6d1",
  2267 => x"3f8053fe",
  2268 => x"eb397351",
  2269 => x"f7cd3ffe",
  2270 => x"9039617b",
  2271 => x"327081ff",
  2272 => x"0655557d",
  2273 => x"802efdf8",
  2274 => x"387a812a",
  2275 => x"74327052",
  2276 => x"54f7b03f",
  2277 => x"7e802efd",
  2278 => x"f038d739",
  2279 => x"81f5d433",
  2280 => x"7c055380",
  2281 => x"527281ff",
  2282 => x"0651f691",
  2283 => x"3f805376",
  2284 => x"a02efdfc",
  2285 => x"387f7829",
  2286 => x"61304157",
  2287 => x"fca1397e",
  2288 => x"87ad3861",
  2289 => x"85eb387d",
  2290 => x"802e80ec",
  2291 => x"38791470",
  2292 => x"337c0770",
  2293 => x"52545680",
  2294 => x"5578752e",
  2295 => x"85387284",
  2296 => x"2a567583",
  2297 => x"2a708106",
  2298 => x"51537280",
  2299 => x"2e843881",
  2300 => x"c0557582",
  2301 => x"2a708106",
  2302 => x"51537280",
  2303 => x"2e853874",
  2304 => x"b0075575",
  2305 => x"812a7081",
  2306 => x"06515372",
  2307 => x"802e8538",
  2308 => x"748c0755",
  2309 => x"75810653",
  2310 => x"72802e85",
  2311 => x"38748307",
  2312 => x"557451f6",
  2313 => x"9e3f7714",
  2314 => x"982b7098",
  2315 => x"2c555376",
  2316 => x"7424ff99",
  2317 => x"38fcb939",
  2318 => x"79147033",
  2319 => x"7c075256",
  2320 => x"f6813f77",
  2321 => x"14982b70",
  2322 => x"982c5559",
  2323 => x"737725fc",
  2324 => x"9f387914",
  2325 => x"70337c07",
  2326 => x"5256f5e7",
  2327 => x"3f771498",
  2328 => x"2b70982c",
  2329 => x"55597674",
  2330 => x"24ce38fc",
  2331 => x"83397d80",
  2332 => x"2e80f038",
  2333 => x"79147033",
  2334 => x"70585455",
  2335 => x"80557875",
  2336 => x"2e853872",
  2337 => x"842a5675",
  2338 => x"832a7081",
  2339 => x"06515372",
  2340 => x"802e8438",
  2341 => x"81c05575",
  2342 => x"822a7081",
  2343 => x"06515372",
  2344 => x"802e8538",
  2345 => x"74b00755",
  2346 => x"75812a70",
  2347 => x"81065153",
  2348 => x"72802e85",
  2349 => x"38748c07",
  2350 => x"55758106",
  2351 => x"5372802e",
  2352 => x"85387483",
  2353 => x"07557409",
  2354 => x"7081ff06",
  2355 => x"5253f4f3",
  2356 => x"3f771498",
  2357 => x"2b70982c",
  2358 => x"55567674",
  2359 => x"24ff9538",
  2360 => x"fb8e3979",
  2361 => x"14703370",
  2362 => x"097081ff",
  2363 => x"06545854",
  2364 => x"55f4d03f",
  2365 => x"7714982b",
  2366 => x"70982c55",
  2367 => x"59737725",
  2368 => x"faee3879",
  2369 => x"14703370",
  2370 => x"097081ff",
  2371 => x"06545854",
  2372 => x"55f4b03f",
  2373 => x"7714982b",
  2374 => x"70982c55",
  2375 => x"59767424",
  2376 => x"c238facc",
  2377 => x"3961802e",
  2378 => x"81ce387d",
  2379 => x"802e80f7",
  2380 => x"38791470",
  2381 => x"33705854",
  2382 => x"55805578",
  2383 => x"752e8538",
  2384 => x"72842a56",
  2385 => x"75832a70",
  2386 => x"81065153",
  2387 => x"72802e84",
  2388 => x"3881c055",
  2389 => x"75822a70",
  2390 => x"81065153",
  2391 => x"72802e85",
  2392 => x"3874b007",
  2393 => x"5575812a",
  2394 => x"70810651",
  2395 => x"5372802e",
  2396 => x"8538748c",
  2397 => x"07557581",
  2398 => x"06537280",
  2399 => x"2e853874",
  2400 => x"83075574",
  2401 => x"097081ff",
  2402 => x"06705357",
  2403 => x"53f3b43f",
  2404 => x"7551f3af",
  2405 => x"3f771498",
  2406 => x"2b70982c",
  2407 => x"55557674",
  2408 => x"24ff8e38",
  2409 => x"f9ca3979",
  2410 => x"14703370",
  2411 => x"097081ff",
  2412 => x"06705559",
  2413 => x"555659f3",
  2414 => x"8a3f7551",
  2415 => x"f3853f77",
  2416 => x"14982b70",
  2417 => x"982c5559",
  2418 => x"737725f9",
  2419 => x"a3387914",
  2420 => x"70337009",
  2421 => x"7081ff06",
  2422 => x"70555955",
  2423 => x"5659f2e3",
  2424 => x"3f7551f2",
  2425 => x"de3f7714",
  2426 => x"982b7098",
  2427 => x"2c555976",
  2428 => x"7424ffb3",
  2429 => x"38f8f939",
  2430 => x"7d802e80",
  2431 => x"f4387914",
  2432 => x"70337058",
  2433 => x"54558055",
  2434 => x"78752e85",
  2435 => x"3872842a",
  2436 => x"5675832a",
  2437 => x"70810651",
  2438 => x"5372802e",
  2439 => x"843881c0",
  2440 => x"5575822a",
  2441 => x"70810651",
  2442 => x"5372802e",
  2443 => x"853874b0",
  2444 => x"07557581",
  2445 => x"2a708106",
  2446 => x"51537280",
  2447 => x"2e853874",
  2448 => x"8c075575",
  2449 => x"81065372",
  2450 => x"802e8538",
  2451 => x"74830755",
  2452 => x"7481ff06",
  2453 => x"705256f1",
  2454 => x"ea3f7551",
  2455 => x"f1e53f77",
  2456 => x"14982b70",
  2457 => x"982c5555",
  2458 => x"767424ff",
  2459 => x"9138f880",
  2460 => x"39791470",
  2461 => x"33705357",
  2462 => x"53f1c83f",
  2463 => x"7551f1c3",
  2464 => x"3f771498",
  2465 => x"2b70982c",
  2466 => x"55597377",
  2467 => x"25f7e138",
  2468 => x"79147033",
  2469 => x"70535753",
  2470 => x"f1a93f75",
  2471 => x"51f1a43f",
  2472 => x"7714982b",
  2473 => x"70982c55",
  2474 => x"59767424",
  2475 => x"c438f7c0",
  2476 => x"397d802e",
  2477 => x"80f23879",
  2478 => x"1470337c",
  2479 => x"07705254",
  2480 => x"56805578",
  2481 => x"752e8538",
  2482 => x"72842a56",
  2483 => x"75832a70",
  2484 => x"81065153",
  2485 => x"72802e84",
  2486 => x"3881c055",
  2487 => x"75822a70",
  2488 => x"81065153",
  2489 => x"72802e85",
  2490 => x"3874b007",
  2491 => x"5575812a",
  2492 => x"70810651",
  2493 => x"5372802e",
  2494 => x"8538748c",
  2495 => x"07557581",
  2496 => x"06537280",
  2497 => x"2e853874",
  2498 => x"83075574",
  2499 => x"097081ff",
  2500 => x"065256f0",
  2501 => x"ae3f7714",
  2502 => x"982b7098",
  2503 => x"2c555376",
  2504 => x"7424ff93",
  2505 => x"38f6c939",
  2506 => x"79147033",
  2507 => x"7c077009",
  2508 => x"7081ff06",
  2509 => x"54555659",
  2510 => x"f0893f77",
  2511 => x"14982b70",
  2512 => x"982c5559",
  2513 => x"737725f6",
  2514 => x"a7387914",
  2515 => x"70337c07",
  2516 => x"70097081",
  2517 => x"ff065455",
  2518 => x"5659efe7",
  2519 => x"3f771498",
  2520 => x"2b70982c",
  2521 => x"55597674",
  2522 => x"24ffbd38",
  2523 => x"f6823961",
  2524 => x"802e81d4",
  2525 => x"387d802e",
  2526 => x"80f93879",
  2527 => x"1470337c",
  2528 => x"07705254",
  2529 => x"56805578",
  2530 => x"752e8538",
  2531 => x"72842a56",
  2532 => x"75832a70",
  2533 => x"81065153",
  2534 => x"72802e84",
  2535 => x"3881c055",
  2536 => x"75822a70",
  2537 => x"81065153",
  2538 => x"72802e85",
  2539 => x"3874b007",
  2540 => x"5575812a",
  2541 => x"70810651",
  2542 => x"5372802e",
  2543 => x"8538748c",
  2544 => x"07557581",
  2545 => x"06537280",
  2546 => x"2e853874",
  2547 => x"83075574",
  2548 => x"097081ff",
  2549 => x"06705354",
  2550 => x"56eee83f",
  2551 => x"7251eee3",
  2552 => x"3f771498",
  2553 => x"2b70982c",
  2554 => x"55567674",
  2555 => x"24ff8c38",
  2556 => x"f4fe3979",
  2557 => x"1470337c",
  2558 => x"07700970",
  2559 => x"81ff0670",
  2560 => x"55535757",
  2561 => x"53eebc3f",
  2562 => x"7251eeb7",
  2563 => x"3f771498",
  2564 => x"2b70982c",
  2565 => x"55597377",
  2566 => x"25f4d538",
  2567 => x"79147033",
  2568 => x"7c077009",
  2569 => x"7081ff06",
  2570 => x"70555357",
  2571 => x"5753ee93",
  2572 => x"3f7251ee",
  2573 => x"8e3f7714",
  2574 => x"982b7098",
  2575 => x"2c555976",
  2576 => x"7424ffaf",
  2577 => x"38f4a939",
  2578 => x"7d802e80",
  2579 => x"f6387914",
  2580 => x"70337c07",
  2581 => x"70525456",
  2582 => x"80557875",
  2583 => x"2e853872",
  2584 => x"842a5675",
  2585 => x"832a7081",
  2586 => x"06515372",
  2587 => x"802e8438",
  2588 => x"81c05575",
  2589 => x"822a7081",
  2590 => x"06515372",
  2591 => x"802e8538",
  2592 => x"74b00755",
  2593 => x"75812a70",
  2594 => x"81065153",
  2595 => x"72802e85",
  2596 => x"38748c07",
  2597 => x"55758106",
  2598 => x"5372802e",
  2599 => x"85387483",
  2600 => x"07557481",
  2601 => x"ff067052",
  2602 => x"56ed983f",
  2603 => x"7551ed93",
  2604 => x"3f771498",
  2605 => x"2b70982c",
  2606 => x"55537674",
  2607 => x"24ff8f38",
  2608 => x"f3ae3979",
  2609 => x"1470337c",
  2610 => x"07705354",
  2611 => x"56ecf43f",
  2612 => x"7251ecef",
  2613 => x"3f771498",
  2614 => x"2b70982c",
  2615 => x"55597377",
  2616 => x"25f38d38",
  2617 => x"79147033",
  2618 => x"7c077053",
  2619 => x"5456ecd3",
  2620 => x"3f7251ec",
  2621 => x"ce3f7714",
  2622 => x"982b7098",
  2623 => x"2c555976",
  2624 => x"7424c038",
  2625 => x"f2ea39f8",
  2626 => x"3d0d7a7d",
  2627 => x"028805af",
  2628 => x"05335a55",
  2629 => x"59807470",
  2630 => x"81055633",
  2631 => x"75585657",
  2632 => x"74772e09",
  2633 => x"81068838",
  2634 => x"76b00c8a",
  2635 => x"3d0d0474",
  2636 => x"53775278",
  2637 => x"51ef923f",
  2638 => x"b00881ff",
  2639 => x"06770570",
  2640 => x"83ffff06",
  2641 => x"77708105",
  2642 => x"59335258",
  2643 => x"5574802e",
  2644 => x"d7387453",
  2645 => x"77527851",
  2646 => x"eeef3fb0",
  2647 => x"0881ff06",
  2648 => x"77057083",
  2649 => x"ffff0677",
  2650 => x"70810559",
  2651 => x"33525855",
  2652 => x"74ffbc38",
  2653 => x"ffb239fe",
  2654 => x"3d0d0293",
  2655 => x"05335382",
  2656 => x"9eb83352",
  2657 => x"829eb408",
  2658 => x"51eebe3f",
  2659 => x"b00881ff",
  2660 => x"06b00c84",
  2661 => x"3d0d04fb",
  2662 => x"3d0d800b",
  2663 => x"81dee852",
  2664 => x"5680c283",
  2665 => x"3f755574",
  2666 => x"105381d0",
  2667 => x"5281f684",
  2668 => x"0851e6c1",
  2669 => x"3fb00887",
  2670 => x"2a708106",
  2671 => x"51547380",
  2672 => x"2e80d138",
  2673 => x"81157081",
  2674 => x"ff067098",
  2675 => x"2b525654",
  2676 => x"738025d3",
  2677 => x"3881def4",
  2678 => x"5180c1cb",
  2679 => x"3f805574",
  2680 => x"105381d0",
  2681 => x"5281f680",
  2682 => x"0851e689",
  2683 => x"3fb00887",
  2684 => x"2a708106",
  2685 => x"51547380",
  2686 => x"2e80cf38",
  2687 => x"81157081",
  2688 => x"ff067098",
  2689 => x"2b525654",
  2690 => x"738025d3",
  2691 => x"3875b00c",
  2692 => x"873d0d04",
  2693 => x"81df8051",
  2694 => x"80c18c3f",
  2695 => x"74528851",
  2696 => x"80c1a73f",
  2697 => x"81df8c51",
  2698 => x"80c0fc3f",
  2699 => x"81167083",
  2700 => x"ffff0681",
  2701 => x"177081ff",
  2702 => x"0670982b",
  2703 => x"52585257",
  2704 => x"54738025",
  2705 => x"fee138ff",
  2706 => x"8c3981df",
  2707 => x"805180c0",
  2708 => x"d63f7452",
  2709 => x"885180c0",
  2710 => x"f13f81df",
  2711 => x"8c5180c0",
  2712 => x"c63f8116",
  2713 => x"7083ffff",
  2714 => x"06811770",
  2715 => x"81ff0670",
  2716 => x"982b5258",
  2717 => x"52575473",
  2718 => x"8025fee3",
  2719 => x"38ff8e39",
  2720 => x"f33d0d7f",
  2721 => x"02840580",
  2722 => x"c3053302",
  2723 => x"880580c6",
  2724 => x"052281df",
  2725 => x"9c545b55",
  2726 => x"5880c08b",
  2727 => x"3f785180",
  2728 => x"c1cf3f81",
  2729 => x"dfa851bf",
  2730 => x"fe3f7352",
  2731 => x"885180c0",
  2732 => x"993f81ce",
  2733 => x"c851bfef",
  2734 => x"3f805776",
  2735 => x"79278191",
  2736 => x"3873108e",
  2737 => x"3d5c5a79",
  2738 => x"53819052",
  2739 => x"7751e4a5",
  2740 => x"3f76882a",
  2741 => x"53905277",
  2742 => x"51e49a3f",
  2743 => x"7681ff06",
  2744 => x"53905277",
  2745 => x"51e48e3f",
  2746 => x"811a5381",
  2747 => x"90527751",
  2748 => x"e4833f80",
  2749 => x"5380e052",
  2750 => x"7751e3f9",
  2751 => x"3fb00887",
  2752 => x"2a810654",
  2753 => x"738a3888",
  2754 => x"18087081",
  2755 => x"ff065d56",
  2756 => x"7b81ff06",
  2757 => x"81d5ac52",
  2758 => x"56bf8c3f",
  2759 => x"75528851",
  2760 => x"bfa83f81",
  2761 => x"e9e051be",
  2762 => x"fe3fe016",
  2763 => x"5480df74",
  2764 => x"27b63876",
  2765 => x"8706701c",
  2766 => x"5755a076",
  2767 => x"3474872e",
  2768 => x"b9388117",
  2769 => x"7083ffff",
  2770 => x"06585578",
  2771 => x"7726fef7",
  2772 => x"3880e00b",
  2773 => x"8c190c8c",
  2774 => x"18087081",
  2775 => x"2a810658",
  2776 => x"5a76f438",
  2777 => x"8f3d0d04",
  2778 => x"76870670",
  2779 => x"1c555575",
  2780 => x"74347487",
  2781 => x"2e098106",
  2782 => x"c9387a51",
  2783 => x"bea93f8a",
  2784 => x"51be8a3f",
  2785 => x"81177083",
  2786 => x"ffff0658",
  2787 => x"55787726",
  2788 => x"feb538ff",
  2789 => x"bc39fb3d",
  2790 => x"0d8151cc",
  2791 => x"aa3fb008",
  2792 => x"81ff0654",
  2793 => x"8251cdd2",
  2794 => x"3fb00881",
  2795 => x"ff065683",
  2796 => x"51cc943f",
  2797 => x"b00883ff",
  2798 => x"ff065573",
  2799 => x"9c3881f6",
  2800 => x"80085474",
  2801 => x"84388180",
  2802 => x"55745375",
  2803 => x"527351fd",
  2804 => x"af3f74b0",
  2805 => x"0c873d0d",
  2806 => x"0481f684",
  2807 => x"0854e439",
  2808 => x"fb3d0d77",
  2809 => x"028405a7",
  2810 => x"05330288",
  2811 => x"05a30533",
  2812 => x"70105658",
  2813 => x"56548190",
  2814 => x"527351e1",
  2815 => x"f83f7351",
  2816 => x"e2a53fb0",
  2817 => x"08802e93",
  2818 => x"38745380",
  2819 => x"d0527351",
  2820 => x"e1e33f80",
  2821 => x"0bb00c87",
  2822 => x"3d0d0481",
  2823 => x"dfc451bd",
  2824 => x"863fff0b",
  2825 => x"b00c873d",
  2826 => x"0d04fc3d",
  2827 => x"0d760284",
  2828 => x"059f0533",
  2829 => x"70108105",
  2830 => x"55565481",
  2831 => x"90527351",
  2832 => x"e1b33f73",
  2833 => x"51e1e03f",
  2834 => x"b008802e",
  2835 => x"a7388053",
  2836 => x"80e05273",
  2837 => x"51e19e3f",
  2838 => x"7351e1cb",
  2839 => x"3fb00880",
  2840 => x"2e923888",
  2841 => x"14087090",
  2842 => x"2b70902c",
  2843 => x"b00c5555",
  2844 => x"863d0d04",
  2845 => x"81dfc451",
  2846 => x"bcad3fff",
  2847 => x"0bb00c86",
  2848 => x"3d0d04fd",
  2849 => x"3d0d9c54",
  2850 => x"81dfcc51",
  2851 => x"bc993f73",
  2852 => x"528851bc",
  2853 => x"b53f7351",
  2854 => x"e1a33fb0",
  2855 => x"0881ff06",
  2856 => x"81f68408",
  2857 => x"5253e0ff",
  2858 => x"3fb00880",
  2859 => x"2eaa3881",
  2860 => x"dfdc51bb",
  2861 => x"f23f7252",
  2862 => x"8851bc8e",
  2863 => x"3f8a51bb",
  2864 => x"cc3f8114",
  2865 => x"7081ff06",
  2866 => x"555380d5",
  2867 => x"7427ffb8",
  2868 => x"3872b00c",
  2869 => x"853d0d04",
  2870 => x"81dfe451",
  2871 => x"bbc93fff",
  2872 => x"0bb00c85",
  2873 => x"3d0d04fe",
  2874 => x"3d0d8151",
  2875 => x"cb8c3fb0",
  2876 => x"0881ff06",
  2877 => x"538251cb",
  2878 => x"813fb008",
  2879 => x"81ff0652",
  2880 => x"7251e184",
  2881 => x"3f7251e0",
  2882 => x"b43fb008",
  2883 => x"81ff0681",
  2884 => x"f6840852",
  2885 => x"53e0903f",
  2886 => x"b008802e",
  2887 => x"883872b0",
  2888 => x"0c843d0d",
  2889 => x"0481dfec",
  2890 => x"51bafc3f",
  2891 => x"ff0bb00c",
  2892 => x"843d0d04",
  2893 => x"fe3d0d02",
  2894 => x"93053302",
  2895 => x"84059705",
  2896 => x"33545271",
  2897 => x"73279338",
  2898 => x"a051bac1",
  2899 => x"3f811270",
  2900 => x"81ff0651",
  2901 => x"52727226",
  2902 => x"ef38843d",
  2903 => x"0d04fe3d",
  2904 => x"0d747081",
  2905 => x"06535371",
  2906 => x"85df3872",
  2907 => x"812a7081",
  2908 => x"06515271",
  2909 => x"85bc3872",
  2910 => x"822a7081",
  2911 => x"06515271",
  2912 => x"85993872",
  2913 => x"832a7081",
  2914 => x"06515271",
  2915 => x"84f63872",
  2916 => x"842a7081",
  2917 => x"06515271",
  2918 => x"84d33872",
  2919 => x"852a7081",
  2920 => x"06515271",
  2921 => x"84b03872",
  2922 => x"862a7081",
  2923 => x"06515271",
  2924 => x"848d3872",
  2925 => x"872a7081",
  2926 => x"06515271",
  2927 => x"83ea3872",
  2928 => x"882a7081",
  2929 => x"06515271",
  2930 => x"83c73872",
  2931 => x"892a7081",
  2932 => x"06515271",
  2933 => x"83a43872",
  2934 => x"8a2a7081",
  2935 => x"06515271",
  2936 => x"83813872",
  2937 => x"8b2a7081",
  2938 => x"06515271",
  2939 => x"82de3872",
  2940 => x"8c2a7081",
  2941 => x"06515271",
  2942 => x"82bb3872",
  2943 => x"8d2a7081",
  2944 => x"06515271",
  2945 => x"82983872",
  2946 => x"8e2a7081",
  2947 => x"06515271",
  2948 => x"81f53872",
  2949 => x"8f2a7081",
  2950 => x"06515271",
  2951 => x"81d23872",
  2952 => x"902a7081",
  2953 => x"06515271",
  2954 => x"81af3872",
  2955 => x"912a7081",
  2956 => x"06515271",
  2957 => x"818c3872",
  2958 => x"922a7081",
  2959 => x"06515271",
  2960 => x"80e93872",
  2961 => x"932a7081",
  2962 => x"06515271",
  2963 => x"80c63872",
  2964 => x"942a7081",
  2965 => x"06515271",
  2966 => x"a5387295",
  2967 => x"2a708106",
  2968 => x"5152718b",
  2969 => x"38807324",
  2970 => x"83f63884",
  2971 => x"3d0d0481",
  2972 => x"dffc51b8",
  2973 => x"b23f7280",
  2974 => x"25f13883",
  2975 => x"e33981e0",
  2976 => x"9851b8a3",
  2977 => x"3f72952a",
  2978 => x"70810651",
  2979 => x"5271802e",
  2980 => x"d438dc39",
  2981 => x"81e0b451",
  2982 => x"b88d3f72",
  2983 => x"942a7081",
  2984 => x"06515271",
  2985 => x"802effb2",
  2986 => x"38d43981",
  2987 => x"e0d051b7",
  2988 => x"f63f7293",
  2989 => x"2a708106",
  2990 => x"51527180",
  2991 => x"2eff9038",
  2992 => x"d33981e0",
  2993 => x"ec51b7df",
  2994 => x"3f72922a",
  2995 => x"70810651",
  2996 => x"5271802e",
  2997 => x"feed38d3",
  2998 => x"3981e18c",
  2999 => x"51b7c83f",
  3000 => x"72912a70",
  3001 => x"81065152",
  3002 => x"71802efe",
  3003 => x"ca38d339",
  3004 => x"81e1ac51",
  3005 => x"b7b13f72",
  3006 => x"902a7081",
  3007 => x"06515271",
  3008 => x"802efea7",
  3009 => x"38d33981",
  3010 => x"e1cc51b7",
  3011 => x"9a3f728f",
  3012 => x"2a708106",
  3013 => x"51527180",
  3014 => x"2efe8438",
  3015 => x"d33981e1",
  3016 => x"ec51b783",
  3017 => x"3f728e2a",
  3018 => x"70810651",
  3019 => x"5271802e",
  3020 => x"fde138d3",
  3021 => x"3981e284",
  3022 => x"51b6ec3f",
  3023 => x"728d2a70",
  3024 => x"81065152",
  3025 => x"71802efd",
  3026 => x"be38d339",
  3027 => x"81e29851",
  3028 => x"b6d53f72",
  3029 => x"8c2a7081",
  3030 => x"06515271",
  3031 => x"802efd9b",
  3032 => x"38d33981",
  3033 => x"e2b851b6",
  3034 => x"be3f728b",
  3035 => x"2a708106",
  3036 => x"51527180",
  3037 => x"2efcf838",
  3038 => x"d33981e2",
  3039 => x"e051b6a7",
  3040 => x"3f728a2a",
  3041 => x"70810651",
  3042 => x"5271802e",
  3043 => x"fcd538d3",
  3044 => x"3981e380",
  3045 => x"51b6903f",
  3046 => x"72892a70",
  3047 => x"81065152",
  3048 => x"71802efc",
  3049 => x"b238d339",
  3050 => x"81e3a051",
  3051 => x"b5f93f72",
  3052 => x"882a7081",
  3053 => x"06515271",
  3054 => x"802efc8f",
  3055 => x"38d33981",
  3056 => x"e3c851b5",
  3057 => x"e23f7287",
  3058 => x"2a708106",
  3059 => x"51527180",
  3060 => x"2efbec38",
  3061 => x"d33981e3",
  3062 => x"e851b5cb",
  3063 => x"3f72862a",
  3064 => x"70810651",
  3065 => x"5271802e",
  3066 => x"fbc938d3",
  3067 => x"3981e488",
  3068 => x"51b5b43f",
  3069 => x"72852a70",
  3070 => x"81065152",
  3071 => x"71802efb",
  3072 => x"a638d339",
  3073 => x"81e4b051",
  3074 => x"b59d3f72",
  3075 => x"842a7081",
  3076 => x"06515271",
  3077 => x"802efb83",
  3078 => x"38d33981",
  3079 => x"e4d051b5",
  3080 => x"863f7283",
  3081 => x"2a708106",
  3082 => x"51527180",
  3083 => x"2efae038",
  3084 => x"d33981e4",
  3085 => x"f051b4ef",
  3086 => x"3f72822a",
  3087 => x"70810651",
  3088 => x"5271802e",
  3089 => x"fabd38d3",
  3090 => x"3981e598",
  3091 => x"51b4d83f",
  3092 => x"72812a70",
  3093 => x"81065152",
  3094 => x"71802efa",
  3095 => x"9a38d339",
  3096 => x"81e5b851",
  3097 => x"b4c13f84",
  3098 => x"3d0d04fd",
  3099 => x"3d0d81e5",
  3100 => x"cc51b4b3",
  3101 => x"3fffaf9b",
  3102 => x"3fb00880",
  3103 => x"2e889a38",
  3104 => x"81e5e851",
  3105 => x"b4a13f81",
  3106 => x"e5f051b4",
  3107 => x"9a3f81f6",
  3108 => x"8c088411",
  3109 => x"08709d2a",
  3110 => x"81065154",
  3111 => x"5472802e",
  3112 => x"87933881",
  3113 => x"cea451b3",
  3114 => x"fe3f81e6",
  3115 => x"8c51b3f7",
  3116 => x"3f81f5cc",
  3117 => x"0880d411",
  3118 => x"085253b5",
  3119 => x"b43f81e6",
  3120 => x"a851b3e3",
  3121 => x"3f81f5cc",
  3122 => x"0880d011",
  3123 => x"085254b5",
  3124 => x"a03f8a51",
  3125 => x"b3b73f81",
  3126 => x"e6c451b3",
  3127 => x"ca3f81e6",
  3128 => x"e851b3c3",
  3129 => x"3f81e7b0",
  3130 => x"51b3bc3f",
  3131 => x"81e7f851",
  3132 => x"b3b53f81",
  3133 => x"f5cc0870",
  3134 => x"085253b4",
  3135 => x"f43fb008",
  3136 => x"81ff0653",
  3137 => x"728c2793",
  3138 => x"38a051b3",
  3139 => x"803f8113",
  3140 => x"7081ff06",
  3141 => x"54548c73",
  3142 => x"26ef3881",
  3143 => x"f5cc0884",
  3144 => x"11085253",
  3145 => x"b4cb3fb0",
  3146 => x"0881ff06",
  3147 => x"53728c27",
  3148 => x"9338a051",
  3149 => x"b2d73f81",
  3150 => x"137081ff",
  3151 => x"0654548c",
  3152 => x"7326ef38",
  3153 => x"81f5cc08",
  3154 => x"88110852",
  3155 => x"53b4a23f",
  3156 => x"b00881ff",
  3157 => x"0653728c",
  3158 => x"279338a0",
  3159 => x"51b2ae3f",
  3160 => x"81137081",
  3161 => x"ff065454",
  3162 => x"8c7326ef",
  3163 => x"3881f5cc",
  3164 => x"088c1108",
  3165 => x"5253b3f9",
  3166 => x"3fb00881",
  3167 => x"ff065372",
  3168 => x"8c279338",
  3169 => x"a051b285",
  3170 => x"3f811370",
  3171 => x"81ff0654",
  3172 => x"548c7326",
  3173 => x"ef3881e8",
  3174 => x"9451b28b",
  3175 => x"3f81f5cc",
  3176 => x"08901108",
  3177 => x"5253b3c9",
  3178 => x"3fb00881",
  3179 => x"ff065372",
  3180 => x"8c279338",
  3181 => x"a051b1d5",
  3182 => x"3f811370",
  3183 => x"81ff0654",
  3184 => x"548c7326",
  3185 => x"ef3881f5",
  3186 => x"cc089411",
  3187 => x"085253b3",
  3188 => x"a03fb008",
  3189 => x"81ff0653",
  3190 => x"728c2793",
  3191 => x"38a051b1",
  3192 => x"ac3f8113",
  3193 => x"7081ff06",
  3194 => x"54548c73",
  3195 => x"26ef3881",
  3196 => x"f5cc0898",
  3197 => x"11085253",
  3198 => x"b2f73fb0",
  3199 => x"0881ff06",
  3200 => x"53728c27",
  3201 => x"9338a051",
  3202 => x"b1833f81",
  3203 => x"137081ff",
  3204 => x"0654548c",
  3205 => x"7326ef38",
  3206 => x"81f5cc08",
  3207 => x"9c110852",
  3208 => x"53b2ce3f",
  3209 => x"b00881ff",
  3210 => x"0653728c",
  3211 => x"279338a0",
  3212 => x"51b0da3f",
  3213 => x"81137081",
  3214 => x"ff065454",
  3215 => x"8c7326ef",
  3216 => x"3881e8b0",
  3217 => x"51b0e03f",
  3218 => x"81f5cc08",
  3219 => x"54810bb0",
  3220 => x"150cb014",
  3221 => x"08537280",
  3222 => x"25f838a0",
  3223 => x"140851b2",
  3224 => x"903fb008",
  3225 => x"81ff0653",
  3226 => x"728c2793",
  3227 => x"38a051b0",
  3228 => x"9c3f8113",
  3229 => x"7081ff06",
  3230 => x"54548c73",
  3231 => x"26ef3881",
  3232 => x"f5cc08a4",
  3233 => x"11085253",
  3234 => x"b1e73fb0",
  3235 => x"0881ff06",
  3236 => x"53728c27",
  3237 => x"9338a051",
  3238 => x"aff33f81",
  3239 => x"137081ff",
  3240 => x"0654548c",
  3241 => x"7326ef38",
  3242 => x"81f5cc08",
  3243 => x"a8110852",
  3244 => x"53b1be3f",
  3245 => x"b00881ff",
  3246 => x"0653728c",
  3247 => x"279338a0",
  3248 => x"51afca3f",
  3249 => x"81137081",
  3250 => x"ff065454",
  3251 => x"8c7326ef",
  3252 => x"3881f5cc",
  3253 => x"08ac1108",
  3254 => x"5253b195",
  3255 => x"3fb00881",
  3256 => x"ff065372",
  3257 => x"8c279338",
  3258 => x"a051afa1",
  3259 => x"3f811370",
  3260 => x"81ff0654",
  3261 => x"548c7326",
  3262 => x"ef3881e8",
  3263 => x"cc51afa7",
  3264 => x"3f81f5cc",
  3265 => x"0880e011",
  3266 => x"085254b0",
  3267 => x"e43f81e8",
  3268 => x"e451af93",
  3269 => x"3f81f5cc",
  3270 => x"0880d811",
  3271 => x"085253b0",
  3272 => x"d03f81e8",
  3273 => x"fc51aeff",
  3274 => x"3f81f5cc",
  3275 => x"08b01108",
  3276 => x"fe0a0652",
  3277 => x"54b0ba3f",
  3278 => x"81f5cc08",
  3279 => x"54800bb0",
  3280 => x"150c81e9",
  3281 => x"9451aedf",
  3282 => x"3f81e9ac",
  3283 => x"51aed83f",
  3284 => x"81f5cc08",
  3285 => x"80c01108",
  3286 => x"5253b095",
  3287 => x"3fb00881",
  3288 => x"ff065372",
  3289 => x"98279338",
  3290 => x"a051aea1",
  3291 => x"3f811370",
  3292 => x"81ff0651",
  3293 => x"53987326",
  3294 => x"ef3881f5",
  3295 => x"cc0880c8",
  3296 => x"11085254",
  3297 => x"afeb3fb0",
  3298 => x"0881ff06",
  3299 => x"53729827",
  3300 => x"9338a051",
  3301 => x"adf73f81",
  3302 => x"137081ff",
  3303 => x"06515398",
  3304 => x"7326ef38",
  3305 => x"81e9c851",
  3306 => x"adfd3f81",
  3307 => x"f5cc0880",
  3308 => x"c4110852",
  3309 => x"54afba3f",
  3310 => x"b00881ff",
  3311 => x"06537298",
  3312 => x"279338a0",
  3313 => x"51adc63f",
  3314 => x"81137081",
  3315 => x"ff065153",
  3316 => x"987326ef",
  3317 => x"3881f5cc",
  3318 => x"0880cc11",
  3319 => x"085254af",
  3320 => x"903fb008",
  3321 => x"81ff0653",
  3322 => x"72982793",
  3323 => x"38a051ad",
  3324 => x"9c3f8113",
  3325 => x"7081ff06",
  3326 => x"51539873",
  3327 => x"26ef388a",
  3328 => x"51ad8a3f",
  3329 => x"81f5cc08",
  3330 => x"b4110881",
  3331 => x"e9e45354",
  3332 => x"54ad943f",
  3333 => x"80732481",
  3334 => x"8a387251",
  3335 => x"aed33fa0",
  3336 => x"51acea3f",
  3337 => x"72862681",
  3338 => x"81387210",
  3339 => x"1081eec8",
  3340 => x"05537208",
  3341 => x"0481c6e4",
  3342 => x"51acec3f",
  3343 => x"81e68c51",
  3344 => x"ace53f81",
  3345 => x"f5cc0880",
  3346 => x"d4110852",
  3347 => x"53aea23f",
  3348 => x"81e6a851",
  3349 => x"acd13f81",
  3350 => x"f5cc0880",
  3351 => x"d0110852",
  3352 => x"54ae8e3f",
  3353 => x"8a51aca5",
  3354 => x"3f81e6c4",
  3355 => x"51acb83f",
  3356 => x"81e6e851",
  3357 => x"acb13f81",
  3358 => x"e7b051ac",
  3359 => x"aa3f81e7",
  3360 => x"f851aca3",
  3361 => x"3f81f5cc",
  3362 => x"08700852",
  3363 => x"53ade23f",
  3364 => x"b00881ff",
  3365 => x"0653f8ec",
  3366 => x"3981ce88",
  3367 => x"51ac883f",
  3368 => x"f7de3981",
  3369 => x"e9f851ab",
  3370 => x"fe3f81f5",
  3371 => x"cc08b811",
  3372 => x"0881ea84",
  3373 => x"535553ab",
  3374 => x"ee3f7352",
  3375 => x"a051ac8a",
  3376 => x"3f7351f1",
  3377 => x"993f8a51",
  3378 => x"abc33f80",
  3379 => x"0bb00c85",
  3380 => x"3d0d0481",
  3381 => x"ea9851ab",
  3382 => x"ce3fcf39",
  3383 => x"81eaa451",
  3384 => x"abc53fc6",
  3385 => x"3981eab0",
  3386 => x"51abbc3f",
  3387 => x"ffbc3981",
  3388 => x"eab451ab",
  3389 => x"b23fffb2",
  3390 => x"3981eac0",
  3391 => x"51aba83f",
  3392 => x"ffa83981",
  3393 => x"eacc51ab",
  3394 => x"9e3fff9e",
  3395 => x"3981ead8",
  3396 => x"51ab943f",
  3397 => x"ff9439fd",
  3398 => x"3d0d81ea",
  3399 => x"e451ab87",
  3400 => x"3fffa5ef",
  3401 => x"3fb00882",
  3402 => x"c63881ea",
  3403 => x"ec51aaf7",
  3404 => x"3f81f5d4",
  3405 => x"3353b352",
  3406 => x"7251d381",
  3407 => x"3f81eaf0",
  3408 => x"51aae43f",
  3409 => x"81f68c08",
  3410 => x"84110870",
  3411 => x"9d2a8106",
  3412 => x"51545472",
  3413 => x"802e81ef",
  3414 => x"3881eaf8",
  3415 => x"51aac83f",
  3416 => x"81eafc51",
  3417 => x"aac13f81",
  3418 => x"f5cc0880",
  3419 => x"d0110852",
  3420 => x"54abfe3f",
  3421 => x"81f5cc08",
  3422 => x"54810bb0",
  3423 => x"150cb014",
  3424 => x"08537280",
  3425 => x"25f83881",
  3426 => x"eb8c51aa",
  3427 => x"9a3f81f5",
  3428 => x"cc08a011",
  3429 => x"085254ab",
  3430 => x"d83f81f5",
  3431 => x"d43353b3",
  3432 => x"527251d2",
  3433 => x"983f81eb",
  3434 => x"9451a9fb",
  3435 => x"3f81f5cc",
  3436 => x"08a41108",
  3437 => x"5254abb9",
  3438 => x"3f81eb9c",
  3439 => x"51a9e83f",
  3440 => x"81f5cc08",
  3441 => x"a8110852",
  3442 => x"53aba63f",
  3443 => x"81f5d433",
  3444 => x"54b35273",
  3445 => x"51d1e63f",
  3446 => x"81eba451",
  3447 => x"a9c93f81",
  3448 => x"f5cc08ac",
  3449 => x"11085253",
  3450 => x"ab873f81",
  3451 => x"ebac51a9",
  3452 => x"b63f81f5",
  3453 => x"cc0880e0",
  3454 => x"11085254",
  3455 => x"aaf33f81",
  3456 => x"f5d43353",
  3457 => x"b3527251",
  3458 => x"d1b33f81",
  3459 => x"ebb451a9",
  3460 => x"963f81f5",
  3461 => x"cc08b011",
  3462 => x"08fe0a06",
  3463 => x"5254aad1",
  3464 => x"3f81f5cc",
  3465 => x"0854800b",
  3466 => x"b0150cb4",
  3467 => x"140881eb",
  3468 => x"bc5253a8",
  3469 => x"f23f7286",
  3470 => x"2680c238",
  3471 => x"72101081",
  3472 => x"eee40553",
  3473 => x"72080481",
  3474 => x"ebc851a8",
  3475 => x"da3f81ea",
  3476 => x"fc51a8d3",
  3477 => x"3f81f5cc",
  3478 => x"0880d011",
  3479 => x"085254aa",
  3480 => x"903f81f5",
  3481 => x"cc085481",
  3482 => x"0bb0150c",
  3483 => x"fe903981",
  3484 => x"eaf851fd",
  3485 => x"b93981ea",
  3486 => x"d851a8ab",
  3487 => x"3f81f5cc",
  3488 => x"08b81108",
  3489 => x"81ebd053",
  3490 => x"5553a89b",
  3491 => x"3f7352a0",
  3492 => x"51a8b73f",
  3493 => x"8a51a7f5",
  3494 => x"3f738106",
  3495 => x"537285df",
  3496 => x"3873812a",
  3497 => x"70810651",
  3498 => x"537285bc",
  3499 => x"3873822a",
  3500 => x"70810651",
  3501 => x"53728599",
  3502 => x"3873832a",
  3503 => x"70810651",
  3504 => x"537284f6",
  3505 => x"3873842a",
  3506 => x"70810651",
  3507 => x"537284d3",
  3508 => x"3873852a",
  3509 => x"70810651",
  3510 => x"537284b0",
  3511 => x"3873862a",
  3512 => x"70810651",
  3513 => x"5372848d",
  3514 => x"3873872a",
  3515 => x"70810651",
  3516 => x"537283ea",
  3517 => x"3873882a",
  3518 => x"70810651",
  3519 => x"537283c7",
  3520 => x"3873892a",
  3521 => x"70810651",
  3522 => x"537283a4",
  3523 => x"38738a2a",
  3524 => x"70810651",
  3525 => x"53728381",
  3526 => x"38738b2a",
  3527 => x"70810651",
  3528 => x"537282de",
  3529 => x"38738c2a",
  3530 => x"70810651",
  3531 => x"537282bb",
  3532 => x"38738d2a",
  3533 => x"70810651",
  3534 => x"53728298",
  3535 => x"38738e2a",
  3536 => x"70810651",
  3537 => x"537281f5",
  3538 => x"38738f2a",
  3539 => x"70810651",
  3540 => x"537281d2",
  3541 => x"3873902a",
  3542 => x"70810651",
  3543 => x"537281af",
  3544 => x"3873912a",
  3545 => x"70810651",
  3546 => x"5372818c",
  3547 => x"3873922a",
  3548 => x"70810651",
  3549 => x"537280e9",
  3550 => x"3873932a",
  3551 => x"70810651",
  3552 => x"537280c6",
  3553 => x"3873942a",
  3554 => x"70810651",
  3555 => x"5372a538",
  3556 => x"73952a70",
  3557 => x"81065153",
  3558 => x"728b3880",
  3559 => x"742483f6",
  3560 => x"38853d0d",
  3561 => x"0481ebe0",
  3562 => x"51a5fc3f",
  3563 => x"738025f1",
  3564 => x"3883e339",
  3565 => x"81ebf051",
  3566 => x"a5ed3f73",
  3567 => x"952a7081",
  3568 => x"06515372",
  3569 => x"802ed438",
  3570 => x"dc3981ec",
  3571 => x"8051a5d7",
  3572 => x"3f73942a",
  3573 => x"70810651",
  3574 => x"5372802e",
  3575 => x"ffb238d4",
  3576 => x"3981ec90",
  3577 => x"51a5c03f",
  3578 => x"73932a70",
  3579 => x"81065153",
  3580 => x"72802eff",
  3581 => x"9038d339",
  3582 => x"81eca051",
  3583 => x"a5a93f73",
  3584 => x"922a7081",
  3585 => x"06515372",
  3586 => x"802efeed",
  3587 => x"38d33981",
  3588 => x"ecb051a5",
  3589 => x"923f7391",
  3590 => x"2a708106",
  3591 => x"51537280",
  3592 => x"2efeca38",
  3593 => x"d33981ec",
  3594 => x"c051a4fb",
  3595 => x"3f73902a",
  3596 => x"70810651",
  3597 => x"5372802e",
  3598 => x"fea738d3",
  3599 => x"3981ecd0",
  3600 => x"51a4e43f",
  3601 => x"738f2a70",
  3602 => x"81065153",
  3603 => x"72802efe",
  3604 => x"8438d339",
  3605 => x"81ece051",
  3606 => x"a4cd3f73",
  3607 => x"8e2a7081",
  3608 => x"06515372",
  3609 => x"802efde1",
  3610 => x"38d33981",
  3611 => x"ecf051a4",
  3612 => x"b63f738d",
  3613 => x"2a708106",
  3614 => x"51537280",
  3615 => x"2efdbe38",
  3616 => x"d33981ec",
  3617 => x"fc51a49f",
  3618 => x"3f738c2a",
  3619 => x"70810651",
  3620 => x"5372802e",
  3621 => x"fd9b38d3",
  3622 => x"3981ed8c",
  3623 => x"51a4883f",
  3624 => x"738b2a70",
  3625 => x"81065153",
  3626 => x"72802efc",
  3627 => x"f838d339",
  3628 => x"81ed9c51",
  3629 => x"a3f13f73",
  3630 => x"8a2a7081",
  3631 => x"06515372",
  3632 => x"802efcd5",
  3633 => x"38d33981",
  3634 => x"edac51a3",
  3635 => x"da3f7389",
  3636 => x"2a708106",
  3637 => x"51537280",
  3638 => x"2efcb238",
  3639 => x"d33981ed",
  3640 => x"bc51a3c3",
  3641 => x"3f73882a",
  3642 => x"70810651",
  3643 => x"5372802e",
  3644 => x"fc8f38d3",
  3645 => x"3981edcc",
  3646 => x"51a3ac3f",
  3647 => x"73872a70",
  3648 => x"81065153",
  3649 => x"72802efb",
  3650 => x"ec38d339",
  3651 => x"81eddc51",
  3652 => x"a3953f73",
  3653 => x"862a7081",
  3654 => x"06515372",
  3655 => x"802efbc9",
  3656 => x"38d33981",
  3657 => x"edec51a2",
  3658 => x"fe3f7385",
  3659 => x"2a708106",
  3660 => x"51537280",
  3661 => x"2efba638",
  3662 => x"d33981ed",
  3663 => x"fc51a2e7",
  3664 => x"3f73842a",
  3665 => x"70810651",
  3666 => x"5372802e",
  3667 => x"fb8338d3",
  3668 => x"3981ee8c",
  3669 => x"51a2d03f",
  3670 => x"73832a70",
  3671 => x"81065153",
  3672 => x"72802efa",
  3673 => x"e038d339",
  3674 => x"81ee9c51",
  3675 => x"a2b93f73",
  3676 => x"822a7081",
  3677 => x"06515372",
  3678 => x"802efabd",
  3679 => x"38d33981",
  3680 => x"eeac51a2",
  3681 => x"a23f7381",
  3682 => x"2a708106",
  3683 => x"51537280",
  3684 => x"2efa9a38",
  3685 => x"d33981ee",
  3686 => x"bc51a28b",
  3687 => x"3f853d0d",
  3688 => x"0481ea98",
  3689 => x"51a2803f",
  3690 => x"f9d33981",
  3691 => x"eaa451a1",
  3692 => x"f63ff9c9",
  3693 => x"3981eab0",
  3694 => x"51a1ec3f",
  3695 => x"f9bf3981",
  3696 => x"eab451a1",
  3697 => x"e23ff9b5",
  3698 => x"3981eac0",
  3699 => x"51a1d83f",
  3700 => x"f9ab3981",
  3701 => x"eacc51a1",
  3702 => x"ce3ff9a1",
  3703 => x"39fe3d0d",
  3704 => x"cafe3f80",
  3705 => x"5281d684",
  3706 => x"51cdc83f",
  3707 => x"829ebc08",
  3708 => x"80d2f70b",
  3709 => x"829ebc0c",
  3710 => x"53f69c3f",
  3711 => x"72829ebc",
  3712 => x"0c843d0d",
  3713 => x"04fd3d0d",
  3714 => x"8151ffaf",
  3715 => x"ba3fb008",
  3716 => x"81ff0654",
  3717 => x"8251ffaf",
  3718 => x"ae3fb008",
  3719 => x"9f2b7407",
  3720 => x"81f5cc08",
  3721 => x"53b4130c",
  3722 => x"73b00c85",
  3723 => x"3d0d04fd",
  3724 => x"3d0d81ef",
  3725 => x"f851a0ef",
  3726 => x"3f81f5c8",
  3727 => x"08841108",
  3728 => x"5254a2ad",
  3729 => x"3f81f088",
  3730 => x"51a0dc3f",
  3731 => x"81f5c808",
  3732 => x"88110852",
  3733 => x"53a29a3f",
  3734 => x"81f09851",
  3735 => x"a0c93f81",
  3736 => x"f5c8088c",
  3737 => x"11085254",
  3738 => x"a2873f81",
  3739 => x"f0a851a0",
  3740 => x"b63f81f5",
  3741 => x"c8089011",
  3742 => x"085253a1",
  3743 => x"f43f81f0",
  3744 => x"b851a0a3",
  3745 => x"3f81f5c8",
  3746 => x"08941108",
  3747 => x"5254a1e1",
  3748 => x"3f81f5c8",
  3749 => x"08700881",
  3750 => x"f0c85355",
  3751 => x"53a0883f",
  3752 => x"73528851",
  3753 => x"a0a43f73",
  3754 => x"81065372",
  3755 => x"802e80c2",
  3756 => x"3881ef80",
  3757 => x"519ff03f",
  3758 => x"73812a70",
  3759 => x"81065153",
  3760 => x"72818738",
  3761 => x"73822a70",
  3762 => x"81065153",
  3763 => x"7280e438",
  3764 => x"73832a70",
  3765 => x"81065153",
  3766 => x"7280c338",
  3767 => x"73842a81",
  3768 => x"065473a6",
  3769 => x"388a519f",
  3770 => x"a43f800b",
  3771 => x"b00c853d",
  3772 => x"0d0481ef",
  3773 => x"90519faf",
  3774 => x"3f73812a",
  3775 => x"70810651",
  3776 => x"5372802e",
  3777 => x"ffbe3880",
  3778 => x"c13981ef",
  3779 => x"a4519f97",
  3780 => x"3f8a519e",
  3781 => x"f83f800b",
  3782 => x"b00c853d",
  3783 => x"0d0481ef",
  3784 => x"bc519f83",
  3785 => x"3f73842a",
  3786 => x"81065473",
  3787 => x"802effb5",
  3788 => x"38d83981",
  3789 => x"efd8519e",
  3790 => x"ee3f7383",
  3791 => x"2a708106",
  3792 => x"51537280",
  3793 => x"2eff9538",
  3794 => x"d53981ef",
  3795 => x"ec519ed7",
  3796 => x"3f73822a",
  3797 => x"70810651",
  3798 => x"5372802e",
  3799 => x"fef238d3",
  3800 => x"39ff3d0d",
  3801 => x"8151ffac",
  3802 => x"de3f81f5",
  3803 => x"c808b008",
  3804 => x"90120c52",
  3805 => x"8251ffac",
  3806 => x"ce3f81f5",
  3807 => x"c808b008",
  3808 => x"94120c52",
  3809 => x"800bb00c",
  3810 => x"833d0d04",
  3811 => x"ff3d0d81",
  3812 => x"f5c80870",
  3813 => x"08535180",
  3814 => x"710c71b0",
  3815 => x"0c833d0d",
  3816 => x"04f93d0d",
  3817 => x"02a60522",
  3818 => x"81f5d833",
  3819 => x"81f70655",
  3820 => x"567381f5",
  3821 => x"d8347353",
  3822 => x"a05281f6",
  3823 => x"800851e0",
  3824 => x"9f3f8057",
  3825 => x"8f5581f5",
  3826 => x"d83381fe",
  3827 => x"06547381",
  3828 => x"f5d83473",
  3829 => x"53a05281",
  3830 => x"f6800851",
  3831 => x"e0823f75",
  3832 => x"752c8106",
  3833 => x"5877802e",
  3834 => x"819e3881",
  3835 => x"f5d83382",
  3836 => x"07547381",
  3837 => x"f5d83473",
  3838 => x"53a05281",
  3839 => x"f6800851",
  3840 => x"dfde3fa0",
  3841 => x"5281f680",
  3842 => x"0851e09e",
  3843 => x"3fb00882",
  3844 => x"2a810654",
  3845 => x"73802e8d",
  3846 => x"3881752b",
  3847 => x"77077083",
  3848 => x"ffff0658",
  3849 => x"5481f5d8",
  3850 => x"33810754",
  3851 => x"7381f5d8",
  3852 => x"347353a0",
  3853 => x"5281f680",
  3854 => x"0851dfa4",
  3855 => x"3f748180",
  3856 => x"0a2981ff",
  3857 => x"0a057098",
  3858 => x"2c565874",
  3859 => x"8025fef6",
  3860 => x"3881f5d8",
  3861 => x"33820754",
  3862 => x"7381f5d8",
  3863 => x"347353a0",
  3864 => x"5281f680",
  3865 => x"0851def8",
  3866 => x"3f81f5d8",
  3867 => x"33880756",
  3868 => x"7581f5d8",
  3869 => x"347553a0",
  3870 => x"5281f680",
  3871 => x"0851dee0",
  3872 => x"3f76b00c",
  3873 => x"893d0d04",
  3874 => x"81f5d833",
  3875 => x"81fd0654",
  3876 => x"fee039fb",
  3877 => x"3d0d029f",
  3878 => x"05335680",
  3879 => x"c05381d0",
  3880 => x"5281f680",
  3881 => x"0851c0cd",
  3882 => x"3fb00887",
  3883 => x"2a810655",
  3884 => x"ff5474a5",
  3885 => x"38818051",
  3886 => x"fde73f82",
  3887 => x"8051fde1",
  3888 => x"3f848351",
  3889 => x"fddb3f86",
  3890 => x"f151fdd5",
  3891 => x"3f75832b",
  3892 => x"88830751",
  3893 => x"fdcb3f74",
  3894 => x"5473b00c",
  3895 => x"873d0d04",
  3896 => x"fc3d0d81",
  3897 => x"51ffa9df",
  3898 => x"3fb00881",
  3899 => x"ff065580",
  3900 => x"c05381d0",
  3901 => x"5281f680",
  3902 => x"0851ffbf",
  3903 => x"f83fb008",
  3904 => x"872a7081",
  3905 => x"06515473",
  3906 => x"802e8838",
  3907 => x"74b00c86",
  3908 => x"3d0d0481",
  3909 => x"8051fd89",
  3910 => x"3f828051",
  3911 => x"fd833f84",
  3912 => x"8351fcfd",
  3913 => x"3f86f151",
  3914 => x"fcf73f74",
  3915 => x"832b8883",
  3916 => x"0751fced",
  3917 => x"3f74b00c",
  3918 => x"863d0d04",
  3919 => x"803d0d81",
  3920 => x"51ffaab6",
  3921 => x"3fb00883",
  3922 => x"ffff0651",
  3923 => x"fcd33fb0",
  3924 => x"0883ffff",
  3925 => x"06b00c82",
  3926 => x"3d0d0480",
  3927 => x"0b829dd8",
  3928 => x"34800bb0",
  3929 => x"0c04fb3d",
  3930 => x"0d8151ff",
  3931 => x"aa8c3fb0",
  3932 => x"08538251",
  3933 => x"ffaa833f",
  3934 => x"b00856b0",
  3935 => x"08833890",
  3936 => x"5672fc06",
  3937 => x"5575812e",
  3938 => x"80f13880",
  3939 => x"54737627",
  3940 => x"aa387383",
  3941 => x"06537280",
  3942 => x"2eae3881",
  3943 => x"d5ac519a",
  3944 => x"863f7470",
  3945 => x"84055608",
  3946 => x"52a0519a",
  3947 => x"9d3fa051",
  3948 => x"99db3f81",
  3949 => x"14547574",
  3950 => x"26d8388a",
  3951 => x"5199ce3f",
  3952 => x"800bb00c",
  3953 => x"873d0d04",
  3954 => x"81f0dc51",
  3955 => x"99d93f74",
  3956 => x"52a05199",
  3957 => x"f53f81f1",
  3958 => x"fc5199cb",
  3959 => x"3f81d5ac",
  3960 => x"5199c43f",
  3961 => x"74708405",
  3962 => x"560852a0",
  3963 => x"5199db3f",
  3964 => x"a0519999",
  3965 => x"3f811454",
  3966 => x"ffbc3981",
  3967 => x"d5ac5199",
  3968 => x"a63f7408",
  3969 => x"52a05199",
  3970 => x"c13f8a51",
  3971 => x"98ff3f80",
  3972 => x"0bb00c87",
  3973 => x"3d0d04fc",
  3974 => x"3d0d8151",
  3975 => x"ffa8db3f",
  3976 => x"b0085282",
  3977 => x"51ffa79f",
  3978 => x"3fb00881",
  3979 => x"ff067256",
  3980 => x"53835472",
  3981 => x"802ea238",
  3982 => x"7351ffa8",
  3983 => x"bd3f8114",
  3984 => x"7081ff06",
  3985 => x"ff157081",
  3986 => x"ff06b008",
  3987 => x"79708405",
  3988 => x"5b0c5652",
  3989 => x"555272e0",
  3990 => x"3872b00c",
  3991 => x"863d0d04",
  3992 => x"803d0d8c",
  3993 => x"5198a63f",
  3994 => x"800bb00c",
  3995 => x"823d0d04",
  3996 => x"803d0d81",
  3997 => x"f6980851",
  3998 => x"f8bb9586",
  3999 => x"a1710c81",
  4000 => x"0bb00c82",
  4001 => x"3d0d0480",
  4002 => x"3d0d8151",
  4003 => x"ffa6b83f",
  4004 => x"b00881ff",
  4005 => x"0651ffb8",
  4006 => x"ec3f800b",
  4007 => x"b00c823d",
  4008 => x"0d04fa3d",
  4009 => x"0d880a57",
  4010 => x"840a5681",
  4011 => x"51ffa697",
  4012 => x"3fb00883",
  4013 => x"ffff0654",
  4014 => x"73833890",
  4015 => x"54805574",
  4016 => x"742780e7",
  4017 => x"38757084",
  4018 => x"05570870",
  4019 => x"902c5253",
  4020 => x"999f3f8a",
  4021 => x"52b00851",
  4022 => x"dcda3f72",
  4023 => x"902b7090",
  4024 => x"2c525399",
  4025 => x"8c3f8a52",
  4026 => x"b00851dc",
  4027 => x"c73f7670",
  4028 => x"84055808",
  4029 => x"70902c52",
  4030 => x"5398f63f",
  4031 => x"8a52b008",
  4032 => x"51dcb13f",
  4033 => x"72902b70",
  4034 => x"902c5253",
  4035 => x"98e33f8a",
  4036 => x"52b00851",
  4037 => x"dc9e3f8a",
  4038 => x"5196f23f",
  4039 => x"81157083",
  4040 => x"ffff0656",
  4041 => x"53737526",
  4042 => x"ff9b3873",
  4043 => x"b00c883d",
  4044 => x"0d04fd3d",
  4045 => x"0d81f5e0",
  4046 => x"088c1108",
  4047 => x"70822b83",
  4048 => x"fffc0681",
  4049 => x"f0e05451",
  4050 => x"545496db",
  4051 => x"3f725288",
  4052 => x"0a51ffab",
  4053 => x"c43fb008",
  4054 => x"54b008fe",
  4055 => x"2ea838b0",
  4056 => x"08ff2e94",
  4057 => x"38725198",
  4058 => x"883f81f0",
  4059 => x"f45196b7",
  4060 => x"3f73b00c",
  4061 => x"853d0d04",
  4062 => x"81f18851",
  4063 => x"96a93f73",
  4064 => x"b00c853d",
  4065 => x"0d0481f1",
  4066 => x"9051969b",
  4067 => x"3f73b00c",
  4068 => x"853d0d04",
  4069 => x"fc3d0d81",
  4070 => x"f5e0088c",
  4071 => x"11087082",
  4072 => x"2b83fffc",
  4073 => x"0681f19c",
  4074 => x"54515555",
  4075 => x"95f93f81",
  4076 => x"f6940888",
  4077 => x"11087080",
  4078 => x"c0078813",
  4079 => x"0c545573",
  4080 => x"52880a51",
  4081 => x"ffade43f",
  4082 => x"b00881f6",
  4083 => x"94088811",
  4084 => x"0870ffbf",
  4085 => x"0688130c",
  4086 => x"555555b0",
  4087 => x"08fe2e80",
  4088 => x"c538b008",
  4089 => x"fe249a38",
  4090 => x"b008fd2e",
  4091 => x"ab387451",
  4092 => x"96ff3f81",
  4093 => x"f1b05195",
  4094 => x"ae3f74b0",
  4095 => x"0c863d0d",
  4096 => x"04b008ff",
  4097 => x"2e098106",
  4098 => x"e53881f1",
  4099 => x"88519597",
  4100 => x"3f74b00c",
  4101 => x"863d0d04",
  4102 => x"81f1c451",
  4103 => x"95893f74",
  4104 => x"b00c863d",
  4105 => x"0d0481f1",
  4106 => x"d45194fb",
  4107 => x"3f74b00c",
  4108 => x"863d0d04",
  4109 => x"fe3d0d88",
  4110 => x"0a53840a",
  4111 => x"0b81f5e0",
  4112 => x"088c1108",
  4113 => x"51525280",
  4114 => x"71279538",
  4115 => x"80737084",
  4116 => x"05550c80",
  4117 => x"72708405",
  4118 => x"540cff11",
  4119 => x"5170ed38",
  4120 => x"800bb00c",
  4121 => x"843d0d04",
  4122 => x"fd3d0d81",
  4123 => x"51ffa2d7",
  4124 => x"3fb00881",
  4125 => x"ff065473",
  4126 => x"802ea438",
  4127 => x"73842690",
  4128 => x"3881f5e0",
  4129 => x"0874710c",
  4130 => x"5373b00c",
  4131 => x"853d0d04",
  4132 => x"81f5e008",
  4133 => x"5380730c",
  4134 => x"73b00c85",
  4135 => x"3d0d0481",
  4136 => x"f1e05194",
  4137 => x"823f81f1",
  4138 => x"f05193fb",
  4139 => x"3f81f5e0",
  4140 => x"08700852",
  4141 => x"5395ba3f",
  4142 => x"81f28051",
  4143 => x"93e93f81",
  4144 => x"f5e00884",
  4145 => x"11085353",
  4146 => x"a05193fe",
  4147 => x"3f81f294",
  4148 => x"5193d43f",
  4149 => x"81f5e008",
  4150 => x"88110853",
  4151 => x"53a05193",
  4152 => x"e93f81f2",
  4153 => x"a85193bf",
  4154 => x"3f81f5e0",
  4155 => x"088c1108",
  4156 => x"525394fd",
  4157 => x"3f8a5193",
  4158 => x"943f73b0",
  4159 => x"0c853d0d",
  4160 => x"04bc0802",
  4161 => x"bc0cf93d",
  4162 => x"0d02bc08",
  4163 => x"fc050c88",
  4164 => x"0a0bbc08",
  4165 => x"f4050cfc",
  4166 => x"3d0d823d",
  4167 => x"bc08f005",
  4168 => x"0c8151ff",
  4169 => x"a1a13fb0",
  4170 => x"0881ff06",
  4171 => x"bc08f805",
  4172 => x"0c8251ff",
  4173 => x"a1913fb0",
  4174 => x"08bc08f0",
  4175 => x"05082383",
  4176 => x"51ffa183",
  4177 => x"3fb008bc",
  4178 => x"08f00508",
  4179 => x"82052384",
  4180 => x"51ffa0f3",
  4181 => x"3fb008bc",
  4182 => x"08f00508",
  4183 => x"84052385",
  4184 => x"51ffa0e3",
  4185 => x"3fb008bc",
  4186 => x"08f00508",
  4187 => x"86052386",
  4188 => x"51ffa0d3",
  4189 => x"3fb008bc",
  4190 => x"08f00508",
  4191 => x"88052387",
  4192 => x"51ffa0c3",
  4193 => x"3fb008bc",
  4194 => x"08f00508",
  4195 => x"8a052388",
  4196 => x"51ffa0b3",
  4197 => x"3fb008bc",
  4198 => x"08f00508",
  4199 => x"8c052389",
  4200 => x"51ffa0a3",
  4201 => x"3fb008bc",
  4202 => x"08f00508",
  4203 => x"8e052380",
  4204 => x"0b81f5e0",
  4205 => x"08708c05",
  4206 => x"0851bc08",
  4207 => x"e4050cbc",
  4208 => x"08ec050c",
  4209 => x"bc08ec05",
  4210 => x"08bc08e4",
  4211 => x"05082781",
  4212 => x"8f38bc08",
  4213 => x"e40508bc",
  4214 => x"08e8050c",
  4215 => x"bc08f805",
  4216 => x"08802e81",
  4217 => x"b638bc08",
  4218 => x"ec050810",
  4219 => x"bc08f005",
  4220 => x"08057022",
  4221 => x"bc08f405",
  4222 => x"08820522",
  4223 => x"71902b07",
  4224 => x"bc08f405",
  4225 => x"080cbc08",
  4226 => x"e4050cbc",
  4227 => x"08f8050c",
  4228 => x"bc08ec05",
  4229 => x"08810570",
  4230 => x"81ff06bc",
  4231 => x"08e4050c",
  4232 => x"bc08f805",
  4233 => x"0c860bbc",
  4234 => x"08ec0508",
  4235 => x"27883880",
  4236 => x"0bbc08e4",
  4237 => x"050cbc08",
  4238 => x"e40508bc",
  4239 => x"08f40508",
  4240 => x"8405bc08",
  4241 => x"e80508ff",
  4242 => x"05bc08e8",
  4243 => x"050cbc08",
  4244 => x"f4050cbc",
  4245 => x"08ec050c",
  4246 => x"bc08e805",
  4247 => x"08ff8738",
  4248 => x"bc08fc05",
  4249 => x"080d800b",
  4250 => x"b00c893d",
  4251 => x"0dbc0c04",
  4252 => x"bc08e405",
  4253 => x"08bc08f4",
  4254 => x"05088405",
  4255 => x"bc08e805",
  4256 => x"08ff05bc",
  4257 => x"08e8050c",
  4258 => x"bc08f405",
  4259 => x"0cbc08ec",
  4260 => x"050cbc08",
  4261 => x"e8050880",
  4262 => x"2ec638bc",
  4263 => x"08ec0508",
  4264 => x"10bc08f0",
  4265 => x"05080570",
  4266 => x"2270902b",
  4267 => x"bc08f405",
  4268 => x"0808fc80",
  4269 => x"80067190",
  4270 => x"2c07bc08",
  4271 => x"f405080c",
  4272 => x"52bc08e4",
  4273 => x"050cbc08",
  4274 => x"f8050c80",
  4275 => x"0bbc08e4",
  4276 => x"050cbc08",
  4277 => x"ec050886",
  4278 => x"26ff9538",
  4279 => x"bc08ec05",
  4280 => x"08810570",
  4281 => x"81ff06bc",
  4282 => x"08f40508",
  4283 => x"8405bc08",
  4284 => x"e80508ff",
  4285 => x"05bc08e8",
  4286 => x"050cbc08",
  4287 => x"f4050cbc",
  4288 => x"08ec050c",
  4289 => x"bc08e405",
  4290 => x"0cbc08e8",
  4291 => x"0508ff8b",
  4292 => x"38fecd39",
  4293 => x"f93d0d81",
  4294 => x"51ff9dab",
  4295 => x"3fb00881",
  4296 => x"ff0681f2",
  4297 => x"b852578e",
  4298 => x"fe3f81f2",
  4299 => x"cc518ef7",
  4300 => x"3ff88080",
  4301 => x"9a805480",
  4302 => x"55737084",
  4303 => x"05550874",
  4304 => x"70840556",
  4305 => x"08545672",
  4306 => x"a0388115",
  4307 => x"7081ff06",
  4308 => x"56538775",
  4309 => x"27e33876",
  4310 => x"812e80c3",
  4311 => x"388a518e",
  4312 => x"ac3f76b0",
  4313 => x"0c893d0d",
  4314 => x"048a518e",
  4315 => x"a03f7251",
  4316 => x"8fff3f8c",
  4317 => x"52b00851",
  4318 => x"d3ba3f81",
  4319 => x"f2e4518e",
  4320 => x"a63f7552",
  4321 => x"a0518ec2",
  4322 => x"3f7551d3",
  4323 => x"d13f8115",
  4324 => x"7081ff06",
  4325 => x"56538775",
  4326 => x"27ff9e38",
  4327 => x"ffb939f8",
  4328 => x"80809a80",
  4329 => x"54805380",
  4330 => x"74708405",
  4331 => x"560c8074",
  4332 => x"70840556",
  4333 => x"0c811370",
  4334 => x"81ff0654",
  4335 => x"55728726",
  4336 => x"ff9b3880",
  4337 => x"74708405",
  4338 => x"560c8074",
  4339 => x"70840556",
  4340 => x"0c811370",
  4341 => x"81ff0654",
  4342 => x"55877327",
  4343 => x"ca38fefd",
  4344 => x"39fb3d0d",
  4345 => x"029f0533",
  4346 => x"79982b70",
  4347 => x"982c5154",
  4348 => x"55810a54",
  4349 => x"805672e8",
  4350 => x"25bd38e8",
  4351 => x"53751081",
  4352 => x"07738180",
  4353 => x"0a298180",
  4354 => x"0a057098",
  4355 => x"2c515456",
  4356 => x"807324e9",
  4357 => x"38807325",
  4358 => x"80c73873",
  4359 => x"812a810a",
  4360 => x"07738180",
  4361 => x"0a2981ff",
  4362 => x"0a057098",
  4363 => x"2c515454",
  4364 => x"728024e7",
  4365 => x"38ab3997",
  4366 => x"73259a38",
  4367 => x"9774812a",
  4368 => x"810a0771",
  4369 => x"81800a29",
  4370 => x"81ff0a05",
  4371 => x"70982c51",
  4372 => x"525553dc",
  4373 => x"39807324",
  4374 => x"ffa33872",
  4375 => x"8024ffbb",
  4376 => x"38745280",
  4377 => x"51ffb4d5",
  4378 => x"3f7381ff",
  4379 => x"0651ffb5",
  4380 => x"d23f7452",
  4381 => x"8151ffb4",
  4382 => x"c43f7388",
  4383 => x"2a7081ff",
  4384 => x"065253ff",
  4385 => x"b5bd3f74",
  4386 => x"528251ff",
  4387 => x"b4af3f73",
  4388 => x"902a7081",
  4389 => x"ff065253",
  4390 => x"ffb5a83f",
  4391 => x"74528351",
  4392 => x"ffb49a3f",
  4393 => x"73982a51",
  4394 => x"ffb5983f",
  4395 => x"74528451",
  4396 => x"ffb48a3f",
  4397 => x"7581ff06",
  4398 => x"51ffb587",
  4399 => x"3f745285",
  4400 => x"51ffb3f9",
  4401 => x"3f75882a",
  4402 => x"7081ff06",
  4403 => x"5253ffb4",
  4404 => x"f23f7452",
  4405 => x"8651ffb3",
  4406 => x"e43f7590",
  4407 => x"2a7081ff",
  4408 => x"065254ff",
  4409 => x"b4dd3f74",
  4410 => x"528751ff",
  4411 => x"b3cf3f75",
  4412 => x"982a51ff",
  4413 => x"b4cd3f87",
  4414 => x"3d0d04f2",
  4415 => x"3d0d0280",
  4416 => x"c3053302",
  4417 => x"840580c7",
  4418 => x"05338180",
  4419 => x"0a712b98",
  4420 => x"2a81f5e0",
  4421 => x"088c1108",
  4422 => x"71084453",
  4423 => x"565c5557",
  4424 => x"80730c80",
  4425 => x"7071725c",
  4426 => x"5a5e5b80",
  4427 => x"56757a27",
  4428 => x"80d73881",
  4429 => x"772783cb",
  4430 => x"387783ff",
  4431 => x"ff068119",
  4432 => x"71101084",
  4433 => x"0a057930",
  4434 => x"7a823270",
  4435 => x"30728025",
  4436 => x"71802507",
  4437 => x"56585841",
  4438 => x"57595c7b",
  4439 => x"802e83d2",
  4440 => x"38821522",
  4441 => x"5372902b",
  4442 => x"70902c54",
  4443 => x"55727b25",
  4444 => x"8338725b",
  4445 => x"7c732583",
  4446 => x"38725d81",
  4447 => x"167081ff",
  4448 => x"06575e79",
  4449 => x"7626ffb1",
  4450 => x"38811970",
  4451 => x"81ff065a",
  4452 => x"5680e579",
  4453 => x"27ff9438",
  4454 => x"987d3590",
  4455 => x"2b70902c",
  4456 => x"7c309871",
  4457 => x"35902b70",
  4458 => x"902c5c5c",
  4459 => x"55565477",
  4460 => x"54777525",
  4461 => x"83387454",
  4462 => x"73902b70",
  4463 => x"902c5d55",
  4464 => x"7b54807c",
  4465 => x"2583d438",
  4466 => x"73902b70",
  4467 => x"902c5f56",
  4468 => x"80705d58",
  4469 => x"80705a56",
  4470 => x"757a2780",
  4471 => x"e4388177",
  4472 => x"27838938",
  4473 => x"7783ffff",
  4474 => x"06811971",
  4475 => x"1010840a",
  4476 => x"0579307a",
  4477 => x"82327030",
  4478 => x"72802571",
  4479 => x"80250753",
  4480 => x"51575357",
  4481 => x"59547380",
  4482 => x"2e83a138",
  4483 => x"82152254",
  4484 => x"73902b70",
  4485 => x"902c719f",
  4486 => x"2c707232",
  4487 => x"7131799f",
  4488 => x"2c707b32",
  4489 => x"71315154",
  4490 => x"51565653",
  4491 => x"72742583",
  4492 => x"38745681",
  4493 => x"197081ff",
  4494 => x"065a5579",
  4495 => x"7926ffa4",
  4496 => x"387d7635",
  4497 => x"982b7098",
  4498 => x"2c53547b",
  4499 => x"51fb923f",
  4500 => x"811c7081",
  4501 => x"ff065d59",
  4502 => x"80e57c27",
  4503 => x"fef63881",
  4504 => x"f5e0087f",
  4505 => x"710c5880",
  4506 => x"5281d684",
  4507 => x"51ffb4c3",
  4508 => x"3f829ebc",
  4509 => x"0880d2f7",
  4510 => x"0b829ebc",
  4511 => x"0c5f8052",
  4512 => x"8051ffb0",
  4513 => x"b83f81f2",
  4514 => x"ec51889b",
  4515 => x"3f7c5189",
  4516 => x"e03f8052",
  4517 => x"8751ffb0",
  4518 => x"a43f81f2",
  4519 => x"f4518887",
  4520 => x"3f7a5189",
  4521 => x"cc3f80d2",
  4522 => x"528051ff",
  4523 => x"b08f3f81",
  4524 => x"f2fc5187",
  4525 => x"f23f7651",
  4526 => x"89b73f80",
  4527 => x"c0528751",
  4528 => x"ffaffa3f",
  4529 => x"81f38451",
  4530 => x"87dd3f79",
  4531 => x"80e62951",
  4532 => x"899f3f7e",
  4533 => x"829ebc0c",
  4534 => x"903d0d04",
  4535 => x"74225372",
  4536 => x"902b7090",
  4537 => x"2c545c72",
  4538 => x"7b258338",
  4539 => x"725b7c73",
  4540 => x"25833872",
  4541 => x"5d811670",
  4542 => x"81ff0657",
  4543 => x"5e757a27",
  4544 => x"fd873877",
  4545 => x"83ffff06",
  4546 => x"81197110",
  4547 => x"10880a05",
  4548 => x"79307a82",
  4549 => x"32703072",
  4550 => x"80257180",
  4551 => x"25075658",
  4552 => x"40415759",
  4553 => x"5473802e",
  4554 => x"ffb23882",
  4555 => x"152253ff",
  4556 => x"ae397422",
  4557 => x"53fcae39",
  4558 => x"74225473",
  4559 => x"902b7090",
  4560 => x"2c719f2c",
  4561 => x"70723271",
  4562 => x"31799f2c",
  4563 => x"707b3271",
  4564 => x"31515451",
  4565 => x"56565372",
  4566 => x"74258338",
  4567 => x"74568119",
  4568 => x"7081ff06",
  4569 => x"5a55787a",
  4570 => x"27fdd638",
  4571 => x"7783ffff",
  4572 => x"06811971",
  4573 => x"1010880a",
  4574 => x"0579307a",
  4575 => x"82327030",
  4576 => x"72802571",
  4577 => x"80250753",
  4578 => x"51575357",
  4579 => x"59547380",
  4580 => x"2effa538",
  4581 => x"82152254",
  4582 => x"ffa13981",
  4583 => x"70902b70",
  4584 => x"902c4057",
  4585 => x"5480705d",
  4586 => x"58fca939",
  4587 => x"742254fc",
  4588 => x"df39fe3d",
  4589 => x"0d8151ff",
  4590 => x"948d3fb0",
  4591 => x"0881ff06",
  4592 => x"538251ff",
  4593 => x"94813fb0",
  4594 => x"0881ff06",
  4595 => x"527251fa",
  4596 => x"aa3f800b",
  4597 => x"b00c843d",
  4598 => x"0d04fd3d",
  4599 => x"0d81f68c",
  4600 => x"08841108",
  4601 => x"55538151",
  4602 => x"ff93dc3f",
  4603 => x"b00881ff",
  4604 => x"0674dfff",
  4605 => x"ff065452",
  4606 => x"71802e87",
  4607 => x"3873a080",
  4608 => x"80075382",
  4609 => x"51ff93bf",
  4610 => x"3fb00881",
  4611 => x"ff0673ef",
  4612 => x"ff0a0655",
  4613 => x"5271802e",
  4614 => x"87387290",
  4615 => x"800a0754",
  4616 => x"8351ff93",
  4617 => x"a23fb008",
  4618 => x"81ff0674",
  4619 => x"f7ff0a06",
  4620 => x"54527180",
  4621 => x"2e873873",
  4622 => x"88800a07",
  4623 => x"538451ff",
  4624 => x"93853fb0",
  4625 => x"0881ff06",
  4626 => x"73fbff0a",
  4627 => x"06555271",
  4628 => x"802e8738",
  4629 => x"7284800a",
  4630 => x"07548551",
  4631 => x"ff92e83f",
  4632 => x"b00881ff",
  4633 => x"0674fdff",
  4634 => x"0a065452",
  4635 => x"71802e87",
  4636 => x"38738280",
  4637 => x"0a075381",
  4638 => x"f68c0873",
  4639 => x"84120c54",
  4640 => x"72b00c85",
  4641 => x"3d0d04fa",
  4642 => x"3d0d880a",
  4643 => x"0b81f5e0",
  4644 => x"088c1108",
  4645 => x"59555681",
  4646 => x"51ff92ab",
  4647 => x"3fb00890",
  4648 => x"2b70902c",
  4649 => x"56538077",
  4650 => x"27993880",
  4651 => x"77545473",
  4652 => x"83ffff06",
  4653 => x"76708405",
  4654 => x"580cff13",
  4655 => x"75155553",
  4656 => x"72ed3880",
  4657 => x"0bb00c88",
  4658 => x"3d0d04fd",
  4659 => x"3d0d0297",
  4660 => x"053381f6",
  4661 => x"8c088411",
  4662 => x"0870b080",
  4663 => x"0a0770ef",
  4664 => x"ff0a0651",
  4665 => x"54555552",
  4666 => x"71802e87",
  4667 => x"3872b080",
  4668 => x"0a075170",
  4669 => x"8e800a07",
  4670 => x"84150c85",
  4671 => x"3d0d04ff",
  4672 => x"85f73f04",
  4673 => x"fb3d0d77",
  4674 => x"79555580",
  4675 => x"56757524",
  4676 => x"ab388074",
  4677 => x"249d3880",
  4678 => x"53735274",
  4679 => x"5180e13f",
  4680 => x"b0085475",
  4681 => x"802e8538",
  4682 => x"b0083054",
  4683 => x"73b00c87",
  4684 => x"3d0d0473",
  4685 => x"30768132",
  4686 => x"5754dc39",
  4687 => x"74305581",
  4688 => x"56738025",
  4689 => x"d238ec39",
  4690 => x"fa3d0d78",
  4691 => x"7a575580",
  4692 => x"57767524",
  4693 => x"a438759f",
  4694 => x"2c548153",
  4695 => x"75743274",
  4696 => x"31527451",
  4697 => x"9b3fb008",
  4698 => x"5476802e",
  4699 => x"8538b008",
  4700 => x"305473b0",
  4701 => x"0c883d0d",
  4702 => x"04743055",
  4703 => x"8157d739",
  4704 => x"fc3d0d76",
  4705 => x"78535481",
  4706 => x"53807473",
  4707 => x"26525572",
  4708 => x"802e9838",
  4709 => x"70802ea9",
  4710 => x"38807224",
  4711 => x"a4387110",
  4712 => x"73107572",
  4713 => x"26535452",
  4714 => x"72ea3873",
  4715 => x"51788338",
  4716 => x"745170b0",
  4717 => x"0c863d0d",
  4718 => x"0472812a",
  4719 => x"72812a53",
  4720 => x"5372802e",
  4721 => x"e6387174",
  4722 => x"26ef3873",
  4723 => x"72317574",
  4724 => x"0774812a",
  4725 => x"74812a55",
  4726 => x"555654e5",
  4727 => x"39101010",
  4728 => x"10101010",
  4729 => x"10101010",
  4730 => x"10101010",
  4731 => x"10101010",
  4732 => x"10101010",
  4733 => x"10101010",
  4734 => x"10101010",
  4735 => x"53510473",
  4736 => x"81ff0673",
  4737 => x"83060981",
  4738 => x"05830510",
  4739 => x"10102b07",
  4740 => x"72fc060c",
  4741 => x"5151043c",
  4742 => x"04727280",
  4743 => x"728106ff",
  4744 => x"05097206",
  4745 => x"05711052",
  4746 => x"720a100a",
  4747 => x"5372ed38",
  4748 => x"51515351",
  4749 => x"04b008b4",
  4750 => x"08b80875",
  4751 => x"758192c8",
  4752 => x"2d5050b0",
  4753 => x"0856b80c",
  4754 => x"b40cb00c",
  4755 => x"5104b008",
  4756 => x"b408b808",
  4757 => x"75758192",
  4758 => x"842d5050",
  4759 => x"b00856b8",
  4760 => x"0cb40cb0",
  4761 => x"0c5104b0",
  4762 => x"08b408b8",
  4763 => x"0897d02d",
  4764 => x"b80cb40c",
  4765 => x"b00c04ff",
  4766 => x"3d0d028f",
  4767 => x"053381f6",
  4768 => x"9c085271",
  4769 => x"0c800bb0",
  4770 => x"0c833d0d",
  4771 => x"04ff3d0d",
  4772 => x"028f0533",
  4773 => x"51829ebc",
  4774 => x"0852712d",
  4775 => x"b00881ff",
  4776 => x"06b00c83",
  4777 => x"3d0d04fe",
  4778 => x"3d0d7470",
  4779 => x"33535371",
  4780 => x"802e9338",
  4781 => x"81137252",
  4782 => x"829ebc08",
  4783 => x"5353712d",
  4784 => x"72335271",
  4785 => x"ef38843d",
  4786 => x"0d04f43d",
  4787 => x"0d7f0284",
  4788 => x"05bb0533",
  4789 => x"5557880b",
  4790 => x"8c3d5b59",
  4791 => x"895381f3",
  4792 => x"b0527951",
  4793 => x"86d93f73",
  4794 => x"792e80ff",
  4795 => x"38785673",
  4796 => x"902e80ec",
  4797 => x"3802a705",
  4798 => x"58768f06",
  4799 => x"54738926",
  4800 => x"80c23875",
  4801 => x"18b01555",
  4802 => x"55737534",
  4803 => x"76842aff",
  4804 => x"177081ff",
  4805 => x"06585557",
  4806 => x"75df3878",
  4807 => x"1a557575",
  4808 => x"34797033",
  4809 => x"55557380",
  4810 => x"2e933881",
  4811 => x"15745282",
  4812 => x"9ebc0857",
  4813 => x"55752d74",
  4814 => x"335473ef",
  4815 => x"3878b00c",
  4816 => x"8e3d0d04",
  4817 => x"7518b715",
  4818 => x"55557375",
  4819 => x"3476842a",
  4820 => x"ff177081",
  4821 => x"ff065855",
  4822 => x"5775ff9d",
  4823 => x"38ffbc39",
  4824 => x"84705759",
  4825 => x"02a70558",
  4826 => x"ff8f3982",
  4827 => x"705759f4",
  4828 => x"39f13d0d",
  4829 => x"618d3d70",
  4830 => x"5b5c5a80",
  4831 => x"7a565776",
  4832 => x"7a248185",
  4833 => x"38781754",
  4834 => x"8a527451",
  4835 => x"84ff3fb0",
  4836 => x"08b00553",
  4837 => x"72743481",
  4838 => x"17578a52",
  4839 => x"745184c8",
  4840 => x"3fb00855",
  4841 => x"b008de38",
  4842 => x"b008779f",
  4843 => x"2a187081",
  4844 => x"2c5a5656",
  4845 => x"8078259e",
  4846 => x"387817ff",
  4847 => x"05557519",
  4848 => x"70335553",
  4849 => x"74337334",
  4850 => x"73753481",
  4851 => x"16ff1656",
  4852 => x"56777624",
  4853 => x"e9387619",
  4854 => x"58807834",
  4855 => x"807a2417",
  4856 => x"7081ff06",
  4857 => x"7c703356",
  4858 => x"57555672",
  4859 => x"802e9338",
  4860 => x"81157352",
  4861 => x"829ebc08",
  4862 => x"5855762d",
  4863 => x"74335372",
  4864 => x"ef3873b0",
  4865 => x"0c913d0d",
  4866 => x"04ad7b34",
  4867 => x"02ad057a",
  4868 => x"30711956",
  4869 => x"56598a52",
  4870 => x"745183f1",
  4871 => x"3fb008b0",
  4872 => x"05537274",
  4873 => x"34811757",
  4874 => x"8a527451",
  4875 => x"83ba3fb0",
  4876 => x"0855b008",
  4877 => x"fecf38fe",
  4878 => x"ef39fd3d",
  4879 => x"0d81f690",
  4880 => x"0876b2e4",
  4881 => x"2994120c",
  4882 => x"54850b98",
  4883 => x"150c9814",
  4884 => x"08708106",
  4885 => x"515372f6",
  4886 => x"38853d0d",
  4887 => x"04803d0d",
  4888 => x"81f69008",
  4889 => x"51870b84",
  4890 => x"120cff0b",
  4891 => x"a4120ca7",
  4892 => x"0ba8120c",
  4893 => x"b2e40b94",
  4894 => x"120c870b",
  4895 => x"98120c82",
  4896 => x"3d0d0480",
  4897 => x"3d0d81f6",
  4898 => x"940851b8",
  4899 => x"0b8c120c",
  4900 => x"830b8812",
  4901 => x"0c823d0d",
  4902 => x"04803d0d",
  4903 => x"81f69408",
  4904 => x"84110881",
  4905 => x"06b00c51",
  4906 => x"823d0d04",
  4907 => x"ff3d0d81",
  4908 => x"f6940852",
  4909 => x"84120870",
  4910 => x"81065151",
  4911 => x"70802ef4",
  4912 => x"38710870",
  4913 => x"81ff06b0",
  4914 => x"0c51833d",
  4915 => x"0d04fe3d",
  4916 => x"0d029305",
  4917 => x"3381f694",
  4918 => x"08535384",
  4919 => x"12087089",
  4920 => x"2a708106",
  4921 => x"51515170",
  4922 => x"f2387272",
  4923 => x"0c843d0d",
  4924 => x"04fe3d0d",
  4925 => x"02930533",
  4926 => x"53728a2e",
  4927 => x"9c3881f6",
  4928 => x"94085284",
  4929 => x"12087089",
  4930 => x"2a708106",
  4931 => x"51515170",
  4932 => x"f2387272",
  4933 => x"0c843d0d",
  4934 => x"0481f694",
  4935 => x"08528412",
  4936 => x"0870892a",
  4937 => x"70810651",
  4938 => x"515170f2",
  4939 => x"388d720c",
  4940 => x"84120870",
  4941 => x"892a7081",
  4942 => x"06515151",
  4943 => x"70c538d2",
  4944 => x"39803d0d",
  4945 => x"81f68808",
  4946 => x"51800b84",
  4947 => x"120c83fe",
  4948 => x"800b8812",
  4949 => x"0c800b82",
  4950 => x"9ec03480",
  4951 => x"0b829ec4",
  4952 => x"34823d0d",
  4953 => x"04fa3d0d",
  4954 => x"02a30533",
  4955 => x"81f68808",
  4956 => x"829ec033",
  4957 => x"7081ff06",
  4958 => x"70101011",
  4959 => x"829ec433",
  4960 => x"7081ff06",
  4961 => x"72902911",
  4962 => x"70882b78",
  4963 => x"07770c53",
  4964 => x"5b5b5555",
  4965 => x"59545473",
  4966 => x"8a2e9838",
  4967 => x"7480cf2e",
  4968 => x"9238738c",
  4969 => x"2ea43881",
  4970 => x"16537282",
  4971 => x"9ec43488",
  4972 => x"3d0d0471",
  4973 => x"a326a338",
  4974 => x"81175271",
  4975 => x"829ec034",
  4976 => x"800b829e",
  4977 => x"c434883d",
  4978 => x"0d048052",
  4979 => x"71882b73",
  4980 => x"0c811252",
  4981 => x"97907226",
  4982 => x"f338800b",
  4983 => x"829ec034",
  4984 => x"800b829e",
  4985 => x"c434df39",
  4986 => x"bc0802bc",
  4987 => x"0cfd3d0d",
  4988 => x"8053bc08",
  4989 => x"8c050852",
  4990 => x"bc088805",
  4991 => x"0851f780",
  4992 => x"3fb00870",
  4993 => x"b00c5485",
  4994 => x"3d0dbc0c",
  4995 => x"04bc0802",
  4996 => x"bc0cfd3d",
  4997 => x"0d8153bc",
  4998 => x"088c0508",
  4999 => x"52bc0888",
  5000 => x"050851f6",
  5001 => x"db3fb008",
  5002 => x"70b00c54",
  5003 => x"853d0dbc",
  5004 => x"0c04803d",
  5005 => x"0d865184",
  5006 => x"963f8151",
  5007 => x"a1d33ffc",
  5008 => x"3d0d7670",
  5009 => x"797b5555",
  5010 => x"55558f72",
  5011 => x"278c3872",
  5012 => x"75078306",
  5013 => x"5170802e",
  5014 => x"a738ff12",
  5015 => x"5271ff2e",
  5016 => x"98387270",
  5017 => x"81055433",
  5018 => x"74708105",
  5019 => x"5634ff12",
  5020 => x"5271ff2e",
  5021 => x"098106ea",
  5022 => x"3874b00c",
  5023 => x"863d0d04",
  5024 => x"74517270",
  5025 => x"84055408",
  5026 => x"71708405",
  5027 => x"530c7270",
  5028 => x"84055408",
  5029 => x"71708405",
  5030 => x"530c7270",
  5031 => x"84055408",
  5032 => x"71708405",
  5033 => x"530c7270",
  5034 => x"84055408",
  5035 => x"71708405",
  5036 => x"530cf012",
  5037 => x"52718f26",
  5038 => x"c9388372",
  5039 => x"27953872",
  5040 => x"70840554",
  5041 => x"08717084",
  5042 => x"05530cfc",
  5043 => x"12527183",
  5044 => x"26ed3870",
  5045 => x"54ff8339",
  5046 => x"fd3d0d75",
  5047 => x"5384d813",
  5048 => x"08802e8a",
  5049 => x"38805372",
  5050 => x"b00c853d",
  5051 => x"0d048180",
  5052 => x"5272518d",
  5053 => x"9b3fb008",
  5054 => x"84d8140c",
  5055 => x"ff53b008",
  5056 => x"802ee438",
  5057 => x"b008549f",
  5058 => x"53807470",
  5059 => x"8405560c",
  5060 => x"ff135380",
  5061 => x"7324ce38",
  5062 => x"80747084",
  5063 => x"05560cff",
  5064 => x"13537280",
  5065 => x"25e338ff",
  5066 => x"bc39fd3d",
  5067 => x"0d757755",
  5068 => x"539f7427",
  5069 => x"8d389673",
  5070 => x"0cff5271",
  5071 => x"b00c853d",
  5072 => x"0d0484d8",
  5073 => x"13085271",
  5074 => x"802e9338",
  5075 => x"73101012",
  5076 => x"70087972",
  5077 => x"0c515271",
  5078 => x"b00c853d",
  5079 => x"0d047251",
  5080 => x"fef63fff",
  5081 => x"52b008d3",
  5082 => x"3884d813",
  5083 => x"08741010",
  5084 => x"1170087a",
  5085 => x"720c5151",
  5086 => x"52dd39f9",
  5087 => x"3d0d797b",
  5088 => x"5856769f",
  5089 => x"2680e838",
  5090 => x"84d81608",
  5091 => x"5473802e",
  5092 => x"aa387610",
  5093 => x"10147008",
  5094 => x"55557380",
  5095 => x"2eba3880",
  5096 => x"5873812e",
  5097 => x"8f3873ff",
  5098 => x"2ea33880",
  5099 => x"750c7651",
  5100 => x"732d8058",
  5101 => x"77b00c89",
  5102 => x"3d0d0475",
  5103 => x"51fe993f",
  5104 => x"ff58b008",
  5105 => x"ef3884d8",
  5106 => x"160854c6",
  5107 => x"3996760c",
  5108 => x"810bb00c",
  5109 => x"893d0d04",
  5110 => x"755181ed",
  5111 => x"3f7653b0",
  5112 => x"08527551",
  5113 => x"81ad3fb0",
  5114 => x"08b00c89",
  5115 => x"3d0d0496",
  5116 => x"760cff0b",
  5117 => x"b00c893d",
  5118 => x"0d04fc3d",
  5119 => x"0d767856",
  5120 => x"53ff5474",
  5121 => x"9f26b138",
  5122 => x"84d81308",
  5123 => x"5271802e",
  5124 => x"ae387410",
  5125 => x"10127008",
  5126 => x"53538154",
  5127 => x"71802e98",
  5128 => x"38825471",
  5129 => x"ff2e9138",
  5130 => x"83547181",
  5131 => x"2e8a3880",
  5132 => x"730c7451",
  5133 => x"712d8054",
  5134 => x"73b00c86",
  5135 => x"3d0d0472",
  5136 => x"51fd953f",
  5137 => x"b008f138",
  5138 => x"84d81308",
  5139 => x"52c439ff",
  5140 => x"3d0d7352",
  5141 => x"81f6a008",
  5142 => x"51fea03f",
  5143 => x"833d0d04",
  5144 => x"fe3d0d75",
  5145 => x"53745281",
  5146 => x"f6a00851",
  5147 => x"fdbc3f84",
  5148 => x"3d0d0480",
  5149 => x"3d0d81f6",
  5150 => x"a00851fc",
  5151 => x"db3f823d",
  5152 => x"0d04ff3d",
  5153 => x"0d735281",
  5154 => x"f6a00851",
  5155 => x"feec3f83",
  5156 => x"3d0d04fc",
  5157 => x"3d0d800b",
  5158 => x"829ecc0c",
  5159 => x"78527751",
  5160 => x"9caa3fb0",
  5161 => x"0854b008",
  5162 => x"ff2e8838",
  5163 => x"73b00c86",
  5164 => x"3d0d0482",
  5165 => x"9ecc0855",
  5166 => x"74802ef0",
  5167 => x"38767571",
  5168 => x"0c5373b0",
  5169 => x"0c863d0d",
  5170 => x"049bfc3f",
  5171 => x"04fc3d0d",
  5172 => x"76707970",
  5173 => x"73078306",
  5174 => x"54545455",
  5175 => x"7080c338",
  5176 => x"71700870",
  5177 => x"0970f7fb",
  5178 => x"fdff1306",
  5179 => x"70f88482",
  5180 => x"81800651",
  5181 => x"51535354",
  5182 => x"70a63884",
  5183 => x"14727470",
  5184 => x"8405560c",
  5185 => x"70087009",
  5186 => x"70f7fbfd",
  5187 => x"ff130670",
  5188 => x"f8848281",
  5189 => x"80065151",
  5190 => x"53535470",
  5191 => x"802edc38",
  5192 => x"73527170",
  5193 => x"81055333",
  5194 => x"51707370",
  5195 => x"81055534",
  5196 => x"70f03874",
  5197 => x"b00c863d",
  5198 => x"0d04fd3d",
  5199 => x"0d757071",
  5200 => x"83065355",
  5201 => x"5270b838",
  5202 => x"71700870",
  5203 => x"09f7fbfd",
  5204 => x"ff120670",
  5205 => x"f8848281",
  5206 => x"80065151",
  5207 => x"5253709d",
  5208 => x"38841370",
  5209 => x"087009f7",
  5210 => x"fbfdff12",
  5211 => x"0670f884",
  5212 => x"82818006",
  5213 => x"51515253",
  5214 => x"70802ee5",
  5215 => x"38725271",
  5216 => x"33517080",
  5217 => x"2e8a3881",
  5218 => x"12703352",
  5219 => x"5270f838",
  5220 => x"717431b0",
  5221 => x"0c853d0d",
  5222 => x"04fa3d0d",
  5223 => x"787a7c70",
  5224 => x"54555552",
  5225 => x"72802e80",
  5226 => x"d9387174",
  5227 => x"07830651",
  5228 => x"70802e80",
  5229 => x"d438ff13",
  5230 => x"5372ff2e",
  5231 => x"b1387133",
  5232 => x"74335651",
  5233 => x"74712e09",
  5234 => x"8106a938",
  5235 => x"72802e81",
  5236 => x"87387081",
  5237 => x"ff065170",
  5238 => x"802e80fc",
  5239 => x"38811281",
  5240 => x"15ff1555",
  5241 => x"555272ff",
  5242 => x"2e098106",
  5243 => x"d1387133",
  5244 => x"74335651",
  5245 => x"7081ff06",
  5246 => x"7581ff06",
  5247 => x"71713151",
  5248 => x"525270b0",
  5249 => x"0c883d0d",
  5250 => x"04717457",
  5251 => x"55837327",
  5252 => x"88387108",
  5253 => x"74082e88",
  5254 => x"38747655",
  5255 => x"52ff9739",
  5256 => x"fc135372",
  5257 => x"802eb138",
  5258 => x"74087009",
  5259 => x"f7fbfdff",
  5260 => x"120670f8",
  5261 => x"84828180",
  5262 => x"06515151",
  5263 => x"709a3884",
  5264 => x"15841757",
  5265 => x"55837327",
  5266 => x"d0387408",
  5267 => x"76082ed0",
  5268 => x"38747655",
  5269 => x"52fedf39",
  5270 => x"800bb00c",
  5271 => x"883d0d04",
  5272 => x"f33d0d60",
  5273 => x"6264725a",
  5274 => x"5a5e5e80",
  5275 => x"5c767081",
  5276 => x"05583381",
  5277 => x"f3bd1133",
  5278 => x"70832a70",
  5279 => x"81065155",
  5280 => x"555672e9",
  5281 => x"3875ad2e",
  5282 => x"82883875",
  5283 => x"ab2e8284",
  5284 => x"38773070",
  5285 => x"79078025",
  5286 => x"79903270",
  5287 => x"30707207",
  5288 => x"80257307",
  5289 => x"53575751",
  5290 => x"5372802e",
  5291 => x"873875b0",
  5292 => x"2e81eb38",
  5293 => x"778a3888",
  5294 => x"5875b02e",
  5295 => x"83388a58",
  5296 => x"810a5a7b",
  5297 => x"8438fe0a",
  5298 => x"5a775279",
  5299 => x"51f6be3f",
  5300 => x"b0087853",
  5301 => x"7a525bf6",
  5302 => x"8f3fb008",
  5303 => x"5a807081",
  5304 => x"f3bd1833",
  5305 => x"70822a70",
  5306 => x"81065156",
  5307 => x"565a5572",
  5308 => x"802e80c1",
  5309 => x"38d01656",
  5310 => x"75782580",
  5311 => x"d7388079",
  5312 => x"24757b26",
  5313 => x"07537293",
  5314 => x"38747a2e",
  5315 => x"80eb387a",
  5316 => x"762580ed",
  5317 => x"3872802e",
  5318 => x"80e738ff",
  5319 => x"77708105",
  5320 => x"59335759",
  5321 => x"81f3bd16",
  5322 => x"3370822a",
  5323 => x"70810651",
  5324 => x"545472c1",
  5325 => x"38738306",
  5326 => x"5372802e",
  5327 => x"97387381",
  5328 => x"06c91755",
  5329 => x"53728538",
  5330 => x"ffa91654",
  5331 => x"73567776",
  5332 => x"24ffab38",
  5333 => x"80792480",
  5334 => x"f0387b80",
  5335 => x"2e843874",
  5336 => x"30557c80",
  5337 => x"2e8c38ff",
  5338 => x"17537883",
  5339 => x"387d5372",
  5340 => x"7d0c74b0",
  5341 => x"0c8f3d0d",
  5342 => x"04815375",
  5343 => x"7b24ff95",
  5344 => x"38817579",
  5345 => x"29177870",
  5346 => x"81055a33",
  5347 => x"585659ff",
  5348 => x"9339815c",
  5349 => x"76708105",
  5350 => x"583356fd",
  5351 => x"f4398077",
  5352 => x"33545472",
  5353 => x"80f82eb2",
  5354 => x"387280d8",
  5355 => x"32703070",
  5356 => x"80257607",
  5357 => x"51515372",
  5358 => x"802efdf8",
  5359 => x"38811733",
  5360 => x"82185856",
  5361 => x"9058fdf8",
  5362 => x"39810a55",
  5363 => x"7b8438fe",
  5364 => x"0a557f53",
  5365 => x"a2730cff",
  5366 => x"89398154",
  5367 => x"cc39fd3d",
  5368 => x"0d775476",
  5369 => x"53755281",
  5370 => x"f6a00851",
  5371 => x"fcf23f85",
  5372 => x"3d0d04f3",
  5373 => x"3d0d6062",
  5374 => x"64725a5a",
  5375 => x"5d5d805e",
  5376 => x"76708105",
  5377 => x"583381f3",
  5378 => x"bd113370",
  5379 => x"832a7081",
  5380 => x"06515555",
  5381 => x"5672e938",
  5382 => x"75ad2e81",
  5383 => x"ff3875ab",
  5384 => x"2e81fb38",
  5385 => x"77307079",
  5386 => x"07802579",
  5387 => x"90327030",
  5388 => x"70720780",
  5389 => x"25730753",
  5390 => x"57575153",
  5391 => x"72802e87",
  5392 => x"3875b02e",
  5393 => x"81e23877",
  5394 => x"8a388858",
  5395 => x"75b02e83",
  5396 => x"388a5877",
  5397 => x"52ff51f3",
  5398 => x"8f3fb008",
  5399 => x"78535aff",
  5400 => x"51f3aa3f",
  5401 => x"b0085b80",
  5402 => x"705a5581",
  5403 => x"f3bd1633",
  5404 => x"70822a70",
  5405 => x"81065154",
  5406 => x"5472802e",
  5407 => x"80c138d0",
  5408 => x"16567578",
  5409 => x"2580d738",
  5410 => x"80792475",
  5411 => x"7b260753",
  5412 => x"72933874",
  5413 => x"7a2e80eb",
  5414 => x"387a7625",
  5415 => x"80ed3872",
  5416 => x"802e80e7",
  5417 => x"38ff7770",
  5418 => x"81055933",
  5419 => x"575981f3",
  5420 => x"bd163370",
  5421 => x"822a7081",
  5422 => x"06515454",
  5423 => x"72c13873",
  5424 => x"83065372",
  5425 => x"802e9738",
  5426 => x"738106c9",
  5427 => x"17555372",
  5428 => x"8538ffa9",
  5429 => x"16547356",
  5430 => x"777624ff",
  5431 => x"ab388079",
  5432 => x"24818938",
  5433 => x"7d802e84",
  5434 => x"38743055",
  5435 => x"7b802e8c",
  5436 => x"38ff1753",
  5437 => x"7883387c",
  5438 => x"53727c0c",
  5439 => x"74b00c8f",
  5440 => x"3d0d0481",
  5441 => x"53757b24",
  5442 => x"ff953881",
  5443 => x"75792917",
  5444 => x"78708105",
  5445 => x"5a335856",
  5446 => x"59ff9339",
  5447 => x"815e7670",
  5448 => x"81055833",
  5449 => x"56fdfd39",
  5450 => x"80773354",
  5451 => x"547280f8",
  5452 => x"2e80c338",
  5453 => x"7280d832",
  5454 => x"70307080",
  5455 => x"25760751",
  5456 => x"51537280",
  5457 => x"2efe8038",
  5458 => x"81173382",
  5459 => x"18585690",
  5460 => x"705358ff",
  5461 => x"51f1913f",
  5462 => x"b0087853",
  5463 => x"5aff51f1",
  5464 => x"ac3fb008",
  5465 => x"5b80705a",
  5466 => x"55fe8039",
  5467 => x"ff605455",
  5468 => x"a2730cfe",
  5469 => x"f7398154",
  5470 => x"ffba39fd",
  5471 => x"3d0d7754",
  5472 => x"76537552",
  5473 => x"81f6a008",
  5474 => x"51fce83f",
  5475 => x"853d0d04",
  5476 => x"f33d0d7f",
  5477 => x"618b1170",
  5478 => x"f8065c55",
  5479 => x"555e7296",
  5480 => x"26833890",
  5481 => x"59807924",
  5482 => x"747a2607",
  5483 => x"53805472",
  5484 => x"742e0981",
  5485 => x"0680cb38",
  5486 => x"7d518bca",
  5487 => x"3f7883f7",
  5488 => x"2680c638",
  5489 => x"78832a70",
  5490 => x"10101081",
  5491 => x"fddc058c",
  5492 => x"11085959",
  5493 => x"5a76782e",
  5494 => x"83b03884",
  5495 => x"1708fc06",
  5496 => x"568c1708",
  5497 => x"88180871",
  5498 => x"8c120c88",
  5499 => x"120c5875",
  5500 => x"17841108",
  5501 => x"81078412",
  5502 => x"0c537d51",
  5503 => x"8b893f88",
  5504 => x"175473b0",
  5505 => x"0c8f3d0d",
  5506 => x"0478892a",
  5507 => x"79832a5b",
  5508 => x"5372802e",
  5509 => x"bf387886",
  5510 => x"2ab8055a",
  5511 => x"847327b4",
  5512 => x"3880db13",
  5513 => x"5a947327",
  5514 => x"ab38788c",
  5515 => x"2a80ee05",
  5516 => x"5a80d473",
  5517 => x"279e3878",
  5518 => x"8f2a80f7",
  5519 => x"055a82d4",
  5520 => x"73279138",
  5521 => x"78922a80",
  5522 => x"fc055a8a",
  5523 => x"d4732784",
  5524 => x"3880fe5a",
  5525 => x"79101010",
  5526 => x"81fddc05",
  5527 => x"8c110858",
  5528 => x"5576752e",
  5529 => x"a3388417",
  5530 => x"08fc0670",
  5531 => x"7a315556",
  5532 => x"738f2488",
  5533 => x"d5387380",
  5534 => x"25fee638",
  5535 => x"8c170857",
  5536 => x"76752e09",
  5537 => x"8106df38",
  5538 => x"811a5a81",
  5539 => x"fdec0857",
  5540 => x"7681fde4",
  5541 => x"2e82c038",
  5542 => x"841708fc",
  5543 => x"06707a31",
  5544 => x"5556738f",
  5545 => x"2481f938",
  5546 => x"81fde40b",
  5547 => x"81fdf00c",
  5548 => x"81fde40b",
  5549 => x"81fdec0c",
  5550 => x"738025fe",
  5551 => x"b23883ff",
  5552 => x"762783df",
  5553 => x"3875892a",
  5554 => x"76832a55",
  5555 => x"5372802e",
  5556 => x"bf387586",
  5557 => x"2ab80554",
  5558 => x"847327b4",
  5559 => x"3880db13",
  5560 => x"54947327",
  5561 => x"ab38758c",
  5562 => x"2a80ee05",
  5563 => x"5480d473",
  5564 => x"279e3875",
  5565 => x"8f2a80f7",
  5566 => x"055482d4",
  5567 => x"73279138",
  5568 => x"75922a80",
  5569 => x"fc05548a",
  5570 => x"d4732784",
  5571 => x"3880fe54",
  5572 => x"73101010",
  5573 => x"81fddc05",
  5574 => x"88110856",
  5575 => x"5874782e",
  5576 => x"86cf3884",
  5577 => x"1508fc06",
  5578 => x"53757327",
  5579 => x"8d388815",
  5580 => x"08557478",
  5581 => x"2e098106",
  5582 => x"ea388c15",
  5583 => x"0881fddc",
  5584 => x"0b840508",
  5585 => x"718c1a0c",
  5586 => x"76881a0c",
  5587 => x"7888130c",
  5588 => x"788c180c",
  5589 => x"5d587953",
  5590 => x"807a2483",
  5591 => x"e6387282",
  5592 => x"2c81712b",
  5593 => x"5c537a7c",
  5594 => x"26819838",
  5595 => x"7b7b0653",
  5596 => x"7282f138",
  5597 => x"79fc0684",
  5598 => x"055a7a10",
  5599 => x"707d0654",
  5600 => x"5b7282e0",
  5601 => x"38841a5a",
  5602 => x"f1398817",
  5603 => x"8c110858",
  5604 => x"5876782e",
  5605 => x"098106fc",
  5606 => x"c238821a",
  5607 => x"5afdec39",
  5608 => x"78177981",
  5609 => x"0784190c",
  5610 => x"7081fdf0",
  5611 => x"0c7081fd",
  5612 => x"ec0c81fd",
  5613 => x"e40b8c12",
  5614 => x"0c8c1108",
  5615 => x"88120c74",
  5616 => x"81078412",
  5617 => x"0c741175",
  5618 => x"710c5153",
  5619 => x"7d5187b7",
  5620 => x"3f881754",
  5621 => x"fcac3981",
  5622 => x"fddc0b84",
  5623 => x"05087a54",
  5624 => x"5c798025",
  5625 => x"fef83882",
  5626 => x"da397a09",
  5627 => x"7c067081",
  5628 => x"fddc0b84",
  5629 => x"050c5c7a",
  5630 => x"105b7a7c",
  5631 => x"2685387a",
  5632 => x"85b83881",
  5633 => x"fddc0b88",
  5634 => x"05087084",
  5635 => x"1208fc06",
  5636 => x"707c317c",
  5637 => x"72268f72",
  5638 => x"25075757",
  5639 => x"5c5d5572",
  5640 => x"802e80db",
  5641 => x"38797a16",
  5642 => x"81fdd408",
  5643 => x"1b90115a",
  5644 => x"55575b81",
  5645 => x"fdd008ff",
  5646 => x"2e8838a0",
  5647 => x"8f13e080",
  5648 => x"06577652",
  5649 => x"7d5186c0",
  5650 => x"3fb00854",
  5651 => x"b008ff2e",
  5652 => x"9038b008",
  5653 => x"76278299",
  5654 => x"387481fd",
  5655 => x"dc2e8291",
  5656 => x"3881fddc",
  5657 => x"0b880508",
  5658 => x"55841508",
  5659 => x"fc06707a",
  5660 => x"317a7226",
  5661 => x"8f722507",
  5662 => x"52555372",
  5663 => x"83e63874",
  5664 => x"79810784",
  5665 => x"170c7916",
  5666 => x"7081fddc",
  5667 => x"0b88050c",
  5668 => x"75810784",
  5669 => x"120c547e",
  5670 => x"525785eb",
  5671 => x"3f881754",
  5672 => x"fae03975",
  5673 => x"832a7054",
  5674 => x"54807424",
  5675 => x"819b3872",
  5676 => x"822c8171",
  5677 => x"2b81fde0",
  5678 => x"08077081",
  5679 => x"fddc0b84",
  5680 => x"050c7510",
  5681 => x"101081fd",
  5682 => x"dc058811",
  5683 => x"08585a5d",
  5684 => x"53778c18",
  5685 => x"0c748818",
  5686 => x"0c768819",
  5687 => x"0c768c16",
  5688 => x"0cfcf339",
  5689 => x"797a1010",
  5690 => x"1081fddc",
  5691 => x"05705759",
  5692 => x"5d8c1508",
  5693 => x"5776752e",
  5694 => x"a3388417",
  5695 => x"08fc0670",
  5696 => x"7a315556",
  5697 => x"738f2483",
  5698 => x"ca387380",
  5699 => x"25848138",
  5700 => x"8c170857",
  5701 => x"76752e09",
  5702 => x"8106df38",
  5703 => x"8815811b",
  5704 => x"70830655",
  5705 => x"5b5572c9",
  5706 => x"387c8306",
  5707 => x"5372802e",
  5708 => x"fdb838ff",
  5709 => x"1df81959",
  5710 => x"5d881808",
  5711 => x"782eea38",
  5712 => x"fdb53983",
  5713 => x"1a53fc96",
  5714 => x"39831470",
  5715 => x"822c8171",
  5716 => x"2b81fde0",
  5717 => x"08077081",
  5718 => x"fddc0b84",
  5719 => x"050c7610",
  5720 => x"101081fd",
  5721 => x"dc058811",
  5722 => x"08595b5e",
  5723 => x"5153fee1",
  5724 => x"3981fda0",
  5725 => x"081758b0",
  5726 => x"08762e81",
  5727 => x"8d3881fd",
  5728 => x"d008ff2e",
  5729 => x"83ec3873",
  5730 => x"76311881",
  5731 => x"fda00c73",
  5732 => x"87067057",
  5733 => x"5372802e",
  5734 => x"88388873",
  5735 => x"31701555",
  5736 => x"5676149f",
  5737 => x"ff06a080",
  5738 => x"71311770",
  5739 => x"547f5357",
  5740 => x"5383d53f",
  5741 => x"b00853b0",
  5742 => x"08ff2e81",
  5743 => x"a03881fd",
  5744 => x"a0081670",
  5745 => x"81fda00c",
  5746 => x"747581fd",
  5747 => x"dc0b8805",
  5748 => x"0c747631",
  5749 => x"18708107",
  5750 => x"51555658",
  5751 => x"7b81fddc",
  5752 => x"2e839c38",
  5753 => x"798f2682",
  5754 => x"cb38810b",
  5755 => x"84150c84",
  5756 => x"1508fc06",
  5757 => x"707a317a",
  5758 => x"72268f72",
  5759 => x"25075255",
  5760 => x"5372802e",
  5761 => x"fcf93880",
  5762 => x"db39b008",
  5763 => x"9fff0653",
  5764 => x"72feeb38",
  5765 => x"7781fda0",
  5766 => x"0c81fddc",
  5767 => x"0b880508",
  5768 => x"7b188107",
  5769 => x"84120c55",
  5770 => x"81fdcc08",
  5771 => x"78278638",
  5772 => x"7781fdcc",
  5773 => x"0c81fdc8",
  5774 => x"087827fc",
  5775 => x"ac387781",
  5776 => x"fdc80c84",
  5777 => x"1508fc06",
  5778 => x"707a317a",
  5779 => x"72268f72",
  5780 => x"25075255",
  5781 => x"5372802e",
  5782 => x"fca53888",
  5783 => x"39807454",
  5784 => x"56fedb39",
  5785 => x"7d51829f",
  5786 => x"3f800bb0",
  5787 => x"0c8f3d0d",
  5788 => x"04735380",
  5789 => x"7424a938",
  5790 => x"72822c81",
  5791 => x"712b81fd",
  5792 => x"e0080770",
  5793 => x"81fddc0b",
  5794 => x"84050c5d",
  5795 => x"53778c18",
  5796 => x"0c748818",
  5797 => x"0c768819",
  5798 => x"0c768c16",
  5799 => x"0cf9b739",
  5800 => x"83147082",
  5801 => x"2c81712b",
  5802 => x"81fde008",
  5803 => x"077081fd",
  5804 => x"dc0b8405",
  5805 => x"0c5e5153",
  5806 => x"d4397b7b",
  5807 => x"065372fc",
  5808 => x"a338841a",
  5809 => x"7b105c5a",
  5810 => x"f139ff1a",
  5811 => x"8111515a",
  5812 => x"f7b93978",
  5813 => x"17798107",
  5814 => x"84190c8c",
  5815 => x"18088819",
  5816 => x"08718c12",
  5817 => x"0c88120c",
  5818 => x"597081fd",
  5819 => x"f00c7081",
  5820 => x"fdec0c81",
  5821 => x"fde40b8c",
  5822 => x"120c8c11",
  5823 => x"0888120c",
  5824 => x"74810784",
  5825 => x"120c7411",
  5826 => x"75710c51",
  5827 => x"53f9bd39",
  5828 => x"75178411",
  5829 => x"08810784",
  5830 => x"120c538c",
  5831 => x"17088818",
  5832 => x"08718c12",
  5833 => x"0c88120c",
  5834 => x"587d5180",
  5835 => x"da3f8817",
  5836 => x"54f5cf39",
  5837 => x"7284150c",
  5838 => x"f41af806",
  5839 => x"70841e08",
  5840 => x"81060784",
  5841 => x"1e0c701d",
  5842 => x"545b850b",
  5843 => x"84140c85",
  5844 => x"0b88140c",
  5845 => x"8f7b27fd",
  5846 => x"cf38881c",
  5847 => x"527d5182",
  5848 => x"903f81fd",
  5849 => x"dc0b8805",
  5850 => x"0881fda0",
  5851 => x"085955fd",
  5852 => x"b7397781",
  5853 => x"fda00c73",
  5854 => x"81fdd00c",
  5855 => x"fc913972",
  5856 => x"84150cfd",
  5857 => x"a3390404",
  5858 => x"fd3d0d80",
  5859 => x"0b829ecc",
  5860 => x"0c765186",
  5861 => x"cb3fb008",
  5862 => x"53b008ff",
  5863 => x"2e883872",
  5864 => x"b00c853d",
  5865 => x"0d04829e",
  5866 => x"cc085473",
  5867 => x"802ef038",
  5868 => x"7574710c",
  5869 => x"5272b00c",
  5870 => x"853d0d04",
  5871 => x"fb3d0d77",
  5872 => x"705256c2",
  5873 => x"3f81fddc",
  5874 => x"0b880508",
  5875 => x"841108fc",
  5876 => x"06707b31",
  5877 => x"9fef05e0",
  5878 => x"8006e080",
  5879 => x"05565653",
  5880 => x"a0807424",
  5881 => x"94388052",
  5882 => x"7551ff9c",
  5883 => x"3f81fde4",
  5884 => x"08155372",
  5885 => x"b0082e8f",
  5886 => x"387551ff",
  5887 => x"8a3f8053",
  5888 => x"72b00c87",
  5889 => x"3d0d0473",
  5890 => x"30527551",
  5891 => x"fefa3fb0",
  5892 => x"08ff2ea8",
  5893 => x"3881fddc",
  5894 => x"0b880508",
  5895 => x"75753181",
  5896 => x"0784120c",
  5897 => x"5381fda0",
  5898 => x"08743181",
  5899 => x"fda00c75",
  5900 => x"51fed43f",
  5901 => x"810bb00c",
  5902 => x"873d0d04",
  5903 => x"80527551",
  5904 => x"fec63f81",
  5905 => x"fddc0b88",
  5906 => x"0508b008",
  5907 => x"71315653",
  5908 => x"8f7525ff",
  5909 => x"a438b008",
  5910 => x"81fdd008",
  5911 => x"3181fda0",
  5912 => x"0c748107",
  5913 => x"84140c75",
  5914 => x"51fe9c3f",
  5915 => x"8053ff90",
  5916 => x"39f63d0d",
  5917 => x"7c7e545b",
  5918 => x"72802e82",
  5919 => x"83387a51",
  5920 => x"fe843ff8",
  5921 => x"13841108",
  5922 => x"70fe0670",
  5923 => x"13841108",
  5924 => x"fc065d58",
  5925 => x"59545881",
  5926 => x"fde40875",
  5927 => x"2e82de38",
  5928 => x"7884160c",
  5929 => x"80738106",
  5930 => x"545a727a",
  5931 => x"2e81d538",
  5932 => x"78158411",
  5933 => x"08810651",
  5934 => x"5372a038",
  5935 => x"78175779",
  5936 => x"81e63888",
  5937 => x"15085372",
  5938 => x"81fde42e",
  5939 => x"82f9388c",
  5940 => x"1508708c",
  5941 => x"150c7388",
  5942 => x"120c5676",
  5943 => x"81078419",
  5944 => x"0c761877",
  5945 => x"710c5379",
  5946 => x"81913883",
  5947 => x"ff772781",
  5948 => x"c8387689",
  5949 => x"2a77832a",
  5950 => x"56537280",
  5951 => x"2ebf3876",
  5952 => x"862ab805",
  5953 => x"55847327",
  5954 => x"b43880db",
  5955 => x"13559473",
  5956 => x"27ab3876",
  5957 => x"8c2a80ee",
  5958 => x"055580d4",
  5959 => x"73279e38",
  5960 => x"768f2a80",
  5961 => x"f7055582",
  5962 => x"d4732791",
  5963 => x"3876922a",
  5964 => x"80fc0555",
  5965 => x"8ad47327",
  5966 => x"843880fe",
  5967 => x"55741010",
  5968 => x"1081fddc",
  5969 => x"05881108",
  5970 => x"55567376",
  5971 => x"2e82b338",
  5972 => x"841408fc",
  5973 => x"06537673",
  5974 => x"278d3888",
  5975 => x"14085473",
  5976 => x"762e0981",
  5977 => x"06ea388c",
  5978 => x"1408708c",
  5979 => x"1a0c7488",
  5980 => x"1a0c7888",
  5981 => x"120c5677",
  5982 => x"8c150c7a",
  5983 => x"51fc883f",
  5984 => x"8c3d0d04",
  5985 => x"77087871",
  5986 => x"31597705",
  5987 => x"88190854",
  5988 => x"577281fd",
  5989 => x"e42e80e0",
  5990 => x"388c1808",
  5991 => x"708c150c",
  5992 => x"7388120c",
  5993 => x"56fe8939",
  5994 => x"8815088c",
  5995 => x"1608708c",
  5996 => x"130c5788",
  5997 => x"170cfea3",
  5998 => x"3976832a",
  5999 => x"70545580",
  6000 => x"75248198",
  6001 => x"3872822c",
  6002 => x"81712b81",
  6003 => x"fde00807",
  6004 => x"81fddc0b",
  6005 => x"84050c53",
  6006 => x"74101010",
  6007 => x"81fddc05",
  6008 => x"88110855",
  6009 => x"56758c19",
  6010 => x"0c738819",
  6011 => x"0c778817",
  6012 => x"0c778c15",
  6013 => x"0cff8439",
  6014 => x"815afdb4",
  6015 => x"39781773",
  6016 => x"81065457",
  6017 => x"72983877",
  6018 => x"08787131",
  6019 => x"5977058c",
  6020 => x"1908881a",
  6021 => x"08718c12",
  6022 => x"0c88120c",
  6023 => x"57577681",
  6024 => x"0784190c",
  6025 => x"7781fddc",
  6026 => x"0b88050c",
  6027 => x"81fdd808",
  6028 => x"7726fec7",
  6029 => x"3881fdd4",
  6030 => x"08527a51",
  6031 => x"fafe3f7a",
  6032 => x"51fac43f",
  6033 => x"feba3981",
  6034 => x"788c150c",
  6035 => x"7888150c",
  6036 => x"738c1a0c",
  6037 => x"73881a0c",
  6038 => x"5afd8039",
  6039 => x"83157082",
  6040 => x"2c81712b",
  6041 => x"81fde008",
  6042 => x"0781fddc",
  6043 => x"0b84050c",
  6044 => x"51537410",
  6045 => x"101081fd",
  6046 => x"dc058811",
  6047 => x"085556fe",
  6048 => x"e4397453",
  6049 => x"807524a7",
  6050 => x"3872822c",
  6051 => x"81712b81",
  6052 => x"fde00807",
  6053 => x"81fddc0b",
  6054 => x"84050c53",
  6055 => x"758c190c",
  6056 => x"7388190c",
  6057 => x"7788170c",
  6058 => x"778c150c",
  6059 => x"fdcd3983",
  6060 => x"1570822c",
  6061 => x"81712b81",
  6062 => x"fde00807",
  6063 => x"81fddc0b",
  6064 => x"84050c51",
  6065 => x"53d63981",
  6066 => x"0bb00c04",
  6067 => x"803d0d72",
  6068 => x"812e8938",
  6069 => x"800bb00c",
  6070 => x"823d0d04",
  6071 => x"7351b23f",
  6072 => x"fe3d0d82",
  6073 => x"9ec80851",
  6074 => x"708a3882",
  6075 => x"9ed07082",
  6076 => x"9ec80c51",
  6077 => x"70751252",
  6078 => x"52ff5370",
  6079 => x"87fb8080",
  6080 => x"26883870",
  6081 => x"829ec80c",
  6082 => x"715372b0",
  6083 => x"0c843d0d",
  6084 => x"0400ff39",
  6085 => x"00000000",
  6086 => x"00000000",
  6087 => x"00000000",
  6088 => x"00000000",
  6089 => x"00cac5ca",
  6090 => x"c5c0c0c0",
  6091 => x"c0c0c0c0",
  6092 => x"c0c0c0cf",
  6093 => x"cfcfcf00",
  6094 => x"00000f0f",
  6095 => x"0f0f8f8f",
  6096 => x"cfcfcfcf",
  6097 => x"cfcf4f0f",
  6098 => x"0f0f0000",
  6099 => x"cfcfcfcf",
  6100 => x"0f0f0f0f",
  6101 => x"0f0f0f0f",
  6102 => x"0f0ffefe",
  6103 => x"fefc0000",
  6104 => x"cfcfcfcf",
  6105 => x"cfcfcfcf",
  6106 => x"cfcfcfcf",
  6107 => x"cfffff7e",
  6108 => x"7e000000",
  6109 => x"00000000",
  6110 => x"00000000",
  6111 => x"00000000",
  6112 => x"00003f3f",
  6113 => x"3f3f0101",
  6114 => x"01010101",
  6115 => x"01010101",
  6116 => x"3f3f3f3f",
  6117 => x"0000383c",
  6118 => x"3e3e3f3f",
  6119 => x"3f3b3b39",
  6120 => x"39383838",
  6121 => x"38383800",
  6122 => x"003f3f3f",
  6123 => x"3f383838",
  6124 => x"38383838",
  6125 => x"38383c3f",
  6126 => x"3f1f0f00",
  6127 => x"003f3f3f",
  6128 => x"3f030303",
  6129 => x"03030303",
  6130 => x"03033f3f",
  6131 => x"3f3e0000",
  6132 => x"00000000",
  6133 => x"00000000",
  6134 => x"00000000",
  6135 => x"00000000",
  6136 => x"00000000",
  6137 => x"00000000",
  6138 => x"00000000",
  6139 => x"00000000",
  6140 => x"00000000",
  6141 => x"00000000",
  6142 => x"00000000",
  6143 => x"00000000",
  6144 => x"00000000",
  6145 => x"00000000",
  6146 => x"00000000",
  6147 => x"00000000",
  6148 => x"00000000",
  6149 => x"00000000",
  6150 => x"00000000",
  6151 => x"00000000",
  6152 => x"00000000",
  6153 => x"00000000",
  6154 => x"00000000",
  6155 => x"00000000",
  6156 => x"8080c0c0",
  6157 => x"e0e06000",
  6158 => x"00000000",
  6159 => x"00000000",
  6160 => x"00000000",
  6161 => x"00000000",
  6162 => x"00000000",
  6163 => x"00000000",
  6164 => x"00000000",
  6165 => x"00000000",
  6166 => x"00000000",
  6167 => x"00000000",
  6168 => x"00000000",
  6169 => x"00000000",
  6170 => x"00000000",
  6171 => x"00000000",
  6172 => x"00000000",
  6173 => x"00000000",
  6174 => x"00000000",
  6175 => x"00000000",
  6176 => x"00000000",
  6177 => x"00000000",
  6178 => x"806098ee",
  6179 => x"77bbddec",
  6180 => x"ee6e0200",
  6181 => x"00000000",
  6182 => x"00e08080",
  6183 => x"e00000e0",
  6184 => x"a0a00000",
  6185 => x"e0000000",
  6186 => x"00e0c000",
  6187 => x"c0e00000",
  6188 => x"e08080e0",
  6189 => x"0000c020",
  6190 => x"20c00000",
  6191 => x"e0000000",
  6192 => x"20e02000",
  6193 => x"0020a060",
  6194 => x"20000000",
  6195 => x"00000000",
  6196 => x"00000000",
  6197 => x"00000000",
  6198 => x"00000000",
  6199 => x"00000000",
  6200 => x"00000000",
  6201 => x"00030007",
  6202 => x"00070701",
  6203 => x"00000000",
  6204 => x"00000000",
  6205 => x"00000300",
  6206 => x"c0030000",
  6207 => x"034242c0",
  6208 => x"00c34242",
  6209 => x"0000c380",
  6210 => x"01c00340",
  6211 => x"c04300c0",
  6212 => x"43408001",
  6213 => x"c20201c0",
  6214 => x"00c38202",
  6215 => x"80c00300",
  6216 => x"00c04342",
  6217 => x"8202c040",
  6218 => x"40800000",
  6219 => x"c0404000",
  6220 => x"80404000",
  6221 => x"00c04040",
  6222 => x"8000c040",
  6223 => x"4000c080",
  6224 => x"00c00000",
  6225 => x"00000000",
  6226 => x"00000000",
  6227 => x"00000000",
  6228 => x"00000000",
  6229 => x"00ff0000",
  6230 => x"0000c645",
  6231 => x"44800785",
  6232 => x"45408007",
  6233 => x"80424700",
  6234 => x"80474000",
  6235 => x"07c14344",
  6236 => x"00c38404",
  6237 => x"c30007c1",
  6238 => x"42418700",
  6239 => x"80404784",
  6240 => x"04c34047",
  6241 => x"8101c640",
  6242 => x"40070505",
  6243 => x"00040502",
  6244 => x"00000704",
  6245 => x"04030007",
  6246 => x"05050007",
  6247 => x"00020700",
  6248 => x"00000000",
  6249 => x"00000000",
  6250 => x"00000000",
  6251 => x"00000000",
  6252 => x"0000ff00",
  6253 => x"00000007",
  6254 => x"01030500",
  6255 => x"03040403",
  6256 => x"00040502",
  6257 => x"00040502",
  6258 => x"00000705",
  6259 => x"05000700",
  6260 => x"02070000",
  6261 => x"07040403",
  6262 => x"00030404",
  6263 => x"03000701",
  6264 => x"03050007",
  6265 => x"01010000",
  6266 => x"00000000",
  6267 => x"00000000",
  6268 => x"00000000",
  6269 => x"00000000",
  6270 => x"00000000",
  6271 => x"71756974",
  6272 => x"00000000",
  6273 => x"68656c70",
  6274 => x"00000000",
  6275 => x"73686f77",
  6276 => x"2042504d",
  6277 => x"20726567",
  6278 => x"69737465",
  6279 => x"72730000",
  6280 => x"62706d00",
  6281 => x"73686f77",
  6282 => x"2044434d",
  6283 => x"20726567",
  6284 => x"69737465",
  6285 => x"72730000",
  6286 => x"64636d00",
  6287 => x"64696167",
  6288 => x"6e6f7365",
  6289 => x"206f7574",
  6290 => x"70757420",
  6291 => x"2b206d6f",
  6292 => x"64652028",
  6293 => x"302d3320",
  6294 => x"73756d20",
  6295 => x"48205629",
  6296 => x"00000000",
  6297 => x"73656c65",
  6298 => x"63740000",
  6299 => x"73797374",
  6300 => x"656d2072",
  6301 => x"65736574",
  6302 => x"00000000",
  6303 => x"72657365",
  6304 => x"74000000",
  6305 => x"73686f77",
  6306 => x"20737973",
  6307 => x"74656d20",
  6308 => x"696e666f",
  6309 => x"203c7665",
  6310 => x"72626f73",
  6311 => x"653e0000",
  6312 => x"73797369",
  6313 => x"6e666f00",
  6314 => x"3c6c6f77",
  6315 => x"65723e20",
  6316 => x"3c757070",
  6317 => x"65723e20",
  6318 => x"73657220",
  6319 => x"44434d20",
  6320 => x"626f756e",
  6321 => x"64730000",
  6322 => x"73686f77",
  6323 => x"2f736574",
  6324 => x"20646562",
  6325 => x"75672072",
  6326 => x"65676973",
  6327 => x"74657273",
  6328 => x"203c7365",
  6329 => x"74206d6f",
  6330 => x"64653e00",
  6331 => x"64656275",
  6332 => x"67000000",
  6333 => x"736f7572",
  6334 => x"63653a20",
  6335 => x"2030203d",
  6336 => x"20696e74",
  6337 => x"2c203120",
  6338 => x"3d206578",
  6339 => x"74000000",
  6340 => x"636c6b00",
  6341 => x"70756c73",
  6342 => x"6520736f",
  6343 => x"75726365",
  6344 => x"3a203020",
  6345 => x"3d207465",
  6346 => x"73746765",
  6347 => x"6e2c2031",
  6348 => x"203d2065",
  6349 => x"78740000",
  6350 => x"6d696372",
  6351 => x"6f000000",
  6352 => x"74657374",
  6353 => x"67656e65",
  6354 => x"7261746f",
  6355 => x"72203c73",
  6356 => x"63616c65",
  6357 => x"723e203c",
  6358 => x"72657374",
  6359 => x"6172743e",
  6360 => x"00000000",
  6361 => x"74657374",
  6362 => x"67656e00",
  6363 => x"3c6d7574",
  6364 => x"655f6e3e",
  6365 => x"203c7273",
  6366 => x"745f6e3e",
  6367 => x"203c6270",
  6368 => x"625f6e3e",
  6369 => x"203c6f73",
  6370 => x"72313e20",
  6371 => x"3c6f7372",
  6372 => x"323e0000",
  6373 => x"64616363",
  6374 => x"6f6e6600",
  6375 => x"3c6d756c",
  6376 => x"7469706c",
  6377 => x"6965723e",
  6378 => x"20696e69",
  6379 => x"7469616c",
  6380 => x"697a6520",
  6381 => x"62756666",
  6382 => x"65720000",
  6383 => x"64616374",
  6384 => x"65737400",
  6385 => x"72657365",
  6386 => x"74204250",
  6387 => x"4d206361",
  6388 => x"6c63756c",
  6389 => x"6174696f",
  6390 => x"6e206572",
  6391 => x"726f7273",
  6392 => x"00000000",
  6393 => x"62706d72",
  6394 => x"65730000",
  6395 => x"72657365",
  6396 => x"74204443",
  6397 => x"4d206572",
  6398 => x"726f7273",
  6399 => x"00000000",
  6400 => x"64636d72",
  6401 => x"65730000",
  6402 => x"73686f77",
  6403 => x"20646562",
  6404 => x"75672062",
  6405 => x"75666665",
  6406 => x"72203c6c",
  6407 => x"656e6774",
  6408 => x"683e0000",
  6409 => x"636c6561",
  6410 => x"72206465",
  6411 => x"62756720",
  6412 => x"62756666",
  6413 => x"65720000",
  6414 => x"62636c65",
  6415 => x"61720000",
  6416 => x"646f776e",
  6417 => x"6c6f6164",
  6418 => x"20646562",
  6419 => x"75672062",
  6420 => x"75666665",
  6421 => x"72202878",
  6422 => x"6d6f6465",
  6423 => x"6d290000",
  6424 => x"62726561",
  6425 => x"64000000",
  6426 => x"75706c6f",
  6427 => x"61642064",
  6428 => x"65627567",
  6429 => x"20627566",
  6430 => x"66657220",
  6431 => x"28786d6f",
  6432 => x"64656d29",
  6433 => x"00000000",
  6434 => x"62777269",
  6435 => x"74650000",
  6436 => x"62756666",
  6437 => x"6572206f",
  6438 => x"6e204c43",
  6439 => x"44203c63",
  6440 => x"683e203c",
  6441 => x"636f6d62",
  6442 => x"3e000000",
  6443 => x"73636f70",
  6444 => x"65000000",
  6445 => x"64656275",
  6446 => x"67207472",
  6447 => x"61636520",
  6448 => x"3c636c65",
  6449 => x"61723e00",
  6450 => x"74726163",
  6451 => x"65000000",
  6452 => x"73657475",
  6453 => x"70206368",
  6454 => x"616e6e65",
  6455 => x"6c207465",
  6456 => x"7374203c",
  6457 => x"63683e20",
  6458 => x"3c76616c",
  6459 => x"302e2e37",
  6460 => x"3e000000",
  6461 => x"63687465",
  6462 => x"73740000",
  6463 => x"72756e6e",
  6464 => x"696e6720",
  6465 => x"6c696768",
  6466 => x"74000000",
  6467 => x"72756e00",
  6468 => x"72756e20",
  6469 => x"64697370",
  6470 => x"6c617920",
  6471 => x"74657374",
  6472 => x"2066756e",
  6473 => x"6374696f",
  6474 => x"6e000000",
  6475 => x"64697370",
  6476 => x"6c617900",
  6477 => x"73657420",
  6478 => x"6261636b",
  6479 => x"6c696768",
  6480 => x"74203c30",
  6481 => x"2e2e3331",
  6482 => x"3e000000",
  6483 => x"6261636b",
  6484 => x"00000000",
  6485 => x"73686f77",
  6486 => x"206c6f67",
  6487 => x"6f206f6e",
  6488 => x"20676c63",
  6489 => x"64000000",
  6490 => x"6c6f676f",
  6491 => x"00000000",
  6492 => x"63686563",
  6493 => x"6b204932",
  6494 => x"43206164",
  6495 => x"64726573",
  6496 => x"73000000",
  6497 => x"69326300",
  6498 => x"72656164",
  6499 => x"20454550",
  6500 => x"524f4d20",
  6501 => x"3c627573",
  6502 => x"3e203c69",
  6503 => x"32635f61",
  6504 => x"6464723e",
  6505 => x"203c6c65",
  6506 => x"6e677468",
  6507 => x"3e000000",
  6508 => x"65657072",
  6509 => x"6f6d0000",
  6510 => x"41444320",
  6511 => x"72656769",
  6512 => x"73746572",
  6513 => x"20747261",
  6514 => x"6e736665",
  6515 => x"72203c76",
  6516 => x"616c7565",
  6517 => x"3e000000",
  6518 => x"61747261",
  6519 => x"6e730000",
  6520 => x"696e6974",
  6521 => x"20414443",
  6522 => x"20726567",
  6523 => x"69737465",
  6524 => x"72730000",
  6525 => x"61696e69",
  6526 => x"74000000",
  6527 => x"72656164",
  6528 => x"20636872",
  6529 => x"6f6e7465",
  6530 => x"6c207265",
  6531 => x"67697374",
  6532 => x"65727300",
  6533 => x"63726561",
  6534 => x"64000000",
  6535 => x"696e6974",
  6536 => x"20636872",
  6537 => x"6f6e7465",
  6538 => x"6c207265",
  6539 => x"67697374",
  6540 => x"65727300",
  6541 => x"63696e69",
  6542 => x"74000000",
  6543 => x"77726974",
  6544 => x"65206368",
  6545 => x"726f6e74",
  6546 => x"656c2072",
  6547 => x"65676973",
  6548 => x"74657220",
  6549 => x"3c726567",
  6550 => x"3e203c76",
  6551 => x"616c7565",
  6552 => x"3e000000",
  6553 => x"63777269",
  6554 => x"74650000",
  6555 => x"616c6961",
  6556 => x"7320666f",
  6557 => x"72207800",
  6558 => x"6d656d00",
  6559 => x"77726974",
  6560 => x"6520776f",
  6561 => x"7264203c",
  6562 => x"61646472",
  6563 => x"3e203c6c",
  6564 => x"656e6774",
  6565 => x"683e203c",
  6566 => x"76616c75",
  6567 => x"65287329",
  6568 => x"3e000000",
  6569 => x"776d656d",
  6570 => x"00000000",
  6571 => x"6558616d",
  6572 => x"696e6520",
  6573 => x"6d656d6f",
  6574 => x"7279203c",
  6575 => x"61646472",
  6576 => x"3e203c6c",
  6577 => x"656e6774",
  6578 => x"683e0000",
  6579 => x"636c6561",
  6580 => x"72207363",
  6581 => x"7265656e",
  6582 => x"00000000",
  6583 => x"636c6561",
  6584 => x"72000000",
  6585 => x"65787465",
  6586 => x"726e616c",
  6587 => x"20636c6f",
  6588 => x"636b2000",
  6589 => x"61637469",
  6590 => x"76650a00",
  6591 => x"73656c65",
  6592 => x"63746564",
  6593 => x"0a000000",
  6594 => x"4e4f5420",
  6595 => x"00000000",
  6596 => x"6d696372",
  6597 => x"6f70756c",
  6598 => x"73652073",
  6599 => x"6f757263",
  6600 => x"653a2000",
  6601 => x"65787465",
  6602 => x"726e616c",
  6603 => x"00000000",
  6604 => x"6265616d",
  6605 => x"20706f73",
  6606 => x"6974696f",
  6607 => x"6e206d6f",
  6608 => x"6e69746f",
  6609 => x"72000000",
  6610 => x"0a0a0000",
  6611 => x"20286f6e",
  6612 => x"2073696d",
  6613 => x"290a0000",
  6614 => x"0a485720",
  6615 => x"73796e74",
  6616 => x"68657369",
  6617 => x"7a65643a",
  6618 => x"20000000",
  6619 => x"0a535720",
  6620 => x"636f6d70",
  6621 => x"696c6564",
  6622 => x"2020203a",
  6623 => x"20536570",
  6624 => x"20203920",
  6625 => x"32303131",
  6626 => x"20203134",
  6627 => x"3a31363a",
  6628 => x"34340000",
  6629 => x"0a737973",
  6630 => x"74656d20",
  6631 => x"636c6f63",
  6632 => x"6b20203a",
  6633 => x"20000000",
  6634 => x"204d487a",
  6635 => x"0a000000",
  6636 => x"44454255",
  6637 => x"47204d4f",
  6638 => x"44450000",
  6639 => x"20282b44",
  6640 => x"56492900",
  6641 => x"20282b64",
  6642 => x"65627567",
  6643 => x"20627566",
  6644 => x"66657220",
  6645 => x"7472616e",
  6646 => x"73666572",
  6647 => x"29000000",
  6648 => x"204f4e0a",
  6649 => x"00000000",
  6650 => x"6265616d",
  6651 => x"20706f73",
  6652 => x"6974696f",
  6653 => x"6e206d6f",
  6654 => x"6e69746f",
  6655 => x"720a0000",
  6656 => x"0a536570",
  6657 => x"20203920",
  6658 => x"32303131",
  6659 => x"20203134",
  6660 => x"3a31363a",
  6661 => x"34340000",
  6662 => x"0a696e69",
  6663 => x"74204144",
  6664 => x"43000000",
  6665 => x"0a696e69",
  6666 => x"7420434c",
  6667 => x"4b000000",
  6668 => x"0a696e69",
  6669 => x"74204441",
  6670 => x"43000000",
  6671 => x"0a696e69",
  6672 => x"74204250",
  6673 => x"4d000000",
  6674 => x"202d2d3e",
  6675 => x"20455252",
  6676 => x"4f520000",
  6677 => x"4552524f",
  6678 => x"523a2074",
  6679 => x"6f6f206d",
  6680 => x"75636820",
  6681 => x"636f6d6d",
  6682 => x"616e6473",
  6683 => x"2e0a0000",
  6684 => x"3e200000",
  6685 => x"636f6d6d",
  6686 => x"616e6420",
  6687 => x"6e6f7420",
  6688 => x"666f756e",
  6689 => x"642e0a00",
  6690 => x"73757070",
  6691 => x"6f727465",
  6692 => x"6420636f",
  6693 => x"6d6d616e",
  6694 => x"64733a0a",
  6695 => x"0a000000",
  6696 => x"202d2000",
  6697 => x"76656e64",
  6698 => x"6f723f20",
  6699 => x"20000000",
  6700 => x"485a4452",
  6701 => x"20202020",
  6702 => x"20000000",
  6703 => x"67616973",
  6704 => x"6c657220",
  6705 => x"20000000",
  6706 => x"4148422f",
  6707 => x"41504220",
  6708 => x"42726964",
  6709 => x"67650000",
  6710 => x"45534120",
  6711 => x"20202020",
  6712 => x"20000000",
  6713 => x"756e6b6e",
  6714 => x"6f776e20",
  6715 => x"64657669",
  6716 => x"63650000",
  6717 => x"4c656f6e",
  6718 => x"32204d65",
  6719 => x"6d6f7279",
  6720 => x"20436f6e",
  6721 => x"74726f6c",
  6722 => x"6c657200",
  6723 => x"47522031",
  6724 => x"302f3130",
  6725 => x"30204d62",
  6726 => x"69742045",
  6727 => x"74686572",
  6728 => x"6e657420",
  6729 => x"4d414300",
  6730 => x"64696666",
  6731 => x"6572656e",
  6732 => x"7469616c",
  6733 => x"20637572",
  6734 => x"72656e74",
  6735 => x"206d6f6e",
  6736 => x"69746f72",
  6737 => x"00000000",
  6738 => x"64656275",
  6739 => x"67207472",
  6740 => x"61636572",
  6741 => x"206d656d",
  6742 => x"6f727900",
  6743 => x"4541444f",
  6744 => x"47533130",
  6745 => x"32206469",
  6746 => x"73706c61",
  6747 => x"79206472",
  6748 => x"69766572",
  6749 => x"00000000",
  6750 => x"64656275",
  6751 => x"67206275",
  6752 => x"66666572",
  6753 => x"20636f6e",
  6754 => x"74726f6c",
  6755 => x"00000000",
  6756 => x"74726967",
  6757 => x"67657220",
  6758 => x"67656e65",
  6759 => x"7261746f",
  6760 => x"72000000",
  6761 => x"64656275",
  6762 => x"6720636f",
  6763 => x"6e736f6c",
  6764 => x"65000000",
  6765 => x"44434d20",
  6766 => x"70686173",
  6767 => x"65207368",
  6768 => x"69667420",
  6769 => x"636f6e74",
  6770 => x"726f6c00",
  6771 => x"5a505520",
  6772 => x"4d656d6f",
  6773 => x"72792077",
  6774 => x"72617070",
  6775 => x"65720000",
  6776 => x"5a505520",
  6777 => x"41484220",
  6778 => x"57726170",
  6779 => x"70657200",
  6780 => x"56474120",
  6781 => x"636f6e74",
  6782 => x"726f6c6c",
  6783 => x"65720000",
  6784 => x"4d6f6475",
  6785 => x"6c617220",
  6786 => x"54696d65",
  6787 => x"7220556e",
  6788 => x"69740000",
  6789 => x"47656e65",
  6790 => x"72616c20",
  6791 => x"50757270",
  6792 => x"6f736520",
  6793 => x"492f4f20",
  6794 => x"706f7274",
  6795 => x"00000000",
  6796 => x"47656e65",
  6797 => x"72696320",
  6798 => x"55415254",
  6799 => x"00000000",
  6800 => x"414d4241",
  6801 => x"20577261",
  6802 => x"70706572",
  6803 => x"20666f72",
  6804 => x"204f4320",
  6805 => x"4932432d",
  6806 => x"6d617374",
  6807 => x"65720000",
  6808 => x"53504920",
  6809 => x"4d656d6f",
  6810 => x"72792043",
  6811 => x"6f6e7472",
  6812 => x"6f6c6c65",
  6813 => x"72000000",
  6814 => x"4475616c",
  6815 => x"2d706f72",
  6816 => x"74204148",
  6817 => x"42205352",
  6818 => x"414d206d",
  6819 => x"6f64756c",
  6820 => x"65000000",
  6821 => x"20206170",
  6822 => x"62736c76",
  6823 => x"00000000",
  6824 => x"76656e64",
  6825 => x"20307800",
  6826 => x"64657620",
  6827 => x"30780000",
  6828 => x"76657220",
  6829 => x"00000000",
  6830 => x"69727120",
  6831 => x"00000000",
  6832 => x"61646472",
  6833 => x"20307800",
  6834 => x"6168626d",
  6835 => x"73740000",
  6836 => x"61686273",
  6837 => x"6c760000",
  6838 => x"000018db",
  6839 => x"0000197f",
  6840 => x"00001973",
  6841 => x"00001967",
  6842 => x"0000195b",
  6843 => x"0000194f",
  6844 => x"00001943",
  6845 => x"00001937",
  6846 => x"0000192b",
  6847 => x"0000191f",
  6848 => x"00001913",
  6849 => x"04580808",
  6850 => x"20ff0000",
  6851 => x"00006b14",
  6852 => x"00006bf4",
  6853 => x"02010305",
  6854 => x"05070501",
  6855 => x"03030505",
  6856 => x"02030104",
  6857 => x"05050505",
  6858 => x"05050505",
  6859 => x"05050101",
  6860 => x"04050404",
  6861 => x"07050505",
  6862 => x"05050505",
  6863 => x"05030405",
  6864 => x"05050505",
  6865 => x"05050505",
  6866 => x"05050505",
  6867 => x"05050503",
  6868 => x"04030505",
  6869 => x"02050504",
  6870 => x"05050405",
  6871 => x"04010204",
  6872 => x"02050404",
  6873 => x"05050404",
  6874 => x"04040507",
  6875 => x"05040404",
  6876 => x"02040500",
  6877 => x"04050200",
  6878 => x"04080303",
  6879 => x"04090003",
  6880 => x"06000000",
  6881 => x"00020204",
  6882 => x"04040400",
  6883 => x"04060003",
  6884 => x"05000000",
  6885 => x"00000404",
  6886 => x"05050204",
  6887 => x"05060305",
  6888 => x"04030705",
  6889 => x"04050303",
  6890 => x"02040502",
  6891 => x"03020405",
  6892 => x"06060604",
  6893 => x"05050505",
  6894 => x"05050504",
  6895 => x"04040404",
  6896 => x"03030303",
  6897 => x"05050505",
  6898 => x"05050505",
  6899 => x"05040404",
  6900 => x"04050404",
  6901 => x"04040404",
  6902 => x"04040503",
  6903 => x"04040404",
  6904 => x"02020303",
  6905 => x"04040404",
  6906 => x"04040405",
  6907 => x"04040404",
  6908 => x"04030303",
  6909 => x"00005f07",
  6910 => x"0007741c",
  6911 => x"771c172e",
  6912 => x"6a3e2b3a",
  6913 => x"06493608",
  6914 => x"36493036",
  6915 => x"49597648",
  6916 => x"073c4281",
  6917 => x"81423c0a",
  6918 => x"041f040a",
  6919 => x"08083e08",
  6920 => x"08806008",
  6921 => x"080840c0",
  6922 => x"300c033e",
  6923 => x"4141413e",
  6924 => x"44427f40",
  6925 => x"40466151",
  6926 => x"49462241",
  6927 => x"49493618",
  6928 => x"14127f10",
  6929 => x"27454545",
  6930 => x"393e4949",
  6931 => x"49300101",
  6932 => x"710d0336",
  6933 => x"49494936",
  6934 => x"06494929",
  6935 => x"1e36d008",
  6936 => x"14224114",
  6937 => x"14141414",
  6938 => x"41221408",
  6939 => x"02510906",
  6940 => x"3c4299a5",
  6941 => x"bd421c7c",
  6942 => x"1211127c",
  6943 => x"7f494949",
  6944 => x"363e4141",
  6945 => x"41227f41",
  6946 => x"41413e7f",
  6947 => x"49494941",
  6948 => x"7f090909",
  6949 => x"013e4149",
  6950 => x"497a7f08",
  6951 => x"08087f41",
  6952 => x"7f414041",
  6953 => x"413f7f08",
  6954 => x"1422417f",
  6955 => x"40404040",
  6956 => x"7f060c06",
  6957 => x"7f7f0608",
  6958 => x"307f3e41",
  6959 => x"41413e7f",
  6960 => x"09090906",
  6961 => x"3e4161c1",
  6962 => x"be7f0919",
  6963 => x"29462649",
  6964 => x"49493201",
  6965 => x"017f0101",
  6966 => x"3f404040",
  6967 => x"3f073840",
  6968 => x"38071f60",
  6969 => x"1f601f63",
  6970 => x"14081463",
  6971 => x"01067806",
  6972 => x"01615149",
  6973 => x"45437f41",
  6974 => x"41030c30",
  6975 => x"c041417f",
  6976 => x"04020102",
  6977 => x"04808080",
  6978 => x"80800102",
  6979 => x"20545454",
  6980 => x"787f4444",
  6981 => x"44383844",
  6982 => x"44443844",
  6983 => x"44447f38",
  6984 => x"54545458",
  6985 => x"087e0901",
  6986 => x"18a4a4a4",
  6987 => x"787f0404",
  6988 => x"787d807d",
  6989 => x"7f102844",
  6990 => x"3f407c04",
  6991 => x"7804787c",
  6992 => x"04047838",
  6993 => x"444438fc",
  6994 => x"24242418",
  6995 => x"18242424",
  6996 => x"fc7c0804",
  6997 => x"04485454",
  6998 => x"24043f44",
  6999 => x"403c4040",
  7000 => x"7c1c2040",
  7001 => x"201c1c60",
  7002 => x"601c6060",
  7003 => x"1c442810",
  7004 => x"28449ca0",
  7005 => x"601c6454",
  7006 => x"544c187e",
  7007 => x"8181ffff",
  7008 => x"81817e18",
  7009 => x"18040810",
  7010 => x"0c143e55",
  7011 => x"55ff8181",
  7012 => x"81ff8060",
  7013 => x"80608060",
  7014 => x"60600060",
  7015 => x"60006060",
  7016 => x"047f0414",
  7017 => x"7f140201",
  7018 => x"01024629",
  7019 => x"1608344a",
  7020 => x"31483000",
  7021 => x"18243e41",
  7022 => x"227f4941",
  7023 => x"03040403",
  7024 => x"03040304",
  7025 => x"04030403",
  7026 => x"183c3c18",
  7027 => x"08080808",
  7028 => x"03010203",
  7029 => x"020e020e",
  7030 => x"060e0048",
  7031 => x"30384438",
  7032 => x"54483844",
  7033 => x"fe44487e",
  7034 => x"49014438",
  7035 => x"28384403",
  7036 => x"147c1403",
  7037 => x"e7e74e55",
  7038 => x"55390101",
  7039 => x"0001011c",
  7040 => x"2a555522",
  7041 => x"1c1d151e",
  7042 => x"18240018",
  7043 => x"24080808",
  7044 => x"18080808",
  7045 => x"3c42bd95",
  7046 => x"a9423c01",
  7047 => x"01010101",
  7048 => x"06090906",
  7049 => x"44445f44",
  7050 => x"44191512",
  7051 => x"15150a02",
  7052 => x"01fc2020",
  7053 => x"1c0e7f01",
  7054 => x"7f011818",
  7055 => x"00804002",
  7056 => x"1f060909",
  7057 => x"06241800",
  7058 => x"2418824f",
  7059 => x"304c62f1",
  7060 => x"824f300c",
  7061 => x"d2b1955f",
  7062 => x"304c62f1",
  7063 => x"30484520",
  7064 => x"60392e38",
  7065 => x"6060382e",
  7066 => x"3960701d",
  7067 => x"131d7072",
  7068 => x"1d121e71",
  7069 => x"701d121d",
  7070 => x"70603b25",
  7071 => x"3b607e11",
  7072 => x"7f49411e",
  7073 => x"2161927c",
  7074 => x"5556447c",
  7075 => x"5655447c",
  7076 => x"5655467d",
  7077 => x"54544545",
  7078 => x"7e44447e",
  7079 => x"45467d46",
  7080 => x"457c4508",
  7081 => x"7f49413e",
  7082 => x"7e091222",
  7083 => x"7d384546",
  7084 => x"44383844",
  7085 => x"46453838",
  7086 => x"46454638",
  7087 => x"3a454546",
  7088 => x"39384544",
  7089 => x"45382214",
  7090 => x"081422bc",
  7091 => x"625a463d",
  7092 => x"3c41423c",
  7093 => x"3c42413c",
  7094 => x"3c42413e",
  7095 => x"3d40403d",
  7096 => x"0608f209",
  7097 => x"067f2222",
  7098 => x"1cfe0989",
  7099 => x"76205556",
  7100 => x"78205655",
  7101 => x"78225555",
  7102 => x"7a235556",
  7103 => x"7b205554",
  7104 => x"79275557",
  7105 => x"78205438",
  7106 => x"54483844",
  7107 => x"c4385556",
  7108 => x"58385655",
  7109 => x"583a5555",
  7110 => x"5a395454",
  7111 => x"59017a7a",
  7112 => x"01027902",
  7113 => x"02780260",
  7114 => x"91927c7b",
  7115 => x"090a7338",
  7116 => x"45463838",
  7117 => x"4645383a",
  7118 => x"45453a3b",
  7119 => x"45463b39",
  7120 => x"44443908",
  7121 => x"082a0808",
  7122 => x"b8644c3a",
  7123 => x"3c41427c",
  7124 => x"3c42417c",
  7125 => x"3a41417a",
  7126 => x"3d40407d",
  7127 => x"986219ff",
  7128 => x"423c9a60",
  7129 => x"1a000000",
  7130 => x"69326320",
  7131 => x"4456490a",
  7132 => x"00000000",
  7133 => x"69326320",
  7134 => x"464d430a",
  7135 => x"00000000",
  7136 => x"61646472",
  7137 => x"6573733a",
  7138 => x"20307800",
  7139 => x"2020202d",
  7140 => x"2d3e2020",
  7141 => x"2041434b",
  7142 => x"0a000000",
  7143 => x"72656164",
  7144 => x"20646174",
  7145 => x"61202800",
  7146 => x"20627974",
  7147 => x"65732920",
  7148 => x"66726f6d",
  7149 => x"20493243",
  7150 => x"2d616464",
  7151 => x"72657373",
  7152 => x"20307800",
  7153 => x"6e6f6163",
  7154 => x"6b200000",
  7155 => x"6368726f",
  7156 => x"6e74656c",
  7157 => x"20726567",
  7158 => x"20307800",
  7159 => x"3a203078",
  7160 => x"00000000",
  7161 => x"206e6163",
  7162 => x"6b000000",
  7163 => x"6572726f",
  7164 => x"7220286e",
  7165 => x"61636b29",
  7166 => x"0a000000",
  7167 => x"0a202063",
  7168 => x"68616e6e",
  7169 => x"656c2033",
  7170 => x"20696e70",
  7171 => x"7574206f",
  7172 => x"76657266",
  7173 => x"6c6f7700",
  7174 => x"0a202063",
  7175 => x"68616e6e",
  7176 => x"656c2032",
  7177 => x"20696e70",
  7178 => x"7574206f",
  7179 => x"76657266",
  7180 => x"6c6f7700",
  7181 => x"0a202063",
  7182 => x"68616e6e",
  7183 => x"656c2031",
  7184 => x"20696e70",
  7185 => x"7574206f",
  7186 => x"76657266",
  7187 => x"6c6f7700",
  7188 => x"0a202063",
  7189 => x"68616e6e",
  7190 => x"656c2030",
  7191 => x"20696e70",
  7192 => x"7574206f",
  7193 => x"76657266",
  7194 => x"6c6f7700",
  7195 => x"0a202063",
  7196 => x"68616e6e",
  7197 => x"656c2033",
  7198 => x"20717561",
  7199 => x"6473756d",
  7200 => x"206f7665",
  7201 => x"72666c6f",
  7202 => x"77000000",
  7203 => x"0a202063",
  7204 => x"68616e6e",
  7205 => x"656c2032",
  7206 => x"20717561",
  7207 => x"6473756d",
  7208 => x"206f7665",
  7209 => x"72666c6f",
  7210 => x"77000000",
  7211 => x"0a202063",
  7212 => x"68616e6e",
  7213 => x"656c2031",
  7214 => x"20717561",
  7215 => x"6473756d",
  7216 => x"206f7665",
  7217 => x"72666c6f",
  7218 => x"77000000",
  7219 => x"0a202063",
  7220 => x"68616e6e",
  7221 => x"656c2030",
  7222 => x"20717561",
  7223 => x"6473756d",
  7224 => x"206f7665",
  7225 => x"72666c6f",
  7226 => x"77000000",
  7227 => x"0a202073",
  7228 => x"756d2073",
  7229 => x"63616c65",
  7230 => x"72206f76",
  7231 => x"6572666c",
  7232 => x"6f770000",
  7233 => x"0a202073",
  7234 => x"756d2076",
  7235 => x"616c7565",
  7236 => x"20637574",
  7237 => x"74656400",
  7238 => x"0a202063",
  7239 => x"68616e6e",
  7240 => x"656c2033",
  7241 => x"20646976",
  7242 => x"6964656e",
  7243 => x"64206375",
  7244 => x"74746564",
  7245 => x"00000000",
  7246 => x"0a202063",
  7247 => x"68616e6e",
  7248 => x"656c2033",
  7249 => x"206e6f69",
  7250 => x"73652063",
  7251 => x"6f6d7065",
  7252 => x"6e736174",
  7253 => x"696f6e20",
  7254 => x"746f2062",
  7255 => x"69670000",
  7256 => x"0a202063",
  7257 => x"68616e6e",
  7258 => x"656c2033",
  7259 => x"206e6f69",
  7260 => x"73652076",
  7261 => x"616c7565",
  7262 => x"20637574",
  7263 => x"74656400",
  7264 => x"0a202063",
  7265 => x"68616e6e",
  7266 => x"656c2032",
  7267 => x"20646976",
  7268 => x"6964656e",
  7269 => x"64206375",
  7270 => x"74746564",
  7271 => x"00000000",
  7272 => x"0a202063",
  7273 => x"68616e6e",
  7274 => x"656c2032",
  7275 => x"206e6f69",
  7276 => x"73652063",
  7277 => x"6f6d7065",
  7278 => x"6e736174",
  7279 => x"696f6e20",
  7280 => x"746f2062",
  7281 => x"69670000",
  7282 => x"0a202063",
  7283 => x"68616e6e",
  7284 => x"656c2032",
  7285 => x"206e6f69",
  7286 => x"73652076",
  7287 => x"616c7565",
  7288 => x"20637574",
  7289 => x"74656400",
  7290 => x"0a202063",
  7291 => x"68616e6e",
  7292 => x"656c2031",
  7293 => x"20646976",
  7294 => x"6964656e",
  7295 => x"64206375",
  7296 => x"74746564",
  7297 => x"00000000",
  7298 => x"0a202063",
  7299 => x"68616e6e",
  7300 => x"656c2031",
  7301 => x"206e6f69",
  7302 => x"73652063",
  7303 => x"6f6d7065",
  7304 => x"6e736174",
  7305 => x"696f6e20",
  7306 => x"746f2062",
  7307 => x"69670000",
  7308 => x"0a202063",
  7309 => x"68616e6e",
  7310 => x"656c2031",
  7311 => x"206e6f69",
  7312 => x"73652076",
  7313 => x"616c7565",
  7314 => x"20637574",
  7315 => x"74656400",
  7316 => x"0a202063",
  7317 => x"68616e6e",
  7318 => x"656c2030",
  7319 => x"20646976",
  7320 => x"6964656e",
  7321 => x"64206375",
  7322 => x"74746564",
  7323 => x"00000000",
  7324 => x"0a202063",
  7325 => x"68616e6e",
  7326 => x"656c2030",
  7327 => x"206e6f69",
  7328 => x"73652063",
  7329 => x"6f6d7065",
  7330 => x"6e736174",
  7331 => x"696f6e20",
  7332 => x"746f2062",
  7333 => x"69670000",
  7334 => x"0a202063",
  7335 => x"68616e6e",
  7336 => x"656c2030",
  7337 => x"206e6f69",
  7338 => x"73652076",
  7339 => x"616c7565",
  7340 => x"20637574",
  7341 => x"74656400",
  7342 => x"0a202073",
  7343 => x"6f667477",
  7344 => x"61726520",
  7345 => x"6572726f",
  7346 => x"72000000",
  7347 => x"0a657874",
  7348 => x"65726e61",
  7349 => x"6c20636c",
  7350 => x"6f636b20",
  7351 => x"20202020",
  7352 => x"2020203a",
  7353 => x"20000000",
  7354 => x"61637469",
  7355 => x"76650000",
  7356 => x"0a6d6963",
  7357 => x"726f7075",
  7358 => x"6c736520",
  7359 => x"736f7572",
  7360 => x"63652020",
  7361 => x"2020203a",
  7362 => x"20000000",
  7363 => x"0a6d6963",
  7364 => x"726f7075",
  7365 => x"6c736520",
  7366 => x"6576656e",
  7367 => x"74206c69",
  7368 => x"6d69743a",
  7369 => x"20000000",
  7370 => x"0a6d6561",
  7371 => x"73757265",
  7372 => x"6d656e74",
  7373 => x"206c656e",
  7374 => x"67746820",
  7375 => x"2020203a",
  7376 => x"20000000",
  7377 => x"0a626561",
  7378 => x"6d20706f",
  7379 => x"73697469",
  7380 => x"6f6e206d",
  7381 => x"6f6e6974",
  7382 => x"6f722072",
  7383 => x"65676973",
  7384 => x"74657273",
  7385 => x"00000000",
  7386 => x"0a202020",
  7387 => x"20202020",
  7388 => x"20202020",
  7389 => x"20202020",
  7390 => x"20202020",
  7391 => x"20202020",
  7392 => x"20636861",
  7393 => x"6e6e656c",
  7394 => x"20302020",
  7395 => x"20636861",
  7396 => x"6e6e656c",
  7397 => x"20312020",
  7398 => x"20636861",
  7399 => x"6e6e656c",
  7400 => x"20322020",
  7401 => x"20636861",
  7402 => x"6e6e656c",
  7403 => x"20330000",
  7404 => x"0a202020",
  7405 => x"20202020",
  7406 => x"20202020",
  7407 => x"20202020",
  7408 => x"20202020",
  7409 => x"20202020",
  7410 => x"202d2d2d",
  7411 => x"2d20686f",
  7412 => x"72697a6f",
  7413 => x"6e74616c",
  7414 => x"202d2d2d",
  7415 => x"2d2d2020",
  7416 => x"202d2d2d",
  7417 => x"2d2d2d20",
  7418 => x"76657274",
  7419 => x"6963616c",
  7420 => x"202d2d2d",
  7421 => x"2d2d0000",
  7422 => x"0a736361",
  7423 => x"6c657220",
  7424 => x"76616c75",
  7425 => x"65732020",
  7426 => x"20202020",
  7427 => x"20202020",
  7428 => x"20000000",
  7429 => x"0a6e6f69",
  7430 => x"73652063",
  7431 => x"6f6d7065",
  7432 => x"6e736174",
  7433 => x"696f6e20",
  7434 => x"20202020",
  7435 => x"20000000",
  7436 => x"0a6d6561",
  7437 => x"73757265",
  7438 => x"6d656e74",
  7439 => x"20202020",
  7440 => x"20202020",
  7441 => x"20202020",
  7442 => x"20000000",
  7443 => x"0a73616d",
  7444 => x"706c6573",
  7445 => x"20286469",
  7446 => x"76292020",
  7447 => x"20202020",
  7448 => x"3a200000",
  7449 => x"0a73756d",
  7450 => x"20636861",
  7451 => x"6e6e656c",
  7452 => x"20736361",
  7453 => x"6c657220",
  7454 => x"3a200000",
  7455 => x"0a73756d",
  7456 => x"20636861",
  7457 => x"6e6e656c",
  7458 => x"20202020",
  7459 => x"20202020",
  7460 => x"3a200000",
  7461 => x"0a0a706f",
  7462 => x"73697469",
  7463 => x"6f6e2063",
  7464 => x"6f6d7075",
  7465 => x"74617469",
  7466 => x"6f6e0000",
  7467 => x"0a202073",
  7468 => x"63616c65",
  7469 => x"72207661",
  7470 => x"6c756573",
  7471 => x"20202020",
  7472 => x"20202020",
  7473 => x"20000000",
  7474 => x"0a20206f",
  7475 => x"66667365",
  7476 => x"74202020",
  7477 => x"20202020",
  7478 => x"20202020",
  7479 => x"20202020",
  7480 => x"20000000",
  7481 => x"0a6f7574",
  7482 => x"70757420",
  7483 => x"73656c65",
  7484 => x"6374203a",
  7485 => x"20000000",
  7486 => x"64697265",
  7487 => x"6374206d",
  7488 => x"6f646500",
  7489 => x"0a63616c",
  7490 => x"63207374",
  7491 => x"61746520",
  7492 => x"2020203a",
  7493 => x"20307800",
  7494 => x"76657274",
  7495 => x"6963616c",
  7496 => x"00000000",
  7497 => x"686f7269",
  7498 => x"7a6f6e74",
  7499 => x"616c0000",
  7500 => x"73756d00",
  7501 => x"6368616e",
  7502 => x"6e656c20",
  7503 => x"33000000",
  7504 => x"6368616e",
  7505 => x"6e656c20",
  7506 => x"32000000",
  7507 => x"6368616e",
  7508 => x"6e656c20",
  7509 => x"31000000",
  7510 => x"6368616e",
  7511 => x"6e656c20",
  7512 => x"30000000",
  7513 => x"636c6b3a",
  7514 => x"20000000",
  7515 => x"494e5400",
  7516 => x"6d70756c",
  7517 => x"733a2000",
  7518 => x"65787400",
  7519 => x"0a6d6561",
  7520 => x"732e206c",
  7521 => x"656e6774",
  7522 => x"683a2000",
  7523 => x"0a636830",
  7524 => x"3a200000",
  7525 => x"6368313a",
  7526 => x"20000000",
  7527 => x"0a636832",
  7528 => x"3a200000",
  7529 => x"6368333a",
  7530 => x"20000000",
  7531 => x"0a73706c",
  7532 => x"3a200000",
  7533 => x"73756d3a",
  7534 => x"20000000",
  7535 => x"0a6f7574",
  7536 => x"7075743a",
  7537 => x"20000000",
  7538 => x"7467656e",
  7539 => x"00000000",
  7540 => x"0a63616c",
  7541 => x"63207374",
  7542 => x"6174653a",
  7543 => x"20000000",
  7544 => x"63683320",
  7545 => x"696e7020",
  7546 => x"6f762020",
  7547 => x"00000000",
  7548 => x"63683220",
  7549 => x"696e7020",
  7550 => x"6f762020",
  7551 => x"00000000",
  7552 => x"63683120",
  7553 => x"696e7020",
  7554 => x"6f762020",
  7555 => x"00000000",
  7556 => x"63683020",
  7557 => x"696e7020",
  7558 => x"6f762020",
  7559 => x"00000000",
  7560 => x"63683320",
  7561 => x"73756d20",
  7562 => x"6f762020",
  7563 => x"00000000",
  7564 => x"63683220",
  7565 => x"73756d20",
  7566 => x"6f762020",
  7567 => x"00000000",
  7568 => x"63683120",
  7569 => x"73756d20",
  7570 => x"6f762020",
  7571 => x"00000000",
  7572 => x"63683020",
  7573 => x"73756d20",
  7574 => x"6f762020",
  7575 => x"00000000",
  7576 => x"73756d20",
  7577 => x"73636c20",
  7578 => x"6f762020",
  7579 => x"00000000",
  7580 => x"73756d20",
  7581 => x"63757420",
  7582 => x"20000000",
  7583 => x"63683320",
  7584 => x"64697620",
  7585 => x"63757420",
  7586 => x"20000000",
  7587 => x"63683320",
  7588 => x"6e736520",
  7589 => x"636d7020",
  7590 => x"20000000",
  7591 => x"63683320",
  7592 => x"6e736520",
  7593 => x"63757420",
  7594 => x"20000000",
  7595 => x"63683220",
  7596 => x"64697620",
  7597 => x"63757420",
  7598 => x"20000000",
  7599 => x"63683220",
  7600 => x"6e736520",
  7601 => x"636d7020",
  7602 => x"20000000",
  7603 => x"63683220",
  7604 => x"6e736520",
  7605 => x"63757420",
  7606 => x"20000000",
  7607 => x"63683120",
  7608 => x"64697620",
  7609 => x"63757420",
  7610 => x"20000000",
  7611 => x"63683120",
  7612 => x"6e736520",
  7613 => x"636d7020",
  7614 => x"20000000",
  7615 => x"63683120",
  7616 => x"6e736520",
  7617 => x"63757420",
  7618 => x"20000000",
  7619 => x"63683020",
  7620 => x"64697620",
  7621 => x"63757420",
  7622 => x"20000000",
  7623 => x"63683020",
  7624 => x"6e736520",
  7625 => x"636d7020",
  7626 => x"20000000",
  7627 => x"63683020",
  7628 => x"6e736520",
  7629 => x"63757420",
  7630 => x"20000000",
  7631 => x"736f6674",
  7632 => x"20657272",
  7633 => x"20200000",
  7634 => x"0000350d",
  7635 => x"00003503",
  7636 => x"000034f9",
  7637 => x"000034ef",
  7638 => x"000034e5",
  7639 => x"000034dc",
  7640 => x"000034d3",
  7641 => x"00003676",
  7642 => x"000039d3",
  7643 => x"000039c9",
  7644 => x"000039bf",
  7645 => x"000039b5",
  7646 => x"000039ab",
  7647 => x"000039a1",
  7648 => x"0a202044",
  7649 => x"434d2061",
  7650 => x"63746976",
  7651 => x"65000000",
  7652 => x"0a202044",
  7653 => x"434d204e",
  7654 => x"4f542061",
  7655 => x"63746976",
  7656 => x"65000000",
  7657 => x"0a202075",
  7658 => x"70706572",
  7659 => x"20626f75",
  7660 => x"6e64206f",
  7661 => x"76657266",
  7662 => x"6c6f7700",
  7663 => x"0a20206c",
  7664 => x"6f776572",
  7665 => x"20626f75",
  7666 => x"6e642075",
  7667 => x"6e646572",
  7668 => x"666c6f77",
  7669 => x"00000000",
  7670 => x"0a202063",
  7671 => x"6f6e6e65",
  7672 => x"6374696f",
  7673 => x"6e206c6f",
  7674 => x"73740000",
  7675 => x"0a202074",
  7676 => x"696d656f",
  7677 => x"75740000",
  7678 => x"0a646174",
  7679 => x"6120696e",
  7680 => x"20202020",
  7681 => x"203a2000",
  7682 => x"0a73756d",
  7683 => x"20696e20",
  7684 => x"20202020",
  7685 => x"203a2000",
  7686 => x"0a617665",
  7687 => x"72616765",
  7688 => x"20202020",
  7689 => x"203a2000",
  7690 => x"0a6c6f77",
  7691 => x"65722062",
  7692 => x"6f756e64",
  7693 => x"203a2000",
  7694 => x"0a757070",
  7695 => x"65722062",
  7696 => x"6f756e64",
  7697 => x"203a2000",
  7698 => x"0a737461",
  7699 => x"74652020",
  7700 => x"20202020",
  7701 => x"203a2030",
  7702 => x"78000000",
  7703 => x"0a307800",
  7704 => x"786d6f64",
  7705 => x"656d2074",
  7706 => x"72616e73",
  7707 => x"6d69742e",
  7708 => x"2e2e0a00",
  7709 => x"20627974",
  7710 => x"65732074",
  7711 => x"72616e73",
  7712 => x"6d697474",
  7713 => x"65640a00",
  7714 => x"63616e63",
  7715 => x"656c0a00",
  7716 => x"72657472",
  7717 => x"79206f75",
  7718 => x"740a0000",
  7719 => x"786d6f64",
  7720 => x"656d2072",
  7721 => x"65636569",
  7722 => x"76652e2e",
  7723 => x"2e0a0000",
  7724 => x"20627974",
  7725 => x"65732072",
  7726 => x"65636569",
  7727 => x"7665640a",
  7728 => x"00000000",
  7729 => x"72782062",
  7730 => x"75666665",
  7731 => x"72206675",
  7732 => x"6c6c0a00",
  7733 => x"74696d65",
  7734 => x"206f7574",
  7735 => x"0a000000",
  7736 => x"64656275",
  7737 => x"67207265",
  7738 => x"67697374",
  7739 => x"65727300",
  7740 => x"0a6d6f64",
  7741 => x"65202020",
  7742 => x"20202020",
  7743 => x"203a2000",
  7744 => x"0a616464",
  7745 => x"72657373",
  7746 => x"20302020",
  7747 => x"203a2030",
  7748 => x"78000000",
  7749 => x"0a616464",
  7750 => x"72657373",
  7751 => x"20312020",
  7752 => x"203a2030",
  7753 => x"78000000",
  7754 => x"0a627566",
  7755 => x"66657220",
  7756 => x"73697a65",
  7757 => x"203a2000",
  7758 => x"0a646562",
  7759 => x"75672074",
  7760 => x"72616365",
  7761 => x"206d656d",
  7762 => x"6f727900",
  7763 => x"0a74696d",
  7764 => x"65207374",
  7765 => x"616d7020",
  7766 => x"20202073",
  7767 => x"74617465",
  7768 => x"00000000",
  7769 => x"20203078",
  7770 => x"00000000",
  7771 => x"6d61783a",
  7772 => x"20000000",
  7773 => x"6d696e3a",
  7774 => x"20000000",
  7775 => x"63683a20",
  7776 => x"00000000",
  7777 => x"73706c3a",
  7778 => x"20000000",
  7779 => x"30622020",
  7780 => x"20202020",
  7781 => x"20202020",
  7782 => x"20202020",
  7783 => x"20202020",
  7784 => x"20202020",
  7785 => x"20202020",
  7786 => x"20202020",
  7787 => x"20200000",
  7788 => x"20202020",
  7789 => x"20202020",
  7790 => x"00000000",
  7791 => x"00202020",
  7792 => x"20202020",
  7793 => x"20202828",
  7794 => x"28282820",
  7795 => x"20202020",
  7796 => x"20202020",
  7797 => x"20202020",
  7798 => x"20202020",
  7799 => x"20881010",
  7800 => x"10101010",
  7801 => x"10101010",
  7802 => x"10101010",
  7803 => x"10040404",
  7804 => x"04040404",
  7805 => x"04040410",
  7806 => x"10101010",
  7807 => x"10104141",
  7808 => x"41414141",
  7809 => x"01010101",
  7810 => x"01010101",
  7811 => x"01010101",
  7812 => x"01010101",
  7813 => x"01010101",
  7814 => x"10101010",
  7815 => x"10104242",
  7816 => x"42424242",
  7817 => x"02020202",
  7818 => x"02020202",
  7819 => x"02020202",
  7820 => x"02020202",
  7821 => x"02020202",
  7822 => x"10101010",
  7823 => x"20000000",
  7824 => x"00000000",
  7825 => x"00000000",
  7826 => x"00000000",
  7827 => x"00000000",
  7828 => x"00000000",
  7829 => x"00000000",
  7830 => x"00000000",
  7831 => x"00000000",
  7832 => x"00000000",
  7833 => x"00000000",
  7834 => x"00000000",
  7835 => x"00000000",
  7836 => x"00000000",
  7837 => x"00000000",
  7838 => x"00000000",
  7839 => x"00000000",
  7840 => x"00000000",
  7841 => x"00000000",
  7842 => x"00000000",
  7843 => x"00000000",
  7844 => x"00000000",
  7845 => x"00000000",
  7846 => x"00000000",
  7847 => x"00000000",
  7848 => x"00000000",
  7849 => x"00000000",
  7850 => x"00000000",
  7851 => x"00000000",
  7852 => x"00000000",
  7853 => x"00000000",
  7854 => x"00000000",
  7855 => x"00000000",
  7856 => x"80000c00",
  7857 => x"00000000",
  7858 => x"80000900",
  7859 => x"80000800",
  7860 => x"00000000",
  7861 => x"00000000",
  7862 => x"ff000000",
  7863 => x"00000000",
  7864 => x"80000b00",
  7865 => x"00ffffff",
  7866 => x"ff00ffff",
  7867 => x"ffff00ff",
  7868 => x"ffffff00",
  7869 => x"00000000",
  7870 => x"00000000",
  7871 => x"80000f00",
  7872 => x"80000a00",
  7873 => x"80000700",
  7874 => x"80000600",
  7875 => x"80000400",
  7876 => x"80000200",
  7877 => x"80000100",
  7878 => x"80000004",
  7879 => x"80000000",
  7880 => x"00007b24",
  7881 => x"00000000",
  7882 => x"00007d8c",
  7883 => x"00007de8",
  7884 => x"00007e44",
  7885 => x"00000000",
  7886 => x"00000000",
  7887 => x"00000000",
  7888 => x"00000000",
  7889 => x"00000000",
  7890 => x"00000000",
  7891 => x"00000000",
  7892 => x"00000000",
  7893 => x"00000000",
  7894 => x"00006838",
  7895 => x"00000000",
  7896 => x"00000000",
  7897 => x"00000000",
  7898 => x"00000000",
  7899 => x"00000000",
  7900 => x"00000000",
  7901 => x"00000000",
  7902 => x"00000000",
  7903 => x"00000000",
  7904 => x"00000000",
  7905 => x"00000000",
  7906 => x"00000000",
  7907 => x"00000000",
  7908 => x"00000000",
  7909 => x"00000000",
  7910 => x"00000000",
  7911 => x"00000000",
  7912 => x"00000000",
  7913 => x"00000000",
  7914 => x"00000000",
  7915 => x"00000000",
  7916 => x"00000000",
  7917 => x"00000000",
  7918 => x"00000000",
  7919 => x"00000000",
  7920 => x"00000000",
  7921 => x"00000000",
  7922 => x"00000000",
  7923 => x"00000001",
  7924 => x"330eabcd",
  7925 => x"1234e66d",
  7926 => x"deec0005",
  7927 => x"000b0000",
  7928 => x"00000000",
  7929 => x"00000000",
  7930 => x"00000000",
  7931 => x"00000000",
  7932 => x"00000000",
  7933 => x"00000000",
  7934 => x"00000000",
  7935 => x"00000000",
  7936 => x"00000000",
  7937 => x"00000000",
  7938 => x"00000000",
  7939 => x"00000000",
  7940 => x"00000000",
  7941 => x"00000000",
  7942 => x"00000000",
  7943 => x"00000000",
  7944 => x"00000000",
  7945 => x"00000000",
  7946 => x"00000000",
  7947 => x"00000000",
  7948 => x"00000000",
  7949 => x"00000000",
  7950 => x"00000000",
  7951 => x"00000000",
  7952 => x"00000000",
  7953 => x"00000000",
  7954 => x"00000000",
  7955 => x"00000000",
  7956 => x"00000000",
  7957 => x"00000000",
  7958 => x"00000000",
  7959 => x"00000000",
  7960 => x"00000000",
  7961 => x"00000000",
  7962 => x"00000000",
  7963 => x"00000000",
  7964 => x"00000000",
  7965 => x"00000000",
  7966 => x"00000000",
  7967 => x"00000000",
  7968 => x"00000000",
  7969 => x"00000000",
  7970 => x"00000000",
  7971 => x"00000000",
  7972 => x"00000000",
  7973 => x"00000000",
  7974 => x"00000000",
  7975 => x"00000000",
  7976 => x"00000000",
  7977 => x"00000000",
  7978 => x"00000000",
  7979 => x"00000000",
  7980 => x"00000000",
  7981 => x"00000000",
  7982 => x"00000000",
  7983 => x"00000000",
  7984 => x"00000000",
  7985 => x"00000000",
  7986 => x"00000000",
  7987 => x"00000000",
  7988 => x"00000000",
  7989 => x"00000000",
  7990 => x"00000000",
  7991 => x"00000000",
  7992 => x"00000000",
  7993 => x"00000000",
  7994 => x"00000000",
  7995 => x"00000000",
  7996 => x"00000000",
  7997 => x"00000000",
  7998 => x"00000000",
  7999 => x"00000000",
  8000 => x"00000000",
  8001 => x"00000000",
  8002 => x"00000000",
  8003 => x"00000000",
  8004 => x"00000000",
  8005 => x"00000000",
  8006 => x"00000000",
  8007 => x"00000000",
  8008 => x"00000000",
  8009 => x"00000000",
  8010 => x"00000000",
  8011 => x"00000000",
  8012 => x"00000000",
  8013 => x"00000000",
  8014 => x"00000000",
  8015 => x"00000000",
  8016 => x"00000000",
  8017 => x"00000000",
  8018 => x"00000000",
  8019 => x"00000000",
  8020 => x"00000000",
  8021 => x"00000000",
  8022 => x"00000000",
  8023 => x"00000000",
  8024 => x"00000000",
  8025 => x"00000000",
  8026 => x"00000000",
  8027 => x"00000000",
  8028 => x"00000000",
  8029 => x"00000000",
  8030 => x"00000000",
  8031 => x"00000000",
  8032 => x"00000000",
  8033 => x"00000000",
  8034 => x"00000000",
  8035 => x"00000000",
  8036 => x"00000000",
  8037 => x"00000000",
  8038 => x"00000000",
  8039 => x"00000000",
  8040 => x"00000000",
  8041 => x"00000000",
  8042 => x"00000000",
  8043 => x"00000000",
  8044 => x"00000000",
  8045 => x"00000000",
  8046 => x"00000000",
  8047 => x"00000000",
  8048 => x"00000000",
  8049 => x"00000000",
  8050 => x"00000000",
  8051 => x"00000000",
  8052 => x"00000000",
  8053 => x"00000000",
  8054 => x"00000000",
  8055 => x"00000000",
  8056 => x"00000000",
  8057 => x"00000000",
  8058 => x"00000000",
  8059 => x"00000000",
  8060 => x"00000000",
  8061 => x"00000000",
  8062 => x"00000000",
  8063 => x"00000000",
  8064 => x"00000000",
  8065 => x"00000000",
  8066 => x"00000000",
  8067 => x"00000000",
  8068 => x"00000000",
  8069 => x"00000000",
  8070 => x"00000000",
  8071 => x"00000000",
  8072 => x"00000000",
  8073 => x"00000000",
  8074 => x"00000000",
  8075 => x"00000000",
  8076 => x"00000000",
  8077 => x"00000000",
  8078 => x"00000000",
  8079 => x"00000000",
  8080 => x"00000000",
  8081 => x"00000000",
  8082 => x"00000000",
  8083 => x"00000000",
  8084 => x"00000000",
  8085 => x"00000000",
  8086 => x"00000000",
  8087 => x"00000000",
  8088 => x"00000000",
  8089 => x"00000000",
  8090 => x"00000000",
  8091 => x"00000000",
  8092 => x"00000000",
  8093 => x"00000000",
  8094 => x"00000000",
  8095 => x"00000000",
  8096 => x"00000000",
  8097 => x"00000000",
  8098 => x"00000000",
  8099 => x"00000000",
  8100 => x"00000000",
  8101 => x"00000000",
  8102 => x"00000000",
  8103 => x"00000000",
  8104 => x"00000000",
  8105 => x"00000000",
  8106 => x"00000000",
  8107 => x"00000000",
  8108 => x"00000000",
  8109 => x"00000000",
  8110 => x"00000000",
  8111 => x"00000000",
  8112 => x"00000000",
  8113 => x"00000000",
  8114 => x"00000000",
  8115 => x"00000000",
  8116 => x"ffffffff",
  8117 => x"00000000",
  8118 => x"00020000",
  8119 => x"00000000",
  8120 => x"00000000",
  8121 => x"00007edc",
  8122 => x"00007edc",
  8123 => x"00007ee4",
  8124 => x"00007ee4",
  8125 => x"00007eec",
  8126 => x"00007eec",
  8127 => x"00007ef4",
  8128 => x"00007ef4",
  8129 => x"00007efc",
  8130 => x"00007efc",
  8131 => x"00007f04",
  8132 => x"00007f04",
  8133 => x"00007f0c",
  8134 => x"00007f0c",
  8135 => x"00007f14",
  8136 => x"00007f14",
  8137 => x"00007f1c",
  8138 => x"00007f1c",
  8139 => x"00007f24",
  8140 => x"00007f24",
  8141 => x"00007f2c",
  8142 => x"00007f2c",
  8143 => x"00007f34",
  8144 => x"00007f34",
  8145 => x"00007f3c",
  8146 => x"00007f3c",
  8147 => x"00007f44",
  8148 => x"00007f44",
  8149 => x"00007f4c",
  8150 => x"00007f4c",
  8151 => x"00007f54",
  8152 => x"00007f54",
  8153 => x"00007f5c",
  8154 => x"00007f5c",
  8155 => x"00007f64",
  8156 => x"00007f64",
  8157 => x"00007f6c",
  8158 => x"00007f6c",
  8159 => x"00007f74",
  8160 => x"00007f74",
  8161 => x"00007f7c",
  8162 => x"00007f7c",
  8163 => x"00007f84",
  8164 => x"00007f84",
  8165 => x"00007f8c",
  8166 => x"00007f8c",
  8167 => x"00007f94",
  8168 => x"00007f94",
  8169 => x"00007f9c",
  8170 => x"00007f9c",
  8171 => x"00007fa4",
  8172 => x"00007fa4",
  8173 => x"00007fac",
  8174 => x"00007fac",
  8175 => x"00007fb4",
  8176 => x"00007fb4",
  8177 => x"00007fbc",
  8178 => x"00007fbc",
  8179 => x"00007fc4",
  8180 => x"00007fc4",
  8181 => x"00007fcc",
  8182 => x"00007fcc",
  8183 => x"00007fd4",
  8184 => x"00007fd4",
  8185 => x"00007fdc",
  8186 => x"00007fdc",
  8187 => x"00007fe4",
  8188 => x"00007fe4",
  8189 => x"00007fec",
  8190 => x"00007fec",
  8191 => x"00007ff4",
  8192 => x"00007ff4",
  8193 => x"00007ffc",
  8194 => x"00007ffc",
  8195 => x"00008004",
  8196 => x"00008004",
  8197 => x"0000800c",
  8198 => x"0000800c",
  8199 => x"00008014",
  8200 => x"00008014",
  8201 => x"0000801c",
  8202 => x"0000801c",
  8203 => x"00008024",
  8204 => x"00008024",
  8205 => x"0000802c",
  8206 => x"0000802c",
  8207 => x"00008034",
  8208 => x"00008034",
  8209 => x"0000803c",
  8210 => x"0000803c",
  8211 => x"00008044",
  8212 => x"00008044",
  8213 => x"0000804c",
  8214 => x"0000804c",
  8215 => x"00008054",
  8216 => x"00008054",
  8217 => x"0000805c",
  8218 => x"0000805c",
  8219 => x"00008064",
  8220 => x"00008064",
  8221 => x"0000806c",
  8222 => x"0000806c",
  8223 => x"00008074",
  8224 => x"00008074",
  8225 => x"0000807c",
  8226 => x"0000807c",
  8227 => x"00008084",
  8228 => x"00008084",
  8229 => x"0000808c",
  8230 => x"0000808c",
  8231 => x"00008094",
  8232 => x"00008094",
  8233 => x"0000809c",
  8234 => x"0000809c",
  8235 => x"000080a4",
  8236 => x"000080a4",
  8237 => x"000080ac",
  8238 => x"000080ac",
  8239 => x"000080b4",
  8240 => x"000080b4",
  8241 => x"000080bc",
  8242 => x"000080bc",
  8243 => x"000080c4",
  8244 => x"000080c4",
  8245 => x"000080cc",
  8246 => x"000080cc",
  8247 => x"000080d4",
  8248 => x"000080d4",
  8249 => x"000080dc",
  8250 => x"000080dc",
  8251 => x"000080e4",
  8252 => x"000080e4",
  8253 => x"000080ec",
  8254 => x"000080ec",
  8255 => x"000080f4",
  8256 => x"000080f4",
  8257 => x"000080fc",
  8258 => x"000080fc",
  8259 => x"00008104",
  8260 => x"00008104",
  8261 => x"0000810c",
  8262 => x"0000810c",
  8263 => x"00008114",
  8264 => x"00008114",
  8265 => x"0000811c",
  8266 => x"0000811c",
  8267 => x"00008124",
  8268 => x"00008124",
  8269 => x"0000812c",
  8270 => x"0000812c",
  8271 => x"00008134",
  8272 => x"00008134",
  8273 => x"0000813c",
  8274 => x"0000813c",
  8275 => x"00008144",
  8276 => x"00008144",
  8277 => x"0000814c",
  8278 => x"0000814c",
  8279 => x"00008154",
  8280 => x"00008154",
  8281 => x"0000815c",
  8282 => x"0000815c",
  8283 => x"00008164",
  8284 => x"00008164",
  8285 => x"0000816c",
  8286 => x"0000816c",
  8287 => x"00008174",
  8288 => x"00008174",
  8289 => x"0000817c",
  8290 => x"0000817c",
  8291 => x"00008184",
  8292 => x"00008184",
  8293 => x"0000818c",
  8294 => x"0000818c",
  8295 => x"00008194",
  8296 => x"00008194",
  8297 => x"0000819c",
  8298 => x"0000819c",
  8299 => x"000081a4",
  8300 => x"000081a4",
  8301 => x"000081ac",
  8302 => x"000081ac",
  8303 => x"000081b4",
  8304 => x"000081b4",
  8305 => x"000081bc",
  8306 => x"000081bc",
  8307 => x"000081c4",
  8308 => x"000081c4",
  8309 => x"000081cc",
  8310 => x"000081cc",
  8311 => x"000081d4",
  8312 => x"000081d4",
  8313 => x"000081dc",
  8314 => x"000081dc",
  8315 => x"000081e4",
  8316 => x"000081e4",
  8317 => x"000081ec",
  8318 => x"000081ec",
  8319 => x"000081f4",
  8320 => x"000081f4",
  8321 => x"000081fc",
  8322 => x"000081fc",
  8323 => x"00008204",
  8324 => x"00008204",
  8325 => x"0000820c",
  8326 => x"0000820c",
  8327 => x"00008214",
  8328 => x"00008214",
  8329 => x"0000821c",
  8330 => x"0000821c",
  8331 => x"00008224",
  8332 => x"00008224",
  8333 => x"0000822c",
  8334 => x"0000822c",
  8335 => x"00008234",
  8336 => x"00008234",
  8337 => x"0000823c",
  8338 => x"0000823c",
  8339 => x"00008244",
  8340 => x"00008244",
  8341 => x"0000824c",
  8342 => x"0000824c",
  8343 => x"00008254",
  8344 => x"00008254",
  8345 => x"0000825c",
  8346 => x"0000825c",
  8347 => x"00008264",
  8348 => x"00008264",
  8349 => x"0000826c",
  8350 => x"0000826c",
  8351 => x"00008274",
  8352 => x"00008274",
  8353 => x"0000827c",
  8354 => x"0000827c",
  8355 => x"00008284",
  8356 => x"00008284",
  8357 => x"0000828c",
  8358 => x"0000828c",
  8359 => x"00008294",
  8360 => x"00008294",
  8361 => x"0000829c",
  8362 => x"0000829c",
  8363 => x"000082a4",
  8364 => x"000082a4",
  8365 => x"000082ac",
  8366 => x"000082ac",
  8367 => x"000082b4",
  8368 => x"000082b4",
  8369 => x"000082bc",
  8370 => x"000082bc",
  8371 => x"000082c4",
  8372 => x"000082c4",
  8373 => x"000082cc",
  8374 => x"000082cc",
  8375 => x"000082d4",
  8376 => x"000082d4",
	others => x"00dead00" -- mask for mem check
	--others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
