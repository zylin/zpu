-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80e3880c",
     3 => x"3a0b0b80",
     4 => x"d2c20400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80d38b2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80e2",
   162 => x"f4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80cd",
   171 => x"ad2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80ce",
   179 => x"df2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80e3840c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"ccac3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80e38408",
   281 => x"802ea438",
   282 => x"80e38808",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80ea",
   286 => x"c40c82a0",
   287 => x"800b80ea",
   288 => x"c80c8290",
   289 => x"800b80ea",
   290 => x"cc0c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"eac40cf8",
   294 => x"80808280",
   295 => x"0b80eac8",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"eacc0c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80eac40c",
   302 => x"80c0a880",
   303 => x"940b80ea",
   304 => x"c80c0b0b",
   305 => x"80d4e00b",
   306 => x"80eacc0c",
   307 => x"04ff3d0d",
   308 => x"80ead033",
   309 => x"5170a738",
   310 => x"80e39008",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"e3900c70",
   315 => x"2d80e390",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80ea",
   319 => x"d034833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80eac008",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"eac0510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404fb3d",
   333 => x"0d775680",
   334 => x"55747627",
   335 => x"81993880",
   336 => x"e3a40854",
   337 => x"bfa9bc0b",
   338 => x"94150c85",
   339 => x"0b98150c",
   340 => x"98140870",
   341 => x"81065153",
   342 => x"72f638bf",
   343 => x"a9bc0b94",
   344 => x"150c850b",
   345 => x"98150c98",
   346 => x"14087081",
   347 => x"06515372",
   348 => x"f638bfa9",
   349 => x"bc0b9415",
   350 => x"0c850b98",
   351 => x"150c9814",
   352 => x"08708106",
   353 => x"515372f6",
   354 => x"38bfa9bc",
   355 => x"0b94150c",
   356 => x"850b9815",
   357 => x"0c981408",
   358 => x"70810651",
   359 => x"5372f638",
   360 => x"bfa9bc0b",
   361 => x"94150c85",
   362 => x"0b98150c",
   363 => x"98140870",
   364 => x"81065153",
   365 => x"72f638bf",
   366 => x"a9bc0b94",
   367 => x"150c850b",
   368 => x"98150c98",
   369 => x"14087081",
   370 => x"06515372",
   371 => x"f6388115",
   372 => x"55757526",
   373 => x"feee3887",
   374 => x"3d0d0480",
   375 => x"3d0d80e3",
   376 => x"a4085187",
   377 => x"0b84120c",
   378 => x"823d0d04",
   379 => x"f83d0d7a",
   380 => x"7c595380",
   381 => x"73565776",
   382 => x"732480de",
   383 => x"38771754",
   384 => x"8a527451",
   385 => x"80c1813f",
   386 => x"8008b005",
   387 => x"53727434",
   388 => x"8117578a",
   389 => x"52745180",
   390 => x"c0c93f80",
   391 => x"08558008",
   392 => x"dc388008",
   393 => x"779f2a18",
   394 => x"70812c5b",
   395 => x"56568079",
   396 => x"259e3877",
   397 => x"17ff0555",
   398 => x"75187033",
   399 => x"55537433",
   400 => x"73347375",
   401 => x"348116ff",
   402 => x"16565678",
   403 => x"7624e938",
   404 => x"76185680",
   405 => x"76348a3d",
   406 => x"0d04ad78",
   407 => x"7081055a",
   408 => x"34723078",
   409 => x"1855558a",
   410 => x"52745180",
   411 => x"c09a3f80",
   412 => x"08b00553",
   413 => x"72743481",
   414 => x"17578a52",
   415 => x"7451bfe3",
   416 => x"3f800855",
   417 => x"8008fef5",
   418 => x"38ff9739",
   419 => x"f93d0d79",
   420 => x"70713370",
   421 => x"81ff0654",
   422 => x"55555570",
   423 => x"802eb138",
   424 => x"80e3a808",
   425 => x"527281ff",
   426 => x"06811555",
   427 => x"53728a2e",
   428 => x"80f53884",
   429 => x"12087082",
   430 => x"2a810652",
   431 => x"5770802e",
   432 => x"f2387272",
   433 => x"0c733370",
   434 => x"81ff0659",
   435 => x"5377d638",
   436 => x"74753352",
   437 => x"5670802e",
   438 => x"80c93870",
   439 => x"80e3a008",
   440 => x"59538116",
   441 => x"80ead833",
   442 => x"7081ff06",
   443 => x"70101011",
   444 => x"80eadc33",
   445 => x"7081ff06",
   446 => x"72902911",
   447 => x"70882b7a",
   448 => x"077f0c53",
   449 => x"59595454",
   450 => x"5856728a",
   451 => x"2ebe3873",
   452 => x"80cf2eb8",
   453 => x"38811553",
   454 => x"7280eadc",
   455 => x"34753353",
   456 => x"72c03889",
   457 => x"3d0d0484",
   458 => x"12087082",
   459 => x"2a810657",
   460 => x"5875802e",
   461 => x"f2388d72",
   462 => x"0c841208",
   463 => x"70822a81",
   464 => x"06525770",
   465 => x"802efeeb",
   466 => x"38fef739",
   467 => x"71a32699",
   468 => x"38811752",
   469 => x"7180ead8",
   470 => x"34800b80",
   471 => x"eadc3475",
   472 => x"335372fe",
   473 => x"fd38ffbb",
   474 => x"39800b80",
   475 => x"ead83480",
   476 => x"0b80eadc",
   477 => x"34e939fd",
   478 => x"3d0d80e3",
   479 => x"9c085480",
   480 => x"d50b8415",
   481 => x"0c80e3a8",
   482 => x"08528412",
   483 => x"08810651",
   484 => x"70802ef6",
   485 => x"38710870",
   486 => x"81ff06f6",
   487 => x"11525451",
   488 => x"70ae268c",
   489 => x"38701010",
   490 => x"80e0f405",
   491 => x"51700804",
   492 => x"84120870",
   493 => x"822a7081",
   494 => x"06515151",
   495 => x"70802ef0",
   496 => x"38ab720c",
   497 => x"728a2eaa",
   498 => x"38841208",
   499 => x"70822a70",
   500 => x"81065151",
   501 => x"5170802e",
   502 => x"f0387272",
   503 => x"0c841208",
   504 => x"70822a81",
   505 => x"06515372",
   506 => x"802ef238",
   507 => x"ad720cff",
   508 => x"99398412",
   509 => x"0870822a",
   510 => x"70810651",
   511 => x"51517080",
   512 => x"2ef0388d",
   513 => x"720c8412",
   514 => x"0870822a",
   515 => x"70810651",
   516 => x"51517080",
   517 => x"2effb238",
   518 => x"c13981ff",
   519 => x"0b84150c",
   520 => x"fee83980",
   521 => x"ff0b8415",
   522 => x"0cfedf39",
   523 => x"bf0b8415",
   524 => x"0cfed739",
   525 => x"9f0b8415",
   526 => x"0cfecf39",
   527 => x"8f0b8415",
   528 => x"0cfec739",
   529 => x"870b8415",
   530 => x"0cfebf39",
   531 => x"830b8415",
   532 => x"0cfeb739",
   533 => x"810b8415",
   534 => x"0cfeaf39",
   535 => x"800b8415",
   536 => x"0cfea739",
   537 => x"d73d0d80",
   538 => x"e3a00855",
   539 => x"800b8416",
   540 => x"0cfe800a",
   541 => x"0b88160c",
   542 => x"800b80ea",
   543 => x"d834800b",
   544 => x"80eadc34",
   545 => x"a63d7053",
   546 => x"80e39808",
   547 => x"8c110853",
   548 => x"555bfad8",
   549 => x"3f80d88c",
   550 => x"0b80d88c",
   551 => x"33555a73",
   552 => x"802e80cc",
   553 => x"3880e3a0",
   554 => x"0874575c",
   555 => x"811a80ea",
   556 => x"d8337081",
   557 => x"ff067010",
   558 => x"101180ea",
   559 => x"dc337081",
   560 => x"ff067290",
   561 => x"29117088",
   562 => x"2b7d0763",
   563 => x"0c445c5c",
   564 => x"42575a5a",
   565 => x"758a2e87",
   566 => x"bc387680",
   567 => x"cf2e87b5",
   568 => x"38811857",
   569 => x"7680eadc",
   570 => x"34793356",
   571 => x"75ffbd38",
   572 => x"7a7b3355",
   573 => x"5a73802e",
   574 => x"80cc3880",
   575 => x"e3a00874",
   576 => x"575b811a",
   577 => x"80ead833",
   578 => x"7081ff06",
   579 => x"70101011",
   580 => x"80eadc33",
   581 => x"7081ff06",
   582 => x"72902911",
   583 => x"70882b7d",
   584 => x"07620c46",
   585 => x"5c5c4457",
   586 => x"5a5a758a",
   587 => x"2e878438",
   588 => x"7680cf2e",
   589 => x"86fd3881",
   590 => x"18597880",
   591 => x"eadc3479",
   592 => x"335675ff",
   593 => x"bd3880d8",
   594 => x"a40b80d8",
   595 => x"a433555a",
   596 => x"73802e80",
   597 => x"cc3880e3",
   598 => x"a0087457",
   599 => x"5b811a80",
   600 => x"ead83370",
   601 => x"81ff0670",
   602 => x"10101180",
   603 => x"eadc3370",
   604 => x"81ff0672",
   605 => x"90291170",
   606 => x"882b7d07",
   607 => x"620c495c",
   608 => x"5c57575a",
   609 => x"5a758a2e",
   610 => x"85ed3876",
   611 => x"80cf2e85",
   612 => x"e6388118",
   613 => x"5d7c80ea",
   614 => x"dc347933",
   615 => x"5675ffbd",
   616 => x"3880e398",
   617 => x"087008a5",
   618 => x"3d5b575a",
   619 => x"8b5380d4",
   620 => x"e4527851",
   621 => x"bdf33f82",
   622 => x"02840581",
   623 => x"89055957",
   624 => x"758f0654",
   625 => x"73892685",
   626 => x"92387618",
   627 => x"b0155555",
   628 => x"73753475",
   629 => x"842aff18",
   630 => x"7081ff06",
   631 => x"595c5676",
   632 => x"df387879",
   633 => x"33555a73",
   634 => x"802e80cc",
   635 => x"3880e3a0",
   636 => x"0874575b",
   637 => x"811a80ea",
   638 => x"d8337081",
   639 => x"ff067010",
   640 => x"101180ea",
   641 => x"dc337081",
   642 => x"ff067290",
   643 => x"29117088",
   644 => x"2b7d0762",
   645 => x"0c455c5c",
   646 => x"5f575a5a",
   647 => x"758a2e87",
   648 => x"f3387680",
   649 => x"cf2e87ec",
   650 => x"38811857",
   651 => x"7680eadc",
   652 => x"34793356",
   653 => x"75ffbd38",
   654 => x"80d8b00b",
   655 => x"80d8b033",
   656 => x"555a7380",
   657 => x"2e80cc38",
   658 => x"80e3a008",
   659 => x"74575b81",
   660 => x"1a80ead8",
   661 => x"337081ff",
   662 => x"06701010",
   663 => x"1180eadc",
   664 => x"337081ff",
   665 => x"06729029",
   666 => x"1170882b",
   667 => x"7d07620c",
   668 => x"475c5c45",
   669 => x"575a5a75",
   670 => x"8a2e87b6",
   671 => x"387680cf",
   672 => x"2e87af38",
   673 => x"81185978",
   674 => x"80eadc34",
   675 => x"79335675",
   676 => x"ffbd3880",
   677 => x"5f890a5c",
   678 => x"ac3d087f",
   679 => x"2e098106",
   680 => x"87ca387e",
   681 => x"a13d0288",
   682 => x"0580fd05",
   683 => x"40415d7c",
   684 => x"bf064362",
   685 => x"85d43880",
   686 => x"d8840b80",
   687 => x"d8843355",
   688 => x"5a73802e",
   689 => x"80cc3880",
   690 => x"e3a00874",
   691 => x"575b811a",
   692 => x"80ead833",
   693 => x"7081ff06",
   694 => x"70101011",
   695 => x"80eadc33",
   696 => x"7081ff06",
   697 => x"72902911",
   698 => x"70882b7d",
   699 => x"07620c47",
   700 => x"5c5c4557",
   701 => x"5a5a758a",
   702 => x"2e848a38",
   703 => x"7680cf2e",
   704 => x"84833881",
   705 => x"18567580",
   706 => x"eadc3479",
   707 => x"335675ff",
   708 => x"bd387b56",
   709 => x"8b5380d4",
   710 => x"e4527f51",
   711 => x"bb8b3f88",
   712 => x"57758f06",
   713 => x"54738926",
   714 => x"83d23876",
   715 => x"1eb01555",
   716 => x"55737534",
   717 => x"75842aff",
   718 => x"187081ff",
   719 => x"06595b56",
   720 => x"76df387f",
   721 => x"6033555a",
   722 => x"73802e85",
   723 => x"bf3880e3",
   724 => x"a0087457",
   725 => x"5b811a80",
   726 => x"ead83370",
   727 => x"81ff0670",
   728 => x"10101180",
   729 => x"eadc3370",
   730 => x"81ff0672",
   731 => x"90291170",
   732 => x"882b7d07",
   733 => x"620c5a5c",
   734 => x"5c44575a",
   735 => x"5a758a2e",
   736 => x"83bf3876",
   737 => x"80cf2e83",
   738 => x"b8388118",
   739 => x"597880ea",
   740 => x"dc347933",
   741 => x"5675ffbd",
   742 => x"3880d8b4",
   743 => x"0b80d8b4",
   744 => x"33555a73",
   745 => x"802e80c7",
   746 => x"38735681",
   747 => x"1a80ead8",
   748 => x"337081ff",
   749 => x"06701010",
   750 => x"1180eadc",
   751 => x"337081ff",
   752 => x"06729029",
   753 => x"1170882b",
   754 => x"7d07620c",
   755 => x"495c5c57",
   756 => x"575a5a75",
   757 => x"8a2e82cb",
   758 => x"387680cf",
   759 => x"2e82c438",
   760 => x"81185574",
   761 => x"80eadc34",
   762 => x"79335675",
   763 => x"ffbd387b",
   764 => x"087c3270",
   765 => x"30710770",
   766 => x"9f2a7081",
   767 => x"ff06b011",
   768 => x"7081ff06",
   769 => x"80ead833",
   770 => x"7081ff06",
   771 => x"70101011",
   772 => x"80eadc33",
   773 => x"7081ff06",
   774 => x"72902911",
   775 => x"70882b77",
   776 => x"07670c4e",
   777 => x"58595c53",
   778 => x"5f465a52",
   779 => x"595b5860",
   780 => x"8a2e83a4",
   781 => x"387680cf",
   782 => x"2e839d38",
   783 => x"81184160",
   784 => x"80eadc34",
   785 => x"791f841d",
   786 => x"811f5f5d",
   787 => x"5f8fff7d",
   788 => x"27fcdc38",
   789 => x"7e800cab",
   790 => x"3d0d0476",
   791 => x"18b71555",
   792 => x"55737534",
   793 => x"75842aff",
   794 => x"187081ff",
   795 => x"06595c56",
   796 => x"76facd38",
   797 => x"faec3974",
   798 => x"a32680f1",
   799 => x"38811955",
   800 => x"7480ead8",
   801 => x"34800b80",
   802 => x"eadc3479",
   803 => x"335675f9",
   804 => x"cc38fa8d",
   805 => x"3974a326",
   806 => x"80c43881",
   807 => x"19567580",
   808 => x"ead83480",
   809 => x"0b80eadc",
   810 => x"34793356",
   811 => x"75f7fd38",
   812 => x"f8be3974",
   813 => x"a3269938",
   814 => x"81195877",
   815 => x"80ead834",
   816 => x"800b80ea",
   817 => x"dc347933",
   818 => x"5675f8b6",
   819 => x"38f8f739",
   820 => x"800b80ea",
   821 => x"d834800b",
   822 => x"80eadc34",
   823 => x"e939800b",
   824 => x"80ead834",
   825 => x"800b80ea",
   826 => x"dc34ffbd",
   827 => x"39800b80",
   828 => x"ead83480",
   829 => x"0b80eadc",
   830 => x"34ff9039",
   831 => x"761eb715",
   832 => x"5555fcad",
   833 => x"3974a326",
   834 => x"80f13881",
   835 => x"19557480",
   836 => x"ead83480",
   837 => x"0b80eadc",
   838 => x"34793356",
   839 => x"75fbaf38",
   840 => x"fbf03974",
   841 => x"a32680c4",
   842 => x"38811958",
   843 => x"7780ead8",
   844 => x"34800b80",
   845 => x"eadc3479",
   846 => x"335675fc",
   847 => x"ee38fdaf",
   848 => x"3974a326",
   849 => x"99388119",
   850 => x"577680ea",
   851 => x"d834800b",
   852 => x"80eadc34",
   853 => x"79335675",
   854 => x"fbfb38fc",
   855 => x"bc39800b",
   856 => x"80ead834",
   857 => x"800b80ea",
   858 => x"dc34e939",
   859 => x"800b80ea",
   860 => x"d834800b",
   861 => x"80eadc34",
   862 => x"ffbd3980",
   863 => x"0b80ead8",
   864 => x"34800b80",
   865 => x"eadc34ff",
   866 => x"903980e3",
   867 => x"a0087c08",
   868 => x"7d327030",
   869 => x"7107709f",
   870 => x"2a7081ff",
   871 => x"06b01170",
   872 => x"81ff0680",
   873 => x"ead83370",
   874 => x"81ff0670",
   875 => x"10101180",
   876 => x"eadc3370",
   877 => x"81ff0672",
   878 => x"90291170",
   879 => x"882b7707",
   880 => x"7d0c4f58",
   881 => x"595d5340",
   882 => x"475b525a",
   883 => x"5c595b60",
   884 => x"8a2e0981",
   885 => x"06fcde38",
   886 => x"75a326a2",
   887 => x"3881195b",
   888 => x"7a80ead8",
   889 => x"34800b80",
   890 => x"eadc3479",
   891 => x"1f841d81",
   892 => x"1f5f5d5f",
   893 => x"8fff7d27",
   894 => x"f9b538fc",
   895 => x"d739800b",
   896 => x"80ead834",
   897 => x"800b80ea",
   898 => x"dc34e039",
   899 => x"80e3a008",
   900 => x"5bfb8639",
   901 => x"74a32680",
   902 => x"c4388119",
   903 => x"567580ea",
   904 => x"d834800b",
   905 => x"80eadc34",
   906 => x"79335675",
   907 => x"f7c638f8",
   908 => x"873974a3",
   909 => x"26993881",
   910 => x"19587780",
   911 => x"ead83480",
   912 => x"0b80eadc",
   913 => x"34793356",
   914 => x"75f88438",
   915 => x"f8c53980",
   916 => x"0b80ead8",
   917 => x"34800b80",
   918 => x"eadc34e9",
   919 => x"39800b80",
   920 => x"ead83480",
   921 => x"0b80eadc",
   922 => x"34ffbd39",
   923 => x"7b7f9f3d",
   924 => x"028c0580",
   925 => x"f105983d",
   926 => x"02940580",
   927 => x"cd054542",
   928 => x"4543445d",
   929 => x"80d8840b",
   930 => x"80d88433",
   931 => x"555a7380",
   932 => x"2e80cc38",
   933 => x"80e3a008",
   934 => x"74575b81",
   935 => x"1a80ead8",
   936 => x"337081ff",
   937 => x"06701010",
   938 => x"1180eadc",
   939 => x"337081ff",
   940 => x"06729029",
   941 => x"1170882b",
   942 => x"7d07620c",
   943 => x"5a5c5c5f",
   944 => x"575a5a75",
   945 => x"8a2e8483",
   946 => x"387680cf",
   947 => x"2e83fc38",
   948 => x"81185776",
   949 => x"80eadc34",
   950 => x"79335675",
   951 => x"ffbd387c",
   952 => x"568b5380",
   953 => x"d4e45260",
   954 => x"51b3be3f",
   955 => x"8857758f",
   956 => x"06547389",
   957 => x"2683cb38",
   958 => x"6117b015",
   959 => x"55557375",
   960 => x"3475842a",
   961 => x"ff187081",
   962 => x"ff06595b",
   963 => x"5676df38",
   964 => x"60613355",
   965 => x"5a73802e",
   966 => x"84e33880",
   967 => x"e3a00874",
   968 => x"575b811a",
   969 => x"80ead833",
   970 => x"7081ff06",
   971 => x"70101011",
   972 => x"80eadc33",
   973 => x"7081ff06",
   974 => x"72902911",
   975 => x"70882b7d",
   976 => x"07620c42",
   977 => x"5c5c5757",
   978 => x"5a5a758a",
   979 => x"2e839a38",
   980 => x"7680cf2e",
   981 => x"83933881",
   982 => x"18597880",
   983 => x"eadc3479",
   984 => x"335675ff",
   985 => x"bd3880ea",
   986 => x"d8337081",
   987 => x"ff067010",
   988 => x"101180ea",
   989 => x"dc337081",
   990 => x"ff067290",
   991 => x"29117088",
   992 => x"2ba00761",
   993 => x"0c41595a",
   994 => x"56575874",
   995 => x"80cf2e84",
   996 => x"a0388117",
   997 => x"567580ea",
   998 => x"dc347c08",
   999 => x"70585ca3",
  1000 => x"5380d4f0",
  1001 => x"527d51b2",
  1002 => x"803fa056",
  1003 => x"7f1677b1",
  1004 => x"06b00756",
  1005 => x"59747934",
  1006 => x"760a100a",
  1007 => x"ff177081",
  1008 => x"ff065859",
  1009 => x"5775e538",
  1010 => x"7d7e3355",
  1011 => x"5a73802e",
  1012 => x"84883880",
  1013 => x"e3a00874",
  1014 => x"575b811a",
  1015 => x"80ead833",
  1016 => x"7081ff06",
  1017 => x"70101011",
  1018 => x"80eadc33",
  1019 => x"7081ff06",
  1020 => x"72902911",
  1021 => x"70882b7d",
  1022 => x"07620c53",
  1023 => x"5c5c5757",
  1024 => x"5a5a758a",
  1025 => x"2e828038",
  1026 => x"7680cf2e",
  1027 => x"81f93881",
  1028 => x"18567580",
  1029 => x"eadc3479",
  1030 => x"335675ff",
  1031 => x"bd3880ea",
  1032 => x"d8337081",
  1033 => x"ff067010",
  1034 => x"101180ea",
  1035 => x"dc337081",
  1036 => x"ff067290",
  1037 => x"29117088",
  1038 => x"2ba00761",
  1039 => x"0c5a5e5a",
  1040 => x"56575879",
  1041 => x"80cf2e83",
  1042 => x"c5388117",
  1043 => x"587780ea",
  1044 => x"dc347c7c",
  1045 => x"2e83d438",
  1046 => x"80d8b80b",
  1047 => x"80d8b833",
  1048 => x"555a7380",
  1049 => x"2e80c738",
  1050 => x"7356811a",
  1051 => x"80ead833",
  1052 => x"7081ff06",
  1053 => x"70101011",
  1054 => x"80eadc33",
  1055 => x"7081ff06",
  1056 => x"72902911",
  1057 => x"70882b7d",
  1058 => x"07620c42",
  1059 => x"5c5c5757",
  1060 => x"5a5a758a",
  1061 => x"2e818d38",
  1062 => x"7680cf2e",
  1063 => x"81863881",
  1064 => x"18577680",
  1065 => x"eadc3479",
  1066 => x"335675ff",
  1067 => x"bd38841d",
  1068 => x"63810544",
  1069 => x"5d9f6327",
  1070 => x"fbca387e",
  1071 => x"800cab3d",
  1072 => x"0d046117",
  1073 => x"b7155555",
  1074 => x"fcb43974",
  1075 => x"a3268180",
  1076 => x"38811956",
  1077 => x"7580ead8",
  1078 => x"34800b80",
  1079 => x"eadc3479",
  1080 => x"335675fb",
  1081 => x"b638fbf7",
  1082 => x"3974a326",
  1083 => x"80f13881",
  1084 => x"19587780",
  1085 => x"ead83480",
  1086 => x"0b80eadc",
  1087 => x"34793356",
  1088 => x"75fc9f38",
  1089 => x"fce03974",
  1090 => x"a326b738",
  1091 => x"81195776",
  1092 => x"80ead834",
  1093 => x"800b80ea",
  1094 => x"dc347933",
  1095 => x"5675fdba",
  1096 => x"38fdfb39",
  1097 => x"74a32680",
  1098 => x"c5388119",
  1099 => x"557480ea",
  1100 => x"d834800b",
  1101 => x"80eadc34",
  1102 => x"79335675",
  1103 => x"feac38fe",
  1104 => x"ed39800b",
  1105 => x"80ead834",
  1106 => x"800b80ea",
  1107 => x"dc34cb39",
  1108 => x"800b80ea",
  1109 => x"d834800b",
  1110 => x"80eadc34",
  1111 => x"ff813980",
  1112 => x"0b80ead8",
  1113 => x"34800b80",
  1114 => x"eadc34ff",
  1115 => x"9039800b",
  1116 => x"80ead834",
  1117 => x"800b80ea",
  1118 => x"dc34ffbc",
  1119 => x"3980e3a0",
  1120 => x"0880ead8",
  1121 => x"337081ff",
  1122 => x"06701010",
  1123 => x"1180eadc",
  1124 => x"337081ff",
  1125 => x"06729029",
  1126 => x"1170882b",
  1127 => x"a007770c",
  1128 => x"425a5b57",
  1129 => x"58595b74",
  1130 => x"80cf2e09",
  1131 => x"8106fbe2",
  1132 => x"3875a326",
  1133 => x"82b83881",
  1134 => x"185b7a80",
  1135 => x"ead83480",
  1136 => x"0b80eadc",
  1137 => x"347c0870",
  1138 => x"585ca353",
  1139 => x"80d4f052",
  1140 => x"7d51add5",
  1141 => x"3fa056fb",
  1142 => x"d33980e3",
  1143 => x"a00880ea",
  1144 => x"d8337081",
  1145 => x"ff067010",
  1146 => x"101180ea",
  1147 => x"dc337081",
  1148 => x"ff067290",
  1149 => x"29117088",
  1150 => x"2ba00777",
  1151 => x"0c5b5f5b",
  1152 => x"5758595b",
  1153 => x"7980cf2e",
  1154 => x"098106fc",
  1155 => x"bd3875a3",
  1156 => x"2681cc38",
  1157 => x"81185776",
  1158 => x"80ead834",
  1159 => x"800b80ea",
  1160 => x"dc347c7c",
  1161 => x"2e098106",
  1162 => x"fcae3880",
  1163 => x"d8c00b80",
  1164 => x"d8c03355",
  1165 => x"5a73802e",
  1166 => x"fcf43873",
  1167 => x"811b80ea",
  1168 => x"d8337081",
  1169 => x"ff067010",
  1170 => x"101180ea",
  1171 => x"dc337081",
  1172 => x"ff067290",
  1173 => x"29117088",
  1174 => x"2b780763",
  1175 => x"0c5b5d5d",
  1176 => x"40585b5b",
  1177 => x"56758a2e",
  1178 => x"80ca3876",
  1179 => x"80cf2e80",
  1180 => x"c3388118",
  1181 => x"597880ea",
  1182 => x"dc347933",
  1183 => x"5675802e",
  1184 => x"fcac3881",
  1185 => x"1a80ead8",
  1186 => x"337081ff",
  1187 => x"06701010",
  1188 => x"1180eadc",
  1189 => x"337081ff",
  1190 => x"06729029",
  1191 => x"1170882b",
  1192 => x"7d07620c",
  1193 => x"5a5c5c5f",
  1194 => x"575a5a75",
  1195 => x"8a2e0981",
  1196 => x"06ffb838",
  1197 => x"74a32699",
  1198 => x"38811956",
  1199 => x"7580ead8",
  1200 => x"34800b80",
  1201 => x"eadc3479",
  1202 => x"335675ff",
  1203 => x"b638fbde",
  1204 => x"39800b80",
  1205 => x"ead83480",
  1206 => x"0b80eadc",
  1207 => x"34e93980",
  1208 => x"0b80ead8",
  1209 => x"34800b80",
  1210 => x"eadc34fe",
  1211 => x"b539800b",
  1212 => x"80ead834",
  1213 => x"800b80ea",
  1214 => x"dc34fdc9",
  1215 => x"39d93d0d",
  1216 => x"80d8c851",
  1217 => x"e7863f80",
  1218 => x"e3940870",
  1219 => x"0880d8d8",
  1220 => x"535d55e6",
  1221 => x"f73fa63d",
  1222 => x"70537c81",
  1223 => x"ffff0652",
  1224 => x"5de5c93f",
  1225 => x"7c51e6e4",
  1226 => x"3f80d8ec",
  1227 => x"51e6dd3f",
  1228 => x"7b8f2a81",
  1229 => x"06a43d5a",
  1230 => x"568b5380",
  1231 => x"d4e45278",
  1232 => x"51aae63f",
  1233 => x"82028405",
  1234 => x"81890559",
  1235 => x"57758f06",
  1236 => x"54738926",
  1237 => x"89b33876",
  1238 => x"18b01555",
  1239 => x"55737534",
  1240 => x"75842aff",
  1241 => x"187081ff",
  1242 => x"06595b56",
  1243 => x"76df3878",
  1244 => x"79335557",
  1245 => x"73802ea9",
  1246 => x"387380e3",
  1247 => x"a8085656",
  1248 => x"81175775",
  1249 => x"8a2e899d",
  1250 => x"38841508",
  1251 => x"70822a81",
  1252 => x"065b5b79",
  1253 => x"802ef238",
  1254 => x"75750c76",
  1255 => x"335675e0",
  1256 => x"38787933",
  1257 => x"555a7380",
  1258 => x"2e80cc38",
  1259 => x"7380e3a0",
  1260 => x"085c5681",
  1261 => x"1a80ead8",
  1262 => x"337081ff",
  1263 => x"06701010",
  1264 => x"1180eadc",
  1265 => x"337081ff",
  1266 => x"06729029",
  1267 => x"1170882b",
  1268 => x"7d07620c",
  1269 => x"535c5c57",
  1270 => x"575a5a75",
  1271 => x"8a2e8986",
  1272 => x"387680cf",
  1273 => x"2e88ff38",
  1274 => x"81185776",
  1275 => x"80eadc34",
  1276 => x"79335675",
  1277 => x"ffbd3880",
  1278 => x"d98051e5",
  1279 => x"8f3f7b90",
  1280 => x"2a8106a1",
  1281 => x"3d5a568b",
  1282 => x"5380d4e4",
  1283 => x"527851a9",
  1284 => x"983f8202",
  1285 => x"840580fd",
  1286 => x"05595775",
  1287 => x"8f065473",
  1288 => x"892688a6",
  1289 => x"387618b0",
  1290 => x"15555573",
  1291 => x"75347584",
  1292 => x"2aff1870",
  1293 => x"81ff0659",
  1294 => x"565676df",
  1295 => x"38787933",
  1296 => x"55577380",
  1297 => x"2ea93880",
  1298 => x"e3a80874",
  1299 => x"57558117",
  1300 => x"57758a2e",
  1301 => x"88bb3884",
  1302 => x"15087082",
  1303 => x"2a810655",
  1304 => x"5873802e",
  1305 => x"f2387575",
  1306 => x"0c763356",
  1307 => x"75e03878",
  1308 => x"7933555a",
  1309 => x"73802e80",
  1310 => x"cc3880e3",
  1311 => x"a0087457",
  1312 => x"5b811a80",
  1313 => x"ead83370",
  1314 => x"81ff0670",
  1315 => x"10101180",
  1316 => x"eadc3370",
  1317 => x"81ff0672",
  1318 => x"90291170",
  1319 => x"882b7d07",
  1320 => x"620c535c",
  1321 => x"5c57575a",
  1322 => x"5a758a2e",
  1323 => x"93a13876",
  1324 => x"80cf2e93",
  1325 => x"9a388118",
  1326 => x"577680ea",
  1327 => x"dc347933",
  1328 => x"5675ffbd",
  1329 => x"3880d994",
  1330 => x"51e3c13f",
  1331 => x"7b952a83",
  1332 => x"06547381",
  1333 => x"2e94fa38",
  1334 => x"81742694",
  1335 => x"ea387382",
  1336 => x"2e94f838",
  1337 => x"73832e88",
  1338 => x"e13880d9",
  1339 => x"a851e39c",
  1340 => x"3f7c527b",
  1341 => x"972a8706",
  1342 => x"83058171",
  1343 => x"2b525ae1",
  1344 => x"eb3f7c51",
  1345 => x"e3863f80",
  1346 => x"d9bc51e2",
  1347 => x"ff3f80d9",
  1348 => x"c451e2f8",
  1349 => x"3f7c527b",
  1350 => x"9a2a8106",
  1351 => x"810551e1",
  1352 => x"cb3f7c51",
  1353 => x"e2e63f80",
  1354 => x"d9d851e2",
  1355 => x"df3f7c52",
  1356 => x"7b9b2a87",
  1357 => x"06830551",
  1358 => x"e1b23f7c",
  1359 => x"51e2cd3f",
  1360 => x"80d9ec51",
  1361 => x"e2c63f7c",
  1362 => x"527b9e2a",
  1363 => x"820751e1",
  1364 => x"9b3f7c51",
  1365 => x"e2b63f80",
  1366 => x"da8051e2",
  1367 => x"af3f7b9f",
  1368 => x"2a9e3d5a",
  1369 => x"568b5380",
  1370 => x"d4e45278",
  1371 => x"51a6ba3f",
  1372 => x"82028405",
  1373 => x"80f10559",
  1374 => x"57758f06",
  1375 => x"54738926",
  1376 => x"90f63876",
  1377 => x"18b01555",
  1378 => x"55737534",
  1379 => x"75842aff",
  1380 => x"187081ff",
  1381 => x"06595d56",
  1382 => x"76df3878",
  1383 => x"79335557",
  1384 => x"73802ea9",
  1385 => x"3880e3a8",
  1386 => x"08745755",
  1387 => x"81175775",
  1388 => x"8a2e8682",
  1389 => x"38841508",
  1390 => x"70822a81",
  1391 => x"06595477",
  1392 => x"802ef238",
  1393 => x"75750c76",
  1394 => x"335675e0",
  1395 => x"38787933",
  1396 => x"555a7380",
  1397 => x"2e80cc38",
  1398 => x"80e3a008",
  1399 => x"74575b81",
  1400 => x"1a80ead8",
  1401 => x"337081ff",
  1402 => x"06701010",
  1403 => x"1180eadc",
  1404 => x"337081ff",
  1405 => x"06729029",
  1406 => x"1170882b",
  1407 => x"7d07620c",
  1408 => x"5a5c5c5f",
  1409 => x"575a5a75",
  1410 => x"8a2e90e1",
  1411 => x"387680cf",
  1412 => x"2e90da38",
  1413 => x"81185776",
  1414 => x"80eadc34",
  1415 => x"79335675",
  1416 => x"ffbd3880",
  1417 => x"e3940884",
  1418 => x"110880da",
  1419 => x"94535658",
  1420 => x"e0da3f7c",
  1421 => x"52749fff",
  1422 => x"0651dfb0",
  1423 => x"3f7c51e0",
  1424 => x"cb3f80da",
  1425 => x"a851e0c4",
  1426 => x"3f7c5274",
  1427 => x"8c2a8706",
  1428 => x"83058171",
  1429 => x"2b525bdf",
  1430 => x"933f7c51",
  1431 => x"e0ae3f74",
  1432 => x"8f2a8106",
  1433 => x"80dabc52",
  1434 => x"5ce0a13f",
  1435 => x"7b9b3d5a",
  1436 => x"568b5380",
  1437 => x"d4e45278",
  1438 => x"51a4ae3f",
  1439 => x"82028405",
  1440 => x"80e50559",
  1441 => x"57758f06",
  1442 => x"54738926",
  1443 => x"8efc3876",
  1444 => x"18b01555",
  1445 => x"55737534",
  1446 => x"75842aff",
  1447 => x"187081ff",
  1448 => x"06595556",
  1449 => x"76df3878",
  1450 => x"79335557",
  1451 => x"73802ea9",
  1452 => x"3880e3a8",
  1453 => x"08745755",
  1454 => x"81175775",
  1455 => x"8a2e849b",
  1456 => x"38841508",
  1457 => x"70822a81",
  1458 => x"06555a73",
  1459 => x"802ef238",
  1460 => x"75750c76",
  1461 => x"335675e0",
  1462 => x"38787933",
  1463 => x"555a7380",
  1464 => x"2e80cc38",
  1465 => x"80e3a008",
  1466 => x"74575b81",
  1467 => x"1a80ead8",
  1468 => x"337081ff",
  1469 => x"06701010",
  1470 => x"1180eadc",
  1471 => x"337081ff",
  1472 => x"06729029",
  1473 => x"1170882b",
  1474 => x"7d07620c",
  1475 => x"535c5c57",
  1476 => x"575a5a75",
  1477 => x"8a2e8e99",
  1478 => x"387680cf",
  1479 => x"2e8e9238",
  1480 => x"81185776",
  1481 => x"80eadc34",
  1482 => x"79335675",
  1483 => x"ffbd387b",
  1484 => x"83f33880",
  1485 => x"e3940890",
  1486 => x"110880da",
  1487 => x"d0535856",
  1488 => x"deca3f76",
  1489 => x"8f3d5a56",
  1490 => x"8b5380d4",
  1491 => x"e4527851",
  1492 => x"a2d73f88",
  1493 => x"028405b5",
  1494 => x"05595775",
  1495 => x"8f065473",
  1496 => x"89268d9d",
  1497 => x"387618b0",
  1498 => x"15555573",
  1499 => x"75347584",
  1500 => x"2aff1870",
  1501 => x"81ff0659",
  1502 => x"5c5676df",
  1503 => x"38787933",
  1504 => x"55577380",
  1505 => x"2ea93880",
  1506 => x"e3a80874",
  1507 => x"57558117",
  1508 => x"57758a2e",
  1509 => x"82ea3884",
  1510 => x"15087082",
  1511 => x"2a81065d",
  1512 => x"5b7b802e",
  1513 => x"f2387575",
  1514 => x"0c763356",
  1515 => x"75e03878",
  1516 => x"7933555a",
  1517 => x"73802e80",
  1518 => x"cc3880e3",
  1519 => x"a0087457",
  1520 => x"5b811a80",
  1521 => x"ead83370",
  1522 => x"81ff0670",
  1523 => x"10101180",
  1524 => x"eadc3370",
  1525 => x"81ff0672",
  1526 => x"90291170",
  1527 => x"882b7d07",
  1528 => x"620c425c",
  1529 => x"5c40575a",
  1530 => x"5a758a2e",
  1531 => x"8ca53876",
  1532 => x"80cf2e8c",
  1533 => x"9e388118",
  1534 => x"597880ea",
  1535 => x"dc347933",
  1536 => x"5675ffbd",
  1537 => x"38a93d0d",
  1538 => x"047618b7",
  1539 => x"15555573",
  1540 => x"75347584",
  1541 => x"2aff1870",
  1542 => x"81ff0659",
  1543 => x"5b5676f6",
  1544 => x"ac38f6cb",
  1545 => x"39841508",
  1546 => x"70822a81",
  1547 => x"06595477",
  1548 => x"802ef238",
  1549 => x"8d750c84",
  1550 => x"15087082",
  1551 => x"2a81065b",
  1552 => x"5b79802e",
  1553 => x"f6c338f6",
  1554 => x"cf397618",
  1555 => x"b7155555",
  1556 => x"73753475",
  1557 => x"842aff18",
  1558 => x"7081ff06",
  1559 => x"59565676",
  1560 => x"f7b938f7",
  1561 => x"d83974a3",
  1562 => x"26993881",
  1563 => x"19567580",
  1564 => x"ead83480",
  1565 => x"0b80eadc",
  1566 => x"34793356",
  1567 => x"75f6b438",
  1568 => x"f6f53980",
  1569 => x"0b80ead8",
  1570 => x"34800b80",
  1571 => x"eadc34e9",
  1572 => x"39841508",
  1573 => x"70822a81",
  1574 => x"065b5b79",
  1575 => x"802ef238",
  1576 => x"8d750c84",
  1577 => x"15087082",
  1578 => x"2a810655",
  1579 => x"5873802e",
  1580 => x"f7a538f7",
  1581 => x"b1398415",
  1582 => x"0870822a",
  1583 => x"8106555a",
  1584 => x"73802ef2",
  1585 => x"388d750c",
  1586 => x"84150870",
  1587 => x"822a8106",
  1588 => x"59547780",
  1589 => x"2ef9de38",
  1590 => x"f9ea3984",
  1591 => x"15087082",
  1592 => x"2a81065c",
  1593 => x"587a802e",
  1594 => x"f2388d75",
  1595 => x"0c841508",
  1596 => x"70822a81",
  1597 => x"06555a73",
  1598 => x"802efbc5",
  1599 => x"38fbd139",
  1600 => x"84150870",
  1601 => x"822a8106",
  1602 => x"59547780",
  1603 => x"2ef2388d",
  1604 => x"750c8415",
  1605 => x"0870822a",
  1606 => x"81065d5b",
  1607 => x"7b802efc",
  1608 => x"f638fd82",
  1609 => x"3980e394",
  1610 => x"08881108",
  1611 => x"80dae453",
  1612 => x"565cdad8",
  1613 => x"3f748706",
  1614 => x"54738626",
  1615 => x"81a53873",
  1616 => x"101080e2",
  1617 => x"b0055978",
  1618 => x"080480da",
  1619 => x"f851dabc",
  1620 => x"3f80d9a8",
  1621 => x"51dab53f",
  1622 => x"7c527b97",
  1623 => x"2a870683",
  1624 => x"0581712b",
  1625 => x"525ad984",
  1626 => x"3f7c51da",
  1627 => x"9f3f80d9",
  1628 => x"bc51da98",
  1629 => x"3f80d9c4",
  1630 => x"51da913f",
  1631 => x"7c527b9a",
  1632 => x"2a810681",
  1633 => x"0551d8e4",
  1634 => x"3f7c51d9",
  1635 => x"ff3f80d9",
  1636 => x"d851d9f8",
  1637 => x"3f7c527b",
  1638 => x"9b2a8706",
  1639 => x"830551d8",
  1640 => x"cb3f7c51",
  1641 => x"d9e63f80",
  1642 => x"d9ec51d9",
  1643 => x"df3f7c52",
  1644 => x"7b9e2a82",
  1645 => x"0751d8b4",
  1646 => x"3f7c51d9",
  1647 => x"cf3f80da",
  1648 => x"8051d9c8",
  1649 => x"3f7b9f2a",
  1650 => x"9e3d5a56",
  1651 => x"8b5380d4",
  1652 => x"e4527851",
  1653 => x"9dd33f82",
  1654 => x"02840580",
  1655 => x"f1055957",
  1656 => x"f7973980",
  1657 => x"db8051d9",
  1658 => x"a33f80db",
  1659 => x"8851d99c",
  1660 => x"3f80db90",
  1661 => x"51d9953f",
  1662 => x"74832a83",
  1663 => x"06547381",
  1664 => x"2e90e238",
  1665 => x"8174268a",
  1666 => x"e6387382",
  1667 => x"2e90ea38",
  1668 => x"73832e90",
  1669 => x"c63880db",
  1670 => x"a451d8f0",
  1671 => x"3f80dba8",
  1672 => x"51d8e93f",
  1673 => x"74852a87",
  1674 => x"06547381",
  1675 => x"2e90c038",
  1676 => x"8174268a",
  1677 => x"b0387382",
  1678 => x"2e90c838",
  1679 => x"73832e90",
  1680 => x"903880db",
  1681 => x"bc51d8c4",
  1682 => x"3f74902a",
  1683 => x"87065473",
  1684 => x"85268c38",
  1685 => x"73101080",
  1686 => x"e2cc0554",
  1687 => x"73080480",
  1688 => x"db8051d8",
  1689 => x"a73f80db",
  1690 => x"d051d8a0",
  1691 => x"3f7c5274",
  1692 => x"932a8306",
  1693 => x"820751d6",
  1694 => x"f33f7c51",
  1695 => x"d88e3f80",
  1696 => x"dbe451d8",
  1697 => x"873f7c52",
  1698 => x"74942a8f",
  1699 => x"0651d6dc",
  1700 => x"3f7c51d7",
  1701 => x"f73f80db",
  1702 => x"f851d7f0",
  1703 => x"3f7c5274",
  1704 => x"982a8106",
  1705 => x"810551d6",
  1706 => x"c33f7c51",
  1707 => x"d7de3f80",
  1708 => x"dc8c51d7",
  1709 => x"d73f7c52",
  1710 => x"749e2a82",
  1711 => x"0751d6ac",
  1712 => x"3f7c51d7",
  1713 => x"c73f80dc",
  1714 => x"a051d7c0",
  1715 => x"3f749f2a",
  1716 => x"983d5a56",
  1717 => x"8b5380d4",
  1718 => x"e4527851",
  1719 => x"9bcb3f82",
  1720 => x"02840580",
  1721 => x"d9055957",
  1722 => x"758f0654",
  1723 => x"73892687",
  1724 => x"d4387618",
  1725 => x"b0155555",
  1726 => x"73753475",
  1727 => x"842aff18",
  1728 => x"7081ff06",
  1729 => x"595e5676",
  1730 => x"df387879",
  1731 => x"33555773",
  1732 => x"802ea938",
  1733 => x"80e3a808",
  1734 => x"74575581",
  1735 => x"1757758a",
  1736 => x"2e84e638",
  1737 => x"84150870",
  1738 => x"822a8106",
  1739 => x"555d7380",
  1740 => x"2ef23875",
  1741 => x"750c7633",
  1742 => x"5675e038",
  1743 => x"78793355",
  1744 => x"5a73802e",
  1745 => x"80cc3880",
  1746 => x"e3a00874",
  1747 => x"575b811a",
  1748 => x"80ead833",
  1749 => x"7081ff06",
  1750 => x"70101011",
  1751 => x"80eadc33",
  1752 => x"7081ff06",
  1753 => x"72902911",
  1754 => x"70882b7d",
  1755 => x"07620c42",
  1756 => x"5c5c4057",
  1757 => x"5a5a758a",
  1758 => x"2e878338",
  1759 => x"7680cf2e",
  1760 => x"86fc3881",
  1761 => x"18597880",
  1762 => x"eadc3479",
  1763 => x"335675ff",
  1764 => x"bd3880e3",
  1765 => x"94089411",
  1766 => x"0880dcb4",
  1767 => x"535856d5",
  1768 => x"eb3f7695",
  1769 => x"3d5a568b",
  1770 => x"5380d4e4",
  1771 => x"52785199",
  1772 => x"f83f8802",
  1773 => x"840580cd",
  1774 => x"05595775",
  1775 => x"8f065473",
  1776 => x"89268693",
  1777 => x"387618b0",
  1778 => x"15555573",
  1779 => x"75347584",
  1780 => x"2aff1870",
  1781 => x"81ff0659",
  1782 => x"5c5676df",
  1783 => x"38787933",
  1784 => x"55577380",
  1785 => x"2ea93880",
  1786 => x"e3a80874",
  1787 => x"57558117",
  1788 => x"57758a2e",
  1789 => x"83b83884",
  1790 => x"15087082",
  1791 => x"2a81065d",
  1792 => x"5b7b802e",
  1793 => x"f2387575",
  1794 => x"0c763356",
  1795 => x"75e03878",
  1796 => x"7933555a",
  1797 => x"73802e80",
  1798 => x"cc3880e3",
  1799 => x"a0087457",
  1800 => x"5b811a80",
  1801 => x"ead83370",
  1802 => x"81ff0670",
  1803 => x"10101180",
  1804 => x"eadc3370",
  1805 => x"81ff0672",
  1806 => x"90291170",
  1807 => x"882b7d07",
  1808 => x"620c425c",
  1809 => x"5c40575a",
  1810 => x"5a758a2e",
  1811 => x"85923876",
  1812 => x"80cf2e85",
  1813 => x"8b388118",
  1814 => x"597880ea",
  1815 => x"dc347933",
  1816 => x"5675ffbd",
  1817 => x"3880e394",
  1818 => x"08981108",
  1819 => x"80dcc853",
  1820 => x"5856d498",
  1821 => x"3f76923d",
  1822 => x"5a568b53",
  1823 => x"80d4e452",
  1824 => x"785198a5",
  1825 => x"3f880284",
  1826 => x"0580c105",
  1827 => x"5957758f",
  1828 => x"06547389",
  1829 => x"2684b738",
  1830 => x"7618b015",
  1831 => x"55557375",
  1832 => x"3475842a",
  1833 => x"ff187081",
  1834 => x"ff06595b",
  1835 => x"5676df38",
  1836 => x"78793355",
  1837 => x"5773802e",
  1838 => x"a93880e3",
  1839 => x"a8087457",
  1840 => x"55811757",
  1841 => x"758a2e82",
  1842 => x"8a388415",
  1843 => x"0870822a",
  1844 => x"81065d5a",
  1845 => x"7b802ef2",
  1846 => x"3875750c",
  1847 => x"76335675",
  1848 => x"e0387879",
  1849 => x"33555a73",
  1850 => x"802ef4c7",
  1851 => x"3880e3a0",
  1852 => x"0874811c",
  1853 => x"80ead833",
  1854 => x"7081ff06",
  1855 => x"70101011",
  1856 => x"80eadc33",
  1857 => x"7081ff06",
  1858 => x"72902911",
  1859 => x"70882b78",
  1860 => x"07790c44",
  1861 => x"5e5e4259",
  1862 => x"5c5c575b",
  1863 => x"758a2e80",
  1864 => x"ca387680",
  1865 => x"cf2e80c3",
  1866 => x"38811859",
  1867 => x"7880eadc",
  1868 => x"34793356",
  1869 => x"75802ef3",
  1870 => x"fa38811a",
  1871 => x"80ead833",
  1872 => x"7081ff06",
  1873 => x"70101011",
  1874 => x"80eadc33",
  1875 => x"7081ff06",
  1876 => x"72902911",
  1877 => x"70882b7d",
  1878 => x"07620c42",
  1879 => x"5c5c4057",
  1880 => x"5a5a758a",
  1881 => x"2e098106",
  1882 => x"ffb83874",
  1883 => x"a32683ab",
  1884 => x"38811955",
  1885 => x"7480ead8",
  1886 => x"34800b80",
  1887 => x"eadc3479",
  1888 => x"335675ff",
  1889 => x"b538f3ab",
  1890 => x"39841508",
  1891 => x"70822a81",
  1892 => x"06595a77",
  1893 => x"802ef238",
  1894 => x"8d750c84",
  1895 => x"15087082",
  1896 => x"2a810655",
  1897 => x"5d73802e",
  1898 => x"fafa38fb",
  1899 => x"86398415",
  1900 => x"0870822a",
  1901 => x"81065954",
  1902 => x"77802ef2",
  1903 => x"388d750c",
  1904 => x"84150870",
  1905 => x"822a8106",
  1906 => x"5d5b7b80",
  1907 => x"2efca838",
  1908 => x"fcb43984",
  1909 => x"15087082",
  1910 => x"2a810659",
  1911 => x"5477802e",
  1912 => x"f2388d75",
  1913 => x"0c841508",
  1914 => x"70822a81",
  1915 => x"065d5a7b",
  1916 => x"802efdd6",
  1917 => x"38fde239",
  1918 => x"7618b715",
  1919 => x"5555ef89",
  1920 => x"397618b7",
  1921 => x"155555f2",
  1922 => x"e2397618",
  1923 => x"b7155555",
  1924 => x"f1833974",
  1925 => x"a326819e",
  1926 => x"38811955",
  1927 => x"7480ead8",
  1928 => x"34800b80",
  1929 => x"eadc3479",
  1930 => x"335675f3",
  1931 => x"9438f3d5",
  1932 => x"3974a326",
  1933 => x"80f13881",
  1934 => x"19567580",
  1935 => x"ead83480",
  1936 => x"0b80eadc",
  1937 => x"34793356",
  1938 => x"75f1a038",
  1939 => x"f1e13974",
  1940 => x"a32680c4",
  1941 => x"38811956",
  1942 => x"7580ead8",
  1943 => x"34800b80",
  1944 => x"eadc3479",
  1945 => x"335675ec",
  1946 => x"9838ecd9",
  1947 => x"3974a326",
  1948 => x"99388119",
  1949 => x"567580ea",
  1950 => x"d834800b",
  1951 => x"80eadc34",
  1952 => x"79335675",
  1953 => x"eed938ef",
  1954 => x"9a39800b",
  1955 => x"80ead834",
  1956 => x"800b80ea",
  1957 => x"dc34e939",
  1958 => x"800b80ea",
  1959 => x"d834800b",
  1960 => x"80eadc34",
  1961 => x"ffbd3980",
  1962 => x"0b80ead8",
  1963 => x"34800b80",
  1964 => x"eadc34ff",
  1965 => x"9039800b",
  1966 => x"80ead834",
  1967 => x"800b80ea",
  1968 => x"dc34fee3",
  1969 => x"397618b7",
  1970 => x"155555f8",
  1971 => x"ab397618",
  1972 => x"b7155555",
  1973 => x"fbc83976",
  1974 => x"18b71555",
  1975 => x"55f9ec39",
  1976 => x"74a32680",
  1977 => x"d3388119",
  1978 => x"557480ea",
  1979 => x"d834800b",
  1980 => x"80eadc34",
  1981 => x"79335675",
  1982 => x"faa738fa",
  1983 => x"e83974a3",
  1984 => x"26a83881",
  1985 => x"19557480",
  1986 => x"ead83480",
  1987 => x"0b80eadc",
  1988 => x"34793356",
  1989 => x"75f8b738",
  1990 => x"f8f83980",
  1991 => x"0b80ead8",
  1992 => x"34800b80",
  1993 => x"eadc34fc",
  1994 => x"d639800b",
  1995 => x"80ead834",
  1996 => x"800b80ea",
  1997 => x"dc34da39",
  1998 => x"800b80ea",
  1999 => x"d834800b",
  2000 => x"80eadc34",
  2001 => x"ffae3980",
  2002 => x"dcdc51ce",
  2003 => x"bf3ff481",
  2004 => x"3980dce4",
  2005 => x"51ceb53f",
  2006 => x"f3f73980",
  2007 => x"dcec51ce",
  2008 => x"ab3ff3ed",
  2009 => x"3980dcf4",
  2010 => x"51cea13f",
  2011 => x"f5d43980",
  2012 => x"dcfc51ce",
  2013 => x"973ff59e",
  2014 => x"3980dd80",
  2015 => x"51f4e839",
  2016 => x"80dd8451",
  2017 => x"f4e13980",
  2018 => x"dd8851f4",
  2019 => x"da3980dd",
  2020 => x"8c51f4d3",
  2021 => x"3980dd90",
  2022 => x"51cdf13f",
  2023 => x"80dbd051",
  2024 => x"cdea3f7c",
  2025 => x"5274932a",
  2026 => x"83068207",
  2027 => x"51ccbd3f",
  2028 => x"7c51cdd8",
  2029 => x"3f80dbe4",
  2030 => x"51cdd13f",
  2031 => x"7c527494",
  2032 => x"2a8f0651",
  2033 => x"cca63f7c",
  2034 => x"51cdc13f",
  2035 => x"80dbf851",
  2036 => x"cdba3f7c",
  2037 => x"5274982a",
  2038 => x"81068105",
  2039 => x"51cc8d3f",
  2040 => x"7c51cda8",
  2041 => x"3f80dc8c",
  2042 => x"51cda13f",
  2043 => x"7c52749e",
  2044 => x"2a820751",
  2045 => x"cbf63f7c",
  2046 => x"51cd913f",
  2047 => x"80dca051",
  2048 => x"cd8a3f74",
  2049 => x"9f2a983d",
  2050 => x"5a568b53",
  2051 => x"80d4e452",
  2052 => x"78519195",
  2053 => x"3f820284",
  2054 => x"0580d905",
  2055 => x"5957f5c8",
  2056 => x"3980dda0",
  2057 => x"51cce53f",
  2058 => x"80dbd051",
  2059 => x"ccde3f7c",
  2060 => x"5274932a",
  2061 => x"83068207",
  2062 => x"51cbb13f",
  2063 => x"7c51cccc",
  2064 => x"3f80dbe4",
  2065 => x"51ccc53f",
  2066 => x"7c527494",
  2067 => x"2a8f0651",
  2068 => x"cb9a3f7c",
  2069 => x"51ccb53f",
  2070 => x"80dbf851",
  2071 => x"ccae3f7c",
  2072 => x"5274982a",
  2073 => x"81068105",
  2074 => x"51cb813f",
  2075 => x"7c51cc9c",
  2076 => x"3f80dc8c",
  2077 => x"51cc953f",
  2078 => x"7c52749e",
  2079 => x"2a820751",
  2080 => x"caea3f7c",
  2081 => x"51cc853f",
  2082 => x"80dca051",
  2083 => x"cbfe3f74",
  2084 => x"9f2a983d",
  2085 => x"5a568b53",
  2086 => x"80d4e452",
  2087 => x"78519089",
  2088 => x"3f820284",
  2089 => x"0580d905",
  2090 => x"5957f4bc",
  2091 => x"3980ddac",
  2092 => x"51cbd93f",
  2093 => x"80dbd051",
  2094 => x"cbd23f7c",
  2095 => x"5274932a",
  2096 => x"83068207",
  2097 => x"51caa53f",
  2098 => x"7c51cbc0",
  2099 => x"3f80dbe4",
  2100 => x"51cbb93f",
  2101 => x"7c527494",
  2102 => x"2a8f0651",
  2103 => x"ca8e3f7c",
  2104 => x"51cba93f",
  2105 => x"80dbf851",
  2106 => x"cba23f7c",
  2107 => x"5274982a",
  2108 => x"81068105",
  2109 => x"51c9f53f",
  2110 => x"7c51cb90",
  2111 => x"3f80dc8c",
  2112 => x"51cb893f",
  2113 => x"7c52749e",
  2114 => x"2a820751",
  2115 => x"c9de3f7c",
  2116 => x"51caf93f",
  2117 => x"80dca051",
  2118 => x"caf23f74",
  2119 => x"9f2a983d",
  2120 => x"5a568b53",
  2121 => x"80d4e452",
  2122 => x"78518efd",
  2123 => x"3f820284",
  2124 => x"0580d905",
  2125 => x"5957f3b0",
  2126 => x"3980ddbc",
  2127 => x"51cacd3f",
  2128 => x"80dbd051",
  2129 => x"cac63f7c",
  2130 => x"5274932a",
  2131 => x"83068207",
  2132 => x"51c9993f",
  2133 => x"7c51cab4",
  2134 => x"3f80dbe4",
  2135 => x"51caad3f",
  2136 => x"7c527494",
  2137 => x"2a8f0651",
  2138 => x"c9823f7c",
  2139 => x"51ca9d3f",
  2140 => x"80dbf851",
  2141 => x"ca963f7c",
  2142 => x"5274982a",
  2143 => x"81068105",
  2144 => x"51c8e93f",
  2145 => x"7c51ca84",
  2146 => x"3f80dc8c",
  2147 => x"51c9fd3f",
  2148 => x"7c52749e",
  2149 => x"2a820751",
  2150 => x"c8d23f7c",
  2151 => x"51c9ed3f",
  2152 => x"80dca051",
  2153 => x"c9e63f74",
  2154 => x"9f2a983d",
  2155 => x"5a568b53",
  2156 => x"80d4e452",
  2157 => x"78518df1",
  2158 => x"3f820284",
  2159 => x"0580d905",
  2160 => x"5957f2a4",
  2161 => x"3980ddc8",
  2162 => x"51c9c13f",
  2163 => x"80dbd051",
  2164 => x"c9ba3f7c",
  2165 => x"5274932a",
  2166 => x"83068207",
  2167 => x"51c88d3f",
  2168 => x"7c51c9a8",
  2169 => x"3f80dbe4",
  2170 => x"51c9a13f",
  2171 => x"7c527494",
  2172 => x"2a8f0651",
  2173 => x"c7f63f7c",
  2174 => x"51c9913f",
  2175 => x"80dbf851",
  2176 => x"c98a3f7c",
  2177 => x"5274982a",
  2178 => x"81068105",
  2179 => x"51c7dd3f",
  2180 => x"7c51c8f8",
  2181 => x"3f80dc8c",
  2182 => x"51c8f13f",
  2183 => x"7c52749e",
  2184 => x"2a820751",
  2185 => x"c7c63f7c",
  2186 => x"51c8e13f",
  2187 => x"80dca051",
  2188 => x"c8da3f74",
  2189 => x"9f2a983d",
  2190 => x"5a568b53",
  2191 => x"80d4e452",
  2192 => x"78518ce5",
  2193 => x"3f820284",
  2194 => x"0580d905",
  2195 => x"5957f198",
  2196 => x"3980ddd0",
  2197 => x"51c8b53f",
  2198 => x"efe83980",
  2199 => x"ddd451c8",
  2200 => x"ab3fefb2",
  2201 => x"3980ddd8",
  2202 => x"51c8a13f",
  2203 => x"efa83980",
  2204 => x"dddc51c8",
  2205 => x"973fefca",
  2206 => x"3980dde4",
  2207 => x"51c88d3f",
  2208 => x"ef943980",
  2209 => x"dd8451c8",
  2210 => x"833fefb6",
  2211 => x"39e93d0d",
  2212 => x"80e39408",
  2213 => x"84110870",
  2214 => x"9fff0651",
  2215 => x"54548a54",
  2216 => x"bb732783",
  2217 => x"388f5472",
  2218 => x"5287e851",
  2219 => x"87b53f80",
  2220 => x"08fd0574",
  2221 => x"297083ff",
  2222 => x"ff065a55",
  2223 => x"80705d5e",
  2224 => x"f17e5e5a",
  2225 => x"8f0b80e3",
  2226 => x"98087a30",
  2227 => x"56595b8c",
  2228 => x"18085673",
  2229 => x"76249638",
  2230 => x"800b8419",
  2231 => x"0c770857",
  2232 => x"76ed3877",
  2233 => x"08577680",
  2234 => x"2ef338e3",
  2235 => x"397b307c",
  2236 => x"07708025",
  2237 => x"7e813207",
  2238 => x"54547280",
  2239 => x"2e80fb38",
  2240 => x"8c180855",
  2241 => x"74792480",
  2242 => x"f1388057",
  2243 => x"890a558f",
  2244 => x"ff567408",
  2245 => x"75327030",
  2246 => x"70720770",
  2247 => x"9f2a7a05",
  2248 => x"8419ff1b",
  2249 => x"5b595a51",
  2250 => x"54547580",
  2251 => x"25e43876",
  2252 => x"83ffff06",
  2253 => x"7c813254",
  2254 => x"54739238",
  2255 => x"81707406",
  2256 => x"57557580",
  2257 => x"2e873874",
  2258 => x"8c19085b",
  2259 => x"5c73802e",
  2260 => x"92388170",
  2261 => x"7d065654",
  2262 => x"74802e87",
  2263 => x"38738c19",
  2264 => x"085c5d80",
  2265 => x"0b88190c",
  2266 => x"77085776",
  2267 => x"feff3877",
  2268 => x"08577680",
  2269 => x"2ef238fe",
  2270 => x"f439739f",
  2271 => x"2a537c80",
  2272 => x"2e82b138",
  2273 => x"81707406",
  2274 => x"5a557880",
  2275 => x"2e82a538",
  2276 => x"7a7a3156",
  2277 => x"9e762582",
  2278 => x"9f38759f",
  2279 => x"2a167076",
  2280 => x"2c7c7131",
  2281 => x"778c1c08",
  2282 => x"70733153",
  2283 => x"5b52525f",
  2284 => x"54807425",
  2285 => x"9938ff14",
  2286 => x"54800b84",
  2287 => x"190c7708",
  2288 => x"5372ee38",
  2289 => x"77085372",
  2290 => x"802ef338",
  2291 => x"e439800b",
  2292 => x"80e3a008",
  2293 => x"56547388",
  2294 => x"2b750c81",
  2295 => x"14549790",
  2296 => x"7426f338",
  2297 => x"800b80ea",
  2298 => x"d834800b",
  2299 => x"80eadc34",
  2300 => x"80d88451",
  2301 => x"c5963f7d",
  2302 => x"802e81ca",
  2303 => x"3880dff0",
  2304 => x"51c5893f",
  2305 => x"80d88451",
  2306 => x"c5823f7b",
  2307 => x"802e81c4",
  2308 => x"3880dffc",
  2309 => x"51c4f53f",
  2310 => x"80d88451",
  2311 => x"c4ee3f7c",
  2312 => x"802e81a9",
  2313 => x"3880debc",
  2314 => x"51c4e13f",
  2315 => x"80dec851",
  2316 => x"c4da3f94",
  2317 => x"3d70537a",
  2318 => x"525cc3b0",
  2319 => x"3f7b51c4",
  2320 => x"cb3f80de",
  2321 => x"d851c4c4",
  2322 => x"3f7b527a",
  2323 => x"51c39d3f",
  2324 => x"7b51c4b8",
  2325 => x"3f80d884",
  2326 => x"51c4b13f",
  2327 => x"80dee851",
  2328 => x"c4aa3f7b",
  2329 => x"527551c3",
  2330 => x"833f7b51",
  2331 => x"c49e3f80",
  2332 => x"def851c4",
  2333 => x"973f7b52",
  2334 => x"759f2a16",
  2335 => x"70812c52",
  2336 => x"5bc2e93f",
  2337 => x"7b51c484",
  2338 => x"3f80d884",
  2339 => x"51c3fd3f",
  2340 => x"80dfb851",
  2341 => x"c3f63f7b",
  2342 => x"5280e398",
  2343 => x"088c1108",
  2344 => x"525ac2c8",
  2345 => x"3f7b51c3",
  2346 => x"e33f7d81",
  2347 => x"ff06800c",
  2348 => x"993d0d04",
  2349 => x"7a7a3156",
  2350 => x"a80b8c19",
  2351 => x"08707231",
  2352 => x"525854fd",
  2353 => x"ec3980e0",
  2354 => x"8851feb5",
  2355 => x"3980dfd0",
  2356 => x"51fed639",
  2357 => x"80e09851",
  2358 => x"febb39f7",
  2359 => x"3d0d800b",
  2360 => x"80e39c08",
  2361 => x"7008810a",
  2362 => x"0680ead4",
  2363 => x"0c5355c1",
  2364 => x"ea3f80e3",
  2365 => x"a80853b6",
  2366 => x"0b8c140c",
  2367 => x"830b8814",
  2368 => x"0c80e3a0",
  2369 => x"08758412",
  2370 => x"0c52fe80",
  2371 => x"0a0b8813",
  2372 => x"0c7480ea",
  2373 => x"d8347480",
  2374 => x"eadc3480",
  2375 => x"e3940853",
  2376 => x"fac98e86",
  2377 => x"8c730c72",
  2378 => x"0870842a",
  2379 => x"81065154",
  2380 => x"73f53880",
  2381 => x"e0a851c2",
  2382 => x"d33f80ea",
  2383 => x"d408802e",
  2384 => x"829a3880",
  2385 => x"e0b051c2",
  2386 => x"c33f80e0",
  2387 => x"c051c2bc",
  2388 => x"3f890a52",
  2389 => x"83ffff53",
  2390 => x"71720c84",
  2391 => x"12ff1454",
  2392 => x"52728025",
  2393 => x"f33880d7",
  2394 => x"d451c2a0",
  2395 => x"3fdb8e3f",
  2396 => x"8551ffbf",
  2397 => x"bd3ffa95",
  2398 => x"3f8551ff",
  2399 => x"bfb43f80",
  2400 => x"0b80e3a0",
  2401 => x"08555372",
  2402 => x"882b740c",
  2403 => x"81135397",
  2404 => x"907326f3",
  2405 => x"38800b80",
  2406 => x"ead83480",
  2407 => x"0b80eadc",
  2408 => x"347451c5",
  2409 => x"bf3f80e3",
  2410 => x"9c087008",
  2411 => x"70872a81",
  2412 => x"06515553",
  2413 => x"73802e8b",
  2414 => x"3880e398",
  2415 => x"0852800b",
  2416 => x"84130c72",
  2417 => x"0870842a",
  2418 => x"81065154",
  2419 => x"73802e8b",
  2420 => x"3880e398",
  2421 => x"0852800b",
  2422 => x"88130c72",
  2423 => x"0870852a",
  2424 => x"81065154",
  2425 => x"73802ebc",
  2426 => x"3880e394",
  2427 => x"0853fac9",
  2428 => x"8e868c73",
  2429 => x"0c720870",
  2430 => x"842a8106",
  2431 => x"515271f5",
  2432 => x"38f98a3f",
  2433 => x"8551ffbe",
  2434 => x"a93f890a",
  2435 => x"5283ffff",
  2436 => x"5371720c",
  2437 => x"8412ff14",
  2438 => x"54527280",
  2439 => x"25f33880",
  2440 => x"e39c0853",
  2441 => x"72087086",
  2442 => x"2a810654",
  2443 => x"5272802e",
  2444 => x"feef3880",
  2445 => x"0b80e3a0",
  2446 => x"08555372",
  2447 => x"882b740c",
  2448 => x"81135397",
  2449 => x"907326f3",
  2450 => x"38800b80",
  2451 => x"ead83480",
  2452 => x"0b80eadc",
  2453 => x"34748132",
  2454 => x"55fec639",
  2455 => x"80e0e451",
  2456 => x"fde5398c",
  2457 => x"08028c0c",
  2458 => x"fd3d0d80",
  2459 => x"538c088c",
  2460 => x"0508528c",
  2461 => x"08880508",
  2462 => x"5182de3f",
  2463 => x"80087080",
  2464 => x"0c54853d",
  2465 => x"0d8c0c04",
  2466 => x"8c08028c",
  2467 => x"0cfd3d0d",
  2468 => x"81538c08",
  2469 => x"8c050852",
  2470 => x"8c088805",
  2471 => x"085182b9",
  2472 => x"3f800870",
  2473 => x"800c5485",
  2474 => x"3d0d8c0c",
  2475 => x"048c0802",
  2476 => x"8c0cf93d",
  2477 => x"0d800b8c",
  2478 => x"08fc050c",
  2479 => x"8c088805",
  2480 => x"088025ab",
  2481 => x"388c0888",
  2482 => x"0508308c",
  2483 => x"0888050c",
  2484 => x"800b8c08",
  2485 => x"f4050c8c",
  2486 => x"08fc0508",
  2487 => x"8838810b",
  2488 => x"8c08f405",
  2489 => x"0c8c08f4",
  2490 => x"05088c08",
  2491 => x"fc050c8c",
  2492 => x"088c0508",
  2493 => x"8025ab38",
  2494 => x"8c088c05",
  2495 => x"08308c08",
  2496 => x"8c050c80",
  2497 => x"0b8c08f0",
  2498 => x"050c8c08",
  2499 => x"fc050888",
  2500 => x"38810b8c",
  2501 => x"08f0050c",
  2502 => x"8c08f005",
  2503 => x"088c08fc",
  2504 => x"050c8053",
  2505 => x"8c088c05",
  2506 => x"08528c08",
  2507 => x"88050851",
  2508 => x"81a73f80",
  2509 => x"08708c08",
  2510 => x"f8050c54",
  2511 => x"8c08fc05",
  2512 => x"08802e8c",
  2513 => x"388c08f8",
  2514 => x"0508308c",
  2515 => x"08f8050c",
  2516 => x"8c08f805",
  2517 => x"0870800c",
  2518 => x"54893d0d",
  2519 => x"8c0c048c",
  2520 => x"08028c0c",
  2521 => x"fb3d0d80",
  2522 => x"0b8c08fc",
  2523 => x"050c8c08",
  2524 => x"88050880",
  2525 => x"2593388c",
  2526 => x"08880508",
  2527 => x"308c0888",
  2528 => x"050c810b",
  2529 => x"8c08fc05",
  2530 => x"0c8c088c",
  2531 => x"05088025",
  2532 => x"8c388c08",
  2533 => x"8c050830",
  2534 => x"8c088c05",
  2535 => x"0c81538c",
  2536 => x"088c0508",
  2537 => x"528c0888",
  2538 => x"050851ad",
  2539 => x"3f800870",
  2540 => x"8c08f805",
  2541 => x"0c548c08",
  2542 => x"fc050880",
  2543 => x"2e8c388c",
  2544 => x"08f80508",
  2545 => x"308c08f8",
  2546 => x"050c8c08",
  2547 => x"f8050870",
  2548 => x"800c5487",
  2549 => x"3d0d8c0c",
  2550 => x"048c0802",
  2551 => x"8c0cfd3d",
  2552 => x"0d810b8c",
  2553 => x"08fc050c",
  2554 => x"800b8c08",
  2555 => x"f8050c8c",
  2556 => x"088c0508",
  2557 => x"8c088805",
  2558 => x"0827ac38",
  2559 => x"8c08fc05",
  2560 => x"08802ea3",
  2561 => x"38800b8c",
  2562 => x"088c0508",
  2563 => x"2499388c",
  2564 => x"088c0508",
  2565 => x"108c088c",
  2566 => x"050c8c08",
  2567 => x"fc050810",
  2568 => x"8c08fc05",
  2569 => x"0cc9398c",
  2570 => x"08fc0508",
  2571 => x"802e80c9",
  2572 => x"388c088c",
  2573 => x"05088c08",
  2574 => x"88050826",
  2575 => x"a1388c08",
  2576 => x"8805088c",
  2577 => x"088c0508",
  2578 => x"318c0888",
  2579 => x"050c8c08",
  2580 => x"f805088c",
  2581 => x"08fc0508",
  2582 => x"078c08f8",
  2583 => x"050c8c08",
  2584 => x"fc050881",
  2585 => x"2a8c08fc",
  2586 => x"050c8c08",
  2587 => x"8c050881",
  2588 => x"2a8c088c",
  2589 => x"050cffaf",
  2590 => x"398c0890",
  2591 => x"0508802e",
  2592 => x"8f388c08",
  2593 => x"88050870",
  2594 => x"8c08f405",
  2595 => x"0c518d39",
  2596 => x"8c08f805",
  2597 => x"08708c08",
  2598 => x"f4050c51",
  2599 => x"8c08f405",
  2600 => x"08800c85",
  2601 => x"3d0d8c0c",
  2602 => x"04fc3d0d",
  2603 => x"7670797b",
  2604 => x"55555555",
  2605 => x"8f72278c",
  2606 => x"38727507",
  2607 => x"83065170",
  2608 => x"802ea738",
  2609 => x"ff125271",
  2610 => x"ff2e9838",
  2611 => x"72708105",
  2612 => x"54337470",
  2613 => x"81055634",
  2614 => x"ff125271",
  2615 => x"ff2e0981",
  2616 => x"06ea3874",
  2617 => x"800c863d",
  2618 => x"0d047451",
  2619 => x"72708405",
  2620 => x"54087170",
  2621 => x"8405530c",
  2622 => x"72708405",
  2623 => x"54087170",
  2624 => x"8405530c",
  2625 => x"72708405",
  2626 => x"54087170",
  2627 => x"8405530c",
  2628 => x"72708405",
  2629 => x"54087170",
  2630 => x"8405530c",
  2631 => x"f0125271",
  2632 => x"8f26c938",
  2633 => x"83722795",
  2634 => x"38727084",
  2635 => x"05540871",
  2636 => x"70840553",
  2637 => x"0cfc1252",
  2638 => x"718326ed",
  2639 => x"387054ff",
  2640 => x"8339fd3d",
  2641 => x"0d800b80",
  2642 => x"e3880854",
  2643 => x"5472812e",
  2644 => x"9c387380",
  2645 => x"eae00cff",
  2646 => x"b6863fff",
  2647 => x"b5a23f80",
  2648 => x"e3ac5281",
  2649 => x"51f6f43f",
  2650 => x"800851a2",
  2651 => x"3f7280ea",
  2652 => x"e00cffb5",
  2653 => x"eb3fffb5",
  2654 => x"873f80e3",
  2655 => x"ac528151",
  2656 => x"f6d93f80",
  2657 => x"0851873f",
  2658 => x"00ff3900",
  2659 => x"ff39f73d",
  2660 => x"0d7b80e3",
  2661 => x"b00882c8",
  2662 => x"11085a54",
  2663 => x"5a77802e",
  2664 => x"80da3881",
  2665 => x"88188419",
  2666 => x"08ff0581",
  2667 => x"712b5955",
  2668 => x"59807424",
  2669 => x"80ea3880",
  2670 => x"7424b538",
  2671 => x"73822b78",
  2672 => x"11880556",
  2673 => x"56818019",
  2674 => x"08770653",
  2675 => x"72802eb6",
  2676 => x"38781670",
  2677 => x"08535379",
  2678 => x"51740853",
  2679 => x"722dff14",
  2680 => x"fc17fc17",
  2681 => x"79812c5a",
  2682 => x"57575473",
  2683 => x"8025d638",
  2684 => x"77085877",
  2685 => x"ffad3880",
  2686 => x"e3b00853",
  2687 => x"bc1308a5",
  2688 => x"387951ff",
  2689 => x"833f7408",
  2690 => x"53722dff",
  2691 => x"14fc17fc",
  2692 => x"1779812c",
  2693 => x"5a575754",
  2694 => x"738025ff",
  2695 => x"a838d139",
  2696 => x"8057ff93",
  2697 => x"397251bc",
  2698 => x"13085372",
  2699 => x"2d7951fe",
  2700 => x"d73fff3d",
  2701 => x"0d80eab4",
  2702 => x"0bfc0570",
  2703 => x"08525270",
  2704 => x"ff2e9138",
  2705 => x"702dfc12",
  2706 => x"70085252",
  2707 => x"70ff2e09",
  2708 => x"8106f138",
  2709 => x"833d0d04",
  2710 => x"04ffb4f1",
  2711 => x"3f040000",
  2712 => x"00000040",
  2713 => x"30782020",
  2714 => x"20202020",
  2715 => x"20200000",
  2716 => x"30622020",
  2717 => x"20202020",
  2718 => x"20202020",
  2719 => x"20202020",
  2720 => x"20202020",
  2721 => x"20202020",
  2722 => x"20202020",
  2723 => x"20202020",
  2724 => x"20200000",
  2725 => x"0a677265",
  2726 => x"74682072",
  2727 => x"65676973",
  2728 => x"74657273",
  2729 => x"3a000000",
  2730 => x"0a636f6e",
  2731 => x"74726f6c",
  2732 => x"3a202020",
  2733 => x"20202000",
  2734 => x"0a737461",
  2735 => x"7475733a",
  2736 => x"20202020",
  2737 => x"20202000",
  2738 => x"0a6d6163",
  2739 => x"5f6d7362",
  2740 => x"3a202020",
  2741 => x"20202000",
  2742 => x"0a6d6163",
  2743 => x"5f6c7362",
  2744 => x"3a202020",
  2745 => x"20202000",
  2746 => x"0a6d6469",
  2747 => x"6f5f636f",
  2748 => x"6e74726f",
  2749 => x"6c3a2000",
  2750 => x"0a74785f",
  2751 => x"706f696e",
  2752 => x"7465723a",
  2753 => x"20202000",
  2754 => x"0a72785f",
  2755 => x"706f696e",
  2756 => x"7465723a",
  2757 => x"20202000",
  2758 => x"0a656463",
  2759 => x"6c5f6970",
  2760 => x"3a202020",
  2761 => x"20202000",
  2762 => x"0a686173",
  2763 => x"685f6d73",
  2764 => x"623a2020",
  2765 => x"20202000",
  2766 => x"0a686173",
  2767 => x"685f6c73",
  2768 => x"623a2020",
  2769 => x"20202000",
  2770 => x"0a6d6469",
  2771 => x"6f207068",
  2772 => x"79207265",
  2773 => x"67697374",
  2774 => x"65727300",
  2775 => x"0a206d64",
  2776 => x"696f2070",
  2777 => x"68793a20",
  2778 => x"00000000",
  2779 => x"0a202072",
  2780 => x"65673a20",
  2781 => x"00000000",
  2782 => x"2d3e2000",
  2783 => x"0a677265",
  2784 => x"74682d3e",
  2785 => x"636f6e74",
  2786 => x"726f6c20",
  2787 => x"3a000000",
  2788 => x"0a677265",
  2789 => x"74682d3e",
  2790 => x"73746174",
  2791 => x"75732020",
  2792 => x"3a000000",
  2793 => x"0a646573",
  2794 => x"63722d3e",
  2795 => x"636f6e74",
  2796 => x"726f6c20",
  2797 => x"3a000000",
  2798 => x"77726974",
  2799 => x"65206164",
  2800 => x"64726573",
  2801 => x"733a2000",
  2802 => x"20206c65",
  2803 => x"6e677468",
  2804 => x"3a200000",
  2805 => x"0a0a0000",
  2806 => x"72656164",
  2807 => x"20206164",
  2808 => x"64726573",
  2809 => x"733a2000",
  2810 => x"20206578",
  2811 => x"70656374",
  2812 => x"3a200000",
  2813 => x"2020676f",
  2814 => x"743a2000",
  2815 => x"20657272",
  2816 => x"6f720000",
  2817 => x"0a000000",
  2818 => x"206f6b00",
  2819 => x"70686173",
  2820 => x"65207368",
  2821 => x"69667420",
  2822 => x"202d2020",
  2823 => x"76616c75",
  2824 => x"653a2000",
  2825 => x"20207374",
  2826 => x"61747573",
  2827 => x"3a200000",
  2828 => x"20202020",
  2829 => x"20000000",
  2830 => x"4641494c",
  2831 => x"00000000",
  2832 => x"6f6b2020",
  2833 => x"00000000",
  2834 => x"44445220",
  2835 => x"6d656d6f",
  2836 => x"72792069",
  2837 => x"6e666f00",
  2838 => x"0a0a6175",
  2839 => x"746f2074",
  2840 => x"5f524552",
  2841 => x"45534820",
  2842 => x"3a000000",
  2843 => x"0a636c6f",
  2844 => x"636b2065",
  2845 => x"6e61626c",
  2846 => x"6520203a",
  2847 => x"00000000",
  2848 => x"0a696e69",
  2849 => x"74616c69",
  2850 => x"7a652020",
  2851 => x"2020203a",
  2852 => x"00000000",
  2853 => x"0a636f6c",
  2854 => x"756d6e20",
  2855 => x"73697a65",
  2856 => x"2020203a",
  2857 => x"00000000",
  2858 => x"0a62616e",
  2859 => x"6b73697a",
  2860 => x"65202020",
  2861 => x"2020203a",
  2862 => x"00000000",
  2863 => x"4d627974",
  2864 => x"65000000",
  2865 => x"0a745f52",
  2866 => x"43442020",
  2867 => x"20202020",
  2868 => x"2020203a",
  2869 => x"00000000",
  2870 => x"0a745f52",
  2871 => x"46432020",
  2872 => x"20202020",
  2873 => x"2020203a",
  2874 => x"00000000",
  2875 => x"0a745f52",
  2876 => x"50202020",
  2877 => x"20202020",
  2878 => x"2020203a",
  2879 => x"00000000",
  2880 => x"0a726566",
  2881 => x"72657368",
  2882 => x"20656e2e",
  2883 => x"2020203a",
  2884 => x"00000000",
  2885 => x"0a0a4444",
  2886 => x"52206672",
  2887 => x"65717565",
  2888 => x"6e637920",
  2889 => x"3a000000",
  2890 => x"0a444452",
  2891 => x"20646174",
  2892 => x"61207769",
  2893 => x"6474683a",
  2894 => x"00000000",
  2895 => x"0a6d6f62",
  2896 => x"696c6520",
  2897 => x"73757070",
  2898 => x"6f72743a",
  2899 => x"00000000",
  2900 => x"0a0a7374",
  2901 => x"61747573",
  2902 => x"20726561",
  2903 => x"64202020",
  2904 => x"3a000000",
  2905 => x"0a0a7365",
  2906 => x"6c662072",
  2907 => x"65667265",
  2908 => x"73682020",
  2909 => x"3a000000",
  2910 => x"34303639",
  2911 => x"00000000",
  2912 => x"756e6b6e",
  2913 => x"6f776e00",
  2914 => x"20617272",
  2915 => x"61790000",
  2916 => x"0a74656d",
  2917 => x"702d636f",
  2918 => x"6d702072",
  2919 => x"6566723a",
  2920 => x"00000000",
  2921 => x"c2b04300",
  2922 => x"0a647269",
  2923 => x"76652073",
  2924 => x"7472656e",
  2925 => x"6774683a",
  2926 => x"00000000",
  2927 => x"0a706f77",
  2928 => x"65722073",
  2929 => x"6176696e",
  2930 => x"6720203a",
  2931 => x"00000000",
  2932 => x"0a745f58",
  2933 => x"50202020",
  2934 => x"20202020",
  2935 => x"2020203a",
  2936 => x"00000000",
  2937 => x"0a745f58",
  2938 => x"53522020",
  2939 => x"20202020",
  2940 => x"2020203a",
  2941 => x"00000000",
  2942 => x"0a745f43",
  2943 => x"4b452020",
  2944 => x"20202020",
  2945 => x"2020203a",
  2946 => x"00000000",
  2947 => x"0a434153",
  2948 => x"206c6174",
  2949 => x"656e6379",
  2950 => x"2020203a",
  2951 => x"00000000",
  2952 => x"0a6d6f62",
  2953 => x"696c6520",
  2954 => x"656e6162",
  2955 => x"6c65643a",
  2956 => x"00000000",
  2957 => x"0a0a7068",
  2958 => x"7920636f",
  2959 => x"6e666967",
  2960 => x"20302020",
  2961 => x"3a000000",
  2962 => x"0a0a7068",
  2963 => x"7920636f",
  2964 => x"6e666967",
  2965 => x"20312020",
  2966 => x"3a000000",
  2967 => x"20353132",
  2968 => x"00000000",
  2969 => x"31303234",
  2970 => x"00000000",
  2971 => x"32303438",
  2972 => x"00000000",
  2973 => x"66756c6c",
  2974 => x"00000000",
  2975 => x"37300000",
  2976 => x"312f3800",
  2977 => x"312f3400",
  2978 => x"312f3200",
  2979 => x"312f3100",
  2980 => x"64656570",
  2981 => x"20706f77",
  2982 => x"65722064",
  2983 => x"6f776e00",
  2984 => x"636c6f63",
  2985 => x"6b207374",
  2986 => x"6f700000",
  2987 => x"73656c66",
  2988 => x"20726566",
  2989 => x"72657368",
  2990 => x"00000000",
  2991 => x"706f7765",
  2992 => x"7220646f",
  2993 => x"776e0000",
  2994 => x"6e6f6e65",
  2995 => x"00000000",
  2996 => x"332f3400",
  2997 => x"38350000",
  2998 => x"34350000",
  2999 => x"68616c66",
  3000 => x"00000000",
  3001 => x"31350000",
  3002 => x"61646472",
  3003 => x"6573733a",
  3004 => x"20000000",
  3005 => x"20646174",
  3006 => x"613a2000",
  3007 => x"0a0a4443",
  3008 => x"4d207068",
  3009 => x"61736520",
  3010 => x"73686966",
  3011 => x"74207465",
  3012 => x"7374696e",
  3013 => x"67000000",
  3014 => x"0a696e69",
  3015 => x"7469616c",
  3016 => x"3a200000",
  3017 => x"09000000",
  3018 => x"20202020",
  3019 => x"00000000",
  3020 => x"6c6f7720",
  3021 => x"666f756e",
  3022 => x"64000000",
  3023 => x"68696768",
  3024 => x"20666f75",
  3025 => x"6e640000",
  3026 => x"0a6c6f77",
  3027 => x"3a202020",
  3028 => x"20202020",
  3029 => x"20200000",
  3030 => x"0a686967",
  3031 => x"683a2020",
  3032 => x"20202020",
  3033 => x"20200000",
  3034 => x"0a646966",
  3035 => x"663a2020",
  3036 => x"20202020",
  3037 => x"20200000",
  3038 => x"0a646966",
  3039 => x"662f323a",
  3040 => x"20202020",
  3041 => x"20200000",
  3042 => x"0a6d696e",
  3043 => x"5f657272",
  3044 => x"3a202020",
  3045 => x"20200000",
  3046 => x"0a6d696e",
  3047 => x"5f657272",
  3048 => x"5f706f73",
  3049 => x"3a200000",
  3050 => x"676f206d",
  3051 => x"696e5f65",
  3052 => x"72726f72",
  3053 => x"00000000",
  3054 => x"0a66696e",
  3055 => x"616c3a20",
  3056 => x"20202020",
  3057 => x"20200000",
  3058 => x"676f207a",
  3059 => x"65726f00",
  3060 => x"68696768",
  3061 => x"204e4f54",
  3062 => x"20666f75",
  3063 => x"6e640000",
  3064 => x"6c6f7720",
  3065 => x"4e4f5420",
  3066 => x"666f756e",
  3067 => x"64000000",
  3068 => x"64617461",
  3069 => x"2076616c",
  3070 => x"69640000",
  3071 => x"6c6f7720",
  3072 => x"20666f75",
  3073 => x"6e640000",
  3074 => x"64617461",
  3075 => x"204e4f54",
  3076 => x"2076616c",
  3077 => x"69640000",
  3078 => x"6c6f7720",
  3079 => x"204e4f54",
  3080 => x"20666f75",
  3081 => x"6e640000",
  3082 => x"74657374",
  3083 => x"2e632000",
  3084 => x"286f6e20",
  3085 => x"73696d75",
  3086 => x"6c61746f",
  3087 => x"72290a00",
  3088 => x"636f6d70",
  3089 => x"696c6564",
  3090 => x"3a204f63",
  3091 => x"74203236",
  3092 => x"20323031",
  3093 => x"30202031",
  3094 => x"343a3430",
  3095 => x"3a35340a",
  3096 => x"00000000",
  3097 => x"286f6e20",
  3098 => x"68617264",
  3099 => x"77617265",
  3100 => x"290a0000",
  3101 => x"0000078a",
  3102 => x"000007b0",
  3103 => x"000007b0",
  3104 => x"0000078a",
  3105 => x"000007b0",
  3106 => x"000007b0",
  3107 => x"000007b0",
  3108 => x"000007b0",
  3109 => x"000007b0",
  3110 => x"000007b0",
  3111 => x"000007b0",
  3112 => x"000007b0",
  3113 => x"000007b0",
  3114 => x"000007b0",
  3115 => x"000007b0",
  3116 => x"000007b0",
  3117 => x"000007b0",
  3118 => x"000007b0",
  3119 => x"000007b0",
  3120 => x"000007b0",
  3121 => x"000007b0",
  3122 => x"000007b0",
  3123 => x"000007b0",
  3124 => x"000007b0",
  3125 => x"000007b0",
  3126 => x"000007b0",
  3127 => x"000007b0",
  3128 => x"000007b0",
  3129 => x"000007b0",
  3130 => x"000007b0",
  3131 => x"000007b0",
  3132 => x"000007b0",
  3133 => x"000007b0",
  3134 => x"000007b0",
  3135 => x"000007b0",
  3136 => x"000007b0",
  3137 => x"000007b0",
  3138 => x"000007b0",
  3139 => x"0000085c",
  3140 => x"00000854",
  3141 => x"0000084c",
  3142 => x"00000844",
  3143 => x"0000083c",
  3144 => x"00000834",
  3145 => x"0000082c",
  3146 => x"00000823",
  3147 => x"0000081a",
  3148 => x"00001f8e",
  3149 => x"00001f87",
  3150 => x"00001f80",
  3151 => x"000019e3",
  3152 => x"000019e3",
  3153 => x"00001f79",
  3154 => x"00001f79",
  3155 => x"000021c5",
  3156 => x"00002139",
  3157 => x"000020ad",
  3158 => x"00001a5f",
  3159 => x"00002021",
  3160 => x"00001f95",
  3161 => x"64756d6d",
  3162 => x"792e6578",
  3163 => x"65000000",
  3164 => x"43000000",
  3165 => x"00ffffff",
  3166 => x"ff00ffff",
  3167 => x"ffff00ff",
  3168 => x"ffffff00",
  3169 => x"00000000",
  3170 => x"00000000",
  3171 => x"00000000",
  3172 => x"0000353c",
  3173 => x"fff00000",
  3174 => x"80000e00",
  3175 => x"80000800",
  3176 => x"80000600",
  3177 => x"80000200",
  3178 => x"80000100",
  3179 => x"00003164",
  3180 => x"000031b4",
  3181 => x"00000000",
  3182 => x"0000341c",
  3183 => x"00003478",
  3184 => x"000034d4",
  3185 => x"00000000",
  3186 => x"00000000",
  3187 => x"00000000",
  3188 => x"00000000",
  3189 => x"00000000",
  3190 => x"00000000",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00003170",
  3195 => x"00000000",
  3196 => x"00000000",
  3197 => x"00000000",
  3198 => x"00000000",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000001",
  3224 => x"330eabcd",
  3225 => x"1234e66d",
  3226 => x"deec0005",
  3227 => x"000b0000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000000",
  3246 => x"00000000",
  3247 => x"00000000",
  3248 => x"00000000",
  3249 => x"00000000",
  3250 => x"00000000",
  3251 => x"00000000",
  3252 => x"00000000",
  3253 => x"00000000",
  3254 => x"00000000",
  3255 => x"00000000",
  3256 => x"00000000",
  3257 => x"00000000",
  3258 => x"00000000",
  3259 => x"00000000",
  3260 => x"00000000",
  3261 => x"00000000",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00000000",
  3265 => x"00000000",
  3266 => x"00000000",
  3267 => x"00000000",
  3268 => x"00000000",
  3269 => x"00000000",
  3270 => x"00000000",
  3271 => x"00000000",
  3272 => x"00000000",
  3273 => x"00000000",
  3274 => x"00000000",
  3275 => x"00000000",
  3276 => x"00000000",
  3277 => x"00000000",
  3278 => x"00000000",
  3279 => x"00000000",
  3280 => x"00000000",
  3281 => x"00000000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"00000000",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00000000",
  3288 => x"00000000",
  3289 => x"00000000",
  3290 => x"00000000",
  3291 => x"00000000",
  3292 => x"00000000",
  3293 => x"00000000",
  3294 => x"00000000",
  3295 => x"00000000",
  3296 => x"00000000",
  3297 => x"00000000",
  3298 => x"00000000",
  3299 => x"00000000",
  3300 => x"00000000",
  3301 => x"00000000",
  3302 => x"00000000",
  3303 => x"00000000",
  3304 => x"00000000",
  3305 => x"00000000",
  3306 => x"00000000",
  3307 => x"00000000",
  3308 => x"00000000",
  3309 => x"00000000",
  3310 => x"00000000",
  3311 => x"00000000",
  3312 => x"00000000",
  3313 => x"00000000",
  3314 => x"00000000",
  3315 => x"00000000",
  3316 => x"00000000",
  3317 => x"00000000",
  3318 => x"00000000",
  3319 => x"00000000",
  3320 => x"00000000",
  3321 => x"00000000",
  3322 => x"00000000",
  3323 => x"00000000",
  3324 => x"00000000",
  3325 => x"00000000",
  3326 => x"00000000",
  3327 => x"00000000",
  3328 => x"00000000",
  3329 => x"00000000",
  3330 => x"00000000",
  3331 => x"00000000",
  3332 => x"00000000",
  3333 => x"00000000",
  3334 => x"00000000",
  3335 => x"00000000",
  3336 => x"00000000",
  3337 => x"00000000",
  3338 => x"00000000",
  3339 => x"00000000",
  3340 => x"00000000",
  3341 => x"00000000",
  3342 => x"00000000",
  3343 => x"00000000",
  3344 => x"00000000",
  3345 => x"00000000",
  3346 => x"00000000",
  3347 => x"00000000",
  3348 => x"00000000",
  3349 => x"00000000",
  3350 => x"00000000",
  3351 => x"00000000",
  3352 => x"00000000",
  3353 => x"00000000",
  3354 => x"00000000",
  3355 => x"00000000",
  3356 => x"00000000",
  3357 => x"00000000",
  3358 => x"00000000",
  3359 => x"00000000",
  3360 => x"00000000",
  3361 => x"00000000",
  3362 => x"00000000",
  3363 => x"00000000",
  3364 => x"00000000",
  3365 => x"00000000",
  3366 => x"00000000",
  3367 => x"00000000",
  3368 => x"00000000",
  3369 => x"00000000",
  3370 => x"00000000",
  3371 => x"00000000",
  3372 => x"00000000",
  3373 => x"00000000",
  3374 => x"00000000",
  3375 => x"00000000",
  3376 => x"00000000",
  3377 => x"00000000",
  3378 => x"00000000",
  3379 => x"00000000",
  3380 => x"00000000",
  3381 => x"00000000",
  3382 => x"00000000",
  3383 => x"00000000",
  3384 => x"00000000",
  3385 => x"00000000",
  3386 => x"00000000",
  3387 => x"00000000",
  3388 => x"00000000",
  3389 => x"00000000",
  3390 => x"00000000",
  3391 => x"00000000",
  3392 => x"00000000",
  3393 => x"00000000",
  3394 => x"00000000",
  3395 => x"00000000",
  3396 => x"00000000",
  3397 => x"00000000",
  3398 => x"00000000",
  3399 => x"00000000",
  3400 => x"00000000",
  3401 => x"00000000",
  3402 => x"00000000",
  3403 => x"00000000",
  3404 => x"ffffffff",
  3405 => x"00000000",
  3406 => x"ffffffff",
  3407 => x"00000000",
  3408 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
