-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b80db",
     1 => x"cb040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b80de",
     9 => x"b2040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b80dd",
    73 => x"e4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b80ddc7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b81ab",
   162 => x"f4738306",
   163 => x"10100508",
   164 => x"060b0b80",
   165 => x"ddca0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b80de",
   169 => x"99040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b80de",
   177 => x"80040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"81ac840c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053370",
   258 => x"525280db",
   259 => x"bb3f7151",
   260 => x"80dca93f",
   261 => x"71b00c83",
   262 => x"3d0d04fd",
   263 => x"3d0d8a51",
   264 => x"80d6b63f",
   265 => x"a6e53f96",
   266 => x"d353818d",
   267 => x"e852818d",
   268 => x"fc51a6ea",
   269 => x"3fa3c353",
   270 => x"818e8052",
   271 => x"818ea451",
   272 => x"a6dc3fa6",
   273 => x"d553818e",
   274 => x"ac52818e",
   275 => x"bc51a6ce",
   276 => x"3f9fe053",
   277 => x"818ec452",
   278 => x"818fbc51",
   279 => x"a6c03fa1",
   280 => x"c353818e",
   281 => x"e052818f",
   282 => x"8051a6b2",
   283 => x"3fa2a453",
   284 => x"818f8852",
   285 => x"818fa851",
   286 => x"a6a43f9f",
   287 => x"ac53818f",
   288 => x"b052818f",
   289 => x"c451a696",
   290 => x"3fa4db53",
   291 => x"818fcc52",
   292 => x"818fe851",
   293 => x"a6883fa6",
   294 => x"ec53818f",
   295 => x"f0528190",
   296 => x"9451a5fa",
   297 => x"3fa7ad53",
   298 => x"81909c52",
   299 => x"8190c451",
   300 => x"a5ec3fa8",
   301 => x"d5538190",
   302 => x"cc528190",
   303 => x"ec51a5de",
   304 => x"3fa6bc53",
   305 => x"8190f052",
   306 => x"81918c51",
   307 => x"a5d03fa9",
   308 => x"b0538191",
   309 => x"94528191",
   310 => x"a451a5c2",
   311 => x"3fabde53",
   312 => x"8191a852",
   313 => x"8191c451",
   314 => x"a5b43fa6",
   315 => x"82538191",
   316 => x"cc528191",
   317 => x"e451a5a6",
   318 => x"3fabe653",
   319 => x"8191ec52",
   320 => x"81928051",
   321 => x"a5983f8d",
   322 => x"cc538192",
   323 => x"88528192",
   324 => x"9c51a58a",
   325 => x"3f90d653",
   326 => x"8192a052",
   327 => x"8192c851",
   328 => x"a4fc3fa6",
   329 => x"9e538192",
   330 => x"d0528192",
   331 => x"f051a4ee",
   332 => x"3f95fa53",
   333 => x"8192f852",
   334 => x"81938c51",
   335 => x"a4e03f8b",
   336 => x"d0538193",
   337 => x"94528193",
   338 => x"a051a4d2",
   339 => x"3f8cf553",
   340 => x"8193a452",
   341 => x"8193cc51",
   342 => x"a4c43f8b",
   343 => x"d0538193",
   344 => x"d452819a",
   345 => x"f851a4b6",
   346 => x"3f8dbb53",
   347 => x"8193e452",
   348 => x"8193f451",
   349 => x"a4a83f8b",
   350 => x"c5538194",
   351 => x"8852818d",
   352 => x"d851a49a",
   353 => x"3fb5f453",
   354 => x"81948852",
   355 => x"818de051",
   356 => x"a48c3faa",
   357 => x"df3fa4d2",
   358 => x"3f810b81",
   359 => x"cf943480",
   360 => x"d7ce3fb0",
   361 => x"089038a4",
   362 => x"cf3f81cf",
   363 => x"94335473",
   364 => x"ee38853d",
   365 => x"0d0480d7",
   366 => x"ca3fb008",
   367 => x"81ff0651",
   368 => x"a5a43fdb",
   369 => x"39800b81",
   370 => x"cf943480",
   371 => x"0bb00c04",
   372 => x"fb3d0d81",
   373 => x"51a8eb3f",
   374 => x"b0085382",
   375 => x"51a8e33f",
   376 => x"b00856b0",
   377 => x"08833890",
   378 => x"5672fc06",
   379 => x"5475812e",
   380 => x"80fb3880",
   381 => x"55747627",
   382 => x"ad387483",
   383 => x"06537280",
   384 => x"2eb23881",
   385 => x"9ff45180",
   386 => x"d2e93f73",
   387 => x"70840555",
   388 => x"0852a051",
   389 => x"80d2ff3f",
   390 => x"a05180d2",
   391 => x"bc3f8115",
   392 => x"55757526",
   393 => x"d5388a51",
   394 => x"80d2ae3f",
   395 => x"800bb00c",
   396 => x"873d0d04",
   397 => x"8193fc51",
   398 => x"80d2b83f",
   399 => x"7352a051",
   400 => x"80d2d33f",
   401 => x"819ae451",
   402 => x"80d2a83f",
   403 => x"819ff451",
   404 => x"80d2a03f",
   405 => x"73708405",
   406 => x"550852a0",
   407 => x"5180d2b6",
   408 => x"3fa05180",
   409 => x"d1f33f81",
   410 => x"1555ffb5",
   411 => x"397308b0",
   412 => x"0c873d0d",
   413 => x"04fc3d0d",
   414 => x"8151a7c6",
   415 => x"3fb00852",
   416 => x"8251a68c",
   417 => x"3fb00881",
   418 => x"ff067256",
   419 => x"53835472",
   420 => x"802ea138",
   421 => x"7351a7aa",
   422 => x"3f811470",
   423 => x"81ff06ff",
   424 => x"157081ff",
   425 => x"06b00879",
   426 => x"7084055b",
   427 => x"0c565255",
   428 => x"5272e138",
   429 => x"72b00c86",
   430 => x"3d0d0480",
   431 => x"3d0d8c51",
   432 => x"80d1963f",
   433 => x"800bb00c",
   434 => x"823d0d04",
   435 => x"fb3d0d80",
   436 => x"0b819480",
   437 => x"525680d1",
   438 => x"9a3f7555",
   439 => x"741081fe",
   440 => x"065381d0",
   441 => x"5281ac8c",
   442 => x"0851b7b9",
   443 => x"3fb00898",
   444 => x"2b548074",
   445 => x"24a23881",
   446 => x"948c5180",
   447 => x"d0f53f74",
   448 => x"52885180",
   449 => x"d1903f81",
   450 => x"94985180",
   451 => x"d0e53f81",
   452 => x"167083ff",
   453 => x"ff065754",
   454 => x"81157081",
   455 => x"ff067098",
   456 => x"2b525654",
   457 => x"738025ff",
   458 => x"b33875b0",
   459 => x"0c873d0d",
   460 => x"04f33d0d",
   461 => x"7f028405",
   462 => x"80c30533",
   463 => x"02880580",
   464 => x"c6052281",
   465 => x"94a8545b",
   466 => x"555880d0",
   467 => x"a63f7851",
   468 => x"80d1ea3f",
   469 => x"8194b451",
   470 => x"80d0983f",
   471 => x"73528851",
   472 => x"80d0b33f",
   473 => x"8194d051",
   474 => x"80d0883f",
   475 => x"80577679",
   476 => x"27819c38",
   477 => x"73108e3d",
   478 => x"5d5a7981",
   479 => x"ff065381",
   480 => x"90527751",
   481 => x"b69f3f76",
   482 => x"882a5390",
   483 => x"527751b6",
   484 => x"943f7681",
   485 => x"ff065390",
   486 => x"527751b6",
   487 => x"883f811a",
   488 => x"7081ff06",
   489 => x"54558190",
   490 => x"527751b5",
   491 => x"f83f8053",
   492 => x"80e05277",
   493 => x"51b5ee3f",
   494 => x"b008982b",
   495 => x"54807424",
   496 => x"8a388818",
   497 => x"087081ff",
   498 => x"065c567a",
   499 => x"81ff0681",
   500 => x"9ff45256",
   501 => x"80cf9c3f",
   502 => x"75528851",
   503 => x"80cfb73f",
   504 => x"8197f051",
   505 => x"80cf8c3f",
   506 => x"e0165480",
   507 => x"df7427b6",
   508 => x"38768706",
   509 => x"701d5755",
   510 => x"a0763474",
   511 => x"872eb938",
   512 => x"81177083",
   513 => x"ffff0658",
   514 => x"55787726",
   515 => x"feec3880",
   516 => x"e00b8c19",
   517 => x"0c8c1808",
   518 => x"70812a81",
   519 => x"06585a76",
   520 => x"f4388f3d",
   521 => x"0d047687",
   522 => x"06701d55",
   523 => x"55757434",
   524 => x"74872e09",
   525 => x"8106c938",
   526 => x"7b5180ce",
   527 => x"b63f8a51",
   528 => x"80ce963f",
   529 => x"81177083",
   530 => x"ffff0658",
   531 => x"55787726",
   532 => x"fea838ff",
   533 => x"ba39fb3d",
   534 => x"0d8151a2",
   535 => x"b33fb008",
   536 => x"81ff0654",
   537 => x"8251a3da",
   538 => x"3fb00881",
   539 => x"ff065683",
   540 => x"51a29d3f",
   541 => x"b00883ff",
   542 => x"ff065573",
   543 => x"9c3881ac",
   544 => x"8c085474",
   545 => x"84388180",
   546 => x"55745375",
   547 => x"527351fd",
   548 => x"a03f74b0",
   549 => x"0c873d0d",
   550 => x"0481ac90",
   551 => x"0854e439",
   552 => x"f83d0d02",
   553 => x"aa052281",
   554 => x"abe83381",
   555 => x"f7065858",
   556 => x"7681abe8",
   557 => x"3481ac8c",
   558 => x"085580c0",
   559 => x"53819052",
   560 => x"7451b3e1",
   561 => x"3f7451b4",
   562 => x"8e3fb008",
   563 => x"81ff0654",
   564 => x"73802e83",
   565 => x"fc387653",
   566 => x"80d05274",
   567 => x"51b3c63f",
   568 => x"80598f57",
   569 => x"81abe833",
   570 => x"81fe0654",
   571 => x"7381abe8",
   572 => x"3481ac8c",
   573 => x"08745755",
   574 => x"80c05381",
   575 => x"90527451",
   576 => x"b3a33f74",
   577 => x"51b3d03f",
   578 => x"b00881ff",
   579 => x"06547380",
   580 => x"2e83b338",
   581 => x"755380d0",
   582 => x"527451b3",
   583 => x"883f7777",
   584 => x"2c810655",
   585 => x"74802e83",
   586 => x"923881ab",
   587 => x"e8338207",
   588 => x"547381ab",
   589 => x"e83481ac",
   590 => x"8c087457",
   591 => x"5580c053",
   592 => x"81905274",
   593 => x"51b2de3f",
   594 => x"7451b38b",
   595 => x"3fb00881",
   596 => x"ff065473",
   597 => x"802e82d8",
   598 => x"38755380",
   599 => x"d0527451",
   600 => x"b2c33f81",
   601 => x"ac8c0855",
   602 => x"80c15381",
   603 => x"90527451",
   604 => x"b2b33f74",
   605 => x"51b2e03f",
   606 => x"b00881ff",
   607 => x"06567580",
   608 => x"2e828138",
   609 => x"805380e0",
   610 => x"527451b2",
   611 => x"983f7451",
   612 => x"b2c53fb0",
   613 => x"0881ff06",
   614 => x"5473802e",
   615 => x"81e63888",
   616 => x"15087090",
   617 => x"2b70902c",
   618 => x"56565673",
   619 => x"822a8106",
   620 => x"5473802e",
   621 => x"8d388177",
   622 => x"2b790770",
   623 => x"83ffff06",
   624 => x"5a5681ab",
   625 => x"e8338107",
   626 => x"547381ab",
   627 => x"e83481ac",
   628 => x"8c087457",
   629 => x"5580c053",
   630 => x"81905274",
   631 => x"51b1c63f",
   632 => x"7451b1f3",
   633 => x"3fb00881",
   634 => x"ff065473",
   635 => x"802e81a1",
   636 => x"38755380",
   637 => x"d0527451",
   638 => x"b1ab3f76",
   639 => x"81800a29",
   640 => x"81ff0a05",
   641 => x"70982c58",
   642 => x"56768025",
   643 => x"fdd63881",
   644 => x"abe83382",
   645 => x"07577681",
   646 => x"abe83481",
   647 => x"ac8c0855",
   648 => x"80c05381",
   649 => x"90527451",
   650 => x"b0fb3f74",
   651 => x"51b1a83f",
   652 => x"b00881ff",
   653 => x"06587780",
   654 => x"2e81b438",
   655 => x"765380d0",
   656 => x"527451b0",
   657 => x"e03f81ab",
   658 => x"e8338807",
   659 => x"577681ab",
   660 => x"e83481ac",
   661 => x"8c085580",
   662 => x"c0538190",
   663 => x"527451b0",
   664 => x"c43f7451",
   665 => x"b0f13fb0",
   666 => x"0881ff06",
   667 => x"5877802e",
   668 => x"80ee3876",
   669 => x"5380d052",
   670 => x"7451b0a9",
   671 => x"3f78b00c",
   672 => x"8a3d0d04",
   673 => x"8194d451",
   674 => x"80c9e83f",
   675 => x"ff54fe9b",
   676 => x"398194d4",
   677 => x"5180c9db",
   678 => x"3f768180",
   679 => x"0a2981ff",
   680 => x"0a057098",
   681 => x"2c585676",
   682 => x"8025fcb8",
   683 => x"38fee039",
   684 => x"8194d451",
   685 => x"80c9bc3f",
   686 => x"fda93981",
   687 => x"abe83381",
   688 => x"fd0654fc",
   689 => x"ec398194",
   690 => x"d45180c9",
   691 => x"a63ffcce",
   692 => x"398194d4",
   693 => x"5180c99b",
   694 => x"3f80598f",
   695 => x"57fc8539",
   696 => x"8194d451",
   697 => x"80c98c3f",
   698 => x"78b00c8a",
   699 => x"3d0d0481",
   700 => x"94d45180",
   701 => x"c8fd3ffe",
   702 => x"cd39803d",
   703 => x"0d828180",
   704 => x"51fb9d3f",
   705 => x"82828051",
   706 => x"fb963f82",
   707 => x"848151fb",
   708 => x"8f3f8286",
   709 => x"f151fb88",
   710 => x"3f8288b8",
   711 => x"51fb813f",
   712 => x"800bb00c",
   713 => x"823d0d04",
   714 => x"fe3d0d02",
   715 => x"93053302",
   716 => x"84059705",
   717 => x"33545271",
   718 => x"73279438",
   719 => x"a05180c8",
   720 => x"983f8112",
   721 => x"7081ff06",
   722 => x"51527272",
   723 => x"26ee3884",
   724 => x"3d0d04fd",
   725 => x"3d0d8195",
   726 => x"8c5180c8",
   727 => x"963f8195",
   728 => x"ac5180c8",
   729 => x"8e3f8195",
   730 => x"f45180c8",
   731 => x"863f8196",
   732 => x"bc5180c7",
   733 => x"fe3f81ab",
   734 => x"e4087008",
   735 => x"525380c9",
   736 => x"bc3fb008",
   737 => x"81ff0653",
   738 => x"728c2794",
   739 => x"38a05180",
   740 => x"c7c73f81",
   741 => x"137081ff",
   742 => x"0654548c",
   743 => x"7326ee38",
   744 => x"81abe408",
   745 => x"84110852",
   746 => x"5380c991",
   747 => x"3fb00881",
   748 => x"ff065372",
   749 => x"8c279438",
   750 => x"a05180c7",
   751 => x"9c3f8113",
   752 => x"7081ff06",
   753 => x"54548c73",
   754 => x"26ee3881",
   755 => x"abe40888",
   756 => x"11085253",
   757 => x"80c8e63f",
   758 => x"b00881ff",
   759 => x"0653728c",
   760 => x"279438a0",
   761 => x"5180c6f1",
   762 => x"3f811370",
   763 => x"81ff0654",
   764 => x"548c7326",
   765 => x"ee3881ab",
   766 => x"e4088c11",
   767 => x"08525380",
   768 => x"c8bb3fb0",
   769 => x"0881ff06",
   770 => x"53728c27",
   771 => x"9438a051",
   772 => x"80c6c63f",
   773 => x"81137081",
   774 => x"ff065454",
   775 => x"8c7326ee",
   776 => x"388196d8",
   777 => x"5180c6cb",
   778 => x"3f81abe4",
   779 => x"08901108",
   780 => x"525380c8",
   781 => x"883fb008",
   782 => x"81ff0653",
   783 => x"728c2794",
   784 => x"38a05180",
   785 => x"c6933f81",
   786 => x"137081ff",
   787 => x"0654548c",
   788 => x"7326ee38",
   789 => x"81abe408",
   790 => x"94110852",
   791 => x"5380c7dd",
   792 => x"3fb00881",
   793 => x"ff065372",
   794 => x"8c279438",
   795 => x"a05180c5",
   796 => x"e83f8113",
   797 => x"7081ff06",
   798 => x"54548c73",
   799 => x"26ee3881",
   800 => x"abe40898",
   801 => x"11085253",
   802 => x"80c7b23f",
   803 => x"b00881ff",
   804 => x"0653728c",
   805 => x"279438a0",
   806 => x"5180c5bd",
   807 => x"3f811370",
   808 => x"81ff0654",
   809 => x"548c7326",
   810 => x"ee3881ab",
   811 => x"e4089c11",
   812 => x"08525380",
   813 => x"c7873fb0",
   814 => x"0881ff06",
   815 => x"53728c27",
   816 => x"9438a051",
   817 => x"80c5923f",
   818 => x"81137081",
   819 => x"ff065454",
   820 => x"8c7326ee",
   821 => x"388196f4",
   822 => x"5180c597",
   823 => x"3f81abe4",
   824 => x"0854810b",
   825 => x"b0150cb0",
   826 => x"14085372",
   827 => x"8025f838",
   828 => x"a0140851",
   829 => x"80c6c63f",
   830 => x"b00881ff",
   831 => x"0653728c",
   832 => x"279438a0",
   833 => x"5180c4d1",
   834 => x"3f811370",
   835 => x"81ff0654",
   836 => x"548c7326",
   837 => x"ee3881ab",
   838 => x"e408a411",
   839 => x"08525380",
   840 => x"c69b3fb0",
   841 => x"0881ff06",
   842 => x"53728c27",
   843 => x"9438a051",
   844 => x"80c4a63f",
   845 => x"81137081",
   846 => x"ff065454",
   847 => x"8c7326ee",
   848 => x"3881abe4",
   849 => x"08a81108",
   850 => x"525380c5",
   851 => x"f03fb008",
   852 => x"81ff0653",
   853 => x"728c2794",
   854 => x"38a05180",
   855 => x"c3fb3f81",
   856 => x"137081ff",
   857 => x"0654548c",
   858 => x"7326ee38",
   859 => x"81abe408",
   860 => x"ac110852",
   861 => x"5380c5c5",
   862 => x"3fb00881",
   863 => x"ff065372",
   864 => x"8c279438",
   865 => x"a05180c3",
   866 => x"d03f8113",
   867 => x"7081ff06",
   868 => x"54548c73",
   869 => x"26ee3881",
   870 => x"97905180",
   871 => x"c3d53f81",
   872 => x"abe408b0",
   873 => x"1108fe0a",
   874 => x"06525480",
   875 => x"c58f3f81",
   876 => x"abe40854",
   877 => x"800bb015",
   878 => x"0c8197a4",
   879 => x"5180c3b3",
   880 => x"3f8197bc",
   881 => x"5180c3ab",
   882 => x"3f81abe4",
   883 => x"0880c011",
   884 => x"08525380",
   885 => x"c4e73fb0",
   886 => x"0881ff06",
   887 => x"53729827",
   888 => x"9438a051",
   889 => x"80c2f23f",
   890 => x"81137081",
   891 => x"ff065153",
   892 => x"987326ee",
   893 => x"3881abe4",
   894 => x"0880c811",
   895 => x"08525480",
   896 => x"c4bb3fb0",
   897 => x"0881ff06",
   898 => x"53729827",
   899 => x"9438a051",
   900 => x"80c2c63f",
   901 => x"81137081",
   902 => x"ff065153",
   903 => x"987326ee",
   904 => x"388197d8",
   905 => x"5180c2cb",
   906 => x"3f81abe4",
   907 => x"0880c411",
   908 => x"08525480",
   909 => x"c4873fb0",
   910 => x"0881ff06",
   911 => x"53729827",
   912 => x"9438a051",
   913 => x"80c2923f",
   914 => x"81137081",
   915 => x"ff065153",
   916 => x"987326ee",
   917 => x"3881abe4",
   918 => x"0880cc11",
   919 => x"08525480",
   920 => x"c3db3fb0",
   921 => x"0881ff06",
   922 => x"53729827",
   923 => x"9438a051",
   924 => x"80c1e63f",
   925 => x"81137081",
   926 => x"ff065153",
   927 => x"987326ee",
   928 => x"388a5180",
   929 => x"c1d33f81",
   930 => x"abe408b4",
   931 => x"11087081",
   932 => x"ff068197",
   933 => x"f4545255",
   934 => x"5380c1d7",
   935 => x"3f725180",
   936 => x"c39b3fa0",
   937 => x"5180c1b1",
   938 => x"3f728626",
   939 => x"94387210",
   940 => x"10819cb4",
   941 => x"05547308",
   942 => x"04819888",
   943 => x"5180c1b3",
   944 => x"3f81abe4",
   945 => x"08b81108",
   946 => x"7081ff06",
   947 => x"81989454",
   948 => x"52545480",
   949 => x"c19d3f73",
   950 => x"52885180",
   951 => x"c1b83f73",
   952 => x"81065372",
   953 => x"80f23873",
   954 => x"812a7081",
   955 => x"06515372",
   956 => x"80ce3873",
   957 => x"822a7081",
   958 => x"06515372",
   959 => x"ae387383",
   960 => x"2a810654",
   961 => x"738f388a",
   962 => x"5180c0cd",
   963 => x"3f800bb0",
   964 => x"0c853d0d",
   965 => x"048198a8",
   966 => x"5180c0d7",
   967 => x"3f8a5180",
   968 => x"c0b73f80",
   969 => x"0bb00c85",
   970 => x"3d0d0481",
   971 => x"98bc5180",
   972 => x"c0c13f73",
   973 => x"832a8106",
   974 => x"5473802e",
   975 => x"ca38d639",
   976 => x"8198dc51",
   977 => x"80c0ac3f",
   978 => x"73822a70",
   979 => x"81065153",
   980 => x"72802eff",
   981 => x"a938d439",
   982 => x"8198f451",
   983 => x"80c0943f",
   984 => x"73812a70",
   985 => x"81065153",
   986 => x"72802eff",
   987 => x"8638d139",
   988 => x"81998851",
   989 => x"bffd3ffe",
   990 => x"c8398199",
   991 => x"9451bff3",
   992 => x"3ffebe39",
   993 => x"8199a051",
   994 => x"bfe93ffe",
   995 => x"b4398199",
   996 => x"a451bfdf",
   997 => x"3ffeaa39",
   998 => x"8199b051",
   999 => x"bfd53ffe",
  1000 => x"a0398199",
  1001 => x"bc51bfcb",
  1002 => x"3ffe9639",
  1003 => x"fe3d0d88",
  1004 => x"0a53840a",
  1005 => x"0b81abe0",
  1006 => x"088c1108",
  1007 => x"51525280",
  1008 => x"71279538",
  1009 => x"80737084",
  1010 => x"05550c80",
  1011 => x"72708405",
  1012 => x"540cff11",
  1013 => x"5170ed38",
  1014 => x"800bb00c",
  1015 => x"843d0d04",
  1016 => x"fa3d0d88",
  1017 => x"0a57840a",
  1018 => x"56815193",
  1019 => x"a33fb008",
  1020 => x"83ffff06",
  1021 => x"54738338",
  1022 => x"90548055",
  1023 => x"74742781",
  1024 => x"bb387508",
  1025 => x"70902c52",
  1026 => x"5380c0b1",
  1027 => x"3fb00881",
  1028 => x"ff065271",
  1029 => x"8a279338",
  1030 => x"a051bebd",
  1031 => x"3f811270",
  1032 => x"81ff0651",
  1033 => x"528a7226",
  1034 => x"ef387290",
  1035 => x"2b70902c",
  1036 => x"525280c0",
  1037 => x"883fb008",
  1038 => x"81ff0652",
  1039 => x"718a2793",
  1040 => x"38a051be",
  1041 => x"943f8112",
  1042 => x"7081ff06",
  1043 => x"53538a72",
  1044 => x"26ef3876",
  1045 => x"0870902c",
  1046 => x"5253bfe1",
  1047 => x"3fb00881",
  1048 => x"ff065271",
  1049 => x"8a279338",
  1050 => x"a051bded",
  1051 => x"3f811270",
  1052 => x"81ff0651",
  1053 => x"528a7226",
  1054 => x"ef387290",
  1055 => x"2b70902c",
  1056 => x"5252bfb9",
  1057 => x"3fb00881",
  1058 => x"ff065271",
  1059 => x"8a279338",
  1060 => x"a051bdc5",
  1061 => x"3f811270",
  1062 => x"81ff0653",
  1063 => x"538a7226",
  1064 => x"ef388a51",
  1065 => x"bdb33f84",
  1066 => x"17841781",
  1067 => x"177083ff",
  1068 => x"ff065854",
  1069 => x"57577375",
  1070 => x"26fec738",
  1071 => x"73b00c88",
  1072 => x"3d0d04fd",
  1073 => x"3d0d81ab",
  1074 => x"e0088c11",
  1075 => x"0870822b",
  1076 => x"83fffc06",
  1077 => x"8199c854",
  1078 => x"515454bd",
  1079 => x"963f7252",
  1080 => x"880a5195",
  1081 => x"af3fb008",
  1082 => x"54b008fe",
  1083 => x"2ea838b0",
  1084 => x"08ff2e94",
  1085 => x"387251be",
  1086 => x"c43f8199",
  1087 => x"dc51bcf3",
  1088 => x"3f73b00c",
  1089 => x"853d0d04",
  1090 => x"8199f051",
  1091 => x"bce53f73",
  1092 => x"b00c853d",
  1093 => x"0d048199",
  1094 => x"f851bcd7",
  1095 => x"3f73b00c",
  1096 => x"853d0d04",
  1097 => x"fc3d0d81",
  1098 => x"abe0088c",
  1099 => x"11087082",
  1100 => x"2b83fffc",
  1101 => x"06819a84",
  1102 => x"54515555",
  1103 => x"bcb53f81",
  1104 => x"aca00888",
  1105 => x"11087080",
  1106 => x"c0078813",
  1107 => x"0c545573",
  1108 => x"52880a51",
  1109 => x"97c03fb0",
  1110 => x"0881aca0",
  1111 => x"08881108",
  1112 => x"70ffbf06",
  1113 => x"88130c55",
  1114 => x"5555b008",
  1115 => x"fe2e80c5",
  1116 => x"38b008fe",
  1117 => x"249a38b0",
  1118 => x"08fd2eab",
  1119 => x"387451bd",
  1120 => x"bc3f819a",
  1121 => x"9851bbeb",
  1122 => x"3f74b00c",
  1123 => x"863d0d04",
  1124 => x"b008ff2e",
  1125 => x"098106e5",
  1126 => x"388199f0",
  1127 => x"51bbd43f",
  1128 => x"74b00c86",
  1129 => x"3d0d0481",
  1130 => x"9aac51bb",
  1131 => x"c63f74b0",
  1132 => x"0c863d0d",
  1133 => x"04819abc",
  1134 => x"51bbb83f",
  1135 => x"74b00c86",
  1136 => x"3d0d04fd",
  1137 => x"3d0d8151",
  1138 => x"8fc63fb0",
  1139 => x"0881ff06",
  1140 => x"5473802e",
  1141 => x"a4387384",
  1142 => x"26903881",
  1143 => x"abe00874",
  1144 => x"710c5373",
  1145 => x"b00c853d",
  1146 => x"0d0481ab",
  1147 => x"e0085380",
  1148 => x"730c73b0",
  1149 => x"0c853d0d",
  1150 => x"04819ac8",
  1151 => x"51baf43f",
  1152 => x"819ad851",
  1153 => x"baed3f81",
  1154 => x"abe00870",
  1155 => x"085253bc",
  1156 => x"ac3f819a",
  1157 => x"e851badb",
  1158 => x"3f81abe0",
  1159 => x"08841108",
  1160 => x"5353a051",
  1161 => x"baf03f81",
  1162 => x"9afc51ba",
  1163 => x"c63f81ab",
  1164 => x"e0088811",
  1165 => x"085353a0",
  1166 => x"51badb3f",
  1167 => x"819b9051",
  1168 => x"bab13f81",
  1169 => x"abe0088c",
  1170 => x"11085253",
  1171 => x"bbef3f8a",
  1172 => x"51ba863f",
  1173 => x"73b00c85",
  1174 => x"3d0d04f6",
  1175 => x"3d0d880a",
  1176 => x"5681518e",
  1177 => x"ab3fb008",
  1178 => x"8b3d2382",
  1179 => x"518ea13f",
  1180 => x"b0080284",
  1181 => x"05a60523",
  1182 => x"83518e94",
  1183 => x"3fb0088c",
  1184 => x"3d238451",
  1185 => x"8e8a3fb0",
  1186 => x"08893d23",
  1187 => x"85518e80",
  1188 => x"3fb00802",
  1189 => x"84059e05",
  1190 => x"2386518d",
  1191 => x"f33fb008",
  1192 => x"8a3d2380",
  1193 => x"0b81abe0",
  1194 => x"088c1108",
  1195 => x"51535574",
  1196 => x"7227b838",
  1197 => x"71548c3d",
  1198 => x"751005f8",
  1199 => x"11227090",
  1200 => x"2bf01322",
  1201 => x"70848080",
  1202 => x"2972902c",
  1203 => x"057a0c52",
  1204 => x"55588116",
  1205 => x"7081ff06",
  1206 => x"52545274",
  1207 => x"822e9438",
  1208 => x"718417ff",
  1209 => x"16565755",
  1210 => x"73cc3880",
  1211 => x"0bb00c8c",
  1212 => x"3d0d0480",
  1213 => x"0b8417ff",
  1214 => x"16565755",
  1215 => x"73ffb738",
  1216 => x"ea39fe3d",
  1217 => x"0d81518d",
  1218 => x"873fb008",
  1219 => x"81ff0681",
  1220 => x"abdc0871",
  1221 => x"88120c53",
  1222 => x"b00c843d",
  1223 => x"0d04803d",
  1224 => x"0d81518e",
  1225 => x"9d3fb008",
  1226 => x"83ffff06",
  1227 => x"51eaf13f",
  1228 => x"b00883ff",
  1229 => x"ff06b00c",
  1230 => x"823d0d04",
  1231 => x"803d0d81",
  1232 => x"518ccd3f",
  1233 => x"b00881ff",
  1234 => x"06519b83",
  1235 => x"3f800bb0",
  1236 => x"0c823d0d",
  1237 => x"04803d0d",
  1238 => x"81aca408",
  1239 => x"51f8bb95",
  1240 => x"86a1710c",
  1241 => x"810bb00c",
  1242 => x"823d0d04",
  1243 => x"fc3d0d81",
  1244 => x"518c9d3f",
  1245 => x"b00881ff",
  1246 => x"06548251",
  1247 => x"8c923fb0",
  1248 => x"0881ff06",
  1249 => x"81ac9808",
  1250 => x"84110870",
  1251 => x"fe8f0a06",
  1252 => x"77982b07",
  1253 => x"51545653",
  1254 => x"72802e86",
  1255 => x"3871810a",
  1256 => x"07527184",
  1257 => x"160c71b0",
  1258 => x"0c863d0d",
  1259 => x"04fd3d0d",
  1260 => x"81ac9808",
  1261 => x"84110855",
  1262 => x"5381518b",
  1263 => x"d33fb008",
  1264 => x"81ff0674",
  1265 => x"dfffff06",
  1266 => x"54527180",
  1267 => x"2e873873",
  1268 => x"a0808007",
  1269 => x"5382518b",
  1270 => x"b73fb008",
  1271 => x"81ff0673",
  1272 => x"efff0a06",
  1273 => x"55527180",
  1274 => x"2e873872",
  1275 => x"90800a07",
  1276 => x"5483518b",
  1277 => x"9b3fb008",
  1278 => x"81ff0674",
  1279 => x"f7ff0a06",
  1280 => x"54527180",
  1281 => x"2e873873",
  1282 => x"88800a07",
  1283 => x"5384518a",
  1284 => x"ff3fb008",
  1285 => x"81ff0673",
  1286 => x"fbff0a06",
  1287 => x"55527180",
  1288 => x"2e873872",
  1289 => x"84800a07",
  1290 => x"5485518a",
  1291 => x"e33fb008",
  1292 => x"81ff0674",
  1293 => x"fdff0a06",
  1294 => x"54527180",
  1295 => x"2e873873",
  1296 => x"82800a07",
  1297 => x"5381ac98",
  1298 => x"08738412",
  1299 => x"0c5472b0",
  1300 => x"0c853d0d",
  1301 => x"04fc3d0d",
  1302 => x"81ac9808",
  1303 => x"7008819b",
  1304 => x"a0535555",
  1305 => x"b68d3f73",
  1306 => x"9e2a8106",
  1307 => x"5271802e",
  1308 => x"b638819b",
  1309 => x"b051b5fb",
  1310 => x"3f81518a",
  1311 => x"933fb008",
  1312 => x"81ff0681",
  1313 => x"ac980884",
  1314 => x"110870fd",
  1315 => x"0a065656",
  1316 => x"56527180",
  1317 => x"2e863873",
  1318 => x"820a0753",
  1319 => x"7284160c",
  1320 => x"72b00c86",
  1321 => x"3d0d0481",
  1322 => x"9bb851b5",
  1323 => x"c63fc339",
  1324 => x"fc3d0d81",
  1325 => x"bbf00852",
  1326 => x"f881c08e",
  1327 => x"80539f0b",
  1328 => x"81ac9808",
  1329 => x"55557180",
  1330 => x"2e80e038",
  1331 => x"7281ff06",
  1332 => x"84150c81",
  1333 => x"bbf43370",
  1334 => x"81ff0651",
  1335 => x"5271802e",
  1336 => x"a438729f",
  1337 => x"2a731007",
  1338 => x"5374802e",
  1339 => x"a338ff15",
  1340 => x"7381ff06",
  1341 => x"84160c81",
  1342 => x"bbf43370",
  1343 => x"81ff0651",
  1344 => x"535571de",
  1345 => x"3872812a",
  1346 => x"739f2b07",
  1347 => x"5374df38",
  1348 => x"800bb00c",
  1349 => x"863d0d04",
  1350 => x"72812a73",
  1351 => x"9f2b0753",
  1352 => x"80fd51b7",
  1353 => x"e13f81ac",
  1354 => x"98085472",
  1355 => x"81ff0684",
  1356 => x"150c81bb",
  1357 => x"f4337081",
  1358 => x"ff065354",
  1359 => x"71802ed8",
  1360 => x"38729f2a",
  1361 => x"73100753",
  1362 => x"80fd51b7",
  1363 => x"b93f81ac",
  1364 => x"980854d7",
  1365 => x"39f73d0d",
  1366 => x"853d5496",
  1367 => x"53819bc0",
  1368 => x"527351bb",
  1369 => x"b13f9ea0",
  1370 => x"3f815188",
  1371 => x"a33f8052",
  1372 => x"80519cf1",
  1373 => x"3f735380",
  1374 => x"5281a0c0",
  1375 => x"51afdc3f",
  1376 => x"80528151",
  1377 => x"9cdf3f73",
  1378 => x"53825281",
  1379 => x"a0c051af",
  1380 => x"ca3f8052",
  1381 => x"82519ccd",
  1382 => x"3f735381",
  1383 => x"5281a0c0",
  1384 => x"51afb83f",
  1385 => x"80528451",
  1386 => x"9cbb3f73",
  1387 => x"53845281",
  1388 => x"a0c051af",
  1389 => x"a63f8052",
  1390 => x"85519ca9",
  1391 => x"3f735390",
  1392 => x"5281a0c0",
  1393 => x"51af943f",
  1394 => x"80528651",
  1395 => x"9c973f73",
  1396 => x"53835281",
  1397 => x"a0c051af",
  1398 => x"823f8b3d",
  1399 => x"0d04fef5",
  1400 => x"3f800bb0",
  1401 => x"0c04fc3d",
  1402 => x"0d9d9d3f",
  1403 => x"8187f054",
  1404 => x"80558452",
  1405 => x"74519bed",
  1406 => x"3f805373",
  1407 => x"70810555",
  1408 => x"33519ce7",
  1409 => x"3f811370",
  1410 => x"81ff0651",
  1411 => x"5380dc73",
  1412 => x"27e93881",
  1413 => x"157081ff",
  1414 => x"06565387",
  1415 => x"7527d338",
  1416 => x"800bb00c",
  1417 => x"863d0d04",
  1418 => x"fc3d0d81",
  1419 => x"ac980870",
  1420 => x"08810a06",
  1421 => x"81bbf00c",
  1422 => x"53b5ee3f",
  1423 => x"b69c3f81",
  1424 => x"bbf00880",
  1425 => x"dec35452",
  1426 => x"71843888",
  1427 => x"80537281",
  1428 => x"cf980c71",
  1429 => x"802e82aa",
  1430 => x"388194d0",
  1431 => x"51b2943f",
  1432 => x"8c51b1f5",
  1433 => x"3f819bc0",
  1434 => x"51b2883f",
  1435 => x"81bbf008",
  1436 => x"802e818f",
  1437 => x"38819bd8",
  1438 => x"51b1f83f",
  1439 => x"81bbf008",
  1440 => x"802e81ed",
  1441 => x"3881ac98",
  1442 => x"08841108",
  1443 => x"54548052",
  1444 => x"72fe8f0a",
  1445 => x"0672982b",
  1446 => x"07708416",
  1447 => x"0c811370",
  1448 => x"81ff0654",
  1449 => x"56538f72",
  1450 => x"27e638f8",
  1451 => x"81c08e80",
  1452 => x"539f5581",
  1453 => x"bbf00880",
  1454 => x"2e818c38",
  1455 => x"7281ff06",
  1456 => x"84150c81",
  1457 => x"bbf43370",
  1458 => x"81ff0651",
  1459 => x"5271802e",
  1460 => x"a438729f",
  1461 => x"2a731007",
  1462 => x"5374802e",
  1463 => x"a338ff15",
  1464 => x"7381ff06",
  1465 => x"84160c81",
  1466 => x"bbf43370",
  1467 => x"81ff0651",
  1468 => x"535571de",
  1469 => x"3872812a",
  1470 => x"739f2b07",
  1471 => x"5374df38",
  1472 => x"b8873f81",
  1473 => x"9be451b0",
  1474 => x"ea3f819c",
  1475 => x"8851b0e3",
  1476 => x"3fb451b2",
  1477 => x"a83f819c",
  1478 => x"9851b0d7",
  1479 => x"3f819ca0",
  1480 => x"51b0d03f",
  1481 => x"819cac51",
  1482 => x"b0c93f81",
  1483 => x"bbf008fe",
  1484 => x"d438be39",
  1485 => x"72812a73",
  1486 => x"9f2b0753",
  1487 => x"80fd51b3",
  1488 => x"c53f81ac",
  1489 => x"98085472",
  1490 => x"81ff0684",
  1491 => x"150c81bb",
  1492 => x"f4337081",
  1493 => x"ff065552",
  1494 => x"73802ed8",
  1495 => x"38729f2a",
  1496 => x"73100753",
  1497 => x"80fd51b3",
  1498 => x"9d3f81ac",
  1499 => x"980854d7",
  1500 => x"39d9a83f",
  1501 => x"81ac9808",
  1502 => x"84110854",
  1503 => x"548052fe",
  1504 => x"8f39b594",
  1505 => x"3f96e63f",
  1506 => x"fdcf3980",
  1507 => x"0b81cf8c",
  1508 => x"34800b81",
  1509 => x"cf883480",
  1510 => x"0b81cf90",
  1511 => x"0c04fc3d",
  1512 => x"0d765281",
  1513 => x"cf883370",
  1514 => x"10101071",
  1515 => x"100581bb",
  1516 => x"f8055254",
  1517 => x"bbee3f77",
  1518 => x"5281cf88",
  1519 => x"33709029",
  1520 => x"71317010",
  1521 => x"1081beb8",
  1522 => x"05535555",
  1523 => x"bbd63f81",
  1524 => x"cf883370",
  1525 => x"101081cd",
  1526 => x"b8057a71",
  1527 => x"0c548105",
  1528 => x"537281cf",
  1529 => x"8834863d",
  1530 => x"0d04803d",
  1531 => x"0d819ce0",
  1532 => x"51af803f",
  1533 => x"823d0d04",
  1534 => x"fe3d0d81",
  1535 => x"cf900853",
  1536 => x"72853884",
  1537 => x"3d0d0472",
  1538 => x"2db00853",
  1539 => x"800b81cf",
  1540 => x"900cb008",
  1541 => x"8c38819c",
  1542 => x"e051aed7",
  1543 => x"3f843d0d",
  1544 => x"04819ff4",
  1545 => x"51aecc3f",
  1546 => x"7283ffff",
  1547 => x"26aa3881",
  1548 => x"ff732796",
  1549 => x"38725290",
  1550 => x"51aedb3f",
  1551 => x"8a51ae99",
  1552 => x"3f819ce0",
  1553 => x"51aeac3f",
  1554 => x"d4397252",
  1555 => x"8851aec6",
  1556 => x"3f8a51ae",
  1557 => x"843fea39",
  1558 => x"7252a051",
  1559 => x"aeb83f8a",
  1560 => x"51adf63f",
  1561 => x"dc39fa3d",
  1562 => x"0d02a305",
  1563 => x"3356758d",
  1564 => x"2e80f438",
  1565 => x"75883270",
  1566 => x"307780ff",
  1567 => x"32703072",
  1568 => x"80257180",
  1569 => x"25075451",
  1570 => x"56585574",
  1571 => x"95389f76",
  1572 => x"278c3881",
  1573 => x"cf8c3355",
  1574 => x"80ce7527",
  1575 => x"ae38883d",
  1576 => x"0d0481cf",
  1577 => x"8c335675",
  1578 => x"802ef338",
  1579 => x"8851ada9",
  1580 => x"3fa051ad",
  1581 => x"a43f8851",
  1582 => x"ad9f3f81",
  1583 => x"cf8c33ff",
  1584 => x"05577681",
  1585 => x"cf8c3488",
  1586 => x"3d0d0475",
  1587 => x"51ad8a3f",
  1588 => x"81cf8c33",
  1589 => x"81115557",
  1590 => x"7381cf8c",
  1591 => x"347581ce",
  1592 => x"b8183488",
  1593 => x"3d0d048a",
  1594 => x"51acee3f",
  1595 => x"81cf8c33",
  1596 => x"81115654",
  1597 => x"7481cf8c",
  1598 => x"34800b81",
  1599 => x"ceb81534",
  1600 => x"8056800b",
  1601 => x"81ceb817",
  1602 => x"33565474",
  1603 => x"a02e8338",
  1604 => x"81547480",
  1605 => x"2e903873",
  1606 => x"802e8b38",
  1607 => x"81167081",
  1608 => x"ff065757",
  1609 => x"dd397580",
  1610 => x"2ebf3880",
  1611 => x"0b81cf88",
  1612 => x"33555574",
  1613 => x"7427ab38",
  1614 => x"73577410",
  1615 => x"10107510",
  1616 => x"05765481",
  1617 => x"ceb85381",
  1618 => x"bbf80551",
  1619 => x"baa23fb0",
  1620 => x"08802ea6",
  1621 => x"38811570",
  1622 => x"81ff0656",
  1623 => x"54767526",
  1624 => x"d938819c",
  1625 => x"e451ac8b",
  1626 => x"3f819ce0",
  1627 => x"51ac843f",
  1628 => x"800b81cf",
  1629 => x"8c34883d",
  1630 => x"0d047410",
  1631 => x"1081cdb8",
  1632 => x"05700881",
  1633 => x"cf900c56",
  1634 => x"800b81cf",
  1635 => x"8c34e739",
  1636 => x"f73d0d02",
  1637 => x"af053359",
  1638 => x"800b81ce",
  1639 => x"b83381ce",
  1640 => x"b8595556",
  1641 => x"73a02e09",
  1642 => x"81069638",
  1643 => x"81167081",
  1644 => x"ff0681ce",
  1645 => x"b8117033",
  1646 => x"53595754",
  1647 => x"73a02eec",
  1648 => x"38805877",
  1649 => x"792780ea",
  1650 => x"38807733",
  1651 => x"56547474",
  1652 => x"2e833881",
  1653 => x"5474a02e",
  1654 => x"9a387380",
  1655 => x"c53874a0",
  1656 => x"2e913881",
  1657 => x"187081ff",
  1658 => x"06595578",
  1659 => x"7826da38",
  1660 => x"80c03981",
  1661 => x"167081ff",
  1662 => x"0681ceb8",
  1663 => x"11703357",
  1664 => x"52575773",
  1665 => x"a02e0981",
  1666 => x"06d93881",
  1667 => x"167081ff",
  1668 => x"0681ceb8",
  1669 => x"11703357",
  1670 => x"52575773",
  1671 => x"a02ed438",
  1672 => x"c2398116",
  1673 => x"7081ff06",
  1674 => x"81ceb811",
  1675 => x"595755ff",
  1676 => x"98398a53",
  1677 => x"8b3dfc05",
  1678 => x"527651bc",
  1679 => x"f83f8b3d",
  1680 => x"0d04f73d",
  1681 => x"0d02af05",
  1682 => x"3359800b",
  1683 => x"81ceb833",
  1684 => x"81ceb859",
  1685 => x"555673a0",
  1686 => x"2e098106",
  1687 => x"96388116",
  1688 => x"7081ff06",
  1689 => x"81ceb811",
  1690 => x"70335359",
  1691 => x"575473a0",
  1692 => x"2eec3880",
  1693 => x"58777927",
  1694 => x"80ea3880",
  1695 => x"77335654",
  1696 => x"74742e83",
  1697 => x"38815474",
  1698 => x"a02e9a38",
  1699 => x"7380c538",
  1700 => x"74a02e91",
  1701 => x"38811870",
  1702 => x"81ff0659",
  1703 => x"55787826",
  1704 => x"da3880c0",
  1705 => x"39811670",
  1706 => x"81ff0681",
  1707 => x"ceb81170",
  1708 => x"33575257",
  1709 => x"5773a02e",
  1710 => x"098106d9",
  1711 => x"38811670",
  1712 => x"81ff0681",
  1713 => x"ceb81170",
  1714 => x"33575257",
  1715 => x"5773a02e",
  1716 => x"d438c239",
  1717 => x"81167081",
  1718 => x"ff0681ce",
  1719 => x"b8115957",
  1720 => x"55ff9839",
  1721 => x"90538b3d",
  1722 => x"fc055276",
  1723 => x"51bee33f",
  1724 => x"8b3d0d04",
  1725 => x"fc3d0d8a",
  1726 => x"51a8de3f",
  1727 => x"819cf851",
  1728 => x"a8f13f80",
  1729 => x"0b81cf88",
  1730 => x"33535372",
  1731 => x"722780f5",
  1732 => x"38721010",
  1733 => x"10731005",
  1734 => x"81bbf805",
  1735 => x"705254a8",
  1736 => x"d23f7284",
  1737 => x"2b707431",
  1738 => x"822b81be",
  1739 => x"b8113351",
  1740 => x"53557180",
  1741 => x"2eb73873",
  1742 => x"51b5d63f",
  1743 => x"b00881ff",
  1744 => x"06527189",
  1745 => x"269338a0",
  1746 => x"51a88e3f",
  1747 => x"81127081",
  1748 => x"ff065354",
  1749 => x"897227ef",
  1750 => x"38819d90",
  1751 => x"51a8943f",
  1752 => x"74733182",
  1753 => x"2b81beb8",
  1754 => x"0551a887",
  1755 => x"3f8a51a7",
  1756 => x"e83f8113",
  1757 => x"7081ff06",
  1758 => x"81cf8833",
  1759 => x"54545571",
  1760 => x"7326ff8d",
  1761 => x"388a51a7",
  1762 => x"d03f81cf",
  1763 => x"8833b00c",
  1764 => x"863d0d04",
  1765 => x"f53d0d7d",
  1766 => x"598a5481",
  1767 => x"028405ba",
  1768 => x"0522575c",
  1769 => x"80e45380",
  1770 => x"52abc53f",
  1771 => x"b008722e",
  1772 => x"09810683",
  1773 => x"38815272",
  1774 => x"802eb138",
  1775 => x"71802e91",
  1776 => x"3880e451",
  1777 => x"aac03fff",
  1778 => x"137081ff",
  1779 => x"065452d7",
  1780 => x"3972802e",
  1781 => x"9738abab",
  1782 => x"3fb00881",
  1783 => x"ff065271",
  1784 => x"952e829a",
  1785 => x"387180c3",
  1786 => x"2e81ec38",
  1787 => x"ff147081",
  1788 => x"ff065553",
  1789 => x"73ffad38",
  1790 => x"75802e81",
  1791 => x"cc388a7c",
  1792 => x"095c5a81",
  1793 => x"51ab9e3f",
  1794 => x"7b51ab99",
  1795 => x"3f7a51ab",
  1796 => x"943f8070",
  1797 => x"55578180",
  1798 => x"55ff1570",
  1799 => x"81ff0656",
  1800 => x"529a5375",
  1801 => x"802e9138",
  1802 => x"78708105",
  1803 => x"5a33ff17",
  1804 => x"7083ffff",
  1805 => x"06585353",
  1806 => x"7251aae9",
  1807 => x"3f77802e",
  1808 => x"81a93872",
  1809 => x"882b7432",
  1810 => x"53875472",
  1811 => x"902b5280",
  1812 => x"72248188",
  1813 => x"38721083",
  1814 => x"fffe0653",
  1815 => x"ff145473",
  1816 => x"8025e838",
  1817 => x"7283ffff",
  1818 => x"065474ff",
  1819 => x"ac387780",
  1820 => x"2e818338",
  1821 => x"73882a51",
  1822 => x"aaab3f73",
  1823 => x"81ff0651",
  1824 => x"aaa33fa9",
  1825 => x"eb3fb008",
  1826 => x"fa38a9f7",
  1827 => x"3fb00881",
  1828 => x"ff065271",
  1829 => x"862e80eb",
  1830 => x"3871982e",
  1831 => x"80f038ff",
  1832 => x"1a7081ff",
  1833 => x"065b5479",
  1834 => x"fed938fe",
  1835 => x"5271b00c",
  1836 => x"8d3d0d04",
  1837 => x"a9ba3fb0",
  1838 => x"08fa38a9",
  1839 => x"c63fb008",
  1840 => x"81ff0652",
  1841 => x"71862ee5",
  1842 => x"388451a9",
  1843 => x"d83fa9a0",
  1844 => x"3fb008e0",
  1845 => x"38e53981",
  1846 => x"58fe9d39",
  1847 => x"7210a0a1",
  1848 => x"327083ff",
  1849 => x"ff065452",
  1850 => x"fef23972",
  1851 => x"177081ff",
  1852 => x"065852fe",
  1853 => x"f5397651",
  1854 => x"a9ab3fff",
  1855 => x"86398058",
  1856 => x"fdf63981",
  1857 => x"1c7081ff",
  1858 => x"065d55fd",
  1859 => x"eb39ff0b",
  1860 => x"b00c8d3d",
  1861 => x"0d04f63d",
  1862 => x"0d7c7e5b",
  1863 => x"5980c357",
  1864 => x"8a55815b",
  1865 => x"805880e4",
  1866 => x"53805477",
  1867 => x"7a2482aa",
  1868 => x"387651a8",
  1869 => x"f03f8052",
  1870 => x"a8b63fb0",
  1871 => x"08722e09",
  1872 => x"81068338",
  1873 => x"81527280",
  1874 => x"2e81e638",
  1875 => x"71802e91",
  1876 => x"3880e451",
  1877 => x"a7b03fff",
  1878 => x"137081ff",
  1879 => x"065452d6",
  1880 => x"3972802e",
  1881 => x"81cb38a8",
  1882 => x"9a3fb008",
  1883 => x"81ff0652",
  1884 => x"71842e82",
  1885 => x"81387184",
  1886 => x"2481ca38",
  1887 => x"71812e09",
  1888 => x"810681ad",
  1889 => x"388657a7",
  1890 => x"fa3fb008",
  1891 => x"81ff0653",
  1892 => x"7a732e83",
  1893 => x"389557a7",
  1894 => x"ea3fb008",
  1895 => x"097081ff",
  1896 => x"0657527a",
  1897 => x"762e8338",
  1898 => x"95578053",
  1899 => x"a7d53f78",
  1900 => x"1356b008",
  1901 => x"76348113",
  1902 => x"7081ff06",
  1903 => x"70982b58",
  1904 => x"54527580",
  1905 => x"25e63880",
  1906 => x"56781670",
  1907 => x"3370882b",
  1908 => x"76325253",
  1909 => x"53875472",
  1910 => x"902b5280",
  1911 => x"72248187",
  1912 => x"38721083",
  1913 => x"fffe0653",
  1914 => x"ff145473",
  1915 => x"8025e838",
  1916 => x"7283ffff",
  1917 => x"06811770",
  1918 => x"81ff0670",
  1919 => x"982b5658",
  1920 => x"53547280",
  1921 => x"25c338a6",
  1922 => x"fa3fb008",
  1923 => x"81ff0674",
  1924 => x"882a5753",
  1925 => x"72762e83",
  1926 => x"389557a6",
  1927 => x"e63fb008",
  1928 => x"81ff0674",
  1929 => x"81ff0653",
  1930 => x"5675722e",
  1931 => x"80d43895",
  1932 => x"57ff1570",
  1933 => x"81ff0656",
  1934 => x"5274fdea",
  1935 => x"38fe0bb0",
  1936 => x"0c8c3d0d",
  1937 => x"0471982e",
  1938 => x"098106e5",
  1939 => x"388651a6",
  1940 => x"d43fff0b",
  1941 => x"b00c8c3d",
  1942 => x"0d049851",
  1943 => x"a6c73ffd",
  1944 => x"0bb00c8c",
  1945 => x"3d0d0472",
  1946 => x"10a0a132",
  1947 => x"7083ffff",
  1948 => x"065452fe",
  1949 => x"f3398651",
  1950 => x"a6ab3f77",
  1951 => x"b00c8c3d",
  1952 => x"0d047686",
  1953 => x"2e098106",
  1954 => x"ffa73877",
  1955 => x"84808029",
  1956 => x"82800a05",
  1957 => x"70902c81",
  1958 => x"801b811e",
  1959 => x"7081ff06",
  1960 => x"5f575b59",
  1961 => x"5374fcfe",
  1962 => x"38ff9239",
  1963 => x"fe3d0d02",
  1964 => x"93053302",
  1965 => x"84059705",
  1966 => x"33545271",
  1967 => x"812e9238",
  1968 => x"7180d52e",
  1969 => x"bb38819d",
  1970 => x"9451a1a7",
  1971 => x"3f843d0d",
  1972 => x"04819da0",
  1973 => x"51a19c3f",
  1974 => x"72912e81",
  1975 => x"d9387291",
  1976 => x"24b53872",
  1977 => x"8c2e81e4",
  1978 => x"38728c24",
  1979 => x"80dc3872",
  1980 => x"862e81b7",
  1981 => x"38819dac",
  1982 => x"51a0f83f",
  1983 => x"843d0d04",
  1984 => x"819dbc51",
  1985 => x"a0ed3f72",
  1986 => x"8726ea38",
  1987 => x"72101081",
  1988 => x"a0a00552",
  1989 => x"71080472",
  1990 => x"a82e81a5",
  1991 => x"3872a824",
  1992 => x"9438729a",
  1993 => x"2e098106",
  1994 => x"cc38819d",
  1995 => x"c851a0c3",
  1996 => x"3f843d0d",
  1997 => x"047280e1",
  1998 => x"2e098106",
  1999 => x"ffb73881",
  2000 => x"9de451a0",
  2001 => x"ae3f843d",
  2002 => x"0d04728f",
  2003 => x"2e098106",
  2004 => x"ffa33881",
  2005 => x"9df451a0",
  2006 => x"9a3f843d",
  2007 => x"0d04819e",
  2008 => x"9051a08f",
  2009 => x"3f843d0d",
  2010 => x"04819bc0",
  2011 => x"51a0843f",
  2012 => x"843d0d04",
  2013 => x"819ea851",
  2014 => x"9ff93f84",
  2015 => x"3d0d0481",
  2016 => x"9ebc519f",
  2017 => x"ee3f843d",
  2018 => x"0d04819e",
  2019 => x"cc519fe3",
  2020 => x"3f843d0d",
  2021 => x"04819ee4",
  2022 => x"519fd83f",
  2023 => x"843d0d04",
  2024 => x"819ef851",
  2025 => x"9fcd3f84",
  2026 => x"3d0d0481",
  2027 => x"9f88519f",
  2028 => x"c23f843d",
  2029 => x"0d04819f",
  2030 => x"98519fb7",
  2031 => x"3f843d0d",
  2032 => x"04819fac",
  2033 => x"519fac3f",
  2034 => x"843d0d04",
  2035 => x"819fcc51",
  2036 => x"9fa13f84",
  2037 => x"3d0d04f7",
  2038 => x"3d0d02b3",
  2039 => x"05337c70",
  2040 => x"08c08080",
  2041 => x"0659545a",
  2042 => x"80567583",
  2043 => x"2b7707bf",
  2044 => x"e0800770",
  2045 => x"70840552",
  2046 => x"0871088c",
  2047 => x"2abffe80",
  2048 => x"06790771",
  2049 => x"982a728c",
  2050 => x"2a9fff06",
  2051 => x"73852a70",
  2052 => x"8f06759f",
  2053 => x"06565158",
  2054 => x"5d585255",
  2055 => x"58748d38",
  2056 => x"8116568f",
  2057 => x"7627c338",
  2058 => x"8b3d0d04",
  2059 => x"819fdc51",
  2060 => x"9ec13f75",
  2061 => x"51a0863f",
  2062 => x"8452b008",
  2063 => x"51d5e93f",
  2064 => x"819fe851",
  2065 => x"9ead3f74",
  2066 => x"5288519e",
  2067 => x"c93f8452",
  2068 => x"b00851d5",
  2069 => x"d33f819f",
  2070 => x"f0519e97",
  2071 => x"3f785290",
  2072 => x"519eb33f",
  2073 => x"8652b008",
  2074 => x"51d5bd3f",
  2075 => x"819ff851",
  2076 => x"9e813f72",
  2077 => x"519fc63f",
  2078 => x"8452b008",
  2079 => x"51d5a93f",
  2080 => x"81a08051",
  2081 => x"9ded3f73",
  2082 => x"519fb23f",
  2083 => x"8452b008",
  2084 => x"51d5953f",
  2085 => x"81a08851",
  2086 => x"9dd93f77",
  2087 => x"52a0519d",
  2088 => x"f53f8a52",
  2089 => x"b00851d4",
  2090 => x"ff3f7992",
  2091 => x"388a519d",
  2092 => x"a83f8116",
  2093 => x"568f7627",
  2094 => x"feb038fe",
  2095 => x"eb397881",
  2096 => x"ff065274",
  2097 => x"51fbe53f",
  2098 => x"8a519d8d",
  2099 => x"3fe439f8",
  2100 => x"3d0d02ab",
  2101 => x"05335980",
  2102 => x"5675852b",
  2103 => x"e09011e0",
  2104 => x"80120870",
  2105 => x"982a718c",
  2106 => x"2a9fff06",
  2107 => x"72852a70",
  2108 => x"8f06749f",
  2109 => x"06555158",
  2110 => x"5b535659",
  2111 => x"5574802e",
  2112 => x"81a13875",
  2113 => x"bf2681a9",
  2114 => x"3881a090",
  2115 => x"519ce43f",
  2116 => x"75519ea9",
  2117 => x"3f8652b0",
  2118 => x"0851d48c",
  2119 => x"3f819fe8",
  2120 => x"519cd03f",
  2121 => x"74528851",
  2122 => x"9cec3f84",
  2123 => x"52b00851",
  2124 => x"d3f63f81",
  2125 => x"9ff0519c",
  2126 => x"ba3f7652",
  2127 => x"90519cd6",
  2128 => x"3f8652b0",
  2129 => x"0851d3e0",
  2130 => x"3f819ff8",
  2131 => x"519ca43f",
  2132 => x"72519de9",
  2133 => x"3f8452b0",
  2134 => x"0851d3cc",
  2135 => x"3f81a080",
  2136 => x"519c903f",
  2137 => x"73519dd5",
  2138 => x"3f8452b0",
  2139 => x"0851d3b8",
  2140 => x"3f81a088",
  2141 => x"519bfc3f",
  2142 => x"7708c080",
  2143 => x"800652a0",
  2144 => x"519c933f",
  2145 => x"8a52b008",
  2146 => x"51d39d3f",
  2147 => x"7881ac38",
  2148 => x"8a519bc5",
  2149 => x"3f805374",
  2150 => x"812e81d9",
  2151 => x"3876862e",
  2152 => x"81b53881",
  2153 => x"165680ff",
  2154 => x"7627fead",
  2155 => x"388a3d0d",
  2156 => x"0481a098",
  2157 => x"519bbc3f",
  2158 => x"c016519d",
  2159 => x"803f8652",
  2160 => x"b00851d2",
  2161 => x"e33f819f",
  2162 => x"e8519ba7",
  2163 => x"3f745288",
  2164 => x"519bc33f",
  2165 => x"8452b008",
  2166 => x"51d2cd3f",
  2167 => x"819ff051",
  2168 => x"9b913f76",
  2169 => x"5290519b",
  2170 => x"ad3f8652",
  2171 => x"b00851d2",
  2172 => x"b73f819f",
  2173 => x"f8519afb",
  2174 => x"3f72519c",
  2175 => x"c03f8452",
  2176 => x"b00851d2",
  2177 => x"a33f81a0",
  2178 => x"80519ae7",
  2179 => x"3f73519c",
  2180 => x"ac3f8452",
  2181 => x"b00851d2",
  2182 => x"8f3f81a0",
  2183 => x"88519ad3",
  2184 => x"3f7708c0",
  2185 => x"80800652",
  2186 => x"a0519aea",
  2187 => x"3f8a52b0",
  2188 => x"0851d1f4",
  2189 => x"3f78802e",
  2190 => x"fed63876",
  2191 => x"81ff0652",
  2192 => x"7451f8e8",
  2193 => x"3f8a519a",
  2194 => x"903f8053",
  2195 => x"74812e09",
  2196 => x"8106fec9",
  2197 => x"389f3972",
  2198 => x"81065776",
  2199 => x"802efec3",
  2200 => x"38785277",
  2201 => x"51faf03f",
  2202 => x"81165680",
  2203 => x"ff7627fc",
  2204 => x"e838feb9",
  2205 => x"39745376",
  2206 => x"862e0981",
  2207 => x"06fea438",
  2208 => x"d639803d",
  2209 => x"0d81ac90",
  2210 => x"08519971",
  2211 => x"0c81800b",
  2212 => x"84120c81",
  2213 => x"ac8c0851",
  2214 => x"99710c81",
  2215 => x"800b8412",
  2216 => x"0c823d0d",
  2217 => x"04fe3d0d",
  2218 => x"74028405",
  2219 => x"97053302",
  2220 => x"88059b05",
  2221 => x"3388130c",
  2222 => x"8c120c53",
  2223 => x"8c130870",
  2224 => x"812a8106",
  2225 => x"515271f4",
  2226 => x"388c1308",
  2227 => x"7081ff06",
  2228 => x"b00c5184",
  2229 => x"3d0d0480",
  2230 => x"3d0d728c",
  2231 => x"11087087",
  2232 => x"2a813281",
  2233 => x"06b00c51",
  2234 => x"51823d0d",
  2235 => x"04fe3d0d",
  2236 => x"ff903f81",
  2237 => x"ec538190",
  2238 => x"5281ac90",
  2239 => x"0851ffa5",
  2240 => x"3f9d5390",
  2241 => x"5281ac90",
  2242 => x"0851ff99",
  2243 => x"3f80c553",
  2244 => x"80d05281",
  2245 => x"ac900851",
  2246 => x"ff8b3f81",
  2247 => x"ec538190",
  2248 => x"5281ac90",
  2249 => x"0851fefd",
  2250 => x"3fa15390",
  2251 => x"5281ac90",
  2252 => x"0851fef1",
  2253 => x"3f895380",
  2254 => x"d05281ac",
  2255 => x"900851fe",
  2256 => x"e43f81ec",
  2257 => x"53819052",
  2258 => x"81ac9008",
  2259 => x"51fed63f",
  2260 => x"b3539052",
  2261 => x"81ac9008",
  2262 => x"51feca3f",
  2263 => x"885380d0",
  2264 => x"5281ac90",
  2265 => x"0851febd",
  2266 => x"3f81ec53",
  2267 => x"81905281",
  2268 => x"ac900851",
  2269 => x"feaf3fb4",
  2270 => x"53905281",
  2271 => x"ac900851",
  2272 => x"fea33f96",
  2273 => x"5380d052",
  2274 => x"81ac9008",
  2275 => x"51fe963f",
  2276 => x"81ec5381",
  2277 => x"905281ac",
  2278 => x"900851fe",
  2279 => x"883fb653",
  2280 => x"905281ac",
  2281 => x"900851fd",
  2282 => x"fc3f80e0",
  2283 => x"5380d052",
  2284 => x"81ac9008",
  2285 => x"51fdee3f",
  2286 => x"81ec5381",
  2287 => x"905281ac",
  2288 => x"900851fd",
  2289 => x"e03f80c9",
  2290 => x"53905281",
  2291 => x"ac900851",
  2292 => x"fdd33f81",
  2293 => x"c05380d0",
  2294 => x"5281ac90",
  2295 => x"0851fdc5",
  2296 => x"3f843d0d",
  2297 => x"04fd3d0d",
  2298 => x"02970533",
  2299 => x"0284059b",
  2300 => x"05337181",
  2301 => x"b00781bf",
  2302 => x"06535454",
  2303 => x"f8808098",
  2304 => x"8071710c",
  2305 => x"73842a90",
  2306 => x"07710c73",
  2307 => x"8f06710c",
  2308 => x"527281ab",
  2309 => x"ec347381",
  2310 => x"abf03485",
  2311 => x"3d0d04fd",
  2312 => x"3d0d0297",
  2313 => x"053381ab",
  2314 => x"f0335473",
  2315 => x"05870602",
  2316 => x"84059a05",
  2317 => x"2281abec",
  2318 => x"33547305",
  2319 => x"7081ff06",
  2320 => x"7281b007",
  2321 => x"54515454",
  2322 => x"f8808098",
  2323 => x"8071710c",
  2324 => x"73842a90",
  2325 => x"07710c73",
  2326 => x"8f06710c",
  2327 => x"527281ab",
  2328 => x"ec347381",
  2329 => x"abf03485",
  2330 => x"3d0d04ff",
  2331 => x"3d0d028f",
  2332 => x"0533f880",
  2333 => x"8098840c",
  2334 => x"81abec33",
  2335 => x"81055170",
  2336 => x"81abec34",
  2337 => x"833d0d04",
  2338 => x"ff3d0d80",
  2339 => x"c00bf880",
  2340 => x"8098800c",
  2341 => x"81a10bf8",
  2342 => x"80809880",
  2343 => x"0c81c00b",
  2344 => x"f8808098",
  2345 => x"800c81a4",
  2346 => x"0bf88080",
  2347 => x"98800c81",
  2348 => x"a60bf880",
  2349 => x"8098800c",
  2350 => x"81a20bf8",
  2351 => x"80809880",
  2352 => x"0caf0bf8",
  2353 => x"80809880",
  2354 => x"0ca50bf8",
  2355 => x"80809880",
  2356 => x"0c81810b",
  2357 => x"f8808098",
  2358 => x"800c9d0b",
  2359 => x"f8808098",
  2360 => x"800c81fa",
  2361 => x"0bf88080",
  2362 => x"98800c80",
  2363 => x"0bf88080",
  2364 => x"98800c80",
  2365 => x"527181b0",
  2366 => x"0781bf06",
  2367 => x"f8808098",
  2368 => x"800c900b",
  2369 => x"f8808098",
  2370 => x"800c800b",
  2371 => x"f8808098",
  2372 => x"800c8051",
  2373 => x"800bf880",
  2374 => x"8098840c",
  2375 => x"81117081",
  2376 => x"ff065151",
  2377 => x"80e57127",
  2378 => x"eb388112",
  2379 => x"7081ff06",
  2380 => x"53518772",
  2381 => x"27ffbe38",
  2382 => x"81b00bf8",
  2383 => x"80809880",
  2384 => x"0c900bf8",
  2385 => x"80809880",
  2386 => x"0c800bf8",
  2387 => x"80809880",
  2388 => x"0c800b81",
  2389 => x"abec3480",
  2390 => x"0b81abf0",
  2391 => x"3481af0b",
  2392 => x"f8808098",
  2393 => x"800c833d",
  2394 => x"0d04ed3d",
  2395 => x"0d650284",
  2396 => x"0580db05",
  2397 => x"33028805",
  2398 => x"80df0533",
  2399 => x"5f5a5680",
  2400 => x"7981067a",
  2401 => x"812a8106",
  2402 => x"7b832b81",
  2403 => x"80067c82",
  2404 => x"2a810657",
  2405 => x"5e435f5c",
  2406 => x"81ff4272",
  2407 => x"7c2e0981",
  2408 => x"0683387b",
  2409 => x"42881608",
  2410 => x"5574802e",
  2411 => x"839f3885",
  2412 => x"16335aff",
  2413 => x"537c7a26",
  2414 => x"8e388416",
  2415 => x"3354737d",
  2416 => x"2685387c",
  2417 => x"74315374",
  2418 => x"13703354",
  2419 => x"577281ff",
  2420 => x"06831733",
  2421 => x"70982b81",
  2422 => x"ff0a119b",
  2423 => x"2a810551",
  2424 => x"5a404081",
  2425 => x"53748338",
  2426 => x"74537281",
  2427 => x"ff064380",
  2428 => x"7a81ff06",
  2429 => x"4557ff54",
  2430 => x"7c64268b",
  2431 => x"38841633",
  2432 => x"537c7327",
  2433 => x"83ce3873",
  2434 => x"7481ff06",
  2435 => x"5553805a",
  2436 => x"797324ab",
  2437 => x"38747a2e",
  2438 => x"09810682",
  2439 => x"bb387e98",
  2440 => x"2b81ff0a",
  2441 => x"119b2a82",
  2442 => x"18337171",
  2443 => x"29117081",
  2444 => x"ff067871",
  2445 => x"298c1c08",
  2446 => x"0552435d",
  2447 => x"5758447f",
  2448 => x"63057081",
  2449 => x"ff067063",
  2450 => x"2b7081ff",
  2451 => x"067b622b",
  2452 => x"7081ff06",
  2453 => x"7e832a81",
  2454 => x"065c5557",
  2455 => x"5256455f",
  2456 => x"75802e8f",
  2457 => x"3881abec",
  2458 => x"33640559",
  2459 => x"7880e624",
  2460 => x"8dc6387f",
  2461 => x"78296430",
  2462 => x"5e577b7e",
  2463 => x"2c982b70",
  2464 => x"982c5540",
  2465 => x"73772580",
  2466 => x"fc38ff1f",
  2467 => x"7c81065a",
  2468 => x"537b732e",
  2469 => x"83843860",
  2470 => x"85da3861",
  2471 => x"84a5387d",
  2472 => x"802e81fe",
  2473 => x"38791470",
  2474 => x"33705254",
  2475 => x"56805578",
  2476 => x"752e8538",
  2477 => x"72842a56",
  2478 => x"75832a81",
  2479 => x"06407f80",
  2480 => x"2e843881",
  2481 => x"c0557582",
  2482 => x"2a810640",
  2483 => x"7f802e85",
  2484 => x"3874b007",
  2485 => x"5575812a",
  2486 => x"8106407f",
  2487 => x"802e8538",
  2488 => x"748c0755",
  2489 => x"75810653",
  2490 => x"72802e85",
  2491 => x"38748307",
  2492 => x"557451fa",
  2493 => x"f63f7714",
  2494 => x"982b7098",
  2495 => x"2c555576",
  2496 => x"7424ffa1",
  2497 => x"3862802e",
  2498 => x"9638617f",
  2499 => x"ff055654",
  2500 => x"7b752e81",
  2501 => x"e3387351",
  2502 => x"fad13f60",
  2503 => x"81bd387c",
  2504 => x"528151f9",
  2505 => x"fa3f811c",
  2506 => x"7081ff06",
  2507 => x"5d547e7c",
  2508 => x"26fec738",
  2509 => x"63527e30",
  2510 => x"70982b70",
  2511 => x"982c535c",
  2512 => x"5cf9dc3f",
  2513 => x"635372b0",
  2514 => x"0c953d0d",
  2515 => x"04821633",
  2516 => x"8517335b",
  2517 => x"53fcf639",
  2518 => x"73802eaf",
  2519 => x"38ff1470",
  2520 => x"81ff0655",
  2521 => x"537381ff",
  2522 => x"2ea13874",
  2523 => x"70810556",
  2524 => x"33770570",
  2525 => x"83ffff06",
  2526 => x"ff167081",
  2527 => x"ff065755",
  2528 => x"585a7381",
  2529 => x"ff2e0981",
  2530 => x"06e1387e",
  2531 => x"982b81ff",
  2532 => x"0a119b2a",
  2533 => x"70792919",
  2534 => x"8c190805",
  2535 => x"5c4055fd",
  2536 => x"9e397914",
  2537 => x"70335259",
  2538 => x"f9c13f77",
  2539 => x"14982b70",
  2540 => x"982c5553",
  2541 => x"737725fe",
  2542 => x"cc387914",
  2543 => x"70335259",
  2544 => x"f9a93f77",
  2545 => x"14982b70",
  2546 => x"982c5553",
  2547 => x"767424d2",
  2548 => x"38feb239",
  2549 => x"7c733154",
  2550 => x"fcad3973",
  2551 => x"51f98c3f",
  2552 => x"7c528151",
  2553 => x"f8b93f81",
  2554 => x"1c7081ff",
  2555 => x"065d547e",
  2556 => x"7c26fd86",
  2557 => x"38febd39",
  2558 => x"617b3270",
  2559 => x"81ff0655",
  2560 => x"567d802e",
  2561 => x"fe90387a",
  2562 => x"812a7432",
  2563 => x"705254f8",
  2564 => x"da3f6080",
  2565 => x"2efe8838",
  2566 => x"c2396087",
  2567 => x"8f386185",
  2568 => x"d3387d80",
  2569 => x"2e80e638",
  2570 => x"79147033",
  2571 => x"7c077052",
  2572 => x"54568055",
  2573 => x"78752e85",
  2574 => x"3872842a",
  2575 => x"5675832a",
  2576 => x"81065372",
  2577 => x"802e8438",
  2578 => x"81c05575",
  2579 => x"822a8106",
  2580 => x"5372802e",
  2581 => x"853874b0",
  2582 => x"07557581",
  2583 => x"2a810653",
  2584 => x"72802e85",
  2585 => x"38748c07",
  2586 => x"55758106",
  2587 => x"407f802e",
  2588 => x"85387483",
  2589 => x"07557451",
  2590 => x"f7f13f77",
  2591 => x"14982b70",
  2592 => x"982c5553",
  2593 => x"767424ff",
  2594 => x"9f38fcf9",
  2595 => x"39791470",
  2596 => x"337c0752",
  2597 => x"55f7d43f",
  2598 => x"7714982b",
  2599 => x"70982c55",
  2600 => x"59737725",
  2601 => x"fcdf3879",
  2602 => x"1470337c",
  2603 => x"075255f7",
  2604 => x"ba3f7714",
  2605 => x"982b7098",
  2606 => x"2c555976",
  2607 => x"7424ce38",
  2608 => x"fcc3397d",
  2609 => x"802e80ea",
  2610 => x"38791470",
  2611 => x"33705854",
  2612 => x"55805578",
  2613 => x"752e8538",
  2614 => x"72842a56",
  2615 => x"75832a81",
  2616 => x"06537280",
  2617 => x"2e843881",
  2618 => x"c0557582",
  2619 => x"2a810653",
  2620 => x"72802e85",
  2621 => x"3874b007",
  2622 => x"5575812a",
  2623 => x"81065372",
  2624 => x"802e8538",
  2625 => x"748c0755",
  2626 => x"75810640",
  2627 => x"7f802e85",
  2628 => x"38748307",
  2629 => x"55740970",
  2630 => x"81ff0652",
  2631 => x"53f6cc3f",
  2632 => x"7714982b",
  2633 => x"70982c55",
  2634 => x"56767424",
  2635 => x"ff9b38fb",
  2636 => x"d4397914",
  2637 => x"70337009",
  2638 => x"7081ff06",
  2639 => x"54585440",
  2640 => x"f6a93f77",
  2641 => x"14982b70",
  2642 => x"982c5559",
  2643 => x"737725fb",
  2644 => x"b4387914",
  2645 => x"70337009",
  2646 => x"7081ff06",
  2647 => x"54585440",
  2648 => x"f6893f77",
  2649 => x"14982b70",
  2650 => x"982c5559",
  2651 => x"767424c2",
  2652 => x"38fb9239",
  2653 => x"61802e81",
  2654 => x"c8387d80",
  2655 => x"2e80f138",
  2656 => x"79147033",
  2657 => x"70585455",
  2658 => x"80557875",
  2659 => x"2e853872",
  2660 => x"842a5675",
  2661 => x"832a8106",
  2662 => x"407f802e",
  2663 => x"843881c0",
  2664 => x"5575822a",
  2665 => x"8106407f",
  2666 => x"802e8538",
  2667 => x"74b00755",
  2668 => x"75812a81",
  2669 => x"06407f80",
  2670 => x"2e853874",
  2671 => x"8c075575",
  2672 => x"81065372",
  2673 => x"802e8538",
  2674 => x"74830755",
  2675 => x"74097081",
  2676 => x"ff067053",
  2677 => x"4156f593",
  2678 => x"3f7f51f5",
  2679 => x"8e3f7714",
  2680 => x"982b7098",
  2681 => x"2c555376",
  2682 => x"7424ff94",
  2683 => x"38fa9639",
  2684 => x"79147033",
  2685 => x"70097081",
  2686 => x"ff067055",
  2687 => x"59554155",
  2688 => x"f4e93f75",
  2689 => x"51f4e43f",
  2690 => x"7714982b",
  2691 => x"70982c55",
  2692 => x"59737725",
  2693 => x"f9ef3879",
  2694 => x"14703370",
  2695 => x"097081ff",
  2696 => x"06705559",
  2697 => x"554155f4",
  2698 => x"c23f7551",
  2699 => x"f4bd3f77",
  2700 => x"14982b70",
  2701 => x"982c5559",
  2702 => x"767424ff",
  2703 => x"b338f9c5",
  2704 => x"397d802e",
  2705 => x"80ee3879",
  2706 => x"14703370",
  2707 => x"58545580",
  2708 => x"5578752e",
  2709 => x"85387284",
  2710 => x"2a567583",
  2711 => x"2a810653",
  2712 => x"72802e84",
  2713 => x"3881c055",
  2714 => x"75822a81",
  2715 => x"06537280",
  2716 => x"2e853874",
  2717 => x"b0075575",
  2718 => x"812a8106",
  2719 => x"5372802e",
  2720 => x"8538748c",
  2721 => x"07557581",
  2722 => x"06407f80",
  2723 => x"2e853874",
  2724 => x"83075574",
  2725 => x"81ff0670",
  2726 => x"5256f3cf",
  2727 => x"3f7551f3",
  2728 => x"ca3f7714",
  2729 => x"982b7098",
  2730 => x"2c555376",
  2731 => x"7424ff97",
  2732 => x"38f8d239",
  2733 => x"79147033",
  2734 => x"70535740",
  2735 => x"f3ad3f75",
  2736 => x"51f3a83f",
  2737 => x"7714982b",
  2738 => x"70982c55",
  2739 => x"59737725",
  2740 => x"f8b33879",
  2741 => x"14703370",
  2742 => x"535740f3",
  2743 => x"8e3f7551",
  2744 => x"f3893f77",
  2745 => x"14982b70",
  2746 => x"982c5559",
  2747 => x"767424c4",
  2748 => x"38f89239",
  2749 => x"7d802e80",
  2750 => x"ec387914",
  2751 => x"70337c07",
  2752 => x"70525456",
  2753 => x"80557875",
  2754 => x"2e853872",
  2755 => x"842a5675",
  2756 => x"832a8106",
  2757 => x"5372802e",
  2758 => x"843881c0",
  2759 => x"5575822a",
  2760 => x"81065372",
  2761 => x"802e8538",
  2762 => x"74b00755",
  2763 => x"75812a81",
  2764 => x"06537280",
  2765 => x"2e853874",
  2766 => x"8c075575",
  2767 => x"8106407f",
  2768 => x"802e8538",
  2769 => x"74830755",
  2770 => x"74097081",
  2771 => x"ff065253",
  2772 => x"f2993f77",
  2773 => x"14982b70",
  2774 => x"982c5556",
  2775 => x"767424ff",
  2776 => x"9938f7a1",
  2777 => x"39791470",
  2778 => x"337c0770",
  2779 => x"097081ff",
  2780 => x"06545541",
  2781 => x"56f1f43f",
  2782 => x"7714982b",
  2783 => x"70982c55",
  2784 => x"59737725",
  2785 => x"f6ff3879",
  2786 => x"1470337c",
  2787 => x"07700970",
  2788 => x"81ff0654",
  2789 => x"554156f1",
  2790 => x"d23f7714",
  2791 => x"982b7098",
  2792 => x"2c555976",
  2793 => x"7424ffbd",
  2794 => x"38f6da39",
  2795 => x"61802e80",
  2796 => x"f9387d80",
  2797 => x"2e81e838",
  2798 => x"79147033",
  2799 => x"7c077052",
  2800 => x"54568055",
  2801 => x"78752e85",
  2802 => x"3872842a",
  2803 => x"5675832a",
  2804 => x"81065372",
  2805 => x"802e8438",
  2806 => x"81c05575",
  2807 => x"822a8106",
  2808 => x"5372802e",
  2809 => x"853874b0",
  2810 => x"07557581",
  2811 => x"2a810653",
  2812 => x"72802e85",
  2813 => x"38748c07",
  2814 => x"55758106",
  2815 => x"407f802e",
  2816 => x"85387483",
  2817 => x"07557409",
  2818 => x"7081ff06",
  2819 => x"70535456",
  2820 => x"f0d93f72",
  2821 => x"51f0d43f",
  2822 => x"7714982b",
  2823 => x"70982c55",
  2824 => x"40767424",
  2825 => x"ff9238f5",
  2826 => x"dc397d80",
  2827 => x"2e81c538",
  2828 => x"79147033",
  2829 => x"7c077052",
  2830 => x"54568055",
  2831 => x"78752e85",
  2832 => x"3872842a",
  2833 => x"5675832a",
  2834 => x"81065372",
  2835 => x"802e8438",
  2836 => x"81c05575",
  2837 => x"822a8106",
  2838 => x"5372802e",
  2839 => x"853874b0",
  2840 => x"07557581",
  2841 => x"2a810653",
  2842 => x"72802e85",
  2843 => x"38748c07",
  2844 => x"55758106",
  2845 => x"407f802e",
  2846 => x"85387483",
  2847 => x"07557481",
  2848 => x"ff067052",
  2849 => x"53efe43f",
  2850 => x"7251efdf",
  2851 => x"3f771498",
  2852 => x"2b70982c",
  2853 => x"55567674",
  2854 => x"24ff9538",
  2855 => x"f4e73979",
  2856 => x"1470337c",
  2857 => x"07700970",
  2858 => x"81ff0670",
  2859 => x"55564256",
  2860 => x"59efb83f",
  2861 => x"7251efb3",
  2862 => x"3f771498",
  2863 => x"2b70982c",
  2864 => x"55597377",
  2865 => x"25f4be38",
  2866 => x"79147033",
  2867 => x"7c077009",
  2868 => x"7081ff06",
  2869 => x"70555642",
  2870 => x"5659ef8f",
  2871 => x"3f7251ef",
  2872 => x"8a3f7714",
  2873 => x"982b7098",
  2874 => x"2c555976",
  2875 => x"7424ffaf",
  2876 => x"38f49239",
  2877 => x"79147033",
  2878 => x"7c077053",
  2879 => x"5455eeeb",
  2880 => x"3f7251ee",
  2881 => x"e63f7714",
  2882 => x"982b7098",
  2883 => x"2c555973",
  2884 => x"7725f3f1",
  2885 => x"38791470",
  2886 => x"337c0770",
  2887 => x"535455ee",
  2888 => x"ca3f7251",
  2889 => x"eec53f77",
  2890 => x"14982b70",
  2891 => x"982c5559",
  2892 => x"767424c0",
  2893 => x"38f3ce39",
  2894 => x"81abf033",
  2895 => x"7f055680",
  2896 => x"527581ff",
  2897 => x"0651ed9d",
  2898 => x"3f80537c",
  2899 => x"a02ef3f6",
  2900 => x"387f7829",
  2901 => x"64305e57",
  2902 => x"f2a039f8",
  2903 => x"3d0d7a7d",
  2904 => x"028805af",
  2905 => x"05335a55",
  2906 => x"59807470",
  2907 => x"81055633",
  2908 => x"75585657",
  2909 => x"74772e09",
  2910 => x"81068838",
  2911 => x"76b00c8a",
  2912 => x"3d0d0474",
  2913 => x"53775278",
  2914 => x"51efdf3f",
  2915 => x"b00881ff",
  2916 => x"06770570",
  2917 => x"83ffff06",
  2918 => x"77708105",
  2919 => x"59335258",
  2920 => x"5574802e",
  2921 => x"d7387453",
  2922 => x"77527851",
  2923 => x"efbc3fb0",
  2924 => x"0881ff06",
  2925 => x"77057083",
  2926 => x"ffff0677",
  2927 => x"70810559",
  2928 => x"33525855",
  2929 => x"74ffbc38",
  2930 => x"ffb239d0",
  2931 => x"db3f04fb",
  2932 => x"3d0d7779",
  2933 => x"55558056",
  2934 => x"757524ab",
  2935 => x"38807424",
  2936 => x"9d388053",
  2937 => x"73527451",
  2938 => x"80e13fb0",
  2939 => x"08547580",
  2940 => x"2e8538b0",
  2941 => x"08305473",
  2942 => x"b00c873d",
  2943 => x"0d047330",
  2944 => x"76813257",
  2945 => x"54dc3974",
  2946 => x"30558156",
  2947 => x"738025d2",
  2948 => x"38ec39fa",
  2949 => x"3d0d787a",
  2950 => x"57558057",
  2951 => x"767524a4",
  2952 => x"38759f2c",
  2953 => x"54815375",
  2954 => x"74327431",
  2955 => x"5274519b",
  2956 => x"3fb00854",
  2957 => x"76802e85",
  2958 => x"38b00830",
  2959 => x"5473b00c",
  2960 => x"883d0d04",
  2961 => x"74305581",
  2962 => x"57d739fc",
  2963 => x"3d0d7678",
  2964 => x"53548153",
  2965 => x"80747326",
  2966 => x"52557280",
  2967 => x"2e983870",
  2968 => x"802ea938",
  2969 => x"807224a4",
  2970 => x"38711073",
  2971 => x"10757226",
  2972 => x"53545272",
  2973 => x"ea387351",
  2974 => x"78833874",
  2975 => x"5170b00c",
  2976 => x"863d0d04",
  2977 => x"72812a72",
  2978 => x"812a5353",
  2979 => x"72802ee6",
  2980 => x"38717426",
  2981 => x"ef387372",
  2982 => x"31757407",
  2983 => x"74812a74",
  2984 => x"812a5555",
  2985 => x"5654e539",
  2986 => x"10101010",
  2987 => x"10101010",
  2988 => x"10101010",
  2989 => x"10101010",
  2990 => x"10101010",
  2991 => x"10101010",
  2992 => x"10101010",
  2993 => x"10101053",
  2994 => x"51047381",
  2995 => x"ff067383",
  2996 => x"06098105",
  2997 => x"83051010",
  2998 => x"102b0772",
  2999 => x"fc060c51",
  3000 => x"51043c04",
  3001 => x"72728072",
  3002 => x"8106ff05",
  3003 => x"09720605",
  3004 => x"71105272",
  3005 => x"0a100a53",
  3006 => x"72ed3851",
  3007 => x"51535104",
  3008 => x"b008b408",
  3009 => x"b8087575",
  3010 => x"80dc932d",
  3011 => x"5050b008",
  3012 => x"56b80cb4",
  3013 => x"0cb00c51",
  3014 => x"04b008b4",
  3015 => x"08b80875",
  3016 => x"7580dbcf",
  3017 => x"2d5050b0",
  3018 => x"0856b80c",
  3019 => x"b40cb00c",
  3020 => x"5104b008",
  3021 => x"b408b808",
  3022 => x"8187eb2d",
  3023 => x"b80cb40c",
  3024 => x"b00c04ff",
  3025 => x"3d0d028f",
  3026 => x"053381ac",
  3027 => x"a8085271",
  3028 => x"0c800bb0",
  3029 => x"0c833d0d",
  3030 => x"04ff3d0d",
  3031 => x"028f0533",
  3032 => x"5181cf98",
  3033 => x"0852712d",
  3034 => x"b00881ff",
  3035 => x"06b00c83",
  3036 => x"3d0d04fe",
  3037 => x"3d0d7470",
  3038 => x"33535371",
  3039 => x"802e9338",
  3040 => x"81137252",
  3041 => x"81cf9808",
  3042 => x"5353712d",
  3043 => x"72335271",
  3044 => x"ef38843d",
  3045 => x"0d04f43d",
  3046 => x"0d7f0284",
  3047 => x"05bb0533",
  3048 => x"5557880b",
  3049 => x"8c3d5b59",
  3050 => x"895381a9",
  3051 => x"c8527951",
  3052 => x"86e43f73",
  3053 => x"792e80ff",
  3054 => x"38785673",
  3055 => x"902e80ec",
  3056 => x"3802a705",
  3057 => x"58768f06",
  3058 => x"54738926",
  3059 => x"80c23875",
  3060 => x"18b01555",
  3061 => x"55737534",
  3062 => x"76842aff",
  3063 => x"177081ff",
  3064 => x"06585557",
  3065 => x"75df3878",
  3066 => x"1a557575",
  3067 => x"34797033",
  3068 => x"55557380",
  3069 => x"2e933881",
  3070 => x"15745281",
  3071 => x"cf980857",
  3072 => x"55752d74",
  3073 => x"335473ef",
  3074 => x"3878b00c",
  3075 => x"8e3d0d04",
  3076 => x"7518b715",
  3077 => x"55557375",
  3078 => x"3476842a",
  3079 => x"ff177081",
  3080 => x"ff065855",
  3081 => x"5775ff9d",
  3082 => x"38ffbc39",
  3083 => x"84705759",
  3084 => x"02a70558",
  3085 => x"ff8f3982",
  3086 => x"705759f4",
  3087 => x"39f13d0d",
  3088 => x"618d3d70",
  3089 => x"5b5c5a80",
  3090 => x"7a565776",
  3091 => x"7a248185",
  3092 => x"38781754",
  3093 => x"8a527451",
  3094 => x"858a3fb0",
  3095 => x"08b00553",
  3096 => x"72743481",
  3097 => x"17578a52",
  3098 => x"745184d3",
  3099 => x"3fb00855",
  3100 => x"b008de38",
  3101 => x"b008779f",
  3102 => x"2a187081",
  3103 => x"2c5a5656",
  3104 => x"8078259e",
  3105 => x"387817ff",
  3106 => x"05557519",
  3107 => x"70335553",
  3108 => x"74337334",
  3109 => x"73753481",
  3110 => x"16ff1656",
  3111 => x"56777624",
  3112 => x"e9387619",
  3113 => x"58807834",
  3114 => x"807a2417",
  3115 => x"7081ff06",
  3116 => x"7c703356",
  3117 => x"57555672",
  3118 => x"802e9338",
  3119 => x"81157352",
  3120 => x"81cf9808",
  3121 => x"5855762d",
  3122 => x"74335372",
  3123 => x"ef3873b0",
  3124 => x"0c913d0d",
  3125 => x"04ad7b34",
  3126 => x"02ad057a",
  3127 => x"30711956",
  3128 => x"56598a52",
  3129 => x"745183fc",
  3130 => x"3fb008b0",
  3131 => x"05537274",
  3132 => x"34811757",
  3133 => x"8a527451",
  3134 => x"83c53fb0",
  3135 => x"0855b008",
  3136 => x"fecf38fe",
  3137 => x"ef39fd3d",
  3138 => x"0d81ac9c",
  3139 => x"0876b2e4",
  3140 => x"2994120c",
  3141 => x"54850b98",
  3142 => x"150c9814",
  3143 => x"08708106",
  3144 => x"515372f6",
  3145 => x"38853d0d",
  3146 => x"04803d0d",
  3147 => x"81ac9c08",
  3148 => x"51870b84",
  3149 => x"120cff0b",
  3150 => x"b4120ca7",
  3151 => x"0bb8120c",
  3152 => x"87e80ba4",
  3153 => x"120ca70b",
  3154 => x"a8120cb2",
  3155 => x"e40b9412",
  3156 => x"0c870b98",
  3157 => x"120c823d",
  3158 => x"0d04803d",
  3159 => x"0d81aca0",
  3160 => x"0851b80b",
  3161 => x"8c120c83",
  3162 => x"0b88120c",
  3163 => x"823d0d04",
  3164 => x"803d0d81",
  3165 => x"aca00884",
  3166 => x"11088106",
  3167 => x"b00c5182",
  3168 => x"3d0d04ff",
  3169 => x"3d0d81ac",
  3170 => x"a0085284",
  3171 => x"12087081",
  3172 => x"06515170",
  3173 => x"802ef438",
  3174 => x"71087081",
  3175 => x"ff06b00c",
  3176 => x"51833d0d",
  3177 => x"04fe3d0d",
  3178 => x"02930533",
  3179 => x"81aca008",
  3180 => x"53538412",
  3181 => x"0870892a",
  3182 => x"70810651",
  3183 => x"515170f2",
  3184 => x"3872720c",
  3185 => x"843d0d04",
  3186 => x"fe3d0d02",
  3187 => x"93053353",
  3188 => x"728a2e9c",
  3189 => x"3881aca0",
  3190 => x"08528412",
  3191 => x"0870892a",
  3192 => x"70810651",
  3193 => x"515170f2",
  3194 => x"3872720c",
  3195 => x"843d0d04",
  3196 => x"81aca008",
  3197 => x"52841208",
  3198 => x"70892a70",
  3199 => x"81065151",
  3200 => x"5170f238",
  3201 => x"8d720c84",
  3202 => x"12087089",
  3203 => x"2a708106",
  3204 => x"51515170",
  3205 => x"c538d239",
  3206 => x"803d0d81",
  3207 => x"ac940851",
  3208 => x"800b8412",
  3209 => x"0c83fe80",
  3210 => x"0b88120c",
  3211 => x"800b81cf",
  3212 => x"9c34800b",
  3213 => x"81cfa034",
  3214 => x"823d0d04",
  3215 => x"fa3d0d02",
  3216 => x"a3053381",
  3217 => x"ac940881",
  3218 => x"cf9c3370",
  3219 => x"81ff0670",
  3220 => x"10101181",
  3221 => x"cfa03370",
  3222 => x"81ff0672",
  3223 => x"90291170",
  3224 => x"882b7807",
  3225 => x"770c535b",
  3226 => x"5b555559",
  3227 => x"5454738a",
  3228 => x"2e983874",
  3229 => x"80cf2e92",
  3230 => x"38738c2e",
  3231 => x"a4388116",
  3232 => x"537281cf",
  3233 => x"a034883d",
  3234 => x"0d0471a3",
  3235 => x"26a33881",
  3236 => x"17527181",
  3237 => x"cf9c3480",
  3238 => x"0b81cfa0",
  3239 => x"34883d0d",
  3240 => x"04805271",
  3241 => x"882b730c",
  3242 => x"81125297",
  3243 => x"907226f3",
  3244 => x"38800b81",
  3245 => x"cf9c3480",
  3246 => x"0b81cfa0",
  3247 => x"34df39bc",
  3248 => x"0802bc0c",
  3249 => x"fd3d0d80",
  3250 => x"53bc088c",
  3251 => x"050852bc",
  3252 => x"08880508",
  3253 => x"51f6f43f",
  3254 => x"b00870b0",
  3255 => x"0c54853d",
  3256 => x"0dbc0c04",
  3257 => x"bc0802bc",
  3258 => x"0cfd3d0d",
  3259 => x"8153bc08",
  3260 => x"8c050852",
  3261 => x"bc088805",
  3262 => x"0851f6cf",
  3263 => x"3fb00870",
  3264 => x"b00c5485",
  3265 => x"3d0dbc0c",
  3266 => x"04803d0d",
  3267 => x"86518496",
  3268 => x"3f8151a1",
  3269 => x"d33ffc3d",
  3270 => x"0d767079",
  3271 => x"7b555555",
  3272 => x"558f7227",
  3273 => x"8c387275",
  3274 => x"07830651",
  3275 => x"70802ea7",
  3276 => x"38ff1252",
  3277 => x"71ff2e98",
  3278 => x"38727081",
  3279 => x"05543374",
  3280 => x"70810556",
  3281 => x"34ff1252",
  3282 => x"71ff2e09",
  3283 => x"8106ea38",
  3284 => x"74b00c86",
  3285 => x"3d0d0474",
  3286 => x"51727084",
  3287 => x"05540871",
  3288 => x"70840553",
  3289 => x"0c727084",
  3290 => x"05540871",
  3291 => x"70840553",
  3292 => x"0c727084",
  3293 => x"05540871",
  3294 => x"70840553",
  3295 => x"0c727084",
  3296 => x"05540871",
  3297 => x"70840553",
  3298 => x"0cf01252",
  3299 => x"718f26c9",
  3300 => x"38837227",
  3301 => x"95387270",
  3302 => x"84055408",
  3303 => x"71708405",
  3304 => x"530cfc12",
  3305 => x"52718326",
  3306 => x"ed387054",
  3307 => x"ff8339fd",
  3308 => x"3d0d7553",
  3309 => x"84d81308",
  3310 => x"802e8a38",
  3311 => x"805372b0",
  3312 => x"0c853d0d",
  3313 => x"04818052",
  3314 => x"72518d9b",
  3315 => x"3fb00884",
  3316 => x"d8140cff",
  3317 => x"53b00880",
  3318 => x"2ee438b0",
  3319 => x"08549f53",
  3320 => x"80747084",
  3321 => x"05560cff",
  3322 => x"13538073",
  3323 => x"24ce3880",
  3324 => x"74708405",
  3325 => x"560cff13",
  3326 => x"53728025",
  3327 => x"e338ffbc",
  3328 => x"39fd3d0d",
  3329 => x"75775553",
  3330 => x"9f74278d",
  3331 => x"3896730c",
  3332 => x"ff5271b0",
  3333 => x"0c853d0d",
  3334 => x"0484d813",
  3335 => x"08527180",
  3336 => x"2e933873",
  3337 => x"10101270",
  3338 => x"0879720c",
  3339 => x"515271b0",
  3340 => x"0c853d0d",
  3341 => x"047251fe",
  3342 => x"f63fff52",
  3343 => x"b008d338",
  3344 => x"84d81308",
  3345 => x"74101011",
  3346 => x"70087a72",
  3347 => x"0c515152",
  3348 => x"dd39f93d",
  3349 => x"0d797b58",
  3350 => x"56769f26",
  3351 => x"80e83884",
  3352 => x"d8160854",
  3353 => x"73802eaa",
  3354 => x"38761010",
  3355 => x"14700855",
  3356 => x"5573802e",
  3357 => x"ba388058",
  3358 => x"73812e8f",
  3359 => x"3873ff2e",
  3360 => x"a3388075",
  3361 => x"0c765173",
  3362 => x"2d805877",
  3363 => x"b00c893d",
  3364 => x"0d047551",
  3365 => x"fe993fff",
  3366 => x"58b008ef",
  3367 => x"3884d816",
  3368 => x"0854c639",
  3369 => x"96760c81",
  3370 => x"0bb00c89",
  3371 => x"3d0d0475",
  3372 => x"5181ed3f",
  3373 => x"7653b008",
  3374 => x"52755181",
  3375 => x"ad3fb008",
  3376 => x"b00c893d",
  3377 => x"0d049676",
  3378 => x"0cff0bb0",
  3379 => x"0c893d0d",
  3380 => x"04fc3d0d",
  3381 => x"76785653",
  3382 => x"ff54749f",
  3383 => x"26b13884",
  3384 => x"d8130852",
  3385 => x"71802eae",
  3386 => x"38741010",
  3387 => x"12700853",
  3388 => x"53815471",
  3389 => x"802e9838",
  3390 => x"825471ff",
  3391 => x"2e913883",
  3392 => x"5471812e",
  3393 => x"8a388073",
  3394 => x"0c745171",
  3395 => x"2d805473",
  3396 => x"b00c863d",
  3397 => x"0d047251",
  3398 => x"fd953fb0",
  3399 => x"08f13884",
  3400 => x"d8130852",
  3401 => x"c439ff3d",
  3402 => x"0d735281",
  3403 => x"acac0851",
  3404 => x"fea03f83",
  3405 => x"3d0d04fe",
  3406 => x"3d0d7553",
  3407 => x"745281ac",
  3408 => x"ac0851fd",
  3409 => x"bc3f843d",
  3410 => x"0d04803d",
  3411 => x"0d81acac",
  3412 => x"0851fcdb",
  3413 => x"3f823d0d",
  3414 => x"04ff3d0d",
  3415 => x"735281ac",
  3416 => x"ac0851fe",
  3417 => x"ec3f833d",
  3418 => x"0d04fc3d",
  3419 => x"0d800b81",
  3420 => x"cfa80c78",
  3421 => x"5277519c",
  3422 => x"aa3fb008",
  3423 => x"54b008ff",
  3424 => x"2e883873",
  3425 => x"b00c863d",
  3426 => x"0d0481cf",
  3427 => x"a8085574",
  3428 => x"802ef038",
  3429 => x"7675710c",
  3430 => x"5373b00c",
  3431 => x"863d0d04",
  3432 => x"9bfc3f04",
  3433 => x"fc3d0d76",
  3434 => x"70797073",
  3435 => x"07830654",
  3436 => x"54545570",
  3437 => x"80c33871",
  3438 => x"70087009",
  3439 => x"70f7fbfd",
  3440 => x"ff130670",
  3441 => x"f8848281",
  3442 => x"80065151",
  3443 => x"53535470",
  3444 => x"a6388414",
  3445 => x"72747084",
  3446 => x"05560c70",
  3447 => x"08700970",
  3448 => x"f7fbfdff",
  3449 => x"130670f8",
  3450 => x"84828180",
  3451 => x"06515153",
  3452 => x"53547080",
  3453 => x"2edc3873",
  3454 => x"52717081",
  3455 => x"05533351",
  3456 => x"70737081",
  3457 => x"05553470",
  3458 => x"f03874b0",
  3459 => x"0c863d0d",
  3460 => x"04fd3d0d",
  3461 => x"75707183",
  3462 => x"06535552",
  3463 => x"70b83871",
  3464 => x"70087009",
  3465 => x"f7fbfdff",
  3466 => x"120670f8",
  3467 => x"84828180",
  3468 => x"06515152",
  3469 => x"53709d38",
  3470 => x"84137008",
  3471 => x"7009f7fb",
  3472 => x"fdff1206",
  3473 => x"70f88482",
  3474 => x"81800651",
  3475 => x"51525370",
  3476 => x"802ee538",
  3477 => x"72527133",
  3478 => x"5170802e",
  3479 => x"8a388112",
  3480 => x"70335252",
  3481 => x"70f83871",
  3482 => x"7431b00c",
  3483 => x"853d0d04",
  3484 => x"fa3d0d78",
  3485 => x"7a7c7054",
  3486 => x"55555272",
  3487 => x"802e80d9",
  3488 => x"38717407",
  3489 => x"83065170",
  3490 => x"802e80d4",
  3491 => x"38ff1353",
  3492 => x"72ff2eb1",
  3493 => x"38713374",
  3494 => x"33565174",
  3495 => x"712e0981",
  3496 => x"06a93872",
  3497 => x"802e8187",
  3498 => x"387081ff",
  3499 => x"06517080",
  3500 => x"2e80fc38",
  3501 => x"81128115",
  3502 => x"ff155555",
  3503 => x"5272ff2e",
  3504 => x"098106d1",
  3505 => x"38713374",
  3506 => x"33565170",
  3507 => x"81ff0675",
  3508 => x"81ff0671",
  3509 => x"71315152",
  3510 => x"5270b00c",
  3511 => x"883d0d04",
  3512 => x"71745755",
  3513 => x"83732788",
  3514 => x"38710874",
  3515 => x"082e8838",
  3516 => x"74765552",
  3517 => x"ff9739fc",
  3518 => x"13537280",
  3519 => x"2eb13874",
  3520 => x"087009f7",
  3521 => x"fbfdff12",
  3522 => x"0670f884",
  3523 => x"82818006",
  3524 => x"51515170",
  3525 => x"9a388415",
  3526 => x"84175755",
  3527 => x"837327d0",
  3528 => x"38740876",
  3529 => x"082ed038",
  3530 => x"74765552",
  3531 => x"fedf3980",
  3532 => x"0bb00c88",
  3533 => x"3d0d04f3",
  3534 => x"3d0d6062",
  3535 => x"64725a5a",
  3536 => x"5e5e805c",
  3537 => x"76708105",
  3538 => x"583381a9",
  3539 => x"d5113370",
  3540 => x"832a7081",
  3541 => x"06515555",
  3542 => x"5672e938",
  3543 => x"75ad2e82",
  3544 => x"883875ab",
  3545 => x"2e828438",
  3546 => x"77307079",
  3547 => x"07802579",
  3548 => x"90327030",
  3549 => x"70720780",
  3550 => x"25730753",
  3551 => x"57575153",
  3552 => x"72802e87",
  3553 => x"3875b02e",
  3554 => x"81eb3877",
  3555 => x"8a388858",
  3556 => x"75b02e83",
  3557 => x"388a5881",
  3558 => x"0a5a7b84",
  3559 => x"38fe0a5a",
  3560 => x"77527951",
  3561 => x"f6be3fb0",
  3562 => x"0878537a",
  3563 => x"525bf68f",
  3564 => x"3fb0085a",
  3565 => x"807081a9",
  3566 => x"d5183370",
  3567 => x"822a7081",
  3568 => x"06515656",
  3569 => x"5a557280",
  3570 => x"2e80c138",
  3571 => x"d0165675",
  3572 => x"782580d7",
  3573 => x"38807924",
  3574 => x"757b2607",
  3575 => x"53729338",
  3576 => x"747a2e80",
  3577 => x"eb387a76",
  3578 => x"2580ed38",
  3579 => x"72802e80",
  3580 => x"e738ff77",
  3581 => x"70810559",
  3582 => x"33575981",
  3583 => x"a9d51633",
  3584 => x"70822a70",
  3585 => x"81065154",
  3586 => x"5472c138",
  3587 => x"73830653",
  3588 => x"72802e97",
  3589 => x"38738106",
  3590 => x"c9175553",
  3591 => x"728538ff",
  3592 => x"a9165473",
  3593 => x"56777624",
  3594 => x"ffab3880",
  3595 => x"792480f0",
  3596 => x"387b802e",
  3597 => x"84387430",
  3598 => x"557c802e",
  3599 => x"8c38ff17",
  3600 => x"53788338",
  3601 => x"7d53727d",
  3602 => x"0c74b00c",
  3603 => x"8f3d0d04",
  3604 => x"8153757b",
  3605 => x"24ff9538",
  3606 => x"81757929",
  3607 => x"17787081",
  3608 => x"055a3358",
  3609 => x"5659ff93",
  3610 => x"39815c76",
  3611 => x"70810558",
  3612 => x"3356fdf4",
  3613 => x"39807733",
  3614 => x"54547280",
  3615 => x"f82eb238",
  3616 => x"7280d832",
  3617 => x"70307080",
  3618 => x"25760751",
  3619 => x"51537280",
  3620 => x"2efdf838",
  3621 => x"81173382",
  3622 => x"18585690",
  3623 => x"58fdf839",
  3624 => x"810a557b",
  3625 => x"8438fe0a",
  3626 => x"557f53a2",
  3627 => x"730cff89",
  3628 => x"398154cc",
  3629 => x"39fd3d0d",
  3630 => x"77547653",
  3631 => x"755281ac",
  3632 => x"ac0851fc",
  3633 => x"f23f853d",
  3634 => x"0d04f33d",
  3635 => x"0d606264",
  3636 => x"725a5a5d",
  3637 => x"5d805e76",
  3638 => x"70810558",
  3639 => x"3381a9d5",
  3640 => x"11337083",
  3641 => x"2a708106",
  3642 => x"51555556",
  3643 => x"72e93875",
  3644 => x"ad2e81ff",
  3645 => x"3875ab2e",
  3646 => x"81fb3877",
  3647 => x"30707907",
  3648 => x"80257990",
  3649 => x"32703070",
  3650 => x"72078025",
  3651 => x"73075357",
  3652 => x"57515372",
  3653 => x"802e8738",
  3654 => x"75b02e81",
  3655 => x"e238778a",
  3656 => x"38885875",
  3657 => x"b02e8338",
  3658 => x"8a587752",
  3659 => x"ff51f38f",
  3660 => x"3fb00878",
  3661 => x"535aff51",
  3662 => x"f3aa3fb0",
  3663 => x"085b8070",
  3664 => x"5a5581a9",
  3665 => x"d5163370",
  3666 => x"822a7081",
  3667 => x"06515454",
  3668 => x"72802e80",
  3669 => x"c138d016",
  3670 => x"56757825",
  3671 => x"80d73880",
  3672 => x"7924757b",
  3673 => x"26075372",
  3674 => x"9338747a",
  3675 => x"2e80eb38",
  3676 => x"7a762580",
  3677 => x"ed387280",
  3678 => x"2e80e738",
  3679 => x"ff777081",
  3680 => x"05593357",
  3681 => x"5981a9d5",
  3682 => x"16337082",
  3683 => x"2a708106",
  3684 => x"51545472",
  3685 => x"c1387383",
  3686 => x"06537280",
  3687 => x"2e973873",
  3688 => x"8106c917",
  3689 => x"55537285",
  3690 => x"38ffa916",
  3691 => x"54735677",
  3692 => x"7624ffab",
  3693 => x"38807924",
  3694 => x"8189387d",
  3695 => x"802e8438",
  3696 => x"7430557b",
  3697 => x"802e8c38",
  3698 => x"ff175378",
  3699 => x"83387c53",
  3700 => x"727c0c74",
  3701 => x"b00c8f3d",
  3702 => x"0d048153",
  3703 => x"757b24ff",
  3704 => x"95388175",
  3705 => x"79291778",
  3706 => x"7081055a",
  3707 => x"33585659",
  3708 => x"ff933981",
  3709 => x"5e767081",
  3710 => x"05583356",
  3711 => x"fdfd3980",
  3712 => x"77335454",
  3713 => x"7280f82e",
  3714 => x"80c33872",
  3715 => x"80d83270",
  3716 => x"30708025",
  3717 => x"76075151",
  3718 => x"5372802e",
  3719 => x"fe803881",
  3720 => x"17338218",
  3721 => x"58569070",
  3722 => x"5358ff51",
  3723 => x"f1913fb0",
  3724 => x"0878535a",
  3725 => x"ff51f1ac",
  3726 => x"3fb0085b",
  3727 => x"80705a55",
  3728 => x"fe8039ff",
  3729 => x"605455a2",
  3730 => x"730cfef7",
  3731 => x"398154ff",
  3732 => x"ba39fd3d",
  3733 => x"0d775476",
  3734 => x"53755281",
  3735 => x"acac0851",
  3736 => x"fce83f85",
  3737 => x"3d0d04f3",
  3738 => x"3d0d7f61",
  3739 => x"8b1170f8",
  3740 => x"065c5555",
  3741 => x"5e729626",
  3742 => x"83389059",
  3743 => x"80792474",
  3744 => x"7a260753",
  3745 => x"80547274",
  3746 => x"2e098106",
  3747 => x"80cb387d",
  3748 => x"518bca3f",
  3749 => x"7883f726",
  3750 => x"80c63878",
  3751 => x"832a7010",
  3752 => x"101081b3",
  3753 => x"e8058c11",
  3754 => x"0859595a",
  3755 => x"76782e83",
  3756 => x"b0388417",
  3757 => x"08fc0656",
  3758 => x"8c170888",
  3759 => x"1808718c",
  3760 => x"120c8812",
  3761 => x"0c587517",
  3762 => x"84110881",
  3763 => x"0784120c",
  3764 => x"537d518b",
  3765 => x"893f8817",
  3766 => x"5473b00c",
  3767 => x"8f3d0d04",
  3768 => x"78892a79",
  3769 => x"832a5b53",
  3770 => x"72802ebf",
  3771 => x"3878862a",
  3772 => x"b8055a84",
  3773 => x"7327b438",
  3774 => x"80db135a",
  3775 => x"947327ab",
  3776 => x"38788c2a",
  3777 => x"80ee055a",
  3778 => x"80d47327",
  3779 => x"9e38788f",
  3780 => x"2a80f705",
  3781 => x"5a82d473",
  3782 => x"27913878",
  3783 => x"922a80fc",
  3784 => x"055a8ad4",
  3785 => x"73278438",
  3786 => x"80fe5a79",
  3787 => x"10101081",
  3788 => x"b3e8058c",
  3789 => x"11085855",
  3790 => x"76752ea3",
  3791 => x"38841708",
  3792 => x"fc06707a",
  3793 => x"31555673",
  3794 => x"8f2488d5",
  3795 => x"38738025",
  3796 => x"fee6388c",
  3797 => x"17085776",
  3798 => x"752e0981",
  3799 => x"06df3881",
  3800 => x"1a5a81b3",
  3801 => x"f8085776",
  3802 => x"81b3f02e",
  3803 => x"82c03884",
  3804 => x"1708fc06",
  3805 => x"707a3155",
  3806 => x"56738f24",
  3807 => x"81f93881",
  3808 => x"b3f00b81",
  3809 => x"b3fc0c81",
  3810 => x"b3f00b81",
  3811 => x"b3f80c73",
  3812 => x"8025feb2",
  3813 => x"3883ff76",
  3814 => x"2783df38",
  3815 => x"75892a76",
  3816 => x"832a5553",
  3817 => x"72802ebf",
  3818 => x"3875862a",
  3819 => x"b8055484",
  3820 => x"7327b438",
  3821 => x"80db1354",
  3822 => x"947327ab",
  3823 => x"38758c2a",
  3824 => x"80ee0554",
  3825 => x"80d47327",
  3826 => x"9e38758f",
  3827 => x"2a80f705",
  3828 => x"5482d473",
  3829 => x"27913875",
  3830 => x"922a80fc",
  3831 => x"05548ad4",
  3832 => x"73278438",
  3833 => x"80fe5473",
  3834 => x"10101081",
  3835 => x"b3e80588",
  3836 => x"11085658",
  3837 => x"74782e86",
  3838 => x"cf388415",
  3839 => x"08fc0653",
  3840 => x"7573278d",
  3841 => x"38881508",
  3842 => x"5574782e",
  3843 => x"098106ea",
  3844 => x"388c1508",
  3845 => x"81b3e80b",
  3846 => x"84050871",
  3847 => x"8c1a0c76",
  3848 => x"881a0c78",
  3849 => x"88130c78",
  3850 => x"8c180c5d",
  3851 => x"58795380",
  3852 => x"7a2483e6",
  3853 => x"3872822c",
  3854 => x"81712b5c",
  3855 => x"537a7c26",
  3856 => x"8198387b",
  3857 => x"7b065372",
  3858 => x"82f13879",
  3859 => x"fc068405",
  3860 => x"5a7a1070",
  3861 => x"7d06545b",
  3862 => x"7282e038",
  3863 => x"841a5af1",
  3864 => x"3988178c",
  3865 => x"11085858",
  3866 => x"76782e09",
  3867 => x"8106fcc2",
  3868 => x"38821a5a",
  3869 => x"fdec3978",
  3870 => x"17798107",
  3871 => x"84190c70",
  3872 => x"81b3fc0c",
  3873 => x"7081b3f8",
  3874 => x"0c81b3f0",
  3875 => x"0b8c120c",
  3876 => x"8c110888",
  3877 => x"120c7481",
  3878 => x"0784120c",
  3879 => x"74117571",
  3880 => x"0c51537d",
  3881 => x"5187b73f",
  3882 => x"881754fc",
  3883 => x"ac3981b3",
  3884 => x"e80b8405",
  3885 => x"087a545c",
  3886 => x"798025fe",
  3887 => x"f83882da",
  3888 => x"397a097c",
  3889 => x"067081b3",
  3890 => x"e80b8405",
  3891 => x"0c5c7a10",
  3892 => x"5b7a7c26",
  3893 => x"85387a85",
  3894 => x"b83881b3",
  3895 => x"e80b8805",
  3896 => x"08708412",
  3897 => x"08fc0670",
  3898 => x"7c317c72",
  3899 => x"268f7225",
  3900 => x"0757575c",
  3901 => x"5d557280",
  3902 => x"2e80db38",
  3903 => x"797a1681",
  3904 => x"b3e0081b",
  3905 => x"90115a55",
  3906 => x"575b81b3",
  3907 => x"dc08ff2e",
  3908 => x"8838a08f",
  3909 => x"13e08006",
  3910 => x"5776527d",
  3911 => x"5186c03f",
  3912 => x"b00854b0",
  3913 => x"08ff2e90",
  3914 => x"38b00876",
  3915 => x"27829938",
  3916 => x"7481b3e8",
  3917 => x"2e829138",
  3918 => x"81b3e80b",
  3919 => x"88050855",
  3920 => x"841508fc",
  3921 => x"06707a31",
  3922 => x"7a72268f",
  3923 => x"72250752",
  3924 => x"55537283",
  3925 => x"e6387479",
  3926 => x"81078417",
  3927 => x"0c791670",
  3928 => x"81b3e80b",
  3929 => x"88050c75",
  3930 => x"81078412",
  3931 => x"0c547e52",
  3932 => x"5785eb3f",
  3933 => x"881754fa",
  3934 => x"e0397583",
  3935 => x"2a705454",
  3936 => x"80742481",
  3937 => x"9b387282",
  3938 => x"2c81712b",
  3939 => x"81b3ec08",
  3940 => x"077081b3",
  3941 => x"e80b8405",
  3942 => x"0c751010",
  3943 => x"1081b3e8",
  3944 => x"05881108",
  3945 => x"585a5d53",
  3946 => x"778c180c",
  3947 => x"7488180c",
  3948 => x"7688190c",
  3949 => x"768c160c",
  3950 => x"fcf33979",
  3951 => x"7a101010",
  3952 => x"81b3e805",
  3953 => x"7057595d",
  3954 => x"8c150857",
  3955 => x"76752ea3",
  3956 => x"38841708",
  3957 => x"fc06707a",
  3958 => x"31555673",
  3959 => x"8f2483ca",
  3960 => x"38738025",
  3961 => x"8481388c",
  3962 => x"17085776",
  3963 => x"752e0981",
  3964 => x"06df3888",
  3965 => x"15811b70",
  3966 => x"8306555b",
  3967 => x"5572c938",
  3968 => x"7c830653",
  3969 => x"72802efd",
  3970 => x"b838ff1d",
  3971 => x"f819595d",
  3972 => x"88180878",
  3973 => x"2eea38fd",
  3974 => x"b539831a",
  3975 => x"53fc9639",
  3976 => x"83147082",
  3977 => x"2c81712b",
  3978 => x"81b3ec08",
  3979 => x"077081b3",
  3980 => x"e80b8405",
  3981 => x"0c761010",
  3982 => x"1081b3e8",
  3983 => x"05881108",
  3984 => x"595b5e51",
  3985 => x"53fee139",
  3986 => x"81b3ac08",
  3987 => x"1758b008",
  3988 => x"762e818d",
  3989 => x"3881b3dc",
  3990 => x"08ff2e83",
  3991 => x"ec387376",
  3992 => x"311881b3",
  3993 => x"ac0c7387",
  3994 => x"06705753",
  3995 => x"72802e88",
  3996 => x"38887331",
  3997 => x"70155556",
  3998 => x"76149fff",
  3999 => x"06a08071",
  4000 => x"31177054",
  4001 => x"7f535753",
  4002 => x"83d53fb0",
  4003 => x"0853b008",
  4004 => x"ff2e81a0",
  4005 => x"3881b3ac",
  4006 => x"08167081",
  4007 => x"b3ac0c74",
  4008 => x"7581b3e8",
  4009 => x"0b88050c",
  4010 => x"74763118",
  4011 => x"70810751",
  4012 => x"5556587b",
  4013 => x"81b3e82e",
  4014 => x"839c3879",
  4015 => x"8f2682cb",
  4016 => x"38810b84",
  4017 => x"150c8415",
  4018 => x"08fc0670",
  4019 => x"7a317a72",
  4020 => x"268f7225",
  4021 => x"07525553",
  4022 => x"72802efc",
  4023 => x"f93880db",
  4024 => x"39b0089f",
  4025 => x"ff065372",
  4026 => x"feeb3877",
  4027 => x"81b3ac0c",
  4028 => x"81b3e80b",
  4029 => x"8805087b",
  4030 => x"18810784",
  4031 => x"120c5581",
  4032 => x"b3d80878",
  4033 => x"27863877",
  4034 => x"81b3d80c",
  4035 => x"81b3d408",
  4036 => x"7827fcac",
  4037 => x"387781b3",
  4038 => x"d40c8415",
  4039 => x"08fc0670",
  4040 => x"7a317a72",
  4041 => x"268f7225",
  4042 => x"07525553",
  4043 => x"72802efc",
  4044 => x"a5388839",
  4045 => x"80745456",
  4046 => x"fedb397d",
  4047 => x"51829f3f",
  4048 => x"800bb00c",
  4049 => x"8f3d0d04",
  4050 => x"73538074",
  4051 => x"24a93872",
  4052 => x"822c8171",
  4053 => x"2b81b3ec",
  4054 => x"08077081",
  4055 => x"b3e80b84",
  4056 => x"050c5d53",
  4057 => x"778c180c",
  4058 => x"7488180c",
  4059 => x"7688190c",
  4060 => x"768c160c",
  4061 => x"f9b73983",
  4062 => x"1470822c",
  4063 => x"81712b81",
  4064 => x"b3ec0807",
  4065 => x"7081b3e8",
  4066 => x"0b84050c",
  4067 => x"5e5153d4",
  4068 => x"397b7b06",
  4069 => x"5372fca3",
  4070 => x"38841a7b",
  4071 => x"105c5af1",
  4072 => x"39ff1a81",
  4073 => x"11515af7",
  4074 => x"b9397817",
  4075 => x"79810784",
  4076 => x"190c8c18",
  4077 => x"08881908",
  4078 => x"718c120c",
  4079 => x"88120c59",
  4080 => x"7081b3fc",
  4081 => x"0c7081b3",
  4082 => x"f80c81b3",
  4083 => x"f00b8c12",
  4084 => x"0c8c1108",
  4085 => x"88120c74",
  4086 => x"81078412",
  4087 => x"0c741175",
  4088 => x"710c5153",
  4089 => x"f9bd3975",
  4090 => x"17841108",
  4091 => x"81078412",
  4092 => x"0c538c17",
  4093 => x"08881808",
  4094 => x"718c120c",
  4095 => x"88120c58",
  4096 => x"7d5180da",
  4097 => x"3f881754",
  4098 => x"f5cf3972",
  4099 => x"84150cf4",
  4100 => x"1af80670",
  4101 => x"841e0881",
  4102 => x"0607841e",
  4103 => x"0c701d54",
  4104 => x"5b850b84",
  4105 => x"140c850b",
  4106 => x"88140c8f",
  4107 => x"7b27fdcf",
  4108 => x"38881c52",
  4109 => x"7d518290",
  4110 => x"3f81b3e8",
  4111 => x"0b880508",
  4112 => x"81b3ac08",
  4113 => x"5955fdb7",
  4114 => x"397781b3",
  4115 => x"ac0c7381",
  4116 => x"b3dc0cfc",
  4117 => x"91397284",
  4118 => x"150cfda3",
  4119 => x"390404fd",
  4120 => x"3d0d800b",
  4121 => x"81cfa80c",
  4122 => x"765186cb",
  4123 => x"3fb00853",
  4124 => x"b008ff2e",
  4125 => x"883872b0",
  4126 => x"0c853d0d",
  4127 => x"0481cfa8",
  4128 => x"08547380",
  4129 => x"2ef03875",
  4130 => x"74710c52",
  4131 => x"72b00c85",
  4132 => x"3d0d04fb",
  4133 => x"3d0d7770",
  4134 => x"5256c23f",
  4135 => x"81b3e80b",
  4136 => x"88050884",
  4137 => x"1108fc06",
  4138 => x"707b319f",
  4139 => x"ef05e080",
  4140 => x"06e08005",
  4141 => x"565653a0",
  4142 => x"80742494",
  4143 => x"38805275",
  4144 => x"51ff9c3f",
  4145 => x"81b3f008",
  4146 => x"155372b0",
  4147 => x"082e8f38",
  4148 => x"7551ff8a",
  4149 => x"3f805372",
  4150 => x"b00c873d",
  4151 => x"0d047330",
  4152 => x"527551fe",
  4153 => x"fa3fb008",
  4154 => x"ff2ea838",
  4155 => x"81b3e80b",
  4156 => x"88050875",
  4157 => x"75318107",
  4158 => x"84120c53",
  4159 => x"81b3ac08",
  4160 => x"743181b3",
  4161 => x"ac0c7551",
  4162 => x"fed43f81",
  4163 => x"0bb00c87",
  4164 => x"3d0d0480",
  4165 => x"527551fe",
  4166 => x"c63f81b3",
  4167 => x"e80b8805",
  4168 => x"08b00871",
  4169 => x"3156538f",
  4170 => x"7525ffa4",
  4171 => x"38b00881",
  4172 => x"b3dc0831",
  4173 => x"81b3ac0c",
  4174 => x"74810784",
  4175 => x"140c7551",
  4176 => x"fe9c3f80",
  4177 => x"53ff9039",
  4178 => x"f63d0d7c",
  4179 => x"7e545b72",
  4180 => x"802e8283",
  4181 => x"387a51fe",
  4182 => x"843ff813",
  4183 => x"84110870",
  4184 => x"fe067013",
  4185 => x"841108fc",
  4186 => x"065d5859",
  4187 => x"545881b3",
  4188 => x"f008752e",
  4189 => x"82de3878",
  4190 => x"84160c80",
  4191 => x"73810654",
  4192 => x"5a727a2e",
  4193 => x"81d53878",
  4194 => x"15841108",
  4195 => x"81065153",
  4196 => x"72a03878",
  4197 => x"17577981",
  4198 => x"e6388815",
  4199 => x"08537281",
  4200 => x"b3f02e82",
  4201 => x"f9388c15",
  4202 => x"08708c15",
  4203 => x"0c738812",
  4204 => x"0c567681",
  4205 => x"0784190c",
  4206 => x"76187771",
  4207 => x"0c537981",
  4208 => x"913883ff",
  4209 => x"772781c8",
  4210 => x"3876892a",
  4211 => x"77832a56",
  4212 => x"5372802e",
  4213 => x"bf387686",
  4214 => x"2ab80555",
  4215 => x"847327b4",
  4216 => x"3880db13",
  4217 => x"55947327",
  4218 => x"ab38768c",
  4219 => x"2a80ee05",
  4220 => x"5580d473",
  4221 => x"279e3876",
  4222 => x"8f2a80f7",
  4223 => x"055582d4",
  4224 => x"73279138",
  4225 => x"76922a80",
  4226 => x"fc05558a",
  4227 => x"d4732784",
  4228 => x"3880fe55",
  4229 => x"74101010",
  4230 => x"81b3e805",
  4231 => x"88110855",
  4232 => x"5673762e",
  4233 => x"82b33884",
  4234 => x"1408fc06",
  4235 => x"53767327",
  4236 => x"8d388814",
  4237 => x"08547376",
  4238 => x"2e098106",
  4239 => x"ea388c14",
  4240 => x"08708c1a",
  4241 => x"0c74881a",
  4242 => x"0c788812",
  4243 => x"0c56778c",
  4244 => x"150c7a51",
  4245 => x"fc883f8c",
  4246 => x"3d0d0477",
  4247 => x"08787131",
  4248 => x"59770588",
  4249 => x"19085457",
  4250 => x"7281b3f0",
  4251 => x"2e80e038",
  4252 => x"8c180870",
  4253 => x"8c150c73",
  4254 => x"88120c56",
  4255 => x"fe893988",
  4256 => x"15088c16",
  4257 => x"08708c13",
  4258 => x"0c578817",
  4259 => x"0cfea339",
  4260 => x"76832a70",
  4261 => x"54558075",
  4262 => x"24819838",
  4263 => x"72822c81",
  4264 => x"712b81b3",
  4265 => x"ec080781",
  4266 => x"b3e80b84",
  4267 => x"050c5374",
  4268 => x"10101081",
  4269 => x"b3e80588",
  4270 => x"11085556",
  4271 => x"758c190c",
  4272 => x"7388190c",
  4273 => x"7788170c",
  4274 => x"778c150c",
  4275 => x"ff843981",
  4276 => x"5afdb439",
  4277 => x"78177381",
  4278 => x"06545772",
  4279 => x"98387708",
  4280 => x"78713159",
  4281 => x"77058c19",
  4282 => x"08881a08",
  4283 => x"718c120c",
  4284 => x"88120c57",
  4285 => x"57768107",
  4286 => x"84190c77",
  4287 => x"81b3e80b",
  4288 => x"88050c81",
  4289 => x"b3e40877",
  4290 => x"26fec738",
  4291 => x"81b3e008",
  4292 => x"527a51fa",
  4293 => x"fe3f7a51",
  4294 => x"fac43ffe",
  4295 => x"ba398178",
  4296 => x"8c150c78",
  4297 => x"88150c73",
  4298 => x"8c1a0c73",
  4299 => x"881a0c5a",
  4300 => x"fd803983",
  4301 => x"1570822c",
  4302 => x"81712b81",
  4303 => x"b3ec0807",
  4304 => x"81b3e80b",
  4305 => x"84050c51",
  4306 => x"53741010",
  4307 => x"1081b3e8",
  4308 => x"05881108",
  4309 => x"5556fee4",
  4310 => x"39745380",
  4311 => x"7524a738",
  4312 => x"72822c81",
  4313 => x"712b81b3",
  4314 => x"ec080781",
  4315 => x"b3e80b84",
  4316 => x"050c5375",
  4317 => x"8c190c73",
  4318 => x"88190c77",
  4319 => x"88170c77",
  4320 => x"8c150cfd",
  4321 => x"cd398315",
  4322 => x"70822c81",
  4323 => x"712b81b3",
  4324 => x"ec080781",
  4325 => x"b3e80b84",
  4326 => x"050c5153",
  4327 => x"d639810b",
  4328 => x"b00c0480",
  4329 => x"3d0d7281",
  4330 => x"2e893880",
  4331 => x"0bb00c82",
  4332 => x"3d0d0473",
  4333 => x"51b23ffe",
  4334 => x"3d0d81cf",
  4335 => x"a4085170",
  4336 => x"8a3881cf",
  4337 => x"ac7081cf",
  4338 => x"a40c5170",
  4339 => x"75125252",
  4340 => x"ff537087",
  4341 => x"fb808026",
  4342 => x"88387081",
  4343 => x"cfa40c71",
  4344 => x"5372b00c",
  4345 => x"843d0d04",
  4346 => x"00ff3900",
  4347 => x"ff390000",
  4348 => x"00000000",
  4349 => x"00000000",
  4350 => x"00000000",
  4351 => x"00000000",
  4352 => x"00cac5ca",
  4353 => x"c5c0c0c0",
  4354 => x"c0c0c0c0",
  4355 => x"c0c0c0cf",
  4356 => x"cfcfcf00",
  4357 => x"00000f0f",
  4358 => x"0f0f8f8f",
  4359 => x"cfcfcfcf",
  4360 => x"cfcf4f0f",
  4361 => x"0f0f0000",
  4362 => x"cfcfcfcf",
  4363 => x"0f0f0f0f",
  4364 => x"0f0f0f0f",
  4365 => x"0f0ffefe",
  4366 => x"fefc0000",
  4367 => x"cfcfcfcf",
  4368 => x"cfcfcfcf",
  4369 => x"cfcfcfcf",
  4370 => x"cfffff7e",
  4371 => x"7e000000",
  4372 => x"00000000",
  4373 => x"00000000",
  4374 => x"00000000",
  4375 => x"00003f3f",
  4376 => x"3f3f0101",
  4377 => x"01010101",
  4378 => x"01010101",
  4379 => x"3f3f3f3f",
  4380 => x"0000383c",
  4381 => x"3e3e3f3f",
  4382 => x"3f3b3b39",
  4383 => x"39383838",
  4384 => x"38383800",
  4385 => x"003f3f3f",
  4386 => x"3f383838",
  4387 => x"38383838",
  4388 => x"38383c3f",
  4389 => x"3f1f0f00",
  4390 => x"003f3f3f",
  4391 => x"3f030303",
  4392 => x"03030303",
  4393 => x"03033f3f",
  4394 => x"3f3e0000",
  4395 => x"00000000",
  4396 => x"00000000",
  4397 => x"00000000",
  4398 => x"00000000",
  4399 => x"00000000",
  4400 => x"00000000",
  4401 => x"00000000",
  4402 => x"00000000",
  4403 => x"00000000",
  4404 => x"00000000",
  4405 => x"00000000",
  4406 => x"00000000",
  4407 => x"00000000",
  4408 => x"00000000",
  4409 => x"00000000",
  4410 => x"00000000",
  4411 => x"00000000",
  4412 => x"00000000",
  4413 => x"00000000",
  4414 => x"00000000",
  4415 => x"00000000",
  4416 => x"00000000",
  4417 => x"00000000",
  4418 => x"00000000",
  4419 => x"8080c0c0",
  4420 => x"e0e06000",
  4421 => x"00000000",
  4422 => x"00000000",
  4423 => x"00000000",
  4424 => x"00000000",
  4425 => x"00000000",
  4426 => x"00000000",
  4427 => x"00000000",
  4428 => x"00000000",
  4429 => x"00000000",
  4430 => x"00000000",
  4431 => x"00000000",
  4432 => x"00000000",
  4433 => x"00000000",
  4434 => x"00000000",
  4435 => x"00000000",
  4436 => x"00000000",
  4437 => x"00000000",
  4438 => x"00000000",
  4439 => x"00000000",
  4440 => x"00000000",
  4441 => x"806098ee",
  4442 => x"77bbddec",
  4443 => x"ee6e0200",
  4444 => x"00000000",
  4445 => x"00e08080",
  4446 => x"e00000e0",
  4447 => x"a0a00000",
  4448 => x"e0000000",
  4449 => x"00e0c000",
  4450 => x"c0e00000",
  4451 => x"e08080e0",
  4452 => x"0000c020",
  4453 => x"20c00000",
  4454 => x"e0000000",
  4455 => x"20e02000",
  4456 => x"0020a060",
  4457 => x"20000000",
  4458 => x"00000000",
  4459 => x"00000000",
  4460 => x"00000000",
  4461 => x"00000000",
  4462 => x"00000000",
  4463 => x"00000000",
  4464 => x"00030007",
  4465 => x"00070701",
  4466 => x"00000000",
  4467 => x"00000000",
  4468 => x"00000300",
  4469 => x"c0030000",
  4470 => x"034242c0",
  4471 => x"00c34242",
  4472 => x"0000c380",
  4473 => x"01c00340",
  4474 => x"c04300c0",
  4475 => x"43408001",
  4476 => x"c20201c0",
  4477 => x"00c38202",
  4478 => x"80c00300",
  4479 => x"00c04342",
  4480 => x"8202c040",
  4481 => x"40800000",
  4482 => x"c0404000",
  4483 => x"80404000",
  4484 => x"00c04040",
  4485 => x"8000c040",
  4486 => x"4000c080",
  4487 => x"00c00000",
  4488 => x"00000000",
  4489 => x"00000000",
  4490 => x"00000000",
  4491 => x"00000000",
  4492 => x"00ff0000",
  4493 => x"0000c645",
  4494 => x"44800785",
  4495 => x"45408007",
  4496 => x"80424700",
  4497 => x"80474000",
  4498 => x"07c14344",
  4499 => x"00c38404",
  4500 => x"c30007c1",
  4501 => x"42418700",
  4502 => x"80404784",
  4503 => x"04c34047",
  4504 => x"8101c640",
  4505 => x"40070505",
  4506 => x"00040502",
  4507 => x"00000704",
  4508 => x"04030007",
  4509 => x"05050007",
  4510 => x"00020700",
  4511 => x"00000000",
  4512 => x"00000000",
  4513 => x"00000000",
  4514 => x"00000000",
  4515 => x"0000ff00",
  4516 => x"00000007",
  4517 => x"01030500",
  4518 => x"03040403",
  4519 => x"00040502",
  4520 => x"00040502",
  4521 => x"00000705",
  4522 => x"05000700",
  4523 => x"02070000",
  4524 => x"07040403",
  4525 => x"00030404",
  4526 => x"03000701",
  4527 => x"03050007",
  4528 => x"01010000",
  4529 => x"00000000",
  4530 => x"00000000",
  4531 => x"00000000",
  4532 => x"00000000",
  4533 => x"00000000",
  4534 => x"71756974",
  4535 => x"00000000",
  4536 => x"68656c70",
  4537 => x"00000000",
  4538 => x"73686f77",
  4539 => x"2042504d",
  4540 => x"20726567",
  4541 => x"69737465",
  4542 => x"72730000",
  4543 => x"62706d00",
  4544 => x"73686f77",
  4545 => x"2f736574",
  4546 => x"20646562",
  4547 => x"75672072",
  4548 => x"65676973",
  4549 => x"74657273",
  4550 => x"203c7365",
  4551 => x"74206d6f",
  4552 => x"64653e00",
  4553 => x"64656275",
  4554 => x"67000000",
  4555 => x"73797374",
  4556 => x"656d2072",
  4557 => x"65736574",
  4558 => x"00000000",
  4559 => x"72657365",
  4560 => x"74000000",
  4561 => x"73686f77",
  4562 => x"20646562",
  4563 => x"75672062",
  4564 => x"75666665",
  4565 => x"72203c6c",
  4566 => x"656e6774",
  4567 => x"683e0000",
  4568 => x"646f776e",
  4569 => x"6c6f6164",
  4570 => x"20646562",
  4571 => x"75672062",
  4572 => x"75666665",
  4573 => x"72202878",
  4574 => x"6d6f6465",
  4575 => x"6d290000",
  4576 => x"62726561",
  4577 => x"64000000",
  4578 => x"75706c6f",
  4579 => x"61642064",
  4580 => x"65627567",
  4581 => x"20627566",
  4582 => x"66657220",
  4583 => x"28786d6f",
  4584 => x"64656d29",
  4585 => x"00000000",
  4586 => x"62777269",
  4587 => x"74650000",
  4588 => x"636c6561",
  4589 => x"72206465",
  4590 => x"62756720",
  4591 => x"62756666",
  4592 => x"65720000",
  4593 => x"62636c65",
  4594 => x"61720000",
  4595 => x"73657475",
  4596 => x"70206368",
  4597 => x"616e6e65",
  4598 => x"6c207465",
  4599 => x"7374203c",
  4600 => x"70302e2e",
  4601 => x"353e0000",
  4602 => x"63687465",
  4603 => x"73740000",
  4604 => x"74657374",
  4605 => x"67656e65",
  4606 => x"7261746f",
  4607 => x"72203c73",
  4608 => x"63616c65",
  4609 => x"723e203c",
  4610 => x"72657374",
  4611 => x"6172743e",
  4612 => x"00000000",
  4613 => x"74657374",
  4614 => x"67656e00",
  4615 => x"3c6d7574",
  4616 => x"655f6e3e",
  4617 => x"203c7273",
  4618 => x"745f6e3e",
  4619 => x"203c6270",
  4620 => x"625f6e3e",
  4621 => x"203c6f73",
  4622 => x"72313e20",
  4623 => x"3c6f7372",
  4624 => x"323e0000",
  4625 => x"64616363",
  4626 => x"6f6e6600",
  4627 => x"636c6b20",
  4628 => x"3c73656c",
  4629 => x"6563743e",
  4630 => x"2030203d",
  4631 => x"20696e74",
  4632 => x"2c203120",
  4633 => x"3d206578",
  4634 => x"74000000",
  4635 => x"636c6b00",
  4636 => x"73686f77",
  4637 => x"20737973",
  4638 => x"74656d20",
  4639 => x"696e666f",
  4640 => x"203c7665",
  4641 => x"72626f73",
  4642 => x"653e0000",
  4643 => x"73797369",
  4644 => x"6e666f00",
  4645 => x"72756e6e",
  4646 => x"696e6720",
  4647 => x"6c696768",
  4648 => x"74000000",
  4649 => x"72756e00",
  4650 => x"72756e20",
  4651 => x"64697370",
  4652 => x"6c617920",
  4653 => x"74657374",
  4654 => x"2066756e",
  4655 => x"6374696f",
  4656 => x"6e000000",
  4657 => x"64697370",
  4658 => x"6c617900",
  4659 => x"73657420",
  4660 => x"6261636b",
  4661 => x"6c696768",
  4662 => x"74203c30",
  4663 => x"2e2e3331",
  4664 => x"3e000000",
  4665 => x"6261636b",
  4666 => x"00000000",
  4667 => x"73686f77",
  4668 => x"206c6f67",
  4669 => x"6f206f6e",
  4670 => x"20676c63",
  4671 => x"64000000",
  4672 => x"6c6f676f",
  4673 => x"00000000",
  4674 => x"63686563",
  4675 => x"6b204932",
  4676 => x"43206164",
  4677 => x"64726573",
  4678 => x"73000000",
  4679 => x"69326300",
  4680 => x"72656164",
  4681 => x"20454550",
  4682 => x"524f4d20",
  4683 => x"3c627573",
  4684 => x"3e203c69",
  4685 => x"32635f61",
  4686 => x"6464723e",
  4687 => x"203c6c65",
  4688 => x"6e677468",
  4689 => x"3e000000",
  4690 => x"65657072",
  4691 => x"6f6d0000",
  4692 => x"41444320",
  4693 => x"72656769",
  4694 => x"73746572",
  4695 => x"20747261",
  4696 => x"6e736665",
  4697 => x"72203c76",
  4698 => x"616c7565",
  4699 => x"3e000000",
  4700 => x"61747261",
  4701 => x"6e730000",
  4702 => x"696e6974",
  4703 => x"20414443",
  4704 => x"20726567",
  4705 => x"69737465",
  4706 => x"72730000",
  4707 => x"61696e69",
  4708 => x"74000000",
  4709 => x"616c6961",
  4710 => x"7320666f",
  4711 => x"72207800",
  4712 => x"6d656d00",
  4713 => x"77726974",
  4714 => x"6520776f",
  4715 => x"7264203c",
  4716 => x"61646472",
  4717 => x"3e203c6c",
  4718 => x"656e6774",
  4719 => x"683e203c",
  4720 => x"76616c75",
  4721 => x"65287329",
  4722 => x"3e000000",
  4723 => x"776d656d",
  4724 => x"00000000",
  4725 => x"6558616d",
  4726 => x"696e6520",
  4727 => x"6d656d6f",
  4728 => x"72790000",
  4729 => x"636c6561",
  4730 => x"72207363",
  4731 => x"7265656e",
  4732 => x"00000000",
  4733 => x"636c6561",
  4734 => x"72000000",
  4735 => x"0a307800",
  4736 => x"69326320",
  4737 => x"464d430a",
  4738 => x"00000000",
  4739 => x"61646472",
  4740 => x"6573733a",
  4741 => x"20307800",
  4742 => x"2020202d",
  4743 => x"2d3e2020",
  4744 => x"2041434b",
  4745 => x"0a000000",
  4746 => x"72656164",
  4747 => x"20646174",
  4748 => x"61202800",
  4749 => x"20627974",
  4750 => x"65732920",
  4751 => x"66726f6d",
  4752 => x"20493243",
  4753 => x"2d616464",
  4754 => x"72657373",
  4755 => x"20307800",
  4756 => x"0a0a0000",
  4757 => x"6e6f6163",
  4758 => x"6b200000",
  4759 => x"6368726f",
  4760 => x"6e74656c",
  4761 => x"20726567",
  4762 => x"20307800",
  4763 => x"3a203078",
  4764 => x"00000000",
  4765 => x"206e6163",
  4766 => x"6b000000",
  4767 => x"6572726f",
  4768 => x"7220286e",
  4769 => x"61636b29",
  4770 => x"0a000000",
  4771 => x"6265616d",
  4772 => x"20706f73",
  4773 => x"6974696f",
  4774 => x"6e206d6f",
  4775 => x"6e69746f",
  4776 => x"72207265",
  4777 => x"67697374",
  4778 => x"65727300",
  4779 => x"0a202020",
  4780 => x"20202020",
  4781 => x"20202020",
  4782 => x"20202020",
  4783 => x"20202020",
  4784 => x"20202020",
  4785 => x"20636861",
  4786 => x"6e6e656c",
  4787 => x"20302020",
  4788 => x"20636861",
  4789 => x"6e6e656c",
  4790 => x"20312020",
  4791 => x"20636861",
  4792 => x"6e6e656c",
  4793 => x"20322020",
  4794 => x"20636861",
  4795 => x"6e6e656c",
  4796 => x"20330000",
  4797 => x"0a202020",
  4798 => x"20202020",
  4799 => x"20202020",
  4800 => x"20202020",
  4801 => x"20202020",
  4802 => x"20202020",
  4803 => x"202d2d2d",
  4804 => x"2d20686f",
  4805 => x"72697a6f",
  4806 => x"6e74616c",
  4807 => x"202d2d2d",
  4808 => x"2d2d2020",
  4809 => x"202d2d2d",
  4810 => x"2d2d2d20",
  4811 => x"76657274",
  4812 => x"6963616c",
  4813 => x"202d2d2d",
  4814 => x"2d2d0000",
  4815 => x"0a736361",
  4816 => x"6c657220",
  4817 => x"76616c75",
  4818 => x"65732020",
  4819 => x"20202020",
  4820 => x"20202020",
  4821 => x"20000000",
  4822 => x"0a6e6f69",
  4823 => x"73652063",
  4824 => x"6f6d7065",
  4825 => x"6e736174",
  4826 => x"696f6e20",
  4827 => x"20202020",
  4828 => x"20000000",
  4829 => x"0a6d6561",
  4830 => x"73757265",
  4831 => x"6d656e74",
  4832 => x"20202020",
  4833 => x"20202020",
  4834 => x"20202020",
  4835 => x"20000000",
  4836 => x"0a73756d",
  4837 => x"20636861",
  4838 => x"6e6e656c",
  4839 => x"2020203a",
  4840 => x"20000000",
  4841 => x"0a706f73",
  4842 => x"6974696f",
  4843 => x"6e20636f",
  4844 => x"6d707574",
  4845 => x"6174696f",
  4846 => x"6e000000",
  4847 => x"0a202073",
  4848 => x"63616c65",
  4849 => x"72207661",
  4850 => x"6c756573",
  4851 => x"20202020",
  4852 => x"20202020",
  4853 => x"20000000",
  4854 => x"0a20206f",
  4855 => x"66667365",
  4856 => x"74202020",
  4857 => x"20202020",
  4858 => x"20202020",
  4859 => x"20202020",
  4860 => x"20000000",
  4861 => x"0a6f7574",
  4862 => x"70757420",
  4863 => x"73656c65",
  4864 => x"6374203a",
  4865 => x"20000000",
  4866 => x"6368616e",
  4867 => x"6e656c20",
  4868 => x"30000000",
  4869 => x"0a63616c",
  4870 => x"63207374",
  4871 => x"61746520",
  4872 => x"2020203a",
  4873 => x"20307800",
  4874 => x"0a202064",
  4875 => x"69766964",
  4876 => x"656e6420",
  4877 => x"63757474",
  4878 => x"65640000",
  4879 => x"0a20206e",
  4880 => x"6f697365",
  4881 => x"20636f6d",
  4882 => x"70656e73",
  4883 => x"6174696f",
  4884 => x"6e20746f",
  4885 => x"20626967",
  4886 => x"00000000",
  4887 => x"0a20206e",
  4888 => x"6f697365",
  4889 => x"2076616c",
  4890 => x"75652063",
  4891 => x"75747465",
  4892 => x"64000000",
  4893 => x"0a202073",
  4894 => x"756d2076",
  4895 => x"616c7565",
  4896 => x"20637574",
  4897 => x"74656400",
  4898 => x"76657274",
  4899 => x"6963616c",
  4900 => x"00000000",
  4901 => x"686f7269",
  4902 => x"7a6f6e74",
  4903 => x"616c0000",
  4904 => x"73756d00",
  4905 => x"6368616e",
  4906 => x"6e656c20",
  4907 => x"33000000",
  4908 => x"6368616e",
  4909 => x"6e656c20",
  4910 => x"32000000",
  4911 => x"6368616e",
  4912 => x"6e656c20",
  4913 => x"31000000",
  4914 => x"786d6f64",
  4915 => x"656d2074",
  4916 => x"72616e73",
  4917 => x"6d69742e",
  4918 => x"2e2e0a00",
  4919 => x"20627974",
  4920 => x"65732074",
  4921 => x"72616e73",
  4922 => x"6d697474",
  4923 => x"65640a00",
  4924 => x"63616e63",
  4925 => x"656c0a00",
  4926 => x"72657472",
  4927 => x"79206f75",
  4928 => x"740a0000",
  4929 => x"786d6f64",
  4930 => x"656d2072",
  4931 => x"65636569",
  4932 => x"76652e2e",
  4933 => x"2e0a0000",
  4934 => x"20627974",
  4935 => x"65732072",
  4936 => x"65636569",
  4937 => x"7665640a",
  4938 => x"00000000",
  4939 => x"72782062",
  4940 => x"75666665",
  4941 => x"72206675",
  4942 => x"6c6c0a00",
  4943 => x"74696d65",
  4944 => x"206f7574",
  4945 => x"0a000000",
  4946 => x"64656275",
  4947 => x"67207265",
  4948 => x"67697374",
  4949 => x"65727300",
  4950 => x"0a6d6f64",
  4951 => x"65202020",
  4952 => x"20202020",
  4953 => x"203a2000",
  4954 => x"0a616464",
  4955 => x"72657373",
  4956 => x"20302020",
  4957 => x"203a2030",
  4958 => x"78000000",
  4959 => x"0a616464",
  4960 => x"72657373",
  4961 => x"20312020",
  4962 => x"203a2030",
  4963 => x"78000000",
  4964 => x"0a627566",
  4965 => x"66657220",
  4966 => x"73697a65",
  4967 => x"203a2000",
  4968 => x"65787465",
  4969 => x"726e616c",
  4970 => x"20636c6f",
  4971 => x"636b2000",
  4972 => x"61637469",
  4973 => x"76650a00",
  4974 => x"4e4f5420",
  4975 => x"00000000",
  4976 => x"6265616d",
  4977 => x"20706f73",
  4978 => x"6974696f",
  4979 => x"6e206d6f",
  4980 => x"6e69746f",
  4981 => x"72000000",
  4982 => x"20286f6e",
  4983 => x"2073696d",
  4984 => x"290a0000",
  4985 => x"0a636f6d",
  4986 => x"70696c65",
  4987 => x"643a204a",
  4988 => x"756e2032",
  4989 => x"34203230",
  4990 => x"31312020",
  4991 => x"31333a33",
  4992 => x"393a3039",
  4993 => x"00000000",
  4994 => x"0a737973",
  4995 => x"74656d20",
  4996 => x"636c6f63",
  4997 => x"6b3a2000",
  4998 => x"204d487a",
  4999 => x"0a000000",
  5000 => x"44454255",
  5001 => x"47204d4f",
  5002 => x"44450000",
  5003 => x"204f4e0a",
  5004 => x"00000000",
  5005 => x"00000eb9",
  5006 => x"00000fa2",
  5007 => x"00000f98",
  5008 => x"00000f8e",
  5009 => x"00000f84",
  5010 => x"00000f7a",
  5011 => x"00000f70",
  5012 => x"0187fc09",
  5013 => x"026f0000",
  5014 => x"0003fff6",
  5015 => x"00060000",
  5016 => x"3e200000",
  5017 => x"636f6d6d",
  5018 => x"616e6420",
  5019 => x"6e6f7420",
  5020 => x"666f756e",
  5021 => x"642e0a00",
  5022 => x"73757070",
  5023 => x"6f727465",
  5024 => x"6420636f",
  5025 => x"6d6d616e",
  5026 => x"64733a0a",
  5027 => x"0a000000",
  5028 => x"202d2000",
  5029 => x"76656e64",
  5030 => x"6f723f20",
  5031 => x"20000000",
  5032 => x"67616973",
  5033 => x"6c657220",
  5034 => x"20000000",
  5035 => x"756e6b6e",
  5036 => x"6f776e20",
  5037 => x"64657669",
  5038 => x"63650000",
  5039 => x"485a4452",
  5040 => x"20202020",
  5041 => x"20000000",
  5042 => x"47656e65",
  5043 => x"72616c20",
  5044 => x"50757270",
  5045 => x"6f736520",
  5046 => x"492f4f20",
  5047 => x"706f7274",
  5048 => x"00000000",
  5049 => x"56474120",
  5050 => x"636f6e74",
  5051 => x"726f6c6c",
  5052 => x"65720000",
  5053 => x"4475616c",
  5054 => x"2d706f72",
  5055 => x"74204148",
  5056 => x"42205352",
  5057 => x"414d206d",
  5058 => x"6f64756c",
  5059 => x"65000000",
  5060 => x"64656275",
  5061 => x"67206275",
  5062 => x"66666572",
  5063 => x"20636f6e",
  5064 => x"74726f6c",
  5065 => x"00000000",
  5066 => x"74726967",
  5067 => x"67657220",
  5068 => x"67656e65",
  5069 => x"7261746f",
  5070 => x"72000000",
  5071 => x"64656275",
  5072 => x"6720636f",
  5073 => x"6e736f6c",
  5074 => x"65000000",
  5075 => x"44434d20",
  5076 => x"70686173",
  5077 => x"65207368",
  5078 => x"69667420",
  5079 => x"636f6e74",
  5080 => x"726f6c00",
  5081 => x"5a505520",
  5082 => x"4d656d6f",
  5083 => x"72792077",
  5084 => x"72617070",
  5085 => x"65720000",
  5086 => x"5a505520",
  5087 => x"41484220",
  5088 => x"57726170",
  5089 => x"70657200",
  5090 => x"4148422f",
  5091 => x"41504220",
  5092 => x"42726964",
  5093 => x"67650000",
  5094 => x"4d6f6475",
  5095 => x"6c617220",
  5096 => x"54696d65",
  5097 => x"7220556e",
  5098 => x"69740000",
  5099 => x"414d4241",
  5100 => x"20577261",
  5101 => x"70706572",
  5102 => x"20666f72",
  5103 => x"204f4320",
  5104 => x"4932432d",
  5105 => x"6d617374",
  5106 => x"65720000",
  5107 => x"47656e65",
  5108 => x"72696320",
  5109 => x"55415254",
  5110 => x"00000000",
  5111 => x"20206170",
  5112 => x"62736c76",
  5113 => x"00000000",
  5114 => x"76656e64",
  5115 => x"20307800",
  5116 => x"64657620",
  5117 => x"30780000",
  5118 => x"76657220",
  5119 => x"00000000",
  5120 => x"69727120",
  5121 => x"00000000",
  5122 => x"61646472",
  5123 => x"20307800",
  5124 => x"6168626d",
  5125 => x"73740000",
  5126 => x"61686273",
  5127 => x"6c760000",
  5128 => x"00001ef5",
  5129 => x"00001fa0",
  5130 => x"00001f95",
  5131 => x"00001f8a",
  5132 => x"00001f7f",
  5133 => x"00001f74",
  5134 => x"00001f69",
  5135 => x"00001f5e",
  5136 => x"04580808",
  5137 => x"20ff0000",
  5138 => x"00005050",
  5139 => x"00005130",
  5140 => x"02010305",
  5141 => x"05070501",
  5142 => x"03030505",
  5143 => x"02030104",
  5144 => x"05050505",
  5145 => x"05050505",
  5146 => x"05050101",
  5147 => x"04050404",
  5148 => x"07050505",
  5149 => x"05050505",
  5150 => x"05030405",
  5151 => x"05050505",
  5152 => x"05050505",
  5153 => x"05050505",
  5154 => x"05050503",
  5155 => x"04030505",
  5156 => x"02050504",
  5157 => x"05050405",
  5158 => x"04010204",
  5159 => x"02050404",
  5160 => x"05050404",
  5161 => x"04040507",
  5162 => x"05040404",
  5163 => x"02040500",
  5164 => x"04050200",
  5165 => x"04080303",
  5166 => x"04090003",
  5167 => x"06000000",
  5168 => x"00020204",
  5169 => x"04040400",
  5170 => x"04060003",
  5171 => x"05000000",
  5172 => x"00000404",
  5173 => x"05050204",
  5174 => x"05060305",
  5175 => x"04030705",
  5176 => x"04050303",
  5177 => x"02040502",
  5178 => x"03020405",
  5179 => x"06060604",
  5180 => x"05050505",
  5181 => x"05050504",
  5182 => x"04040404",
  5183 => x"03030303",
  5184 => x"05050505",
  5185 => x"05050505",
  5186 => x"05040404",
  5187 => x"04050404",
  5188 => x"04040404",
  5189 => x"04040503",
  5190 => x"04040404",
  5191 => x"02020303",
  5192 => x"04040404",
  5193 => x"04040405",
  5194 => x"04040404",
  5195 => x"04030303",
  5196 => x"00005f07",
  5197 => x"0007741c",
  5198 => x"771c172e",
  5199 => x"6a3e2b3a",
  5200 => x"06493608",
  5201 => x"36493036",
  5202 => x"49597648",
  5203 => x"073c4281",
  5204 => x"81423c0a",
  5205 => x"041f040a",
  5206 => x"08083e08",
  5207 => x"08806008",
  5208 => x"080840c0",
  5209 => x"300c033e",
  5210 => x"4141413e",
  5211 => x"44427f40",
  5212 => x"40466151",
  5213 => x"49462241",
  5214 => x"49493618",
  5215 => x"14127f10",
  5216 => x"27454545",
  5217 => x"393e4949",
  5218 => x"49300101",
  5219 => x"710d0336",
  5220 => x"49494936",
  5221 => x"06494929",
  5222 => x"1e36d008",
  5223 => x"14224114",
  5224 => x"14141414",
  5225 => x"41221408",
  5226 => x"02510906",
  5227 => x"3c4299a5",
  5228 => x"bd421c7c",
  5229 => x"1211127c",
  5230 => x"7f494949",
  5231 => x"363e4141",
  5232 => x"41227f41",
  5233 => x"41413e7f",
  5234 => x"49494941",
  5235 => x"7f090909",
  5236 => x"013e4149",
  5237 => x"497a7f08",
  5238 => x"08087f41",
  5239 => x"7f414041",
  5240 => x"413f7f08",
  5241 => x"1422417f",
  5242 => x"40404040",
  5243 => x"7f060c06",
  5244 => x"7f7f0608",
  5245 => x"307f3e41",
  5246 => x"41413e7f",
  5247 => x"09090906",
  5248 => x"3e4161c1",
  5249 => x"be7f0919",
  5250 => x"29462649",
  5251 => x"49493201",
  5252 => x"017f0101",
  5253 => x"3f404040",
  5254 => x"3f073840",
  5255 => x"38071f60",
  5256 => x"1f601f63",
  5257 => x"14081463",
  5258 => x"01067806",
  5259 => x"01615149",
  5260 => x"45437f41",
  5261 => x"41030c30",
  5262 => x"c041417f",
  5263 => x"04020102",
  5264 => x"04808080",
  5265 => x"80800102",
  5266 => x"20545454",
  5267 => x"787f4444",
  5268 => x"44383844",
  5269 => x"44443844",
  5270 => x"44447f38",
  5271 => x"54545458",
  5272 => x"087e0901",
  5273 => x"18a4a4a4",
  5274 => x"787f0404",
  5275 => x"787d807d",
  5276 => x"7f102844",
  5277 => x"3f407c04",
  5278 => x"7804787c",
  5279 => x"04047838",
  5280 => x"444438fc",
  5281 => x"24242418",
  5282 => x"18242424",
  5283 => x"fc7c0804",
  5284 => x"04485454",
  5285 => x"24043f44",
  5286 => x"403c4040",
  5287 => x"7c1c2040",
  5288 => x"201c1c60",
  5289 => x"601c6060",
  5290 => x"1c442810",
  5291 => x"28449ca0",
  5292 => x"601c6454",
  5293 => x"544c187e",
  5294 => x"8181ffff",
  5295 => x"81817e18",
  5296 => x"18040810",
  5297 => x"0c143e55",
  5298 => x"55ff8181",
  5299 => x"81ff8060",
  5300 => x"80608060",
  5301 => x"60600060",
  5302 => x"60006060",
  5303 => x"047f0414",
  5304 => x"7f140201",
  5305 => x"01024629",
  5306 => x"1608344a",
  5307 => x"31483000",
  5308 => x"18243e41",
  5309 => x"227f4941",
  5310 => x"03040403",
  5311 => x"03040304",
  5312 => x"04030403",
  5313 => x"183c3c18",
  5314 => x"08080808",
  5315 => x"03010203",
  5316 => x"020e020e",
  5317 => x"060e0048",
  5318 => x"30384438",
  5319 => x"54483844",
  5320 => x"fe44487e",
  5321 => x"49014438",
  5322 => x"28384403",
  5323 => x"147c1403",
  5324 => x"e7e74e55",
  5325 => x"55390101",
  5326 => x"0001011c",
  5327 => x"2a555522",
  5328 => x"1c1d151e",
  5329 => x"18240018",
  5330 => x"24080808",
  5331 => x"18080808",
  5332 => x"3c42bd95",
  5333 => x"a9423c01",
  5334 => x"01010101",
  5335 => x"06090906",
  5336 => x"44445f44",
  5337 => x"44191512",
  5338 => x"15150a02",
  5339 => x"01fc2020",
  5340 => x"1c0e7f01",
  5341 => x"7f011818",
  5342 => x"00804002",
  5343 => x"1f060909",
  5344 => x"06241800",
  5345 => x"2418824f",
  5346 => x"304c62f1",
  5347 => x"824f300c",
  5348 => x"d2b1955f",
  5349 => x"304c62f1",
  5350 => x"30484520",
  5351 => x"60392e38",
  5352 => x"6060382e",
  5353 => x"3960701d",
  5354 => x"131d7072",
  5355 => x"1d121e71",
  5356 => x"701d121d",
  5357 => x"70603b25",
  5358 => x"3b607e11",
  5359 => x"7f49411e",
  5360 => x"2161927c",
  5361 => x"5556447c",
  5362 => x"5655447c",
  5363 => x"5655467d",
  5364 => x"54544545",
  5365 => x"7e44447e",
  5366 => x"45467d46",
  5367 => x"457c4508",
  5368 => x"7f49413e",
  5369 => x"7e091222",
  5370 => x"7d384546",
  5371 => x"44383844",
  5372 => x"46453838",
  5373 => x"46454638",
  5374 => x"3a454546",
  5375 => x"39384544",
  5376 => x"45382214",
  5377 => x"081422bc",
  5378 => x"625a463d",
  5379 => x"3c41423c",
  5380 => x"3c42413c",
  5381 => x"3c42413e",
  5382 => x"3d40403d",
  5383 => x"0608f209",
  5384 => x"067f2222",
  5385 => x"1cfe0989",
  5386 => x"76205556",
  5387 => x"78205655",
  5388 => x"78225555",
  5389 => x"7a235556",
  5390 => x"7b205554",
  5391 => x"79275557",
  5392 => x"78205438",
  5393 => x"54483844",
  5394 => x"c4385556",
  5395 => x"58385655",
  5396 => x"583a5555",
  5397 => x"5a395454",
  5398 => x"59017a7a",
  5399 => x"01027902",
  5400 => x"02780260",
  5401 => x"91927c7b",
  5402 => x"090a7338",
  5403 => x"45463838",
  5404 => x"4645383a",
  5405 => x"45453a3b",
  5406 => x"45463b39",
  5407 => x"44443908",
  5408 => x"082a0808",
  5409 => x"b8644c3a",
  5410 => x"3c41427c",
  5411 => x"3c42417c",
  5412 => x"3a41417a",
  5413 => x"3d40407d",
  5414 => x"986219ff",
  5415 => x"423c9a60",
  5416 => x"1a000000",
  5417 => x"30622020",
  5418 => x"20202020",
  5419 => x"20202020",
  5420 => x"20202020",
  5421 => x"20202020",
  5422 => x"20202020",
  5423 => x"20202020",
  5424 => x"20202020",
  5425 => x"20200000",
  5426 => x"20202020",
  5427 => x"20202020",
  5428 => x"00000000",
  5429 => x"00202020",
  5430 => x"20202020",
  5431 => x"20202828",
  5432 => x"28282820",
  5433 => x"20202020",
  5434 => x"20202020",
  5435 => x"20202020",
  5436 => x"20202020",
  5437 => x"20881010",
  5438 => x"10101010",
  5439 => x"10101010",
  5440 => x"10101010",
  5441 => x"10040404",
  5442 => x"04040404",
  5443 => x"04040410",
  5444 => x"10101010",
  5445 => x"10104141",
  5446 => x"41414141",
  5447 => x"01010101",
  5448 => x"01010101",
  5449 => x"01010101",
  5450 => x"01010101",
  5451 => x"01010101",
  5452 => x"10101010",
  5453 => x"10104242",
  5454 => x"42424242",
  5455 => x"02020202",
  5456 => x"02020202",
  5457 => x"02020202",
  5458 => x"02020202",
  5459 => x"02020202",
  5460 => x"10101010",
  5461 => x"20000000",
  5462 => x"00000000",
  5463 => x"00000000",
  5464 => x"00000000",
  5465 => x"00000000",
  5466 => x"00000000",
  5467 => x"00000000",
  5468 => x"00000000",
  5469 => x"00000000",
  5470 => x"00000000",
  5471 => x"00000000",
  5472 => x"00000000",
  5473 => x"00000000",
  5474 => x"00000000",
  5475 => x"00000000",
  5476 => x"00000000",
  5477 => x"00000000",
  5478 => x"00000000",
  5479 => x"00000000",
  5480 => x"00000000",
  5481 => x"00000000",
  5482 => x"00000000",
  5483 => x"00000000",
  5484 => x"00000000",
  5485 => x"00000000",
  5486 => x"00000000",
  5487 => x"00000000",
  5488 => x"00000000",
  5489 => x"00000000",
  5490 => x"00000000",
  5491 => x"00000000",
  5492 => x"00000000",
  5493 => x"00000000",
  5494 => x"43000000",
  5495 => x"80000c00",
  5496 => x"80000b00",
  5497 => x"80000800",
  5498 => x"ff000000",
  5499 => x"00000000",
  5500 => x"00000000",
  5501 => x"00ffffff",
  5502 => x"ff00ffff",
  5503 => x"ffff00ff",
  5504 => x"ffffff00",
  5505 => x"00000000",
  5506 => x"00000000",
  5507 => x"80000a00",
  5508 => x"80000700",
  5509 => x"80000600",
  5510 => x"80000400",
  5511 => x"80000200",
  5512 => x"80000100",
  5513 => x"80000004",
  5514 => x"80000000",
  5515 => x"00005630",
  5516 => x"00000000",
  5517 => x"00005898",
  5518 => x"000058f4",
  5519 => x"00005950",
  5520 => x"00000000",
  5521 => x"00000000",
  5522 => x"00000000",
  5523 => x"00000000",
  5524 => x"00000000",
  5525 => x"00000000",
  5526 => x"00000000",
  5527 => x"00000000",
  5528 => x"00000000",
  5529 => x"000055d8",
  5530 => x"00000000",
  5531 => x"00000000",
  5532 => x"00000000",
  5533 => x"00000000",
  5534 => x"00000000",
  5535 => x"00000000",
  5536 => x"00000000",
  5537 => x"00000000",
  5538 => x"00000000",
  5539 => x"00000000",
  5540 => x"00000000",
  5541 => x"00000000",
  5542 => x"00000000",
  5543 => x"00000000",
  5544 => x"00000000",
  5545 => x"00000000",
  5546 => x"00000000",
  5547 => x"00000000",
  5548 => x"00000000",
  5549 => x"00000000",
  5550 => x"00000000",
  5551 => x"00000000",
  5552 => x"00000000",
  5553 => x"00000000",
  5554 => x"00000000",
  5555 => x"00000000",
  5556 => x"00000000",
  5557 => x"00000000",
  5558 => x"00000001",
  5559 => x"330eabcd",
  5560 => x"1234e66d",
  5561 => x"deec0005",
  5562 => x"000b0000",
  5563 => x"00000000",
  5564 => x"00000000",
  5565 => x"00000000",
  5566 => x"00000000",
  5567 => x"00000000",
  5568 => x"00000000",
  5569 => x"00000000",
  5570 => x"00000000",
  5571 => x"00000000",
  5572 => x"00000000",
  5573 => x"00000000",
  5574 => x"00000000",
  5575 => x"00000000",
  5576 => x"00000000",
  5577 => x"00000000",
  5578 => x"00000000",
  5579 => x"00000000",
  5580 => x"00000000",
  5581 => x"00000000",
  5582 => x"00000000",
  5583 => x"00000000",
  5584 => x"00000000",
  5585 => x"00000000",
  5586 => x"00000000",
  5587 => x"00000000",
  5588 => x"00000000",
  5589 => x"00000000",
  5590 => x"00000000",
  5591 => x"00000000",
  5592 => x"00000000",
  5593 => x"00000000",
  5594 => x"00000000",
  5595 => x"00000000",
  5596 => x"00000000",
  5597 => x"00000000",
  5598 => x"00000000",
  5599 => x"00000000",
  5600 => x"00000000",
  5601 => x"00000000",
  5602 => x"00000000",
  5603 => x"00000000",
  5604 => x"00000000",
  5605 => x"00000000",
  5606 => x"00000000",
  5607 => x"00000000",
  5608 => x"00000000",
  5609 => x"00000000",
  5610 => x"00000000",
  5611 => x"00000000",
  5612 => x"00000000",
  5613 => x"00000000",
  5614 => x"00000000",
  5615 => x"00000000",
  5616 => x"00000000",
  5617 => x"00000000",
  5618 => x"00000000",
  5619 => x"00000000",
  5620 => x"00000000",
  5621 => x"00000000",
  5622 => x"00000000",
  5623 => x"00000000",
  5624 => x"00000000",
  5625 => x"00000000",
  5626 => x"00000000",
  5627 => x"00000000",
  5628 => x"00000000",
  5629 => x"00000000",
  5630 => x"00000000",
  5631 => x"00000000",
  5632 => x"00000000",
  5633 => x"00000000",
  5634 => x"00000000",
  5635 => x"00000000",
  5636 => x"00000000",
  5637 => x"00000000",
  5638 => x"00000000",
  5639 => x"00000000",
  5640 => x"00000000",
  5641 => x"00000000",
  5642 => x"00000000",
  5643 => x"00000000",
  5644 => x"00000000",
  5645 => x"00000000",
  5646 => x"00000000",
  5647 => x"00000000",
  5648 => x"00000000",
  5649 => x"00000000",
  5650 => x"00000000",
  5651 => x"00000000",
  5652 => x"00000000",
  5653 => x"00000000",
  5654 => x"00000000",
  5655 => x"00000000",
  5656 => x"00000000",
  5657 => x"00000000",
  5658 => x"00000000",
  5659 => x"00000000",
  5660 => x"00000000",
  5661 => x"00000000",
  5662 => x"00000000",
  5663 => x"00000000",
  5664 => x"00000000",
  5665 => x"00000000",
  5666 => x"00000000",
  5667 => x"00000000",
  5668 => x"00000000",
  5669 => x"00000000",
  5670 => x"00000000",
  5671 => x"00000000",
  5672 => x"00000000",
  5673 => x"00000000",
  5674 => x"00000000",
  5675 => x"00000000",
  5676 => x"00000000",
  5677 => x"00000000",
  5678 => x"00000000",
  5679 => x"00000000",
  5680 => x"00000000",
  5681 => x"00000000",
  5682 => x"00000000",
  5683 => x"00000000",
  5684 => x"00000000",
  5685 => x"00000000",
  5686 => x"00000000",
  5687 => x"00000000",
  5688 => x"00000000",
  5689 => x"00000000",
  5690 => x"00000000",
  5691 => x"00000000",
  5692 => x"00000000",
  5693 => x"00000000",
  5694 => x"00000000",
  5695 => x"00000000",
  5696 => x"00000000",
  5697 => x"00000000",
  5698 => x"00000000",
  5699 => x"00000000",
  5700 => x"00000000",
  5701 => x"00000000",
  5702 => x"00000000",
  5703 => x"00000000",
  5704 => x"00000000",
  5705 => x"00000000",
  5706 => x"00000000",
  5707 => x"00000000",
  5708 => x"00000000",
  5709 => x"00000000",
  5710 => x"00000000",
  5711 => x"00000000",
  5712 => x"00000000",
  5713 => x"00000000",
  5714 => x"00000000",
  5715 => x"00000000",
  5716 => x"00000000",
  5717 => x"00000000",
  5718 => x"00000000",
  5719 => x"00000000",
  5720 => x"00000000",
  5721 => x"00000000",
  5722 => x"00000000",
  5723 => x"00000000",
  5724 => x"00000000",
  5725 => x"00000000",
  5726 => x"00000000",
  5727 => x"00000000",
  5728 => x"00000000",
  5729 => x"00000000",
  5730 => x"00000000",
  5731 => x"00000000",
  5732 => x"00000000",
  5733 => x"00000000",
  5734 => x"00000000",
  5735 => x"00000000",
  5736 => x"00000000",
  5737 => x"00000000",
  5738 => x"00000000",
  5739 => x"00000000",
  5740 => x"00000000",
  5741 => x"00000000",
  5742 => x"00000000",
  5743 => x"00000000",
  5744 => x"00000000",
  5745 => x"00000000",
  5746 => x"00000000",
  5747 => x"00000000",
  5748 => x"00000000",
  5749 => x"00000000",
  5750 => x"00000000",
  5751 => x"ffffffff",
  5752 => x"00000000",
  5753 => x"00020000",
  5754 => x"00000000",
  5755 => x"00000000",
  5756 => x"000059e8",
  5757 => x"000059e8",
  5758 => x"000059f0",
  5759 => x"000059f0",
  5760 => x"000059f8",
  5761 => x"000059f8",
  5762 => x"00005a00",
  5763 => x"00005a00",
  5764 => x"00005a08",
  5765 => x"00005a08",
  5766 => x"00005a10",
  5767 => x"00005a10",
  5768 => x"00005a18",
  5769 => x"00005a18",
  5770 => x"00005a20",
  5771 => x"00005a20",
  5772 => x"00005a28",
  5773 => x"00005a28",
  5774 => x"00005a30",
  5775 => x"00005a30",
  5776 => x"00005a38",
  5777 => x"00005a38",
  5778 => x"00005a40",
  5779 => x"00005a40",
  5780 => x"00005a48",
  5781 => x"00005a48",
  5782 => x"00005a50",
  5783 => x"00005a50",
  5784 => x"00005a58",
  5785 => x"00005a58",
  5786 => x"00005a60",
  5787 => x"00005a60",
  5788 => x"00005a68",
  5789 => x"00005a68",
  5790 => x"00005a70",
  5791 => x"00005a70",
  5792 => x"00005a78",
  5793 => x"00005a78",
  5794 => x"00005a80",
  5795 => x"00005a80",
  5796 => x"00005a88",
  5797 => x"00005a88",
  5798 => x"00005a90",
  5799 => x"00005a90",
  5800 => x"00005a98",
  5801 => x"00005a98",
  5802 => x"00005aa0",
  5803 => x"00005aa0",
  5804 => x"00005aa8",
  5805 => x"00005aa8",
  5806 => x"00005ab0",
  5807 => x"00005ab0",
  5808 => x"00005ab8",
  5809 => x"00005ab8",
  5810 => x"00005ac0",
  5811 => x"00005ac0",
  5812 => x"00005ac8",
  5813 => x"00005ac8",
  5814 => x"00005ad0",
  5815 => x"00005ad0",
  5816 => x"00005ad8",
  5817 => x"00005ad8",
  5818 => x"00005ae0",
  5819 => x"00005ae0",
  5820 => x"00005ae8",
  5821 => x"00005ae8",
  5822 => x"00005af0",
  5823 => x"00005af0",
  5824 => x"00005af8",
  5825 => x"00005af8",
  5826 => x"00005b00",
  5827 => x"00005b00",
  5828 => x"00005b08",
  5829 => x"00005b08",
  5830 => x"00005b10",
  5831 => x"00005b10",
  5832 => x"00005b18",
  5833 => x"00005b18",
  5834 => x"00005b20",
  5835 => x"00005b20",
  5836 => x"00005b28",
  5837 => x"00005b28",
  5838 => x"00005b30",
  5839 => x"00005b30",
  5840 => x"00005b38",
  5841 => x"00005b38",
  5842 => x"00005b40",
  5843 => x"00005b40",
  5844 => x"00005b48",
  5845 => x"00005b48",
  5846 => x"00005b50",
  5847 => x"00005b50",
  5848 => x"00005b58",
  5849 => x"00005b58",
  5850 => x"00005b60",
  5851 => x"00005b60",
  5852 => x"00005b68",
  5853 => x"00005b68",
  5854 => x"00005b70",
  5855 => x"00005b70",
  5856 => x"00005b78",
  5857 => x"00005b78",
  5858 => x"00005b80",
  5859 => x"00005b80",
  5860 => x"00005b88",
  5861 => x"00005b88",
  5862 => x"00005b90",
  5863 => x"00005b90",
  5864 => x"00005b98",
  5865 => x"00005b98",
  5866 => x"00005ba0",
  5867 => x"00005ba0",
  5868 => x"00005ba8",
  5869 => x"00005ba8",
  5870 => x"00005bb0",
  5871 => x"00005bb0",
  5872 => x"00005bb8",
  5873 => x"00005bb8",
  5874 => x"00005bc0",
  5875 => x"00005bc0",
  5876 => x"00005bc8",
  5877 => x"00005bc8",
  5878 => x"00005bd0",
  5879 => x"00005bd0",
  5880 => x"00005bd8",
  5881 => x"00005bd8",
  5882 => x"00005be0",
  5883 => x"00005be0",
  5884 => x"00005be8",
  5885 => x"00005be8",
  5886 => x"00005bf0",
  5887 => x"00005bf0",
  5888 => x"00005bf8",
  5889 => x"00005bf8",
  5890 => x"00005c00",
  5891 => x"00005c00",
  5892 => x"00005c08",
  5893 => x"00005c08",
  5894 => x"00005c10",
  5895 => x"00005c10",
  5896 => x"00005c18",
  5897 => x"00005c18",
  5898 => x"00005c20",
  5899 => x"00005c20",
  5900 => x"00005c28",
  5901 => x"00005c28",
  5902 => x"00005c30",
  5903 => x"00005c30",
  5904 => x"00005c38",
  5905 => x"00005c38",
  5906 => x"00005c40",
  5907 => x"00005c40",
  5908 => x"00005c48",
  5909 => x"00005c48",
  5910 => x"00005c50",
  5911 => x"00005c50",
  5912 => x"00005c58",
  5913 => x"00005c58",
  5914 => x"00005c60",
  5915 => x"00005c60",
  5916 => x"00005c68",
  5917 => x"00005c68",
  5918 => x"00005c70",
  5919 => x"00005c70",
  5920 => x"00005c78",
  5921 => x"00005c78",
  5922 => x"00005c80",
  5923 => x"00005c80",
  5924 => x"00005c88",
  5925 => x"00005c88",
  5926 => x"00005c90",
  5927 => x"00005c90",
  5928 => x"00005c98",
  5929 => x"00005c98",
  5930 => x"00005ca0",
  5931 => x"00005ca0",
  5932 => x"00005ca8",
  5933 => x"00005ca8",
  5934 => x"00005cb0",
  5935 => x"00005cb0",
  5936 => x"00005cb8",
  5937 => x"00005cb8",
  5938 => x"00005cc0",
  5939 => x"00005cc0",
  5940 => x"00005cc8",
  5941 => x"00005cc8",
  5942 => x"00005cd0",
  5943 => x"00005cd0",
  5944 => x"00005cd8",
  5945 => x"00005cd8",
  5946 => x"00005ce0",
  5947 => x"00005ce0",
  5948 => x"00005ce8",
  5949 => x"00005ce8",
  5950 => x"00005cf0",
  5951 => x"00005cf0",
  5952 => x"00005cf8",
  5953 => x"00005cf8",
  5954 => x"00005d00",
  5955 => x"00005d00",
  5956 => x"00005d08",
  5957 => x"00005d08",
  5958 => x"00005d10",
  5959 => x"00005d10",
  5960 => x"00005d18",
  5961 => x"00005d18",
  5962 => x"00005d20",
  5963 => x"00005d20",
  5964 => x"00005d28",
  5965 => x"00005d28",
  5966 => x"00005d30",
  5967 => x"00005d30",
  5968 => x"00005d38",
  5969 => x"00005d38",
  5970 => x"00005d40",
  5971 => x"00005d40",
  5972 => x"00005d48",
  5973 => x"00005d48",
  5974 => x"00005d50",
  5975 => x"00005d50",
  5976 => x"00005d58",
  5977 => x"00005d58",
  5978 => x"00005d60",
  5979 => x"00005d60",
  5980 => x"00005d68",
  5981 => x"00005d68",
  5982 => x"00005d70",
  5983 => x"00005d70",
  5984 => x"00005d78",
  5985 => x"00005d78",
  5986 => x"00005d80",
  5987 => x"00005d80",
  5988 => x"00005d88",
  5989 => x"00005d88",
  5990 => x"00005d90",
  5991 => x"00005d90",
  5992 => x"00005d98",
  5993 => x"00005d98",
  5994 => x"00005da0",
  5995 => x"00005da0",
  5996 => x"00005da8",
  5997 => x"00005da8",
  5998 => x"00005db0",
  5999 => x"00005db0",
  6000 => x"00005db8",
  6001 => x"00005db8",
  6002 => x"00005dc0",
  6003 => x"00005dc0",
  6004 => x"00005dc8",
  6005 => x"00005dc8",
  6006 => x"00005dd0",
  6007 => x"00005dd0",
  6008 => x"00005dd8",
  6009 => x"00005dd8",
  6010 => x"00005de0",
  6011 => x"00005de0",
	--others => x"aaaaaaaa" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
