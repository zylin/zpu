library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80cfd80c",
3 => x"3a0b0b80",
4 => x"c6d00400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"80c7972d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80cf",
162 => x"c4738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0b8b",
171 => x"9f2d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0b8b",
179 => x"e32d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80cfd40c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"82c53f80",
257 => x"c6d93f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"fe3d0d0b",
281 => x"0b80dfc0",
282 => x"08538413",
283 => x"0870882a",
284 => x"70810651",
285 => x"52527080",
286 => x"2ef03871",
287 => x"81ff0680",
288 => x"0c843d0d",
289 => x"04ff3d0d",
290 => x"0b0b80df",
291 => x"c0085271",
292 => x"0870882a",
293 => x"81327081",
294 => x"06515151",
295 => x"70f13873",
296 => x"720c833d",
297 => x"0d0480cf",
298 => x"d408802e",
299 => x"a43880cf",
300 => x"d808822e",
301 => x"bd388380",
302 => x"800b0b0b",
303 => x"80dfc00c",
304 => x"82a0800b",
305 => x"80dfc40c",
306 => x"8290800b",
307 => x"80dfc80c",
308 => x"04f88080",
309 => x"80a40b0b",
310 => x"0b80dfc0",
311 => x"0cf88080",
312 => x"82800b80",
313 => x"dfc40cf8",
314 => x"80808480",
315 => x"0b80dfc8",
316 => x"0c0480c0",
317 => x"a8808c0b",
318 => x"0b0b80df",
319 => x"c00c80c0",
320 => x"a880940b",
321 => x"80dfc40c",
322 => x"0b0b80cf",
323 => x"8c0b80df",
324 => x"c80c0470",
325 => x"7080dfcc",
326 => x"335170a7",
327 => x"3880cfe0",
328 => x"08700852",
329 => x"5270802e",
330 => x"94388412",
331 => x"80cfe00c",
332 => x"702d80cf",
333 => x"e0087008",
334 => x"525270ee",
335 => x"38810b80",
336 => x"dfcc3450",
337 => x"50040470",
338 => x"0b0b80df",
339 => x"bc08802e",
340 => x"8e380b0b",
341 => x"0b0b800b",
342 => x"802e0981",
343 => x"06833850",
344 => x"040b0b80",
345 => x"dfbc510b",
346 => x"0b0bf594",
347 => x"3f500404",
348 => x"fe3d0d89",
349 => x"5380cf90",
350 => x"5182c13f",
351 => x"80cfa051",
352 => x"82ba3f81",
353 => x"0a0b80df",
354 => x"d80cff0b",
355 => x"80dfdc0c",
356 => x"ff135372",
357 => x"8025de38",
358 => x"72800c84",
359 => x"3d0d04fb",
360 => x"3d0d7779",
361 => x"55558056",
362 => x"757524ab",
363 => x"38807424",
364 => x"9d388053",
365 => x"73527451",
366 => x"80e13f80",
367 => x"08547580",
368 => x"2e853880",
369 => x"08305473",
370 => x"800c873d",
371 => x"0d047330",
372 => x"76813257",
373 => x"54dc3974",
374 => x"30558156",
375 => x"738025d2",
376 => x"38ec39fa",
377 => x"3d0d787a",
378 => x"57558057",
379 => x"767524a4",
380 => x"38759f2c",
381 => x"54815375",
382 => x"74327431",
383 => x"5274519b",
384 => x"3f800854",
385 => x"76802e85",
386 => x"38800830",
387 => x"5473800c",
388 => x"883d0d04",
389 => x"74305581",
390 => x"57d739fc",
391 => x"3d0d7678",
392 => x"53548153",
393 => x"80747326",
394 => x"52557280",
395 => x"2e983870",
396 => x"802eab38",
397 => x"807224a6",
398 => x"38711073",
399 => x"10757226",
400 => x"53545272",
401 => x"ea387351",
402 => x"78833874",
403 => x"5170800c",
404 => x"863d0d04",
405 => x"720a100a",
406 => x"720a100a",
407 => x"53537280",
408 => x"2ee43871",
409 => x"7426ed38",
410 => x"73723175",
411 => x"7407740a",
412 => x"100a740a",
413 => x"100a5555",
414 => x"5654e339",
415 => x"f73d0d7c",
416 => x"70525380",
417 => x"f93f7254",
418 => x"80085580",
419 => x"cfb05681",
420 => x"57800881",
421 => x"055a8b3d",
422 => x"e4115953",
423 => x"8259f413",
424 => x"527b8811",
425 => x"08525381",
426 => x"b23f8008",
427 => x"30708008",
428 => x"079f2c8a",
429 => x"07800c53",
430 => x"8b3d0d04",
431 => x"f63d0d7c",
432 => x"80cfe408",
433 => x"71535553",
434 => x"b53f7255",
435 => x"80085680",
436 => x"cfb05781",
437 => x"58800881",
438 => x"055b8c3d",
439 => x"e4115a53",
440 => x"825af413",
441 => x"52881408",
442 => x"5180f03f",
443 => x"80083070",
444 => x"8008079f",
445 => x"2c8a0780",
446 => x"0c548c3d",
447 => x"0d047070",
448 => x"70707570",
449 => x"71830653",
450 => x"555270b4",
451 => x"38717008",
452 => x"7009f7fb",
453 => x"fdff1206",
454 => x"f8848281",
455 => x"80065452",
456 => x"53719b38",
457 => x"84137008",
458 => x"7009f7fb",
459 => x"fdff1206",
460 => x"f8848281",
461 => x"80065452",
462 => x"5371802e",
463 => x"e7387252",
464 => x"71335372",
465 => x"802e8a38",
466 => x"81127033",
467 => x"545272f8",
468 => x"38717431",
469 => x"800c5050",
470 => x"505004f2",
471 => x"3d0d6062",
472 => x"88110870",
473 => x"58565f5a",
474 => x"73802e81",
475 => x"8c388c1a",
476 => x"2270832a",
477 => x"81328106",
478 => x"56587486",
479 => x"38901a08",
480 => x"91387951",
481 => x"90b73fff",
482 => x"55800880",
483 => x"ec388c1a",
484 => x"22587d08",
485 => x"55807883",
486 => x"ffff0670",
487 => x"0a100a81",
488 => x"06415c57",
489 => x"7e772e80",
490 => x"d7387690",
491 => x"38740884",
492 => x"16088817",
493 => x"57585676",
494 => x"802ef238",
495 => x"76548880",
496 => x"77278438",
497 => x"88805473",
498 => x"5375529c",
499 => x"1a0851a4",
500 => x"1a085877",
501 => x"2d800b80",
502 => x"082582e0",
503 => x"38800816",
504 => x"77800831",
505 => x"7f880508",
506 => x"80083170",
507 => x"6188050c",
508 => x"5b585678",
509 => x"ffb43880",
510 => x"5574800c",
511 => x"903d0d04",
512 => x"7a813281",
513 => x"06774056",
514 => x"75802e81",
515 => x"bd387690",
516 => x"38740884",
517 => x"16088817",
518 => x"57585976",
519 => x"802ef238",
520 => x"881a0878",
521 => x"83ffff06",
522 => x"70892a81",
523 => x"06565956",
524 => x"73802e82",
525 => x"f8387577",
526 => x"278b3877",
527 => x"872a8106",
528 => x"5c7b82b5",
529 => x"38767627",
530 => x"83387656",
531 => x"75537852",
532 => x"79085185",
533 => x"833f881a",
534 => x"08763188",
535 => x"1b0c7908",
536 => x"167a0c76",
537 => x"56751977",
538 => x"77317f88",
539 => x"05087831",
540 => x"70618805",
541 => x"0c415859",
542 => x"7e802efe",
543 => x"fa388c1a",
544 => x"2258ff8a",
545 => x"39787954",
546 => x"7c537b52",
547 => x"5684c93f",
548 => x"881a0879",
549 => x"31881b0c",
550 => x"7908197a",
551 => x"0c7c7631",
552 => x"5d7c8e38",
553 => x"79518ff2",
554 => x"3f800881",
555 => x"8f388008",
556 => x"5f751c77",
557 => x"77317f88",
558 => x"05087831",
559 => x"70618805",
560 => x"0c5d585c",
561 => x"7a802efe",
562 => x"ae387681",
563 => x"83387408",
564 => x"84160888",
565 => x"1757585c",
566 => x"76802ef2",
567 => x"3876538a",
568 => x"527b5182",
569 => x"d33f8008",
570 => x"7c318105",
571 => x"5d800884",
572 => x"3881175d",
573 => x"815f7c59",
574 => x"767d2783",
575 => x"38765994",
576 => x"1a08881b",
577 => x"08115758",
578 => x"807a085c",
579 => x"54901a08",
580 => x"7b278338",
581 => x"81547579",
582 => x"25843873",
583 => x"ba387779",
584 => x"24fee238",
585 => x"77537b52",
586 => x"9c1a0851",
587 => x"a41a0859",
588 => x"782d8008",
589 => x"56800880",
590 => x"24fee238",
591 => x"8c1a2280",
592 => x"c0075e7d",
593 => x"8c1b23ff",
594 => x"5574800c",
595 => x"903d0d04",
596 => x"7effa338",
597 => x"ff873975",
598 => x"537b527a",
599 => x"5182f93f",
600 => x"7908167a",
601 => x"0c79518e",
602 => x"b13f8008",
603 => x"cf387c76",
604 => x"315d7cfe",
605 => x"bc38feac",
606 => x"39901a08",
607 => x"7a087131",
608 => x"78117056",
609 => x"5a575280",
610 => x"cfe40851",
611 => x"84943f80",
612 => x"08802eff",
613 => x"a7388008",
614 => x"901b0c80",
615 => x"08167a0c",
616 => x"77941b0c",
617 => x"76881b0c",
618 => x"7656fd99",
619 => x"39790858",
620 => x"901a0878",
621 => x"27833881",
622 => x"54757727",
623 => x"843873b3",
624 => x"38941a08",
625 => x"54737726",
626 => x"80d33873",
627 => x"5378529c",
628 => x"1a0851a4",
629 => x"1a085877",
630 => x"2d800856",
631 => x"80088024",
632 => x"fd83388c",
633 => x"1a2280c0",
634 => x"075e7d8c",
635 => x"1b23ff55",
636 => x"fed73975",
637 => x"53785277",
638 => x"5181dd3f",
639 => x"7908167a",
640 => x"0c79518d",
641 => x"953f8008",
642 => x"802efcd9",
643 => x"388c1a22",
644 => x"80c0075e",
645 => x"7d8c1b23",
646 => x"ff55fead",
647 => x"39767754",
648 => x"79537852",
649 => x"5681b13f",
650 => x"881a0877",
651 => x"31881b0c",
652 => x"7908177a",
653 => x"0cfcae39",
654 => x"fa3d0d7a",
655 => x"79028805",
656 => x"a7053355",
657 => x"53548374",
658 => x"2780df38",
659 => x"71830651",
660 => x"7080d738",
661 => x"71715755",
662 => x"83517582",
663 => x"802913ff",
664 => x"12525670",
665 => x"8025f338",
666 => x"837427bc",
667 => x"38740876",
668 => x"327009f7",
669 => x"fbfdff12",
670 => x"06f88482",
671 => x"81800651",
672 => x"5170802e",
673 => x"98387451",
674 => x"80527033",
675 => x"5772772e",
676 => x"b9388111",
677 => x"81135351",
678 => x"837227ee",
679 => x"38fc1484",
680 => x"16565473",
681 => x"8326c638",
682 => x"7452ff14",
683 => x"5170ff2e",
684 => x"97387133",
685 => x"5472742e",
686 => x"98388112",
687 => x"ff125252",
688 => x"70ff2e09",
689 => x"8106eb38",
690 => x"80517080",
691 => x"0c883d0d",
692 => x"0471800c",
693 => x"883d0d04",
694 => x"fa3d0d78",
695 => x"7a7c7272",
696 => x"72595755",
697 => x"58565774",
698 => x"7727b238",
699 => x"75155176",
700 => x"7127aa38",
701 => x"707618ff",
702 => x"18535353",
703 => x"70ff2e96",
704 => x"38ff12ff",
705 => x"14545272",
706 => x"337234ff",
707 => x"115170ff",
708 => x"2e098106",
709 => x"ec387680",
710 => x"0c883d0d",
711 => x"048f7627",
712 => x"80e63874",
713 => x"77078306",
714 => x"517080dc",
715 => x"38767552",
716 => x"53707084",
717 => x"05520873",
718 => x"70840555",
719 => x"0c727170",
720 => x"84055308",
721 => x"71708405",
722 => x"530c7170",
723 => x"84055308",
724 => x"71708405",
725 => x"530c7170",
726 => x"84055308",
727 => x"71708405",
728 => x"530cf015",
729 => x"5553738f",
730 => x"26c73883",
731 => x"74279538",
732 => x"70708405",
733 => x"52087370",
734 => x"8405550c",
735 => x"fc145473",
736 => x"8326ed38",
737 => x"72715452",
738 => x"ff145170",
739 => x"ff2eff86",
740 => x"38727081",
741 => x"05543372",
742 => x"70810554",
743 => x"34ff1151",
744 => x"ea39ef3d",
745 => x"0d636567",
746 => x"405d427b",
747 => x"802e8582",
748 => x"386151a9",
749 => x"e73ff81c",
750 => x"70841208",
751 => x"70fc0670",
752 => x"628b0570",
753 => x"f8064159",
754 => x"455c5f41",
755 => x"57967427",
756 => x"82c53880",
757 => x"7b247e7c",
758 => x"26075880",
759 => x"5477742e",
760 => x"09810682",
761 => x"ab38787b",
762 => x"2581fe38",
763 => x"781780d7",
764 => x"a00b8805",
765 => x"085b5679",
766 => x"762e84c5",
767 => x"38841608",
768 => x"70fe0617",
769 => x"84110881",
770 => x"06415555",
771 => x"7e828d38",
772 => x"74fc0658",
773 => x"79762e84",
774 => x"e3387818",
775 => x"5f7e7b25",
776 => x"81ff387c",
777 => x"81065473",
778 => x"82c13876",
779 => x"77083184",
780 => x"1108fc06",
781 => x"56577580",
782 => x"2e913879",
783 => x"762e84f0",
784 => x"38741819",
785 => x"58777b25",
786 => x"84913876",
787 => x"802e829b",
788 => x"38781556",
789 => x"7a762482",
790 => x"92388c17",
791 => x"08881808",
792 => x"718c120c",
793 => x"88120c5e",
794 => x"75598817",
795 => x"61fc055b",
796 => x"5679a426",
797 => x"85ff387b",
798 => x"76595593",
799 => x"7a2780c9",
800 => x"387b7084",
801 => x"055d087c",
802 => x"56760c74",
803 => x"70840556",
804 => x"088c180c",
805 => x"9017589b",
806 => x"7a27ae38",
807 => x"74708405",
808 => x"5608780c",
809 => x"74708405",
810 => x"56089418",
811 => x"0c981758",
812 => x"a37a2795",
813 => x"38747084",
814 => x"05560878",
815 => x"0c747084",
816 => x"0556089c",
817 => x"180ca017",
818 => x"58747084",
819 => x"05560875",
820 => x"5f787084",
821 => x"055a0c77",
822 => x"7e708405",
823 => x"40087170",
824 => x"8405530c",
825 => x"7e08710c",
826 => x"5d787b31",
827 => x"56758f26",
828 => x"80c93884",
829 => x"17088106",
830 => x"79078418",
831 => x"0c781784",
832 => x"11088107",
833 => x"84120c5b",
834 => x"6151a791",
835 => x"3f881754",
836 => x"73800c93",
837 => x"3d0d0490",
838 => x"5bfdb839",
839 => x"7756fe83",
840 => x"398c1608",
841 => x"88170871",
842 => x"8c120c88",
843 => x"120c587e",
844 => x"707c3157",
845 => x"598f7627",
846 => x"ffb9387a",
847 => x"17841808",
848 => x"81067c07",
849 => x"84190c76",
850 => x"81078412",
851 => x"0c761184",
852 => x"11088107",
853 => x"84120c5b",
854 => x"88055261",
855 => x"518fda3f",
856 => x"6151a6b9",
857 => x"3f881754",
858 => x"ffa6397d",
859 => x"52615197",
860 => x"d73f8008",
861 => x"5a800880",
862 => x"2e81ab38",
863 => x"8008f805",
864 => x"60840508",
865 => x"fe066105",
866 => x"58557477",
867 => x"2e83f238",
868 => x"fc195877",
869 => x"a42681b0",
870 => x"387b8008",
871 => x"56579378",
872 => x"2780dc38",
873 => x"7b707084",
874 => x"05520880",
875 => x"08708405",
876 => x"800c0c80",
877 => x"08717084",
878 => x"0553085d",
879 => x"567b7670",
880 => x"8405580c",
881 => x"579b7827",
882 => x"b6387670",
883 => x"84055808",
884 => x"75708405",
885 => x"570c7670",
886 => x"84055808",
887 => x"75708405",
888 => x"570ca378",
889 => x"27993876",
890 => x"70840558",
891 => x"08757084",
892 => x"05570c76",
893 => x"70840558",
894 => x"08757084",
895 => x"05570c76",
896 => x"70840558",
897 => x"08775e75",
898 => x"70840557",
899 => x"0c747d70",
900 => x"84055f08",
901 => x"71708405",
902 => x"530c7d08",
903 => x"710c5f7b",
904 => x"5261518e",
905 => x"943f6151",
906 => x"a4f33f79",
907 => x"800c933d",
908 => x"0d047d52",
909 => x"61519690",
910 => x"3f800880",
911 => x"0c933d0d",
912 => x"04841608",
913 => x"55fbc939",
914 => x"77537b52",
915 => x"800851a2",
916 => x"a53f7b52",
917 => x"61518de1",
918 => x"3fcc398c",
919 => x"16088817",
920 => x"08718c12",
921 => x"0c88120c",
922 => x"5d8c1708",
923 => x"88180871",
924 => x"8c120c88",
925 => x"120c5977",
926 => x"59fbef39",
927 => x"7818901c",
928 => x"40557e75",
929 => x"24fb9c38",
930 => x"7a177080",
931 => x"d7a00b88",
932 => x"050c757c",
933 => x"31810784",
934 => x"120c5684",
935 => x"17088106",
936 => x"7b078418",
937 => x"0c6151a3",
938 => x"f43f8817",
939 => x"54fce139",
940 => x"74181990",
941 => x"1c5e5a7c",
942 => x"7a24fb8f",
943 => x"388c1708",
944 => x"88180871",
945 => x"8c120c88",
946 => x"120c5e88",
947 => x"1761fc05",
948 => x"575975a4",
949 => x"2681b638",
950 => x"7b795955",
951 => x"93762780",
952 => x"c9387b70",
953 => x"84055d08",
954 => x"7c56790c",
955 => x"74708405",
956 => x"56088c18",
957 => x"0c901758",
958 => x"9b7627ae",
959 => x"38747084",
960 => x"05560878",
961 => x"0c747084",
962 => x"05560894",
963 => x"180c9817",
964 => x"58a37627",
965 => x"95387470",
966 => x"84055608",
967 => x"780c7470",
968 => x"84055608",
969 => x"9c180ca0",
970 => x"17587470",
971 => x"84055608",
972 => x"75417870",
973 => x"84055a0c",
974 => x"77607084",
975 => x"05420871",
976 => x"70840553",
977 => x"0c600871",
978 => x"0c5e7a17",
979 => x"7080d7a0",
980 => x"0b88050c",
981 => x"7a7c3181",
982 => x"0784120c",
983 => x"58841708",
984 => x"81067b07",
985 => x"84180c61",
986 => x"51a2b23f",
987 => x"78547380",
988 => x"0c933d0d",
989 => x"0479537b",
990 => x"5275519f",
991 => x"f93ffae9",
992 => x"39841508",
993 => x"fc061960",
994 => x"5859fadd",
995 => x"3975537b",
996 => x"5278519f",
997 => x"e13f7a17",
998 => x"7080d7a0",
999 => x"0b88050c",
1000 => x"7a7c3181",
1001 => x"0784120c",
1002 => x"58841708",
1003 => x"81067b07",
1004 => x"84180c61",
1005 => x"51a1e63f",
1006 => x"7854ffb2",
1007 => x"39fa3d0d",
1008 => x"7880cfe4",
1009 => x"085455b8",
1010 => x"1308802e",
1011 => x"81af388c",
1012 => x"15227083",
1013 => x"ffff0670",
1014 => x"832a8132",
1015 => x"81065555",
1016 => x"5672802e",
1017 => x"80da3873",
1018 => x"842a8132",
1019 => x"810657ff",
1020 => x"537680f2",
1021 => x"3873822a",
1022 => x"81065473",
1023 => x"802eb938",
1024 => x"b0150854",
1025 => x"73802e9c",
1026 => x"3880c015",
1027 => x"5373732e",
1028 => x"8f387352",
1029 => x"80cfe408",
1030 => x"518a9e3f",
1031 => x"8c152256",
1032 => x"76b0160c",
1033 => x"75db0657",
1034 => x"768c1623",
1035 => x"800b8416",
1036 => x"0c901508",
1037 => x"750c7656",
1038 => x"75880754",
1039 => x"738c1623",
1040 => x"90150880",
1041 => x"2ebf388c",
1042 => x"15227081",
1043 => x"06555373",
1044 => x"9c38720a",
1045 => x"100a8106",
1046 => x"56758538",
1047 => x"94150854",
1048 => x"7388160c",
1049 => x"80537280",
1050 => x"0c883d0d",
1051 => x"04800b88",
1052 => x"160c9415",
1053 => x"08309816",
1054 => x"0c8053ea",
1055 => x"39725182",
1056 => x"a63ffecb",
1057 => x"3974518f",
1058 => x"bc3f8c15",
1059 => x"22708106",
1060 => x"55537380",
1061 => x"2effbb38",
1062 => x"d439f83d",
1063 => x"0d7a5776",
1064 => x"802e8197",
1065 => x"3880cfe4",
1066 => x"0854b814",
1067 => x"08802e80",
1068 => x"eb388c17",
1069 => x"2270902b",
1070 => x"70902c70",
1071 => x"832a8132",
1072 => x"81065b5b",
1073 => x"57557780",
1074 => x"cb389017",
1075 => x"08567580",
1076 => x"2e80c138",
1077 => x"76087631",
1078 => x"76780c79",
1079 => x"83065555",
1080 => x"73853894",
1081 => x"17085877",
1082 => x"88180c80",
1083 => x"7525a538",
1084 => x"74537552",
1085 => x"9c170851",
1086 => x"a4170854",
1087 => x"732d800b",
1088 => x"80082580",
1089 => x"c9388008",
1090 => x"16758008",
1091 => x"31565674",
1092 => x"8024dd38",
1093 => x"800b800c",
1094 => x"8a3d0d04",
1095 => x"73518187",
1096 => x"3f8c1722",
1097 => x"70902b70",
1098 => x"902c7083",
1099 => x"2a813281",
1100 => x"065b5b57",
1101 => x"5577dd38",
1102 => x"ff9039a1",
1103 => x"9a5280cf",
1104 => x"e408518c",
1105 => x"d03f8008",
1106 => x"800c8a3d",
1107 => x"0d048c17",
1108 => x"2280c007",
1109 => x"58778c18",
1110 => x"23ff0b80",
1111 => x"0c8a3d0d",
1112 => x"04fa3d0d",
1113 => x"797080dc",
1114 => x"298c1154",
1115 => x"7a535657",
1116 => x"8fd63f80",
1117 => x"08800855",
1118 => x"56800880",
1119 => x"2ea23880",
1120 => x"088c0554",
1121 => x"800b8008",
1122 => x"0c768008",
1123 => x"84050c73",
1124 => x"80088805",
1125 => x"0c745380",
1126 => x"5273519c",
1127 => x"f53f7554",
1128 => x"73800c88",
1129 => x"3d0d0470",
1130 => x"707074a8",
1131 => x"e60bbc12",
1132 => x"0c53810b",
1133 => x"b8140c80",
1134 => x"0b84dc14",
1135 => x"0c830b84",
1136 => x"e0140c84",
1137 => x"e81384e4",
1138 => x"140c8413",
1139 => x"08518070",
1140 => x"720c7084",
1141 => x"130c7088",
1142 => x"130c5284",
1143 => x"0b8c1223",
1144 => x"718e1223",
1145 => x"7190120c",
1146 => x"7194120c",
1147 => x"7198120c",
1148 => x"709c120c",
1149 => x"80c1d50b",
1150 => x"a0120c80",
1151 => x"c2a10ba4",
1152 => x"120c80c3",
1153 => x"9d0ba812",
1154 => x"0c80c3ee",
1155 => x"0bac120c",
1156 => x"88130872",
1157 => x"710c7284",
1158 => x"120c7288",
1159 => x"120c5189",
1160 => x"0b8c1223",
1161 => x"810b8e12",
1162 => x"23719012",
1163 => x"0c719412",
1164 => x"0c719812",
1165 => x"0c709c12",
1166 => x"0c80c1d5",
1167 => x"0ba0120c",
1168 => x"80c2a10b",
1169 => x"a4120c80",
1170 => x"c39d0ba8",
1171 => x"120c80c3",
1172 => x"ee0bac12",
1173 => x"0c8c1308",
1174 => x"72710c72",
1175 => x"84120c72",
1176 => x"88120c51",
1177 => x"8a0b8c12",
1178 => x"23820b8e",
1179 => x"12237190",
1180 => x"120c7194",
1181 => x"120c7198",
1182 => x"120c709c",
1183 => x"120c80c1",
1184 => x"d50ba012",
1185 => x"0c80c2a1",
1186 => x"0ba4120c",
1187 => x"80c39d0b",
1188 => x"a8120c80",
1189 => x"c3ee0bac",
1190 => x"120c5050",
1191 => x"5004f83d",
1192 => x"0d7a80cf",
1193 => x"e408b811",
1194 => x"08575758",
1195 => x"7481ec38",
1196 => x"a8e60bbc",
1197 => x"170c810b",
1198 => x"b8170c74",
1199 => x"84dc170c",
1200 => x"830b84e0",
1201 => x"170c84e8",
1202 => x"1684e417",
1203 => x"0c841608",
1204 => x"75710c75",
1205 => x"84120c75",
1206 => x"88120c59",
1207 => x"840b8c1a",
1208 => x"23748e1a",
1209 => x"2374901a",
1210 => x"0c74941a",
1211 => x"0c74981a",
1212 => x"0c789c1a",
1213 => x"0c80c1d5",
1214 => x"0ba01a0c",
1215 => x"80c2a10b",
1216 => x"a41a0c80",
1217 => x"c39d0ba8",
1218 => x"1a0c80c3",
1219 => x"ee0bac1a",
1220 => x"0c881608",
1221 => x"75710c75",
1222 => x"84120c75",
1223 => x"88120c57",
1224 => x"890b8c18",
1225 => x"23810b8e",
1226 => x"18237490",
1227 => x"180c7494",
1228 => x"180c7498",
1229 => x"180c769c",
1230 => x"180c80c1",
1231 => x"d50ba018",
1232 => x"0c80c2a1",
1233 => x"0ba4180c",
1234 => x"80c39d0b",
1235 => x"a8180c80",
1236 => x"c3ee0bac",
1237 => x"180c8c16",
1238 => x"0875710c",
1239 => x"7584120c",
1240 => x"7588120c",
1241 => x"548a0b8c",
1242 => x"1523820b",
1243 => x"8e152374",
1244 => x"90150c74",
1245 => x"94150c74",
1246 => x"98150c73",
1247 => x"9c150c80",
1248 => x"c1d50ba0",
1249 => x"150c80c2",
1250 => x"a10ba415",
1251 => x"0c80c39d",
1252 => x"0ba8150c",
1253 => x"80c3ee0b",
1254 => x"ac150c84",
1255 => x"dc168811",
1256 => x"08841208",
1257 => x"ff055757",
1258 => x"57807524",
1259 => x"9f388c16",
1260 => x"2270902b",
1261 => x"70902c51",
1262 => x"55597380",
1263 => x"2e80ed38",
1264 => x"80dc16ff",
1265 => x"16565674",
1266 => x"8025e338",
1267 => x"76085574",
1268 => x"802e8f38",
1269 => x"74881108",
1270 => x"841208ff",
1271 => x"05575757",
1272 => x"c83982fc",
1273 => x"5277518a",
1274 => x"df3f8008",
1275 => x"80085556",
1276 => x"8008802e",
1277 => x"a3388008",
1278 => x"8c057580",
1279 => x"080c5484",
1280 => x"0b800884",
1281 => x"050c7380",
1282 => x"0888050c",
1283 => x"82f05374",
1284 => x"52735197",
1285 => x"fd3f7554",
1286 => x"7374780c",
1287 => x"5573ffb4",
1288 => x"388c780c",
1289 => x"800b800c",
1290 => x"8a3d0d04",
1291 => x"810b8c17",
1292 => x"2373760c",
1293 => x"7388170c",
1294 => x"7384170c",
1295 => x"7390170c",
1296 => x"7394170c",
1297 => x"7398170c",
1298 => x"ff0b8e17",
1299 => x"2373b017",
1300 => x"0c73b417",
1301 => x"0c7380c4",
1302 => x"170c7380",
1303 => x"c8170c75",
1304 => x"800c8a3d",
1305 => x"0d047070",
1306 => x"a19a5273",
1307 => x"5186a63f",
1308 => x"50500470",
1309 => x"70a19a52",
1310 => x"80cfe408",
1311 => x"5186963f",
1312 => x"505004fb",
1313 => x"3d0d7770",
1314 => x"52569890",
1315 => x"3f80d7a0",
1316 => x"0b880508",
1317 => x"841108fc",
1318 => x"06707b31",
1319 => x"9fef05e0",
1320 => x"8006e080",
1321 => x"05525555",
1322 => x"a0807524",
1323 => x"94388052",
1324 => x"755197ea",
1325 => x"3f80d7a8",
1326 => x"08145372",
1327 => x"80082e8f",
1328 => x"38755197",
1329 => x"d83f8053",
1330 => x"72800c87",
1331 => x"3d0d0474",
1332 => x"30527551",
1333 => x"97c83f80",
1334 => x"08ff2ea8",
1335 => x"3880d7a0",
1336 => x"0b880508",
1337 => x"74763181",
1338 => x"0784120c",
1339 => x"5380d6e4",
1340 => x"08753180",
1341 => x"d6e40c75",
1342 => x"5197a23f",
1343 => x"810b800c",
1344 => x"873d0d04",
1345 => x"80527551",
1346 => x"97943f80",
1347 => x"d7a00b88",
1348 => x"05088008",
1349 => x"71315454",
1350 => x"8f7325ff",
1351 => x"a4388008",
1352 => x"80d79408",
1353 => x"3180d6e4",
1354 => x"0c728107",
1355 => x"84150c75",
1356 => x"5196ea3f",
1357 => x"8053ff90",
1358 => x"39f73d0d",
1359 => x"7b7d545a",
1360 => x"72802e82",
1361 => x"83387951",
1362 => x"96d23ff8",
1363 => x"13841108",
1364 => x"70fe0670",
1365 => x"13841108",
1366 => x"fc065c57",
1367 => x"58545780",
1368 => x"d7a80874",
1369 => x"2e82de38",
1370 => x"7784150c",
1371 => x"80738106",
1372 => x"56597479",
1373 => x"2e81d538",
1374 => x"77148411",
1375 => x"08810656",
1376 => x"5374a038",
1377 => x"77165678",
1378 => x"81e63888",
1379 => x"14085574",
1380 => x"80d7a82e",
1381 => x"82f9388c",
1382 => x"1408708c",
1383 => x"170c7588",
1384 => x"120c5875",
1385 => x"81078418",
1386 => x"0c751776",
1387 => x"710c5478",
1388 => x"81913883",
1389 => x"ff762781",
1390 => x"c8387589",
1391 => x"2a76832a",
1392 => x"54547380",
1393 => x"2ebf3875",
1394 => x"862ab805",
1395 => x"53847427",
1396 => x"b43880db",
1397 => x"14539474",
1398 => x"27ab3875",
1399 => x"8c2a80ee",
1400 => x"055380d4",
1401 => x"74279e38",
1402 => x"758f2a80",
1403 => x"f7055382",
1404 => x"d4742791",
1405 => x"3875922a",
1406 => x"80fc0553",
1407 => x"8ad47427",
1408 => x"843880fe",
1409 => x"53721010",
1410 => x"1080d7a0",
1411 => x"05881108",
1412 => x"55557375",
1413 => x"2e82bf38",
1414 => x"841408fc",
1415 => x"06597579",
1416 => x"278d3888",
1417 => x"14085473",
1418 => x"752e0981",
1419 => x"06ea388c",
1420 => x"1408708c",
1421 => x"190c7488",
1422 => x"190c7788",
1423 => x"120c5576",
1424 => x"8c150c79",
1425 => x"5194d63f",
1426 => x"8b3d0d04",
1427 => x"76087771",
1428 => x"31587605",
1429 => x"88180856",
1430 => x"567480d7",
1431 => x"a82e80e0",
1432 => x"388c1708",
1433 => x"708c170c",
1434 => x"7588120c",
1435 => x"53fe8939",
1436 => x"8814088c",
1437 => x"1508708c",
1438 => x"130c5988",
1439 => x"190cfea3",
1440 => x"3975832a",
1441 => x"70545480",
1442 => x"74248198",
1443 => x"3872822c",
1444 => x"81712b80",
1445 => x"d7a40807",
1446 => x"80d7a00b",
1447 => x"84050c74",
1448 => x"10101080",
1449 => x"d7a00588",
1450 => x"1108718c",
1451 => x"1b0c7088",
1452 => x"1b0c7988",
1453 => x"130c565a",
1454 => x"55768c15",
1455 => x"0cff8439",
1456 => x"8159fdb4",
1457 => x"39771673",
1458 => x"81065455",
1459 => x"72983876",
1460 => x"08777131",
1461 => x"5875058c",
1462 => x"18088819",
1463 => x"08718c12",
1464 => x"0c88120c",
1465 => x"55557481",
1466 => x"0784180c",
1467 => x"7680d7a0",
1468 => x"0b88050c",
1469 => x"80d79c08",
1470 => x"7526fec7",
1471 => x"3880d798",
1472 => x"08527951",
1473 => x"fafd3f79",
1474 => x"5193923f",
1475 => x"feba3981",
1476 => x"778c170c",
1477 => x"7788170c",
1478 => x"758c190c",
1479 => x"7588190c",
1480 => x"59fd8039",
1481 => x"83147082",
1482 => x"2c81712b",
1483 => x"80d7a408",
1484 => x"0780d7a0",
1485 => x"0b84050c",
1486 => x"75101010",
1487 => x"80d7a005",
1488 => x"88110871",
1489 => x"8c1c0c70",
1490 => x"881c0c7a",
1491 => x"88130c57",
1492 => x"5b5653fe",
1493 => x"e4398073",
1494 => x"24a33872",
1495 => x"822c8171",
1496 => x"2b80d7a4",
1497 => x"080780d7",
1498 => x"a00b8405",
1499 => x"0c58748c",
1500 => x"180c7388",
1501 => x"180c7688",
1502 => x"160cfdc3",
1503 => x"39831370",
1504 => x"822c8171",
1505 => x"2b80d7a4",
1506 => x"080780d7",
1507 => x"a00b8405",
1508 => x"0c5953da",
1509 => x"39f93d0d",
1510 => x"797b5853",
1511 => x"800b80cf",
1512 => x"e4085356",
1513 => x"72722ebc",
1514 => x"3884dc13",
1515 => x"5574762e",
1516 => x"b3388815",
1517 => x"08841608",
1518 => x"ff055454",
1519 => x"80732499",
1520 => x"388c1422",
1521 => x"70902b53",
1522 => x"587180d4",
1523 => x"3880dc14",
1524 => x"ff145454",
1525 => x"728025e9",
1526 => x"38740855",
1527 => x"74d43880",
1528 => x"cfe40852",
1529 => x"84dc1255",
1530 => x"74802ead",
1531 => x"38881508",
1532 => x"841608ff",
1533 => x"05545480",
1534 => x"73249838",
1535 => x"8c142270",
1536 => x"902b5358",
1537 => x"71ad3880",
1538 => x"dc14ff14",
1539 => x"54547280",
1540 => x"25ea3874",
1541 => x"085574d5",
1542 => x"3875800c",
1543 => x"893d0d04",
1544 => x"7351762d",
1545 => x"75800807",
1546 => x"80dc15ff",
1547 => x"15555556",
1548 => x"ffa23973",
1549 => x"51762d75",
1550 => x"80080780",
1551 => x"dc15ff15",
1552 => x"555556ca",
1553 => x"39ea3d0d",
1554 => x"688c1122",
1555 => x"700a100a",
1556 => x"81065758",
1557 => x"567480e4",
1558 => x"388e1622",
1559 => x"70902b70",
1560 => x"902c5155",
1561 => x"58807424",
1562 => x"b138983d",
1563 => x"c4055373",
1564 => x"5280cfe4",
1565 => x"08519481",
1566 => x"3f800b80",
1567 => x"08249738",
1568 => x"7983e080",
1569 => x"06547380",
1570 => x"c0802e81",
1571 => x"8f387382",
1572 => x"80802e81",
1573 => x"91388c16",
1574 => x"22577690",
1575 => x"80075473",
1576 => x"8c172388",
1577 => x"805280cf",
1578 => x"e4085181",
1579 => x"9b3f8008",
1580 => x"9d388c16",
1581 => x"22820755",
1582 => x"748c1723",
1583 => x"80c31670",
1584 => x"770c9017",
1585 => x"0c810b94",
1586 => x"170c983d",
1587 => x"0d0480cf",
1588 => x"e408a8e6",
1589 => x"0bbc120c",
1590 => x"588c1622",
1591 => x"81800754",
1592 => x"738c1723",
1593 => x"8008760c",
1594 => x"80089017",
1595 => x"0c88800b",
1596 => x"94170c74",
1597 => x"802ed338",
1598 => x"8e162270",
1599 => x"902b7090",
1600 => x"2c535654",
1601 => x"9afe3f80",
1602 => x"08802eff",
1603 => x"bd388c16",
1604 => x"22810757",
1605 => x"768c1723",
1606 => x"983d0d04",
1607 => x"810b8c17",
1608 => x"225855fe",
1609 => x"f539a816",
1610 => x"0880c39d",
1611 => x"2e098106",
1612 => x"fee4388c",
1613 => x"16228880",
1614 => x"0754738c",
1615 => x"17238880",
1616 => x"0b80cc17",
1617 => x"0cfedc39",
1618 => x"f43d0d7e",
1619 => x"608b1170",
1620 => x"f8065b55",
1621 => x"555d7296",
1622 => x"26833890",
1623 => x"58807824",
1624 => x"74792607",
1625 => x"55805474",
1626 => x"742e0981",
1627 => x"0680ca38",
1628 => x"7c518ea8",
1629 => x"3f7783f7",
1630 => x"2680c538",
1631 => x"77832a70",
1632 => x"10101080",
1633 => x"d7a0058c",
1634 => x"11085858",
1635 => x"5475772e",
1636 => x"81f03884",
1637 => x"1608fc06",
1638 => x"8c170888",
1639 => x"1808718c",
1640 => x"120c8812",
1641 => x"0c5b7605",
1642 => x"84110881",
1643 => x"0784120c",
1644 => x"537c518d",
1645 => x"e83f8816",
1646 => x"5473800c",
1647 => x"8e3d0d04",
1648 => x"77892a78",
1649 => x"832a5854",
1650 => x"73802ebf",
1651 => x"3877862a",
1652 => x"b8055784",
1653 => x"7427b438",
1654 => x"80db1457",
1655 => x"947427ab",
1656 => x"38778c2a",
1657 => x"80ee0557",
1658 => x"80d47427",
1659 => x"9e38778f",
1660 => x"2a80f705",
1661 => x"5782d474",
1662 => x"27913877",
1663 => x"922a80fc",
1664 => x"05578ad4",
1665 => x"74278438",
1666 => x"80fe5776",
1667 => x"10101080",
1668 => x"d7a0058c",
1669 => x"11085653",
1670 => x"74732ea3",
1671 => x"38841508",
1672 => x"fc067079",
1673 => x"31555673",
1674 => x"8f2488e4",
1675 => x"38738025",
1676 => x"88e6388c",
1677 => x"15085574",
1678 => x"732e0981",
1679 => x"06df3881",
1680 => x"175980d7",
1681 => x"b0085675",
1682 => x"80d7a82e",
1683 => x"82cc3884",
1684 => x"1608fc06",
1685 => x"70793155",
1686 => x"55738f24",
1687 => x"bb3880d7",
1688 => x"a80b80d7",
1689 => x"b40c80d7",
1690 => x"a80b80d7",
1691 => x"b00c8074",
1692 => x"2480db38",
1693 => x"74168411",
1694 => x"08810784",
1695 => x"120c53fe",
1696 => x"b0398816",
1697 => x"8c110857",
1698 => x"5975792e",
1699 => x"098106fe",
1700 => x"82388214",
1701 => x"59ffab39",
1702 => x"77167881",
1703 => x"0784180c",
1704 => x"7080d7b4",
1705 => x"0c7080d7",
1706 => x"b00c80d7",
1707 => x"a80b8c12",
1708 => x"0c8c1108",
1709 => x"88120c74",
1710 => x"81078412",
1711 => x"0c740574",
1712 => x"710c5b7c",
1713 => x"518bd63f",
1714 => x"881654fd",
1715 => x"ec3983ff",
1716 => x"75278391",
1717 => x"3874892a",
1718 => x"75832a54",
1719 => x"5473802e",
1720 => x"bf387486",
1721 => x"2ab80553",
1722 => x"847427b4",
1723 => x"3880db14",
1724 => x"53947427",
1725 => x"ab38748c",
1726 => x"2a80ee05",
1727 => x"5380d474",
1728 => x"279e3874",
1729 => x"8f2a80f7",
1730 => x"055382d4",
1731 => x"74279138",
1732 => x"74922a80",
1733 => x"fc05538a",
1734 => x"d4742784",
1735 => x"3880fe53",
1736 => x"72101010",
1737 => x"80d7a005",
1738 => x"88110855",
1739 => x"5773772e",
1740 => x"868b3884",
1741 => x"1408fc06",
1742 => x"5b747b27",
1743 => x"8d388814",
1744 => x"08547377",
1745 => x"2e098106",
1746 => x"ea388c14",
1747 => x"0880d7a0",
1748 => x"0b840508",
1749 => x"718c190c",
1750 => x"7588190c",
1751 => x"7788130c",
1752 => x"5c57758c",
1753 => x"150c7853",
1754 => x"80792483",
1755 => x"98387282",
1756 => x"2c81712b",
1757 => x"5656747b",
1758 => x"2680ca38",
1759 => x"7a750657",
1760 => x"7682a338",
1761 => x"78fc0684",
1762 => x"05597410",
1763 => x"707c0655",
1764 => x"55738292",
1765 => x"38841959",
1766 => x"f13980d7",
1767 => x"a00b8405",
1768 => x"0879545b",
1769 => x"788025c6",
1770 => x"3882da39",
1771 => x"74097b06",
1772 => x"7080d7a0",
1773 => x"0b84050c",
1774 => x"5b741055",
1775 => x"747b2685",
1776 => x"387485bc",
1777 => x"3880d7a0",
1778 => x"0b880508",
1779 => x"70841208",
1780 => x"fc06707b",
1781 => x"317b7226",
1782 => x"8f722507",
1783 => x"5d575c5c",
1784 => x"5578802e",
1785 => x"80d93879",
1786 => x"1580d798",
1787 => x"08199011",
1788 => x"59545680",
1789 => x"d79408ff",
1790 => x"2e8838a0",
1791 => x"8f13e080",
1792 => x"06577652",
1793 => x"7c518996",
1794 => x"3f800854",
1795 => x"8008ff2e",
1796 => x"90388008",
1797 => x"762782a7",
1798 => x"387480d7",
1799 => x"a02e829f",
1800 => x"3880d7a0",
1801 => x"0b880508",
1802 => x"55841508",
1803 => x"fc067079",
1804 => x"31797226",
1805 => x"8f722507",
1806 => x"5d555a7a",
1807 => x"83f23877",
1808 => x"81078416",
1809 => x"0c771570",
1810 => x"80d7a00b",
1811 => x"88050c74",
1812 => x"81078412",
1813 => x"0c567c51",
1814 => x"88c33f88",
1815 => x"15547380",
1816 => x"0c8e3d0d",
1817 => x"0474832a",
1818 => x"70545480",
1819 => x"7424819b",
1820 => x"3872822c",
1821 => x"81712b80",
1822 => x"d7a40807",
1823 => x"7080d7a0",
1824 => x"0b84050c",
1825 => x"75101010",
1826 => x"80d7a005",
1827 => x"88110871",
1828 => x"8c1b0c70",
1829 => x"881b0c79",
1830 => x"88130c57",
1831 => x"555c5575",
1832 => x"8c150cfd",
1833 => x"c1397879",
1834 => x"10101080",
1835 => x"d7a00570",
1836 => x"565b5c8c",
1837 => x"14085675",
1838 => x"742ea338",
1839 => x"841608fc",
1840 => x"06707931",
1841 => x"5853768f",
1842 => x"2483f138",
1843 => x"76802584",
1844 => x"af388c16",
1845 => x"08567574",
1846 => x"2e098106",
1847 => x"df388814",
1848 => x"811a7083",
1849 => x"06555a54",
1850 => x"72c9387b",
1851 => x"83065675",
1852 => x"802efdb8",
1853 => x"38ff1cf8",
1854 => x"1b5b5c88",
1855 => x"1a087a2e",
1856 => x"ea38fdb5",
1857 => x"39831953",
1858 => x"fce43983",
1859 => x"1470822c",
1860 => x"81712b80",
1861 => x"d7a40807",
1862 => x"7080d7a0",
1863 => x"0b84050c",
1864 => x"76101010",
1865 => x"80d7a005",
1866 => x"88110871",
1867 => x"8c1c0c70",
1868 => x"881c0c7a",
1869 => x"88130c58",
1870 => x"535d5653",
1871 => x"fee13980",
1872 => x"d6e40817",
1873 => x"59800876",
1874 => x"2e818b38",
1875 => x"80d79408",
1876 => x"ff2e848e",
1877 => x"38737631",
1878 => x"1980d6e4",
1879 => x"0c738706",
1880 => x"70565372",
1881 => x"802e8838",
1882 => x"88733170",
1883 => x"15555576",
1884 => x"149fff06",
1885 => x"a0807131",
1886 => x"1670547e",
1887 => x"53515386",
1888 => x"9d3f8008",
1889 => x"568008ff",
1890 => x"2e819e38",
1891 => x"80d6e408",
1892 => x"137080d6",
1893 => x"e40c7475",
1894 => x"80d7a00b",
1895 => x"88050c77",
1896 => x"76311581",
1897 => x"07555659",
1898 => x"7a80d7a0",
1899 => x"2e83c038",
1900 => x"798f2682",
1901 => x"ef38810b",
1902 => x"84150c84",
1903 => x"1508fc06",
1904 => x"70793179",
1905 => x"72268f72",
1906 => x"25075d55",
1907 => x"5a7a802e",
1908 => x"fced3880",
1909 => x"db398008",
1910 => x"9fff0655",
1911 => x"74feed38",
1912 => x"7880d6e4",
1913 => x"0c80d7a0",
1914 => x"0b880508",
1915 => x"7a188107",
1916 => x"84120c55",
1917 => x"80d79008",
1918 => x"79278638",
1919 => x"7880d790",
1920 => x"0c80d78c",
1921 => x"087927fc",
1922 => x"a0387880",
1923 => x"d78c0c84",
1924 => x"1508fc06",
1925 => x"70793179",
1926 => x"72268f72",
1927 => x"25075d55",
1928 => x"5a7a802e",
1929 => x"fc993888",
1930 => x"39807457",
1931 => x"53fedd39",
1932 => x"7c5184e9",
1933 => x"3f800b80",
1934 => x"0c8e3d0d",
1935 => x"04807324",
1936 => x"a5387282",
1937 => x"2c81712b",
1938 => x"80d7a408",
1939 => x"077080d7",
1940 => x"a00b8405",
1941 => x"0c5c5a76",
1942 => x"8c170c73",
1943 => x"88170c75",
1944 => x"88180cf9",
1945 => x"fd398313",
1946 => x"70822c81",
1947 => x"712b80d7",
1948 => x"a4080770",
1949 => x"80d7a00b",
1950 => x"84050c5d",
1951 => x"5b53d839",
1952 => x"7a75065c",
1953 => x"7bfc9f38",
1954 => x"84197510",
1955 => x"5659f139",
1956 => x"ff178105",
1957 => x"59f7ab39",
1958 => x"8c150888",
1959 => x"1608718c",
1960 => x"120c8812",
1961 => x"0c597515",
1962 => x"84110881",
1963 => x"0784120c",
1964 => x"587c5183",
1965 => x"e83f8815",
1966 => x"54fba339",
1967 => x"77167881",
1968 => x"0784180c",
1969 => x"8c170888",
1970 => x"1808718c",
1971 => x"120c8812",
1972 => x"0c5c7080",
1973 => x"d7b40c70",
1974 => x"80d7b00c",
1975 => x"80d7a80b",
1976 => x"8c120c8c",
1977 => x"11088812",
1978 => x"0c778107",
1979 => x"84120c77",
1980 => x"0577710c",
1981 => x"557c5183",
1982 => x"a43f8816",
1983 => x"54f5ba39",
1984 => x"72168411",
1985 => x"08810784",
1986 => x"120c588c",
1987 => x"16088817",
1988 => x"08718c12",
1989 => x"0c88120c",
1990 => x"577c5183",
1991 => x"803f8816",
1992 => x"54f59639",
1993 => x"7284150c",
1994 => x"f41af806",
1995 => x"70841d08",
1996 => x"81060784",
1997 => x"1d0c701c",
1998 => x"5556850b",
1999 => x"84150c85",
2000 => x"0b88150c",
2001 => x"8f7627fd",
2002 => x"ab38881b",
2003 => x"527c51eb",
2004 => x"e83f80d7",
2005 => x"a00b8805",
2006 => x"0880d6e4",
2007 => x"085a55fd",
2008 => x"93397880",
2009 => x"d6e40c73",
2010 => x"80d7940c",
2011 => x"fbef3972",
2012 => x"84150cfc",
2013 => x"ff39fb3d",
2014 => x"0d77707a",
2015 => x"7c585553",
2016 => x"568f7527",
2017 => x"80e63872",
2018 => x"76078306",
2019 => x"517080dc",
2020 => x"38757352",
2021 => x"54707084",
2022 => x"05520874",
2023 => x"70840556",
2024 => x"0c737170",
2025 => x"84055308",
2026 => x"71708405",
2027 => x"530c7170",
2028 => x"84055308",
2029 => x"71708405",
2030 => x"530c7170",
2031 => x"84055308",
2032 => x"71708405",
2033 => x"530cf016",
2034 => x"5654748f",
2035 => x"26c73883",
2036 => x"75279538",
2037 => x"70708405",
2038 => x"52087470",
2039 => x"8405560c",
2040 => x"fc155574",
2041 => x"8326ed38",
2042 => x"73715452",
2043 => x"ff155170",
2044 => x"ff2e9838",
2045 => x"72708105",
2046 => x"54337270",
2047 => x"81055434",
2048 => x"ff115170",
2049 => x"ff2e0981",
2050 => x"06ea3875",
2051 => x"800c873d",
2052 => x"0d04fb3d",
2053 => x"0d777a71",
2054 => x"028c05a3",
2055 => x"05335854",
2056 => x"54568373",
2057 => x"2780d438",
2058 => x"75830651",
2059 => x"7080cc38",
2060 => x"74882b75",
2061 => x"07707190",
2062 => x"2b075551",
2063 => x"8f7327a7",
2064 => x"38737270",
2065 => x"8405540c",
2066 => x"71747170",
2067 => x"8405530c",
2068 => x"74717084",
2069 => x"05530c74",
2070 => x"71708405",
2071 => x"530cf014",
2072 => x"5452728f",
2073 => x"26db3883",
2074 => x"73279038",
2075 => x"73727084",
2076 => x"05540cfc",
2077 => x"13537283",
2078 => x"26f238ff",
2079 => x"135170ff",
2080 => x"2e933874",
2081 => x"72708105",
2082 => x"5434ff11",
2083 => x"5170ff2e",
2084 => x"098106ef",
2085 => x"3875800c",
2086 => x"873d0d04",
2087 => x"04047070",
2088 => x"7070800b",
2089 => x"80dfe00c",
2090 => x"765184f3",
2091 => x"3f800853",
2092 => x"8008ff2e",
2093 => x"89387280",
2094 => x"0c505050",
2095 => x"500480df",
2096 => x"e0085473",
2097 => x"802eef38",
2098 => x"7574710c",
2099 => x"5272800c",
2100 => x"50505050",
2101 => x"04f93d0d",
2102 => x"797c557b",
2103 => x"548e1122",
2104 => x"70902b70",
2105 => x"902c5557",
2106 => x"80cfe408",
2107 => x"53585683",
2108 => x"f63f8008",
2109 => x"57800b80",
2110 => x"08249338",
2111 => x"80d01608",
2112 => x"80080580",
2113 => x"d0170c76",
2114 => x"800c893d",
2115 => x"0d048c16",
2116 => x"2283dfff",
2117 => x"0655748c",
2118 => x"17237680",
2119 => x"0c893d0d",
2120 => x"04fa3d0d",
2121 => x"788c1122",
2122 => x"70882a70",
2123 => x"81065157",
2124 => x"585674a9",
2125 => x"388c1622",
2126 => x"83dfff06",
2127 => x"55748c17",
2128 => x"237a5479",
2129 => x"538e1622",
2130 => x"70902b70",
2131 => x"902c5456",
2132 => x"80cfe408",
2133 => x"525681b2",
2134 => x"3f883d0d",
2135 => x"04825480",
2136 => x"538e1622",
2137 => x"70902b70",
2138 => x"902c5456",
2139 => x"80cfe408",
2140 => x"525782bb",
2141 => x"3f8c1622",
2142 => x"83dfff06",
2143 => x"55748c17",
2144 => x"237a5479",
2145 => x"538e1622",
2146 => x"70902b70",
2147 => x"902c5456",
2148 => x"80cfe408",
2149 => x"525680f2",
2150 => x"3f883d0d",
2151 => x"04f93d0d",
2152 => x"797c557b",
2153 => x"548e1122",
2154 => x"70902b70",
2155 => x"902c5557",
2156 => x"80cfe408",
2157 => x"53585681",
2158 => x"f63f8008",
2159 => x"578008ff",
2160 => x"2e99388c",
2161 => x"1622a080",
2162 => x"0755748c",
2163 => x"17238008",
2164 => x"80d0170c",
2165 => x"76800c89",
2166 => x"3d0d048c",
2167 => x"162283df",
2168 => x"ff065574",
2169 => x"8c172376",
2170 => x"800c893d",
2171 => x"0d047070",
2172 => x"70748e11",
2173 => x"2270902b",
2174 => x"70902c55",
2175 => x"51515380",
2176 => x"cfe40851",
2177 => x"bd3f5050",
2178 => x"5004fb3d",
2179 => x"0d800b80",
2180 => x"dfe00c7a",
2181 => x"53795278",
2182 => x"5182ff3f",
2183 => x"80085580",
2184 => x"08ff2e88",
2185 => x"3874800c",
2186 => x"873d0d04",
2187 => x"80dfe008",
2188 => x"5675802e",
2189 => x"f0387776",
2190 => x"710c5474",
2191 => x"800c873d",
2192 => x"0d047070",
2193 => x"7070800b",
2194 => x"80dfe00c",
2195 => x"765184cc",
2196 => x"3f800853",
2197 => x"8008ff2e",
2198 => x"89387280",
2199 => x"0c505050",
2200 => x"500480df",
2201 => x"e0085473",
2202 => x"802eef38",
2203 => x"7574710c",
2204 => x"5272800c",
2205 => x"50505050",
2206 => x"04fc3d0d",
2207 => x"800b80df",
2208 => x"e00c7852",
2209 => x"775187b3",
2210 => x"3f800854",
2211 => x"8008ff2e",
2212 => x"88387380",
2213 => x"0c863d0d",
2214 => x"0480dfe0",
2215 => x"08557480",
2216 => x"2ef03876",
2217 => x"75710c53",
2218 => x"73800c86",
2219 => x"3d0d04fb",
2220 => x"3d0d800b",
2221 => x"80dfe00c",
2222 => x"7a537952",
2223 => x"7851848e",
2224 => x"3f800855",
2225 => x"8008ff2e",
2226 => x"88387480",
2227 => x"0c873d0d",
2228 => x"0480dfe0",
2229 => x"08567580",
2230 => x"2ef03877",
2231 => x"76710c54",
2232 => x"74800c87",
2233 => x"3d0d04fb",
2234 => x"3d0d800b",
2235 => x"80dfe00c",
2236 => x"7a537952",
2237 => x"78518296",
2238 => x"3f800855",
2239 => x"8008ff2e",
2240 => x"88387480",
2241 => x"0c873d0d",
2242 => x"0480dfe0",
2243 => x"08567580",
2244 => x"2ef03877",
2245 => x"76710c54",
2246 => x"74800c87",
2247 => x"3d0d0470",
2248 => x"707080df",
2249 => x"d0088938",
2250 => x"80dfe40b",
2251 => x"80dfd00c",
2252 => x"80dfd008",
2253 => x"75115252",
2254 => x"ff537087",
2255 => x"fb808026",
2256 => x"88387080",
2257 => x"dfd00c71",
2258 => x"5372800c",
2259 => x"50505004",
2260 => x"fd3d0d80",
2261 => x"0b80cfd8",
2262 => x"08545472",
2263 => x"812e9b38",
2264 => x"7380dfd4",
2265 => x"0cc2bf3f",
2266 => x"c1963f80",
2267 => x"dfa85281",
2268 => x"51c3fd3f",
2269 => x"80085186",
2270 => x"c23f7280",
2271 => x"dfd40cc2",
2272 => x"a53fc0fc",
2273 => x"3f80dfa8",
2274 => x"528151c3",
2275 => x"e33f8008",
2276 => x"5186a83f",
2277 => x"00ff3900",
2278 => x"ff39f53d",
2279 => x"0d7e6080",
2280 => x"dfd40870",
2281 => x"5b585b5b",
2282 => x"7580c238",
2283 => x"777a25a1",
2284 => x"38771b70",
2285 => x"337081ff",
2286 => x"06585859",
2287 => x"758a2e98",
2288 => x"387681ff",
2289 => x"0651c1bd",
2290 => x"3f811858",
2291 => x"797824e1",
2292 => x"3879800c",
2293 => x"8d3d0d04",
2294 => x"8d51c1a9",
2295 => x"3f783370",
2296 => x"81ff0652",
2297 => x"57c19e3f",
2298 => x"811858e0",
2299 => x"3979557a",
2300 => x"547d5385",
2301 => x"528d3dfc",
2302 => x"0551c0c6",
2303 => x"3f800856",
2304 => x"85b23f7b",
2305 => x"80080c75",
2306 => x"800c8d3d",
2307 => x"0d04f63d",
2308 => x"0d7d7f80",
2309 => x"dfd40870",
2310 => x"5b585a5a",
2311 => x"7580c138",
2312 => x"777925b3",
2313 => x"38c0b93f",
2314 => x"800881ff",
2315 => x"06708d32",
2316 => x"7030709f",
2317 => x"2a515157",
2318 => x"57768a2e",
2319 => x"80c43875",
2320 => x"802ebf38",
2321 => x"771a5676",
2322 => x"76347651",
2323 => x"c0b73f81",
2324 => x"18587878",
2325 => x"24cf3877",
2326 => x"5675800c",
2327 => x"8c3d0d04",
2328 => x"78557954",
2329 => x"7c538452",
2330 => x"8c3dfc05",
2331 => x"51ffbfd2",
2332 => x"3f800856",
2333 => x"84be3f7a",
2334 => x"80080c75",
2335 => x"800c8c3d",
2336 => x"0d04771a",
2337 => x"598a7934",
2338 => x"8118588d",
2339 => x"51ffbff5",
2340 => x"3f8a51ff",
2341 => x"bfef3f77",
2342 => x"56ffbe39",
2343 => x"fb3d0d80",
2344 => x"dfd40870",
2345 => x"56547388",
2346 => x"3874800c",
2347 => x"873d0d04",
2348 => x"77538352",
2349 => x"873dfc05",
2350 => x"51ffbf86",
2351 => x"3f800854",
2352 => x"83f23f75",
2353 => x"80080c73",
2354 => x"800c873d",
2355 => x"0d04fa3d",
2356 => x"0d80dfd4",
2357 => x"08802ea3",
2358 => x"387a5579",
2359 => x"54785386",
2360 => x"52883dfc",
2361 => x"0551ffbe",
2362 => x"d93f8008",
2363 => x"5683c53f",
2364 => x"7680080c",
2365 => x"75800c88",
2366 => x"3d0d0483",
2367 => x"b73f9d0b",
2368 => x"80080cff",
2369 => x"0b800c88",
2370 => x"3d0d04f7",
2371 => x"3d0d7b7d",
2372 => x"5b59bc53",
2373 => x"80527951",
2374 => x"f5f83f80",
2375 => x"70565798",
2376 => x"56741970",
2377 => x"3370782b",
2378 => x"79078118",
2379 => x"f81a5a58",
2380 => x"59555884",
2381 => x"7524ea38",
2382 => x"767a2384",
2383 => x"19588070",
2384 => x"56579856",
2385 => x"74187033",
2386 => x"70782b79",
2387 => x"078118f8",
2388 => x"1a5a5859",
2389 => x"51548475",
2390 => x"24ea3876",
2391 => x"821b2388",
2392 => x"19588070",
2393 => x"56579856",
2394 => x"74187033",
2395 => x"70782b79",
2396 => x"078118f8",
2397 => x"1a5a5859",
2398 => x"51548475",
2399 => x"24ea3876",
2400 => x"841b0c8c",
2401 => x"19588070",
2402 => x"56579856",
2403 => x"74187033",
2404 => x"70782b79",
2405 => x"078118f8",
2406 => x"1a5a5859",
2407 => x"51548475",
2408 => x"24ea3876",
2409 => x"881b2390",
2410 => x"19588070",
2411 => x"56579856",
2412 => x"74187033",
2413 => x"70782b79",
2414 => x"078118f8",
2415 => x"1a5a5859",
2416 => x"51548475",
2417 => x"24ea3876",
2418 => x"8a1b2394",
2419 => x"19588070",
2420 => x"56579856",
2421 => x"74187033",
2422 => x"70782b79",
2423 => x"078118f8",
2424 => x"1a5a5859",
2425 => x"51548475",
2426 => x"24ea3876",
2427 => x"8c1b2398",
2428 => x"19588070",
2429 => x"56579856",
2430 => x"74187033",
2431 => x"70782b79",
2432 => x"078118f8",
2433 => x"1a5a5859",
2434 => x"51548475",
2435 => x"24ea3876",
2436 => x"8e1b239c",
2437 => x"19588070",
2438 => x"5657b856",
2439 => x"74187033",
2440 => x"70782b79",
2441 => x"078118f8",
2442 => x"1a5a5859",
2443 => x"5a548875",
2444 => x"24ea3876",
2445 => x"901b0c8b",
2446 => x"3d0d04e9",
2447 => x"3d0d6a80",
2448 => x"dfd40857",
2449 => x"57759338",
2450 => x"80c0800b",
2451 => x"84180c75",
2452 => x"ac180c75",
2453 => x"800c993d",
2454 => x"0d04893d",
2455 => x"70556a54",
2456 => x"558a5299",
2457 => x"3dffbc05",
2458 => x"51ffbbd6",
2459 => x"3f800877",
2460 => x"53755256",
2461 => x"fd953fbc",
2462 => x"3f778008",
2463 => x"0c75800c",
2464 => x"993d0d04",
2465 => x"fc3d0d81",
2466 => x"5480dfd4",
2467 => x"08883873",
2468 => x"800c863d",
2469 => x"0d047653",
2470 => x"97b95286",
2471 => x"3dfc0551",
2472 => x"ffbb9f3f",
2473 => x"8008548c",
2474 => x"3f748008",
2475 => x"0c73800c",
2476 => x"863d0d04",
2477 => x"80cfe408",
2478 => x"800c04f7",
2479 => x"3d0d7b80",
2480 => x"cfe40882",
2481 => x"c811085a",
2482 => x"545a7780",
2483 => x"2e80da38",
2484 => x"81881884",
2485 => x"1908ff05",
2486 => x"81712b59",
2487 => x"55598074",
2488 => x"2480ea38",
2489 => x"807424b5",
2490 => x"3873822b",
2491 => x"78118805",
2492 => x"56568180",
2493 => x"19087706",
2494 => x"5372802e",
2495 => x"b6387816",
2496 => x"70085353",
2497 => x"79517408",
2498 => x"53722dff",
2499 => x"14fc17fc",
2500 => x"1779812c",
2501 => x"5a575754",
2502 => x"738025d6",
2503 => x"38770858",
2504 => x"77ffad38",
2505 => x"80cfe408",
2506 => x"53bc1308",
2507 => x"a5387951",
2508 => x"f8e23f74",
2509 => x"0853722d",
2510 => x"ff14fc17",
2511 => x"fc177981",
2512 => x"2c5a5757",
2513 => x"54738025",
2514 => x"ffa838d1",
2515 => x"398057ff",
2516 => x"93397251",
2517 => x"bc130854",
2518 => x"732d7951",
2519 => x"f8b63f70",
2520 => x"7080dfb0",
2521 => x"0bfc0570",
2522 => x"08525270",
2523 => x"ff2e9138",
2524 => x"702dfc12",
2525 => x"70085252",
2526 => x"70ff2e09",
2527 => x"8106f138",
2528 => x"50500404",
2529 => x"ffbb8c3f",
2530 => x"04000000",
2531 => x"00000040",
2532 => x"48656c6c",
2533 => x"6f20776f",
2534 => x"726c6420",
2535 => x"310a0000",
2536 => x"48656c6c",
2537 => x"6f20776f",
2538 => x"726c6420",
2539 => x"320a0000",
2540 => x"0a000000",
2541 => x"43000000",
2542 => x"64756d6d",
2543 => x"792e6578",
2544 => x"65000000",
2545 => x"00ffffff",
2546 => x"ff00ffff",
2547 => x"ffff00ff",
2548 => x"ffffff00",
2549 => x"00000000",
2550 => x"00000000",
2551 => x"00000000",
2552 => x"00002fb8",
2553 => x"000027e8",
2554 => x"00000000",
2555 => x"00002a50",
2556 => x"00002aac",
2557 => x"00002b08",
2558 => x"00000000",
2559 => x"00000000",
2560 => x"00000000",
2561 => x"00000000",
2562 => x"00000000",
2563 => x"00000000",
2564 => x"00000000",
2565 => x"00000000",
2566 => x"00000000",
2567 => x"000027b4",
2568 => x"00000000",
2569 => x"00000000",
2570 => x"00000000",
2571 => x"00000000",
2572 => x"00000000",
2573 => x"00000000",
2574 => x"00000000",
2575 => x"00000000",
2576 => x"00000000",
2577 => x"00000000",
2578 => x"00000000",
2579 => x"00000000",
2580 => x"00000000",
2581 => x"00000000",
2582 => x"00000000",
2583 => x"00000000",
2584 => x"00000000",
2585 => x"00000000",
2586 => x"00000000",
2587 => x"00000000",
2588 => x"00000000",
2589 => x"00000000",
2590 => x"00000000",
2591 => x"00000000",
2592 => x"00000000",
2593 => x"00000000",
2594 => x"00000000",
2595 => x"00000000",
2596 => x"00000001",
2597 => x"330eabcd",
2598 => x"1234e66d",
2599 => x"deec0005",
2600 => x"000b0000",
2601 => x"00000000",
2602 => x"00000000",
2603 => x"00000000",
2604 => x"00000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"00000000",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000000",
2638 => x"00000000",
2639 => x"00000000",
2640 => x"00000000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"ffffffff",
2790 => x"00000000",
2791 => x"00020000",
2792 => x"00000000",
2793 => x"00000000",
2794 => x"00002ba0",
2795 => x"00002ba0",
2796 => x"00002ba8",
2797 => x"00002ba8",
2798 => x"00002bb0",
2799 => x"00002bb0",
2800 => x"00002bb8",
2801 => x"00002bb8",
2802 => x"00002bc0",
2803 => x"00002bc0",
2804 => x"00002bc8",
2805 => x"00002bc8",
2806 => x"00002bd0",
2807 => x"00002bd0",
2808 => x"00002bd8",
2809 => x"00002bd8",
2810 => x"00002be0",
2811 => x"00002be0",
2812 => x"00002be8",
2813 => x"00002be8",
2814 => x"00002bf0",
2815 => x"00002bf0",
2816 => x"00002bf8",
2817 => x"00002bf8",
2818 => x"00002c00",
2819 => x"00002c00",
2820 => x"00002c08",
2821 => x"00002c08",
2822 => x"00002c10",
2823 => x"00002c10",
2824 => x"00002c18",
2825 => x"00002c18",
2826 => x"00002c20",
2827 => x"00002c20",
2828 => x"00002c28",
2829 => x"00002c28",
2830 => x"00002c30",
2831 => x"00002c30",
2832 => x"00002c38",
2833 => x"00002c38",
2834 => x"00002c40",
2835 => x"00002c40",
2836 => x"00002c48",
2837 => x"00002c48",
2838 => x"00002c50",
2839 => x"00002c50",
2840 => x"00002c58",
2841 => x"00002c58",
2842 => x"00002c60",
2843 => x"00002c60",
2844 => x"00002c68",
2845 => x"00002c68",
2846 => x"00002c70",
2847 => x"00002c70",
2848 => x"00002c78",
2849 => x"00002c78",
2850 => x"00002c80",
2851 => x"00002c80",
2852 => x"00002c88",
2853 => x"00002c88",
2854 => x"00002c90",
2855 => x"00002c90",
2856 => x"00002c98",
2857 => x"00002c98",
2858 => x"00002ca0",
2859 => x"00002ca0",
2860 => x"00002ca8",
2861 => x"00002ca8",
2862 => x"00002cb0",
2863 => x"00002cb0",
2864 => x"00002cb8",
2865 => x"00002cb8",
2866 => x"00002cc0",
2867 => x"00002cc0",
2868 => x"00002cc8",
2869 => x"00002cc8",
2870 => x"00002cd0",
2871 => x"00002cd0",
2872 => x"00002cd8",
2873 => x"00002cd8",
2874 => x"00002ce0",
2875 => x"00002ce0",
2876 => x"00002ce8",
2877 => x"00002ce8",
2878 => x"00002cf0",
2879 => x"00002cf0",
2880 => x"00002cf8",
2881 => x"00002cf8",
2882 => x"00002d00",
2883 => x"00002d00",
2884 => x"00002d08",
2885 => x"00002d08",
2886 => x"00002d10",
2887 => x"00002d10",
2888 => x"00002d18",
2889 => x"00002d18",
2890 => x"00002d20",
2891 => x"00002d20",
2892 => x"00002d28",
2893 => x"00002d28",
2894 => x"00002d30",
2895 => x"00002d30",
2896 => x"00002d38",
2897 => x"00002d38",
2898 => x"00002d40",
2899 => x"00002d40",
2900 => x"00002d48",
2901 => x"00002d48",
2902 => x"00002d50",
2903 => x"00002d50",
2904 => x"00002d58",
2905 => x"00002d58",
2906 => x"00002d60",
2907 => x"00002d60",
2908 => x"00002d68",
2909 => x"00002d68",
2910 => x"00002d70",
2911 => x"00002d70",
2912 => x"00002d78",
2913 => x"00002d78",
2914 => x"00002d80",
2915 => x"00002d80",
2916 => x"00002d88",
2917 => x"00002d88",
2918 => x"00002d90",
2919 => x"00002d90",
2920 => x"00002d98",
2921 => x"00002d98",
2922 => x"00002da0",
2923 => x"00002da0",
2924 => x"00002da8",
2925 => x"00002da8",
2926 => x"00002db0",
2927 => x"00002db0",
2928 => x"00002db8",
2929 => x"00002db8",
2930 => x"00002dc0",
2931 => x"00002dc0",
2932 => x"00002dc8",
2933 => x"00002dc8",
2934 => x"00002dd0",
2935 => x"00002dd0",
2936 => x"00002dd8",
2937 => x"00002dd8",
2938 => x"00002de0",
2939 => x"00002de0",
2940 => x"00002de8",
2941 => x"00002de8",
2942 => x"00002df0",
2943 => x"00002df0",
2944 => x"00002df8",
2945 => x"00002df8",
2946 => x"00002e00",
2947 => x"00002e00",
2948 => x"00002e08",
2949 => x"00002e08",
2950 => x"00002e10",
2951 => x"00002e10",
2952 => x"00002e18",
2953 => x"00002e18",
2954 => x"00002e20",
2955 => x"00002e20",
2956 => x"00002e28",
2957 => x"00002e28",
2958 => x"00002e30",
2959 => x"00002e30",
2960 => x"00002e38",
2961 => x"00002e38",
2962 => x"00002e40",
2963 => x"00002e40",
2964 => x"00002e48",
2965 => x"00002e48",
2966 => x"00002e50",
2967 => x"00002e50",
2968 => x"00002e58",
2969 => x"00002e58",
2970 => x"00002e60",
2971 => x"00002e60",
2972 => x"00002e68",
2973 => x"00002e68",
2974 => x"00002e70",
2975 => x"00002e70",
2976 => x"00002e78",
2977 => x"00002e78",
2978 => x"00002e80",
2979 => x"00002e80",
2980 => x"00002e88",
2981 => x"00002e88",
2982 => x"00002e90",
2983 => x"00002e90",
2984 => x"00002e98",
2985 => x"00002e98",
2986 => x"00002ea0",
2987 => x"00002ea0",
2988 => x"00002ea8",
2989 => x"00002ea8",
2990 => x"00002eb0",
2991 => x"00002eb0",
2992 => x"00002eb8",
2993 => x"00002eb8",
2994 => x"00002ec0",
2995 => x"00002ec0",
2996 => x"00002ec8",
2997 => x"00002ec8",
2998 => x"00002ed0",
2999 => x"00002ed0",
3000 => x"00002ed8",
3001 => x"00002ed8",
3002 => x"00002ee0",
3003 => x"00002ee0",
3004 => x"00002ee8",
3005 => x"00002ee8",
3006 => x"00002ef0",
3007 => x"00002ef0",
3008 => x"00002ef8",
3009 => x"00002ef8",
3010 => x"00002f00",
3011 => x"00002f00",
3012 => x"00002f08",
3013 => x"00002f08",
3014 => x"00002f10",
3015 => x"00002f10",
3016 => x"00002f18",
3017 => x"00002f18",
3018 => x"00002f20",
3019 => x"00002f20",
3020 => x"00002f28",
3021 => x"00002f28",
3022 => x"00002f30",
3023 => x"00002f30",
3024 => x"00002f38",
3025 => x"00002f38",
3026 => x"00002f40",
3027 => x"00002f40",
3028 => x"00002f48",
3029 => x"00002f48",
3030 => x"00002f50",
3031 => x"00002f50",
3032 => x"00002f58",
3033 => x"00002f58",
3034 => x"00002f60",
3035 => x"00002f60",
3036 => x"00002f68",
3037 => x"00002f68",
3038 => x"00002f70",
3039 => x"00002f70",
3040 => x"00002f78",
3041 => x"00002f78",
3042 => x"00002f80",
3043 => x"00002f80",
3044 => x"00002f88",
3045 => x"00002f88",
3046 => x"00002f90",
3047 => x"00002f90",
3048 => x"00002f98",
3049 => x"00002f98",
3050 => x"000027b8",
3051 => x"ffffffff",
3052 => x"00000000",
3053 => x"ffffffff",
3054 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
