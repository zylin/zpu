------------------------------------------------------------------------------
----                                                                      ----
----  Single Port RAM that maps to a Xilinx BRAM                          ----
----                                                                      ----
----  http://www.opencores.org/                                           ----
----                                                                      ----
----  Description:                                                        ----
----  This is a program+data memory for the ZPU. It maps to a Xilinx BRAM ----
----                                                                      ----
----  To Do:                                                              ----
----  -                                                                   ----
----                                                                      ----
----  Author:                                                             ----
----    - Salvador E. Tropea, salvador inti.gob.ar                        ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Copyright (c) 2008 Salvador E. Tropea <salvador inti.gob.ar>         ----
---- Copyright (c) 2008 Instituto Nacional de Tecnolog�a Industrial       ----
----                                                                      ----
---- Distributed under the BSD license                                    ----
----                                                                      ----
------------------------------------------------------------------------------
----                                                                      ----
---- Design unit:      SinglePortRAM(Xilinx) (Entity and architecture)    ----
---- File name:        rom_s.in.vhdl (template used)                      ----
---- Note:             None                                               ----
---- Limitations:      None known                                         ----
---- Errors:           None known                                         ----
---- Library:          work                                               ----
---- Dependencies:     IEEE.std_logic_1164                                ----
----                   IEEE.numeric_std                                   ----
---- Target FPGA:      Spartan 3 (XC3S1500-4-FG456)                       ----
---- Language:         VHDL                                               ----
---- Wishbone:         No                                                 ----
---- Synthesis tools:  Xilinx Release 9.2.03i - xst J.39                  ----
---- Simulation tools: GHDL [Sokcho edition] (0.2x)                       ----
---- Text editor:      SETEdit 0.5.x                                      ----
----                                                                      ----
------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity SinglePortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i   : in  std_logic;
      we_i    : in  std_logic;
      re_i    : in  std_logic;
      addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      write_i : in  unsigned(WORD_SIZE-1 downto 0);
      read_o  : out unsigned(WORD_SIZE-1 downto 0);
      busy_o  : out std_logic);
end entity SinglePortRAM;

architecture Xilinx of SinglePortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);
   signal addr_r  : unsigned(BRAM_W-1 downto BYTE_BITS);

   signal ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80f8ec0c",
     3 => x"3a0b0b80",
     4 => x"e7ea0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80e8b72d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80f8",
   162 => x"d8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80ce",
   171 => x"b62d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80cf",
   179 => x"e82d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80f8e80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"83803f80",
   257 => x"e2953f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"ff3d0d0b",
   281 => x"0b8188e0",
   282 => x"08527108",
   283 => x"70882a81",
   284 => x"32708106",
   285 => x"51515170",
   286 => x"f1387372",
   287 => x"0c833d0d",
   288 => x"0480f8e8",
   289 => x"08802ea4",
   290 => x"3880f8ec",
   291 => x"08822ebd",
   292 => x"38838080",
   293 => x"0b0b0b81",
   294 => x"88e00c82",
   295 => x"a0800b81",
   296 => x"88e40c82",
   297 => x"90800b81",
   298 => x"88e80c04",
   299 => x"f8808080",
   300 => x"a40b0b0b",
   301 => x"8188e00c",
   302 => x"f8808082",
   303 => x"800b8188",
   304 => x"e40cf880",
   305 => x"8084800b",
   306 => x"8188e80c",
   307 => x"0480c0a8",
   308 => x"808c0b0b",
   309 => x"0b8188e0",
   310 => x"0c80c0a8",
   311 => x"80940b81",
   312 => x"88e40c0b",
   313 => x"0b80eac8",
   314 => x"0b8188e8",
   315 => x"0c04f23d",
   316 => x"0d608188",
   317 => x"e408565d",
   318 => x"82750c80",
   319 => x"59805a80",
   320 => x"0b8f3d5d",
   321 => x"5b7a1010",
   322 => x"15700871",
   323 => x"08719f2c",
   324 => x"7e852b58",
   325 => x"55557d53",
   326 => x"59579d94",
   327 => x"3f7d7f7a",
   328 => x"72077c72",
   329 => x"07717160",
   330 => x"8105415f",
   331 => x"5d5b5957",
   332 => x"55817b27",
   333 => x"8f38767d",
   334 => x"0c77841e",
   335 => x"0c7c800c",
   336 => x"903d0d04",
   337 => x"8188e408",
   338 => x"55ffba39",
   339 => x"ff3d0d81",
   340 => x"88ec3351",
   341 => x"70a73880",
   342 => x"f8f40870",
   343 => x"08525270",
   344 => x"802e9438",
   345 => x"841280f8",
   346 => x"f40c702d",
   347 => x"80f8f408",
   348 => x"70085252",
   349 => x"70ee3881",
   350 => x"0b8188ec",
   351 => x"34833d0d",
   352 => x"0404803d",
   353 => x"0d0b0b81",
   354 => x"88dc0880",
   355 => x"2e8e380b",
   356 => x"0b0b0b80",
   357 => x"0b802e09",
   358 => x"81068538",
   359 => x"823d0d04",
   360 => x"0b0b8188",
   361 => x"dc510b0b",
   362 => x"0bf4d53f",
   363 => x"823d0d04",
   364 => x"04ff3d0d",
   365 => x"028f0533",
   366 => x"52718a2e",
   367 => x"8a387151",
   368 => x"fd9e3f83",
   369 => x"3d0d048d",
   370 => x"51fd953f",
   371 => x"7151fd90",
   372 => x"3f833d0d",
   373 => x"04ce3d0d",
   374 => x"b53d7070",
   375 => x"84055208",
   376 => x"8bb15c56",
   377 => x"a53d5e5c",
   378 => x"80757081",
   379 => x"05573376",
   380 => x"5b555873",
   381 => x"782e80c1",
   382 => x"388e3d5b",
   383 => x"73a52e09",
   384 => x"810680c5",
   385 => x"38787081",
   386 => x"055a3354",
   387 => x"7380e42e",
   388 => x"81b63873",
   389 => x"80e42480",
   390 => x"c6387380",
   391 => x"e32ea138",
   392 => x"8052a551",
   393 => x"792d8052",
   394 => x"7351792d",
   395 => x"82185878",
   396 => x"7081055a",
   397 => x"335473c4",
   398 => x"3877800c",
   399 => x"b43d0d04",
   400 => x"7b841d83",
   401 => x"1233565d",
   402 => x"57805273",
   403 => x"51792d81",
   404 => x"18797081",
   405 => x"055b3355",
   406 => x"5873ffa0",
   407 => x"38db3973",
   408 => x"80f32e09",
   409 => x"8106ffb8",
   410 => x"387b841d",
   411 => x"7108595d",
   412 => x"56807733",
   413 => x"55567376",
   414 => x"2e8d3881",
   415 => x"16701870",
   416 => x"33575556",
   417 => x"74f538ff",
   418 => x"16558076",
   419 => x"25ffa038",
   420 => x"76708105",
   421 => x"58335480",
   422 => x"52735179",
   423 => x"2d811875",
   424 => x"ff175757",
   425 => x"58807625",
   426 => x"ff853876",
   427 => x"70810558",
   428 => x"33548052",
   429 => x"7351792d",
   430 => x"811875ff",
   431 => x"17575758",
   432 => x"758024cc",
   433 => x"38fee839",
   434 => x"7b841d71",
   435 => x"0870719f",
   436 => x"2c595359",
   437 => x"5d568075",
   438 => x"24819338",
   439 => x"757d7c58",
   440 => x"56548057",
   441 => x"73772e09",
   442 => x"8106b638",
   443 => x"b07b3402",
   444 => x"b505567a",
   445 => x"762e9738",
   446 => x"ff165675",
   447 => x"33757081",
   448 => x"05573481",
   449 => x"17577a76",
   450 => x"2e098106",
   451 => x"eb388075",
   452 => x"34767dff",
   453 => x"12575856",
   454 => x"758024fe",
   455 => x"f338fe8f",
   456 => x"398a5273",
   457 => x"5180c1c0",
   458 => x"3f800880",
   459 => x"eacc0533",
   460 => x"76708105",
   461 => x"58348a52",
   462 => x"7351bffa",
   463 => x"3f800854",
   464 => x"8008802e",
   465 => x"ffad388a",
   466 => x"52735180",
   467 => x"c19a3f80",
   468 => x"0880eacc",
   469 => x"05337670",
   470 => x"81055834",
   471 => x"8a527351",
   472 => x"bfd43f80",
   473 => x"08548008",
   474 => x"ffb738ff",
   475 => x"86397452",
   476 => x"7653b43d",
   477 => x"ffb80551",
   478 => x"978a3fa3",
   479 => x"3d0856fe",
   480 => x"db39803d",
   481 => x"0d80c10b",
   482 => x"81d7b834",
   483 => x"800b81d9",
   484 => x"940c7080",
   485 => x"0c823d0d",
   486 => x"04ff3d0d",
   487 => x"800b81d7",
   488 => x"b8335252",
   489 => x"7080c12e",
   490 => x"99387181",
   491 => x"d9940807",
   492 => x"81d9940c",
   493 => x"80c20b81",
   494 => x"d7bc3470",
   495 => x"800c833d",
   496 => x"0d04810b",
   497 => x"81d99408",
   498 => x"0781d994",
   499 => x"0c80c20b",
   500 => x"81d7bc34",
   501 => x"70800c83",
   502 => x"3d0d04fd",
   503 => x"3d0d7570",
   504 => x"088a0553",
   505 => x"5381d7b8",
   506 => x"33517080",
   507 => x"c12e8b38",
   508 => x"73f33870",
   509 => x"800c853d",
   510 => x"0d04ff12",
   511 => x"7081d7b4",
   512 => x"0831740c",
   513 => x"800c853d",
   514 => x"0d04fc3d",
   515 => x"0d81d7c0",
   516 => x"08557480",
   517 => x"2e8c3876",
   518 => x"7508710c",
   519 => x"81d7c008",
   520 => x"56548c15",
   521 => x"5381d7b4",
   522 => x"08528a51",
   523 => x"8fe73f73",
   524 => x"800c863d",
   525 => x"0d04fb3d",
   526 => x"0d777008",
   527 => x"5656b053",
   528 => x"81d7c008",
   529 => x"52745180",
   530 => x"cdff3f85",
   531 => x"0b8c170c",
   532 => x"850b8c16",
   533 => x"0c750875",
   534 => x"0c81d7c0",
   535 => x"08547380",
   536 => x"2e8a3873",
   537 => x"08750c81",
   538 => x"d7c00854",
   539 => x"8c145381",
   540 => x"d7b40852",
   541 => x"8a518f9d",
   542 => x"3f841508",
   543 => x"ad38860b",
   544 => x"8c160c88",
   545 => x"15528816",
   546 => x"08518ea9",
   547 => x"3f81d7c0",
   548 => x"08700876",
   549 => x"0c548c15",
   550 => x"7054548a",
   551 => x"52730851",
   552 => x"8ef33f73",
   553 => x"800c873d",
   554 => x"0d047508",
   555 => x"54b05373",
   556 => x"52755180",
   557 => x"cd933f73",
   558 => x"800c873d",
   559 => x"0d04d93d",
   560 => x"0d80f980",
   561 => x"0b8188e8",
   562 => x"0cb05180",
   563 => x"c0e43f80",
   564 => x"0881d7b0",
   565 => x"0cb05180",
   566 => x"c0d83f80",
   567 => x"0881d7c0",
   568 => x"0c81d7b0",
   569 => x"0880080c",
   570 => x"800b8008",
   571 => x"84050c82",
   572 => x"0b800888",
   573 => x"050ca80b",
   574 => x"80088c05",
   575 => x"0c9f5380",
   576 => x"ead85280",
   577 => x"08900551",
   578 => x"80ccbe3f",
   579 => x"a13d5e9f",
   580 => x"5380eaf8",
   581 => x"527d5180",
   582 => x"ccaf3f8a",
   583 => x"0b8195f4",
   584 => x"0c80f59c",
   585 => x"51f9ae3f",
   586 => x"80eb9851",
   587 => x"f9a73f80",
   588 => x"f59c51f9",
   589 => x"a03f80f8",
   590 => x"fc08802e",
   591 => x"89d73880",
   592 => x"ebc851f9",
   593 => x"903f80f5",
   594 => x"9c51f989",
   595 => x"3f80f8f8",
   596 => x"085280eb",
   597 => x"f451f8fd",
   598 => x"3f818990",
   599 => x"5180d5da",
   600 => x"3f810b9a",
   601 => x"3d5e5b80",
   602 => x"0b80f8f8",
   603 => x"082582d6",
   604 => x"38903d5f",
   605 => x"80c10b81",
   606 => x"d7b83481",
   607 => x"0b81d994",
   608 => x"0c80c20b",
   609 => x"81d7bc34",
   610 => x"8240835a",
   611 => x"9f5380ec",
   612 => x"a4527c51",
   613 => x"80cbb23f",
   614 => x"8141807d",
   615 => x"537e5256",
   616 => x"8e973f80",
   617 => x"08762e09",
   618 => x"81068338",
   619 => x"81567581",
   620 => x"d9940c7f",
   621 => x"70585675",
   622 => x"8325a238",
   623 => x"75101016",
   624 => x"fd0542a9",
   625 => x"3dffa405",
   626 => x"53835276",
   627 => x"518cc63f",
   628 => x"7f810570",
   629 => x"41705856",
   630 => x"837624e0",
   631 => x"38615475",
   632 => x"53818998",
   633 => x"5281d7cc",
   634 => x"518cba3f",
   635 => x"81d7c008",
   636 => x"70085858",
   637 => x"b0537752",
   638 => x"765180ca",
   639 => x"cc3f850b",
   640 => x"8c190c85",
   641 => x"0b8c180c",
   642 => x"7708770c",
   643 => x"81d7c008",
   644 => x"5675802e",
   645 => x"8a387508",
   646 => x"770c81d7",
   647 => x"c008568c",
   648 => x"165381d7",
   649 => x"b408528a",
   650 => x"518bea3f",
   651 => x"84170887",
   652 => x"eb38860b",
   653 => x"8c180c88",
   654 => x"17528818",
   655 => x"08518af5",
   656 => x"3f81d7c0",
   657 => x"08700878",
   658 => x"0c568c17",
   659 => x"7054598a",
   660 => x"52780851",
   661 => x"8bbf3f80",
   662 => x"c10b81d7",
   663 => x"bc335757",
   664 => x"767626a2",
   665 => x"3880c352",
   666 => x"76518ca3",
   667 => x"3f800861",
   668 => x"2e89e638",
   669 => x"81177081",
   670 => x"ff0681d7",
   671 => x"bc335858",
   672 => x"58757727",
   673 => x"e0387960",
   674 => x"29627054",
   675 => x"71535b59",
   676 => x"b9a43f80",
   677 => x"0840787a",
   678 => x"31708729",
   679 => x"80083180",
   680 => x"088a0581",
   681 => x"d7b83381",
   682 => x"d7b4085e",
   683 => x"5b525a56",
   684 => x"7780c12e",
   685 => x"89d0387b",
   686 => x"f738811b",
   687 => x"5b80f8f8",
   688 => x"087b25fd",
   689 => x"af3881d7",
   690 => x"a85180d2",
   691 => x"ed3f80ec",
   692 => x"c451f681",
   693 => x"3f80f59c",
   694 => x"51f5fa3f",
   695 => x"80ecd451",
   696 => x"f5f33f80",
   697 => x"f59c51f5",
   698 => x"ec3f81d7",
   699 => x"b4085280",
   700 => x"ed8c51f5",
   701 => x"e03f8552",
   702 => x"80eda851",
   703 => x"f5d73f81",
   704 => x"d9940852",
   705 => x"80edc451",
   706 => x"f5cb3f81",
   707 => x"5280eda8",
   708 => x"51f5c23f",
   709 => x"81d7b833",
   710 => x"5280ede0",
   711 => x"51f5b63f",
   712 => x"80c15280",
   713 => x"edfc51f5",
   714 => x"ac3f81d7",
   715 => x"bc335280",
   716 => x"ee9851f5",
   717 => x"a03f80c2",
   718 => x"5280edfc",
   719 => x"51f5963f",
   720 => x"81d7ec08",
   721 => x"5280eeb4",
   722 => x"51f58a3f",
   723 => x"875280ed",
   724 => x"a851f581",
   725 => x"3f8195f4",
   726 => x"085280ee",
   727 => x"d051f4f5",
   728 => x"3f80eeec",
   729 => x"51f4ee3f",
   730 => x"80ef9851",
   731 => x"f4e73f81",
   732 => x"d7c00870",
   733 => x"08535a80",
   734 => x"efa451f4",
   735 => x"d83f80ef",
   736 => x"c051f4d1",
   737 => x"3f81d7c0",
   738 => x"08841108",
   739 => x"535680ef",
   740 => x"f451f4c1",
   741 => x"3f805280",
   742 => x"eda851f4",
   743 => x"b83f81d7",
   744 => x"c0088811",
   745 => x"08535880",
   746 => x"f09051f4",
   747 => x"a83f8252",
   748 => x"80eda851",
   749 => x"f49f3f81",
   750 => x"d7c0088c",
   751 => x"11085357",
   752 => x"80f0ac51",
   753 => x"f48f3f91",
   754 => x"5280eda8",
   755 => x"51f4863f",
   756 => x"81d7c008",
   757 => x"90055280",
   758 => x"f0c851f3",
   759 => x"f83f80f0",
   760 => x"e451f3f1",
   761 => x"3f80f19c",
   762 => x"51f3ea3f",
   763 => x"81d7b008",
   764 => x"7008535f",
   765 => x"80efa451",
   766 => x"f3db3f80",
   767 => x"f1b051f3",
   768 => x"d43f81d7",
   769 => x"b0088411",
   770 => x"08535b80",
   771 => x"eff451f3",
   772 => x"c43f8052",
   773 => x"80eda851",
   774 => x"f3bb3f81",
   775 => x"d7b00888",
   776 => x"1108535c",
   777 => x"80f09051",
   778 => x"f3ab3f81",
   779 => x"5280eda8",
   780 => x"51f3a23f",
   781 => x"81d7b008",
   782 => x"8c110853",
   783 => x"5a80f0ac",
   784 => x"51f3923f",
   785 => x"925280ed",
   786 => x"a851f389",
   787 => x"3f81d7b0",
   788 => x"08900552",
   789 => x"80f0c851",
   790 => x"f2fb3f80",
   791 => x"f0e451f2",
   792 => x"f43f7f52",
   793 => x"80f1f051",
   794 => x"f2eb3f85",
   795 => x"5280eda8",
   796 => x"51f2e23f",
   797 => x"785280f2",
   798 => x"8c51f2d9",
   799 => x"3f8d5280",
   800 => x"eda851f2",
   801 => x"d03f6152",
   802 => x"80f2a851",
   803 => x"f2c73f87",
   804 => x"5280eda8",
   805 => x"51f2be3f",
   806 => x"605280f2",
   807 => x"c451f2b5",
   808 => x"3f815280",
   809 => x"eda851f2",
   810 => x"ac3f7d52",
   811 => x"80f2e051",
   812 => x"f2a33f80",
   813 => x"f2fc51f2",
   814 => x"9c3f7c52",
   815 => x"80f3b451",
   816 => x"f2933f80",
   817 => x"f3d051f2",
   818 => x"8c3f80f5",
   819 => x"9c51f285",
   820 => x"3f81d7a8",
   821 => x"0881d7ac",
   822 => x"08818990",
   823 => x"08818994",
   824 => x"08727131",
   825 => x"70742675",
   826 => x"74317072",
   827 => x"31818988",
   828 => x"0c444481",
   829 => x"898c0c81",
   830 => x"898c0856",
   831 => x"80f48855",
   832 => x"5c595758",
   833 => x"f1cf3f81",
   834 => x"89880856",
   835 => x"80762582",
   836 => x"a43880f8",
   837 => x"f8087071",
   838 => x"9f2c9a3d",
   839 => x"53565681",
   840 => x"89880881",
   841 => x"898c0841",
   842 => x"537f5470",
   843 => x"525a8ef6",
   844 => x"3f66685f",
   845 => x"8188f80c",
   846 => x"7d8188fc",
   847 => x"0c80f8f8",
   848 => x"08709f2c",
   849 => x"58568058",
   850 => x"bd84c078",
   851 => x"55557652",
   852 => x"75537951",
   853 => x"87d23f95",
   854 => x"3d818988",
   855 => x"0881898c",
   856 => x"0841557f",
   857 => x"56676940",
   858 => x"537e5470",
   859 => x"525c8eb6",
   860 => x"3f64665e",
   861 => x"8189800c",
   862 => x"7c818984",
   863 => x"0c80f8f8",
   864 => x"08709f2c",
   865 => x"40588057",
   866 => x"83dceb94",
   867 => x"80775555",
   868 => x"7e527753",
   869 => x"7b518790",
   870 => x"3f64665d",
   871 => x"5b805e8d",
   872 => x"dd7e5555",
   873 => x"81898808",
   874 => x"81898c08",
   875 => x"59527753",
   876 => x"795186f4",
   877 => x"3f666840",
   878 => x"547e557a",
   879 => x"527b53a9",
   880 => x"3dffa805",
   881 => x"518ddf3f",
   882 => x"62645e81",
   883 => x"d7c40c7c",
   884 => x"81d7c80c",
   885 => x"80f49851",
   886 => x"effb3f81",
   887 => x"88fc0852",
   888 => x"80f4c851",
   889 => x"efef3f80",
   890 => x"f4d051ef",
   891 => x"e83f8189",
   892 => x"84085280",
   893 => x"f4c851ef",
   894 => x"dc3f81d7",
   895 => x"c8085280",
   896 => x"f58051ef",
   897 => x"d03f80f5",
   898 => x"9c51efc9",
   899 => x"3f800b80",
   900 => x"0ca93d0d",
   901 => x"0480f5a0",
   902 => x"51f6a839",
   903 => x"770857b0",
   904 => x"53765277",
   905 => x"5180c2a1",
   906 => x"3f80c10b",
   907 => x"81d7bc33",
   908 => x"5757f8ac",
   909 => x"39758a38",
   910 => x"81898c08",
   911 => x"8126fdd2",
   912 => x"3880f5d0",
   913 => x"51ef8e3f",
   914 => x"80f68851",
   915 => x"ef873f80",
   916 => x"f59c51ef",
   917 => x"803f80f8",
   918 => x"f8087071",
   919 => x"9f2c9a3d",
   920 => x"53565681",
   921 => x"89880881",
   922 => x"898c0841",
   923 => x"537f5470",
   924 => x"525a8cb2",
   925 => x"3f66685f",
   926 => x"8188f80c",
   927 => x"7d8188fc",
   928 => x"0c80f8f8",
   929 => x"08709f2c",
   930 => x"58568058",
   931 => x"bd84c078",
   932 => x"55557652",
   933 => x"75537951",
   934 => x"858e3f95",
   935 => x"3d818988",
   936 => x"0881898c",
   937 => x"0841557f",
   938 => x"56676940",
   939 => x"537e5470",
   940 => x"525c8bf2",
   941 => x"3f64665e",
   942 => x"8189800c",
   943 => x"7c818984",
   944 => x"0c80f8f8",
   945 => x"08709f2c",
   946 => x"40588057",
   947 => x"83dceb94",
   948 => x"80775555",
   949 => x"7e527753",
   950 => x"7b5184cc",
   951 => x"3f64665d",
   952 => x"5b805e8d",
   953 => x"dd7e5555",
   954 => x"81898808",
   955 => x"81898c08",
   956 => x"59527753",
   957 => x"795184b0",
   958 => x"3f666840",
   959 => x"547e557a",
   960 => x"527b53a9",
   961 => x"3dffa805",
   962 => x"518b9b3f",
   963 => x"62645e81",
   964 => x"d7c40c7c",
   965 => x"81d7c80c",
   966 => x"80f49851",
   967 => x"edb73f81",
   968 => x"88fc0852",
   969 => x"80f4c851",
   970 => x"edab3f80",
   971 => x"f4d051ed",
   972 => x"a43f8189",
   973 => x"84085280",
   974 => x"f4c851ed",
   975 => x"983f81d7",
   976 => x"c8085280",
   977 => x"f58051ed",
   978 => x"8c3f80f5",
   979 => x"9c51ed85",
   980 => x"3f800b80",
   981 => x"0ca93d0d",
   982 => x"04a93dff",
   983 => x"a0055280",
   984 => x"5180d23f",
   985 => x"9f5380f6",
   986 => x"a8527c51",
   987 => x"bfdb3f7a",
   988 => x"7b81d7b4",
   989 => x"0c811870",
   990 => x"81ff0681",
   991 => x"d7bc3359",
   992 => x"59595af5",
   993 => x"fc39ff16",
   994 => x"707b3160",
   995 => x"0c5c800b",
   996 => x"811c5c5c",
   997 => x"80f8f808",
   998 => x"7b25f3d8",
   999 => x"38f6a739",
  1000 => x"ff3d0d73",
  1001 => x"82327030",
  1002 => x"70720780",
  1003 => x"25800c52",
  1004 => x"52833d0d",
  1005 => x"04fe3d0d",
  1006 => x"74767153",
  1007 => x"54527182",
  1008 => x"2e833883",
  1009 => x"5171812e",
  1010 => x"9a388172",
  1011 => x"269f3871",
  1012 => x"822eb838",
  1013 => x"71842ea9",
  1014 => x"3870730c",
  1015 => x"70800c84",
  1016 => x"3d0d0480",
  1017 => x"e40b81d7",
  1018 => x"b408258b",
  1019 => x"3880730c",
  1020 => x"70800c84",
  1021 => x"3d0d0483",
  1022 => x"730c7080",
  1023 => x"0c843d0d",
  1024 => x"0482730c",
  1025 => x"70800c84",
  1026 => x"3d0d0481",
  1027 => x"730c7080",
  1028 => x"0c843d0d",
  1029 => x"04803d0d",
  1030 => x"74741482",
  1031 => x"05710c80",
  1032 => x"0c823d0d",
  1033 => x"04f73d0d",
  1034 => x"7b7d7f61",
  1035 => x"85127082",
  1036 => x"2b751170",
  1037 => x"74717084",
  1038 => x"05530c5a",
  1039 => x"5a5d5b76",
  1040 => x"0c7980f8",
  1041 => x"180c7986",
  1042 => x"12525758",
  1043 => x"5a5a7676",
  1044 => x"24993876",
  1045 => x"b329822b",
  1046 => x"79115153",
  1047 => x"76737084",
  1048 => x"05550c81",
  1049 => x"14547574",
  1050 => x"25f23876",
  1051 => x"81cc2919",
  1052 => x"fc110881",
  1053 => x"05fc120c",
  1054 => x"7a197008",
  1055 => x"9fa0130c",
  1056 => x"5856850b",
  1057 => x"81d7b40c",
  1058 => x"75800c8b",
  1059 => x"3d0d04fe",
  1060 => x"3d0d0293",
  1061 => x"05335180",
  1062 => x"02840597",
  1063 => x"05335452",
  1064 => x"70732e88",
  1065 => x"3871800c",
  1066 => x"843d0d04",
  1067 => x"7081d7b8",
  1068 => x"34810b80",
  1069 => x"0c843d0d",
  1070 => x"04f83d0d",
  1071 => x"7a7c5956",
  1072 => x"820b8319",
  1073 => x"55557416",
  1074 => x"70337533",
  1075 => x"5b515372",
  1076 => x"792e80c6",
  1077 => x"3880c10b",
  1078 => x"81168116",
  1079 => x"56565782",
  1080 => x"7525e338",
  1081 => x"ffa91770",
  1082 => x"81ff0655",
  1083 => x"59738226",
  1084 => x"83388755",
  1085 => x"81537680",
  1086 => x"d22e9838",
  1087 => x"77527551",
  1088 => x"be963f80",
  1089 => x"53728008",
  1090 => x"25893887",
  1091 => x"1581d7b4",
  1092 => x"0c815372",
  1093 => x"800c8a3d",
  1094 => x"0d047281",
  1095 => x"d7b83482",
  1096 => x"7525ffa2",
  1097 => x"38ffbd39",
  1098 => x"8c08028c",
  1099 => x"0ceb3d0d",
  1100 => x"800b8c08",
  1101 => x"f0050c80",
  1102 => x"0b8c08f4",
  1103 => x"050c8c08",
  1104 => x"8c05088c",
  1105 => x"08900508",
  1106 => x"5654738c",
  1107 => x"08f0050c",
  1108 => x"748c08f4",
  1109 => x"050c8c08",
  1110 => x"f8058c08",
  1111 => x"f0055656",
  1112 => x"88705475",
  1113 => x"53765254",
  1114 => x"bbdf3f80",
  1115 => x"0b8c08e8",
  1116 => x"050c800b",
  1117 => x"8c08ec05",
  1118 => x"0c8c0894",
  1119 => x"05088c08",
  1120 => x"98050856",
  1121 => x"54738c08",
  1122 => x"e8050c74",
  1123 => x"8c08ec05",
  1124 => x"0c8c08f0",
  1125 => x"058c08e8",
  1126 => x"05565688",
  1127 => x"70547553",
  1128 => x"765254bb",
  1129 => x"a43f800b",
  1130 => x"8c08e805",
  1131 => x"0c800b8c",
  1132 => x"08ec050c",
  1133 => x"8c08fc05",
  1134 => x"0883ffff",
  1135 => x"068c08cc",
  1136 => x"050c8c08",
  1137 => x"fc050890",
  1138 => x"2a8c08c4",
  1139 => x"050c8c08",
  1140 => x"f4050883",
  1141 => x"ffff068c",
  1142 => x"08c8050c",
  1143 => x"8c08f405",
  1144 => x"08902a8c",
  1145 => x"08c0050c",
  1146 => x"8c08cc05",
  1147 => x"088c08c8",
  1148 => x"05082970",
  1149 => x"8c08dc05",
  1150 => x"0c8c08cc",
  1151 => x"05088c08",
  1152 => x"c0050829",
  1153 => x"708c08d8",
  1154 => x"050c8c08",
  1155 => x"c405088c",
  1156 => x"08c80508",
  1157 => x"29708c08",
  1158 => x"d4050c8c",
  1159 => x"08c40508",
  1160 => x"8c08c005",
  1161 => x"0829708c",
  1162 => x"08d0050c",
  1163 => x"8c08dc05",
  1164 => x"08902a8c",
  1165 => x"08d80508",
  1166 => x"118c08d8",
  1167 => x"050c8c08",
  1168 => x"d805088c",
  1169 => x"08d40508",
  1170 => x"058c08d8",
  1171 => x"050c5151",
  1172 => x"5151548c",
  1173 => x"08d80508",
  1174 => x"8c08d405",
  1175 => x"08278f38",
  1176 => x"8c08d005",
  1177 => x"08848080",
  1178 => x"058c08d0",
  1179 => x"050c8c08",
  1180 => x"d8050890",
  1181 => x"2a8c08d0",
  1182 => x"0508118c",
  1183 => x"08e0050c",
  1184 => x"8c08d805",
  1185 => x"0883ffff",
  1186 => x"0670902b",
  1187 => x"8c08dc05",
  1188 => x"0883ffff",
  1189 => x"0670128c",
  1190 => x"08e4050c",
  1191 => x"52575154",
  1192 => x"8c08e005",
  1193 => x"088c08e4",
  1194 => x"05085654",
  1195 => x"738c08e8",
  1196 => x"050c748c",
  1197 => x"08ec050c",
  1198 => x"8c08fc05",
  1199 => x"088c08f0",
  1200 => x"0508298c",
  1201 => x"08f80508",
  1202 => x"8c08f405",
  1203 => x"08297012",
  1204 => x"8c08e805",
  1205 => x"08118c08",
  1206 => x"e8050c51",
  1207 => x"55558c08",
  1208 => x"e805088c",
  1209 => x"08ec0508",
  1210 => x"8c088805",
  1211 => x"08585654",
  1212 => x"73760c74",
  1213 => x"84170c8c",
  1214 => x"08880508",
  1215 => x"800c973d",
  1216 => x"0d8c0c04",
  1217 => x"8c08028c",
  1218 => x"0cf63d0d",
  1219 => x"800b8c08",
  1220 => x"f0050c80",
  1221 => x"0b8c08f4",
  1222 => x"050c8c08",
  1223 => x"8c05088c",
  1224 => x"08900508",
  1225 => x"5654738c",
  1226 => x"08f0050c",
  1227 => x"748c08f4",
  1228 => x"050c8c08",
  1229 => x"f8058c08",
  1230 => x"f0055656",
  1231 => x"88705475",
  1232 => x"53765254",
  1233 => x"b8833f80",
  1234 => x"0b8c08f0",
  1235 => x"050c800b",
  1236 => x"8c08f405",
  1237 => x"0c8c08f8",
  1238 => x"0508308c",
  1239 => x"08ec050c",
  1240 => x"8c08fc05",
  1241 => x"08802e8d",
  1242 => x"388c08ec",
  1243 => x"0508ff05",
  1244 => x"8c08ec05",
  1245 => x"0c8c08ec",
  1246 => x"05088c08",
  1247 => x"f0050c8c",
  1248 => x"08fc0508",
  1249 => x"308c08f4",
  1250 => x"050c8c08",
  1251 => x"f005088c",
  1252 => x"08f40508",
  1253 => x"8c088805",
  1254 => x"08585654",
  1255 => x"73760c74",
  1256 => x"84170c8c",
  1257 => x"08880508",
  1258 => x"800c8c3d",
  1259 => x"0d8c0c04",
  1260 => x"8c08028c",
  1261 => x"0cf53d0d",
  1262 => x"8c089405",
  1263 => x"089d388c",
  1264 => x"088c0508",
  1265 => x"8c089005",
  1266 => x"088c0888",
  1267 => x"05085856",
  1268 => x"5473760c",
  1269 => x"7484170c",
  1270 => x"81bf3980",
  1271 => x"0b8c08f0",
  1272 => x"050c800b",
  1273 => x"8c08f405",
  1274 => x"0c8c088c",
  1275 => x"05088c08",
  1276 => x"90050856",
  1277 => x"54738c08",
  1278 => x"f0050c74",
  1279 => x"8c08f405",
  1280 => x"0c8c08f8",
  1281 => x"058c08f0",
  1282 => x"05565688",
  1283 => x"70547553",
  1284 => x"765254b6",
  1285 => x"b43fa00b",
  1286 => x"8c089405",
  1287 => x"08318c08",
  1288 => x"ec050c8c",
  1289 => x"08ec0508",
  1290 => x"80249d38",
  1291 => x"800b8c08",
  1292 => x"f4050c8c",
  1293 => x"08ec0508",
  1294 => x"308c08fc",
  1295 => x"0508712b",
  1296 => x"8c08f005",
  1297 => x"0c54b939",
  1298 => x"8c08fc05",
  1299 => x"088c08ec",
  1300 => x"05082a8c",
  1301 => x"08e8050c",
  1302 => x"8c08fc05",
  1303 => x"088c0894",
  1304 => x"05082b8c",
  1305 => x"08f4050c",
  1306 => x"8c08f805",
  1307 => x"088c0894",
  1308 => x"05082b70",
  1309 => x"8c08e805",
  1310 => x"08078c08",
  1311 => x"f0050c54",
  1312 => x"8c08f005",
  1313 => x"088c08f4",
  1314 => x"05088c08",
  1315 => x"88050858",
  1316 => x"56547376",
  1317 => x"0c748417",
  1318 => x"0c8c0888",
  1319 => x"0508800c",
  1320 => x"8d3d0d8c",
  1321 => x"0c048c08",
  1322 => x"028c0ccc",
  1323 => x"3d0d800b",
  1324 => x"8c08fc05",
  1325 => x"0c800b8c",
  1326 => x"08ec050c",
  1327 => x"800b8c08",
  1328 => x"f0050c8c",
  1329 => x"088c0508",
  1330 => x"8c089005",
  1331 => x"08565473",
  1332 => x"8c08ec05",
  1333 => x"0c748c08",
  1334 => x"f0050c8c",
  1335 => x"08f4058c",
  1336 => x"08ec0556",
  1337 => x"56887054",
  1338 => x"75537652",
  1339 => x"54b4da3f",
  1340 => x"800b8c08",
  1341 => x"e4050c80",
  1342 => x"0b8c08e8",
  1343 => x"050c8c08",
  1344 => x"9405088c",
  1345 => x"08980508",
  1346 => x"5654738c",
  1347 => x"08e4050c",
  1348 => x"748c08e8",
  1349 => x"050c8c08",
  1350 => x"ec058c08",
  1351 => x"e4055656",
  1352 => x"88705475",
  1353 => x"53765254",
  1354 => x"b49f3f8c",
  1355 => x"08f40508",
  1356 => x"8025be38",
  1357 => x"8c08fc05",
  1358 => x"08098c08",
  1359 => x"fc050c8c",
  1360 => x"08d40554",
  1361 => x"8c08f405",
  1362 => x"088c08f8",
  1363 => x"05085755",
  1364 => x"74527553",
  1365 => x"7351fbac",
  1366 => x"3f8c08d4",
  1367 => x"05088c08",
  1368 => x"d8050856",
  1369 => x"54738c08",
  1370 => x"f4050c74",
  1371 => x"8c08f805",
  1372 => x"0c8c08ec",
  1373 => x"05088025",
  1374 => x"be388c08",
  1375 => x"fc050809",
  1376 => x"8c08fc05",
  1377 => x"0c8c08d4",
  1378 => x"05548c08",
  1379 => x"ec05088c",
  1380 => x"08f00508",
  1381 => x"57557452",
  1382 => x"75537351",
  1383 => x"fae63f8c",
  1384 => x"08d40508",
  1385 => x"8c08d805",
  1386 => x"08565473",
  1387 => x"8c08ec05",
  1388 => x"0c748c08",
  1389 => x"f0050c8c",
  1390 => x"08f40508",
  1391 => x"8c08f805",
  1392 => x"08565473",
  1393 => x"8c08d405",
  1394 => x"0c748c08",
  1395 => x"d8050c8c",
  1396 => x"08ec0508",
  1397 => x"8c08f005",
  1398 => x"08565473",
  1399 => x"8c08cc05",
  1400 => x"0c748c08",
  1401 => x"d0050c80",
  1402 => x"0b8c08c8",
  1403 => x"050c800b",
  1404 => x"8c08e405",
  1405 => x"0c800b8c",
  1406 => x"08e8050c",
  1407 => x"8c08d405",
  1408 => x"088c08d8",
  1409 => x"05085654",
  1410 => x"738c08e4",
  1411 => x"050c748c",
  1412 => x"08e8050c",
  1413 => x"800b8c08",
  1414 => x"ffb8050c",
  1415 => x"800b8c08",
  1416 => x"ffbc050c",
  1417 => x"8c08cc05",
  1418 => x"088c08d0",
  1419 => x"05085654",
  1420 => x"738c08ff",
  1421 => x"b8050c74",
  1422 => x"8c08ffbc",
  1423 => x"050c8c08",
  1424 => x"ffbc0508",
  1425 => x"8c08ffac",
  1426 => x"050c8c08",
  1427 => x"ffb80508",
  1428 => x"8c08ffa8",
  1429 => x"050c8c08",
  1430 => x"e805088c",
  1431 => x"08ffa405",
  1432 => x"0c8c08e4",
  1433 => x"05088c08",
  1434 => x"ffa0050c",
  1435 => x"8c08ffa8",
  1436 => x"050891d4",
  1437 => x"388c08ff",
  1438 => x"a005088c",
  1439 => x"08ffac05",
  1440 => x"0827868c",
  1441 => x"388c08ff",
  1442 => x"ac05088c",
  1443 => x"08ff8805",
  1444 => x"0c8c08ff",
  1445 => x"88050883",
  1446 => x"ffff26a0",
  1447 => x"388c08ff",
  1448 => x"88050881",
  1449 => x"ff268b38",
  1450 => x"800b8c08",
  1451 => x"fed8050c",
  1452 => x"a939880b",
  1453 => x"8c08fed8",
  1454 => x"050c9f39",
  1455 => x"8c08ff88",
  1456 => x"0508fe80",
  1457 => x"0a268b38",
  1458 => x"900b8c08",
  1459 => x"fed8050c",
  1460 => x"8939980b",
  1461 => x"8c08fed8",
  1462 => x"050c8c08",
  1463 => x"fed80508",
  1464 => x"8c08ff84",
  1465 => x"050c8c08",
  1466 => x"ff880508",
  1467 => x"8c08ff84",
  1468 => x"05082a80",
  1469 => x"f6c81133",
  1470 => x"8c08ff84",
  1471 => x"050811a0",
  1472 => x"71318c08",
  1473 => x"ff8c050c",
  1474 => x"5151548c",
  1475 => x"08ff8c05",
  1476 => x"08802e80",
  1477 => x"d1388c08",
  1478 => x"ffac0508",
  1479 => x"8c08ff8c",
  1480 => x"05082b8c",
  1481 => x"08ffac05",
  1482 => x"0c8c08ff",
  1483 => x"a005088c",
  1484 => x"08ff8c05",
  1485 => x"082ba00b",
  1486 => x"8c08ff8c",
  1487 => x"0508318c",
  1488 => x"08ffa405",
  1489 => x"08712a70",
  1490 => x"73078c08",
  1491 => x"ffa0050c",
  1492 => x"8c08ffa4",
  1493 => x"05088c08",
  1494 => x"ff8c0508",
  1495 => x"2b8c08ff",
  1496 => x"a4050c51",
  1497 => x"56548c08",
  1498 => x"ffac0508",
  1499 => x"902a8c08",
  1500 => x"ff84050c",
  1501 => x"8c08ffac",
  1502 => x"050883ff",
  1503 => x"ff068c08",
  1504 => x"ff88050c",
  1505 => x"8c08ffa0",
  1506 => x"05088c08",
  1507 => x"ff840508",
  1508 => x"53705254",
  1509 => x"9efb3f80",
  1510 => x"08708c08",
  1511 => x"fef8050c",
  1512 => x"8c08ff84",
  1513 => x"0508538c",
  1514 => x"08ffa005",
  1515 => x"0852549e",
  1516 => x"bb3f8008",
  1517 => x"708c08ff",
  1518 => x"80050c8c",
  1519 => x"08ff8005",
  1520 => x"088c08ff",
  1521 => x"88050829",
  1522 => x"708c08fe",
  1523 => x"f0050c8c",
  1524 => x"08fef805",
  1525 => x"0870902b",
  1526 => x"8c08ffa4",
  1527 => x"0508902a",
  1528 => x"7072078c",
  1529 => x"08fef805",
  1530 => x"0c525851",
  1531 => x"51548c08",
  1532 => x"fef80508",
  1533 => x"8c08fef0",
  1534 => x"05082780",
  1535 => x"e1388c08",
  1536 => x"ff800508",
  1537 => x"ff058c08",
  1538 => x"ff80050c",
  1539 => x"8c08fef8",
  1540 => x"05088c08",
  1541 => x"ffac0508",
  1542 => x"058c08fe",
  1543 => x"f8050c8c",
  1544 => x"08ffac05",
  1545 => x"088c08fe",
  1546 => x"f8050826",
  1547 => x"b1388c08",
  1548 => x"fef80508",
  1549 => x"8c08fef0",
  1550 => x"050827a2",
  1551 => x"388c08ff",
  1552 => x"800508ff",
  1553 => x"058c08ff",
  1554 => x"80050c8c",
  1555 => x"08fef805",
  1556 => x"088c08ff",
  1557 => x"ac050805",
  1558 => x"8c08fef8",
  1559 => x"050c8c08",
  1560 => x"fef80508",
  1561 => x"8c08fef0",
  1562 => x"0508318c",
  1563 => x"08fef805",
  1564 => x"0c8c08fe",
  1565 => x"f805088c",
  1566 => x"08ff8405",
  1567 => x"08537052",
  1568 => x"549d8e3f",
  1569 => x"8008708c",
  1570 => x"08fef405",
  1571 => x"0c8c08ff",
  1572 => x"84050853",
  1573 => x"8c08fef8",
  1574 => x"05085254",
  1575 => x"9cce3f80",
  1576 => x"08708c08",
  1577 => x"fefc050c",
  1578 => x"8c08fefc",
  1579 => x"05088c08",
  1580 => x"ff880508",
  1581 => x"29708c08",
  1582 => x"fef0050c",
  1583 => x"8c08fef4",
  1584 => x"05087090",
  1585 => x"2b8c08ff",
  1586 => x"a4050883",
  1587 => x"ffff0670",
  1588 => x"72078c08",
  1589 => x"fef4050c",
  1590 => x"52585151",
  1591 => x"548c08fe",
  1592 => x"f405088c",
  1593 => x"08fef005",
  1594 => x"082780e1",
  1595 => x"388c08fe",
  1596 => x"fc0508ff",
  1597 => x"058c08fe",
  1598 => x"fc050c8c",
  1599 => x"08fef405",
  1600 => x"088c08ff",
  1601 => x"ac050805",
  1602 => x"8c08fef4",
  1603 => x"050c8c08",
  1604 => x"ffac0508",
  1605 => x"8c08fef4",
  1606 => x"050826b1",
  1607 => x"388c08fe",
  1608 => x"f405088c",
  1609 => x"08fef005",
  1610 => x"0827a238",
  1611 => x"8c08fefc",
  1612 => x"0508ff05",
  1613 => x"8c08fefc",
  1614 => x"050c8c08",
  1615 => x"fef40508",
  1616 => x"8c08ffac",
  1617 => x"0508058c",
  1618 => x"08fef405",
  1619 => x"0c8c08fe",
  1620 => x"f405088c",
  1621 => x"08fef005",
  1622 => x"08318c08",
  1623 => x"fef4050c",
  1624 => x"8c08ff80",
  1625 => x"05087090",
  1626 => x"2b708c08",
  1627 => x"fefc0508",
  1628 => x"078c08ff",
  1629 => x"98050c8c",
  1630 => x"08fef405",
  1631 => x"088c08ff",
  1632 => x"a4050c51",
  1633 => x"54800b8c",
  1634 => x"08ff9405",
  1635 => x"0c8af639",
  1636 => x"8c08ffac",
  1637 => x"05089738",
  1638 => x"8c08ffac",
  1639 => x"05085281",
  1640 => x"519ac93f",
  1641 => x"8008708c",
  1642 => x"08ffac05",
  1643 => x"0c548c08",
  1644 => x"ffac0508",
  1645 => x"8c08fef0",
  1646 => x"050c8c08",
  1647 => x"fef00508",
  1648 => x"83ffff26",
  1649 => x"a0388c08",
  1650 => x"fef00508",
  1651 => x"81ff268b",
  1652 => x"38800b8c",
  1653 => x"08fed405",
  1654 => x"0ca93988",
  1655 => x"0b8c08fe",
  1656 => x"d4050c9f",
  1657 => x"398c08fe",
  1658 => x"f00508fe",
  1659 => x"800a268b",
  1660 => x"38900b8c",
  1661 => x"08fed405",
  1662 => x"0c893998",
  1663 => x"0b8c08fe",
  1664 => x"d4050c8c",
  1665 => x"08fed405",
  1666 => x"088c08fe",
  1667 => x"f4050c8c",
  1668 => x"08fef005",
  1669 => x"088c08fe",
  1670 => x"f405082a",
  1671 => x"80f6c811",
  1672 => x"338c08fe",
  1673 => x"f4050811",
  1674 => x"a071318c",
  1675 => x"08ff8c05",
  1676 => x"0c515154",
  1677 => x"8c08ff8c",
  1678 => x"05089f38",
  1679 => x"8c08ffa0",
  1680 => x"05088c08",
  1681 => x"ffac0508",
  1682 => x"318c08ff",
  1683 => x"a0050c81",
  1684 => x"0b8c08ff",
  1685 => x"94050c85",
  1686 => x"8d39a00b",
  1687 => x"8c08ff8c",
  1688 => x"0508318c",
  1689 => x"08ff9005",
  1690 => x"0c8c08ff",
  1691 => x"ac05088c",
  1692 => x"08ff8c05",
  1693 => x"082b8c08",
  1694 => x"ffac050c",
  1695 => x"8c08ffa0",
  1696 => x"05088c08",
  1697 => x"ff900508",
  1698 => x"2a8c08ff",
  1699 => x"9c050c8c",
  1700 => x"08ffa005",
  1701 => x"088c08ff",
  1702 => x"8c05082b",
  1703 => x"8c08ffa4",
  1704 => x"05088c08",
  1705 => x"ff900508",
  1706 => x"2a707207",
  1707 => x"8c08ffa0",
  1708 => x"050c8c08",
  1709 => x"ffa40508",
  1710 => x"8c08ff8c",
  1711 => x"05082b8c",
  1712 => x"08ffa405",
  1713 => x"0c8c08ff",
  1714 => x"ac050890",
  1715 => x"2a8c08fe",
  1716 => x"f0050c8c",
  1717 => x"08ffac05",
  1718 => x"0883ffff",
  1719 => x"068c08fe",
  1720 => x"f4050c8c",
  1721 => x"08ff9c05",
  1722 => x"088c08fe",
  1723 => x"f0050855",
  1724 => x"70545155",
  1725 => x"55989a3f",
  1726 => x"8008708c",
  1727 => x"08ff8005",
  1728 => x"0c8c08fe",
  1729 => x"f0050853",
  1730 => x"8c08ff9c",
  1731 => x"05085254",
  1732 => x"97da3f80",
  1733 => x"08708c08",
  1734 => x"fef8050c",
  1735 => x"8c08fef8",
  1736 => x"05088c08",
  1737 => x"fef40508",
  1738 => x"29708c08",
  1739 => x"ff88050c",
  1740 => x"8c08ff80",
  1741 => x"05087090",
  1742 => x"2b8c08ff",
  1743 => x"a0050890",
  1744 => x"2a707207",
  1745 => x"8c08ff80",
  1746 => x"050c5258",
  1747 => x"5151548c",
  1748 => x"08ff8005",
  1749 => x"088c08ff",
  1750 => x"88050827",
  1751 => x"80e1388c",
  1752 => x"08fef805",
  1753 => x"08ff058c",
  1754 => x"08fef805",
  1755 => x"0c8c08ff",
  1756 => x"8005088c",
  1757 => x"08ffac05",
  1758 => x"08058c08",
  1759 => x"ff80050c",
  1760 => x"8c08ffac",
  1761 => x"05088c08",
  1762 => x"ff800508",
  1763 => x"26b1388c",
  1764 => x"08ff8005",
  1765 => x"088c08ff",
  1766 => x"88050827",
  1767 => x"a2388c08",
  1768 => x"fef80508",
  1769 => x"ff058c08",
  1770 => x"fef8050c",
  1771 => x"8c08ff80",
  1772 => x"05088c08",
  1773 => x"ffac0508",
  1774 => x"058c08ff",
  1775 => x"80050c8c",
  1776 => x"08ff8005",
  1777 => x"088c08ff",
  1778 => x"88050831",
  1779 => x"8c08ff80",
  1780 => x"050c8c08",
  1781 => x"ff800508",
  1782 => x"8c08fef0",
  1783 => x"05085370",
  1784 => x"525496ad",
  1785 => x"3f800870",
  1786 => x"8c08ff84",
  1787 => x"050c8c08",
  1788 => x"fef00508",
  1789 => x"538c08ff",
  1790 => x"80050852",
  1791 => x"5495ed3f",
  1792 => x"8008708c",
  1793 => x"08fefc05",
  1794 => x"0c8c08fe",
  1795 => x"fc05088c",
  1796 => x"08fef405",
  1797 => x"0829708c",
  1798 => x"08ff8805",
  1799 => x"0c8c08ff",
  1800 => x"84050870",
  1801 => x"902b8c08",
  1802 => x"ffa00508",
  1803 => x"83ffff06",
  1804 => x"7072078c",
  1805 => x"08ff8405",
  1806 => x"0c525851",
  1807 => x"51548c08",
  1808 => x"ff840508",
  1809 => x"8c08ff88",
  1810 => x"05082780",
  1811 => x"e1388c08",
  1812 => x"fefc0508",
  1813 => x"ff058c08",
  1814 => x"fefc050c",
  1815 => x"8c08ff84",
  1816 => x"05088c08",
  1817 => x"ffac0508",
  1818 => x"058c08ff",
  1819 => x"84050c8c",
  1820 => x"08ffac05",
  1821 => x"088c08ff",
  1822 => x"84050826",
  1823 => x"b1388c08",
  1824 => x"ff840508",
  1825 => x"8c08ff88",
  1826 => x"050827a2",
  1827 => x"388c08fe",
  1828 => x"fc0508ff",
  1829 => x"058c08fe",
  1830 => x"fc050c8c",
  1831 => x"08ff8405",
  1832 => x"088c08ff",
  1833 => x"ac050805",
  1834 => x"8c08ff84",
  1835 => x"050c8c08",
  1836 => x"ff840508",
  1837 => x"8c08ff88",
  1838 => x"0508318c",
  1839 => x"08ff8405",
  1840 => x"0c8c08fe",
  1841 => x"f8050870",
  1842 => x"902b708c",
  1843 => x"08fefc05",
  1844 => x"08078c08",
  1845 => x"ff94050c",
  1846 => x"8c08ff84",
  1847 => x"05088c08",
  1848 => x"ffa0050c",
  1849 => x"51548c08",
  1850 => x"ffac0508",
  1851 => x"902a8c08",
  1852 => x"fef0050c",
  1853 => x"8c08ffac",
  1854 => x"050883ff",
  1855 => x"ff068c08",
  1856 => x"fef4050c",
  1857 => x"8c08ffa0",
  1858 => x"05088c08",
  1859 => x"fef00508",
  1860 => x"53705254",
  1861 => x"93fb3f80",
  1862 => x"08708c08",
  1863 => x"ff80050c",
  1864 => x"8c08fef0",
  1865 => x"0508538c",
  1866 => x"08ffa005",
  1867 => x"08525493",
  1868 => x"bb3f8008",
  1869 => x"708c08fe",
  1870 => x"f8050c8c",
  1871 => x"08fef805",
  1872 => x"088c08fe",
  1873 => x"f4050829",
  1874 => x"708c08ff",
  1875 => x"88050c8c",
  1876 => x"08ff8005",
  1877 => x"0870902b",
  1878 => x"8c08ffa4",
  1879 => x"0508902a",
  1880 => x"7072078c",
  1881 => x"08ff8005",
  1882 => x"0c525851",
  1883 => x"51548c08",
  1884 => x"ff800508",
  1885 => x"8c08ff88",
  1886 => x"05082780",
  1887 => x"e1388c08",
  1888 => x"fef80508",
  1889 => x"ff058c08",
  1890 => x"fef8050c",
  1891 => x"8c08ff80",
  1892 => x"05088c08",
  1893 => x"ffac0508",
  1894 => x"058c08ff",
  1895 => x"80050c8c",
  1896 => x"08ffac05",
  1897 => x"088c08ff",
  1898 => x"80050826",
  1899 => x"b1388c08",
  1900 => x"ff800508",
  1901 => x"8c08ff88",
  1902 => x"050827a2",
  1903 => x"388c08fe",
  1904 => x"f80508ff",
  1905 => x"058c08fe",
  1906 => x"f8050c8c",
  1907 => x"08ff8005",
  1908 => x"088c08ff",
  1909 => x"ac050805",
  1910 => x"8c08ff80",
  1911 => x"050c8c08",
  1912 => x"ff800508",
  1913 => x"8c08ff88",
  1914 => x"0508318c",
  1915 => x"08ff8005",
  1916 => x"0c8c08ff",
  1917 => x"8005088c",
  1918 => x"08fef005",
  1919 => x"08537052",
  1920 => x"54928e3f",
  1921 => x"8008708c",
  1922 => x"08ff8405",
  1923 => x"0c8c08fe",
  1924 => x"f0050853",
  1925 => x"8c08ff80",
  1926 => x"05085254",
  1927 => x"91ce3f80",
  1928 => x"08708c08",
  1929 => x"fefc050c",
  1930 => x"8c08fefc",
  1931 => x"05088c08",
  1932 => x"fef40508",
  1933 => x"29708c08",
  1934 => x"ff88050c",
  1935 => x"8c08ff84",
  1936 => x"05087090",
  1937 => x"2b8c08ff",
  1938 => x"a4050883",
  1939 => x"ffff0670",
  1940 => x"72078c08",
  1941 => x"ff84050c",
  1942 => x"52585151",
  1943 => x"548c08ff",
  1944 => x"8405088c",
  1945 => x"08ff8805",
  1946 => x"082780e1",
  1947 => x"388c08fe",
  1948 => x"fc0508ff",
  1949 => x"058c08fe",
  1950 => x"fc050c8c",
  1951 => x"08ff8405",
  1952 => x"088c08ff",
  1953 => x"ac050805",
  1954 => x"8c08ff84",
  1955 => x"050c8c08",
  1956 => x"ffac0508",
  1957 => x"8c08ff84",
  1958 => x"050826b1",
  1959 => x"388c08ff",
  1960 => x"8405088c",
  1961 => x"08ff8805",
  1962 => x"0827a238",
  1963 => x"8c08fefc",
  1964 => x"0508ff05",
  1965 => x"8c08fefc",
  1966 => x"050c8c08",
  1967 => x"ff840508",
  1968 => x"8c08ffac",
  1969 => x"0508058c",
  1970 => x"08ff8405",
  1971 => x"0c8c08ff",
  1972 => x"8405088c",
  1973 => x"08ff8805",
  1974 => x"08318c08",
  1975 => x"ff84050c",
  1976 => x"8c08fef8",
  1977 => x"05087090",
  1978 => x"2b708c08",
  1979 => x"fefc0508",
  1980 => x"078c08ff",
  1981 => x"98050c8c",
  1982 => x"08ff8405",
  1983 => x"088c08ff",
  1984 => x"a4050c51",
  1985 => x"548c08c8",
  1986 => x"0508802e",
  1987 => x"8ea3388c",
  1988 => x"08ffa405",
  1989 => x"088c08ff",
  1990 => x"8c05082a",
  1991 => x"8c08ffb4",
  1992 => x"050c800b",
  1993 => x"8c08ffb0",
  1994 => x"050c8c08",
  1995 => x"c8050856",
  1996 => x"8c08ffb0",
  1997 => x"05088c08",
  1998 => x"ffb40508",
  1999 => x"56547376",
  2000 => x"0c748417",
  2001 => x"0c8dea39",
  2002 => x"8c08ffa0",
  2003 => x"05088c08",
  2004 => x"ffa80508",
  2005 => x"2780d138",
  2006 => x"800b8c08",
  2007 => x"ff98050c",
  2008 => x"800b8c08",
  2009 => x"ff94050c",
  2010 => x"8c08c805",
  2011 => x"08802e8d",
  2012 => x"c0388c08",
  2013 => x"ffa40508",
  2014 => x"8c08ffb4",
  2015 => x"050c8c08",
  2016 => x"ffa00508",
  2017 => x"8c08ffb0",
  2018 => x"050c8c08",
  2019 => x"c8050856",
  2020 => x"8c08ffb0",
  2021 => x"05088c08",
  2022 => x"ffb40508",
  2023 => x"56547376",
  2024 => x"0c748417",
  2025 => x"0c8d8a39",
  2026 => x"8c08ffa8",
  2027 => x"05088c08",
  2028 => x"fef0050c",
  2029 => x"8c08fef0",
  2030 => x"050883ff",
  2031 => x"ff26a038",
  2032 => x"8c08fef0",
  2033 => x"050881ff",
  2034 => x"268b3880",
  2035 => x"0b8c08fe",
  2036 => x"d0050ca9",
  2037 => x"39880b8c",
  2038 => x"08fed005",
  2039 => x"0c9f398c",
  2040 => x"08fef005",
  2041 => x"08fe800a",
  2042 => x"268b3890",
  2043 => x"0b8c08fe",
  2044 => x"d0050c89",
  2045 => x"39980b8c",
  2046 => x"08fed005",
  2047 => x"0c8c08fe",
  2048 => x"d005088c",
  2049 => x"08fef405",
  2050 => x"0c8c08fe",
  2051 => x"f005088c",
  2052 => x"08fef405",
  2053 => x"082a80f6",
  2054 => x"c811338c",
  2055 => x"08fef405",
  2056 => x"0811a071",
  2057 => x"318c08ff",
  2058 => x"8c050c51",
  2059 => x"51548c08",
  2060 => x"ff8c0508",
  2061 => x"81d9388c",
  2062 => x"08ffa005",
  2063 => x"088c08ff",
  2064 => x"a8050826",
  2065 => x"93388c08",
  2066 => x"ffa40508",
  2067 => x"8c08ffac",
  2068 => x"05082784",
  2069 => x"3880e839",
  2070 => x"810b8c08",
  2071 => x"ff98050c",
  2072 => x"8c08ffa4",
  2073 => x"05088c08",
  2074 => x"ffac0508",
  2075 => x"318c08fe",
  2076 => x"f0050c8c",
  2077 => x"08ffa005",
  2078 => x"088c08ff",
  2079 => x"a8050831",
  2080 => x"708c08fe",
  2081 => x"cc050c54",
  2082 => x"8c08ffa4",
  2083 => x"05088c08",
  2084 => x"fef00508",
  2085 => x"278f388c",
  2086 => x"08fecc05",
  2087 => x"08ff058c",
  2088 => x"08fecc05",
  2089 => x"0c8c08fe",
  2090 => x"cc05088c",
  2091 => x"08ffa005",
  2092 => x"0c8c08fe",
  2093 => x"f005088c",
  2094 => x"08ffa405",
  2095 => x"0c893980",
  2096 => x"0b8c08ff",
  2097 => x"98050c80",
  2098 => x"0b8c08ff",
  2099 => x"94050c8c",
  2100 => x"08c80508",
  2101 => x"802e8ad9",
  2102 => x"388c08ff",
  2103 => x"a405088c",
  2104 => x"08ffb405",
  2105 => x"0c8c08ff",
  2106 => x"a005088c",
  2107 => x"08ffb005",
  2108 => x"0c8c08c8",
  2109 => x"0508568c",
  2110 => x"08ffb005",
  2111 => x"088c08ff",
  2112 => x"b4050856",
  2113 => x"5473760c",
  2114 => x"7484170c",
  2115 => x"8aa339a0",
  2116 => x"0b8c08ff",
  2117 => x"8c050831",
  2118 => x"8c08ff90",
  2119 => x"050c8c08",
  2120 => x"ffa80508",
  2121 => x"8c08ff8c",
  2122 => x"05082b8c",
  2123 => x"08ffac05",
  2124 => x"088c08ff",
  2125 => x"9005082a",
  2126 => x"7072078c",
  2127 => x"08ffa805",
  2128 => x"0c8c08ff",
  2129 => x"ac05088c",
  2130 => x"08ff8c05",
  2131 => x"082b8c08",
  2132 => x"ffac050c",
  2133 => x"8c08ffa0",
  2134 => x"05088c08",
  2135 => x"ff900508",
  2136 => x"2a8c08ff",
  2137 => x"9c050c8c",
  2138 => x"08ffa005",
  2139 => x"088c08ff",
  2140 => x"8c05082b",
  2141 => x"8c08ffa4",
  2142 => x"05088c08",
  2143 => x"ff900508",
  2144 => x"2a707207",
  2145 => x"8c08ffa0",
  2146 => x"050c8c08",
  2147 => x"ffa40508",
  2148 => x"8c08ff8c",
  2149 => x"05082b8c",
  2150 => x"08ffa405",
  2151 => x"0c8c08ff",
  2152 => x"a8050890",
  2153 => x"2a8c08fe",
  2154 => x"f8050c8c",
  2155 => x"08ffa805",
  2156 => x"0883ffff",
  2157 => x"068c08fe",
  2158 => x"fc050c8c",
  2159 => x"08ff9c05",
  2160 => x"088c08fe",
  2161 => x"f8050857",
  2162 => x"70565152",
  2163 => x"5255558a",
  2164 => x"c03f8008",
  2165 => x"708c08ff",
  2166 => x"88050c8c",
  2167 => x"08fef805",
  2168 => x"08538c08",
  2169 => x"ff9c0508",
  2170 => x"52548a80",
  2171 => x"3f800870",
  2172 => x"8c08ff80",
  2173 => x"050c8c08",
  2174 => x"ff800508",
  2175 => x"8c08fefc",
  2176 => x"05082970",
  2177 => x"8c08fee8",
  2178 => x"050c8c08",
  2179 => x"ff880508",
  2180 => x"70902b8c",
  2181 => x"08ffa005",
  2182 => x"08902a70",
  2183 => x"72078c08",
  2184 => x"ff88050c",
  2185 => x"52585151",
  2186 => x"548c08ff",
  2187 => x"8805088c",
  2188 => x"08fee805",
  2189 => x"082780e1",
  2190 => x"388c08ff",
  2191 => x"800508ff",
  2192 => x"058c08ff",
  2193 => x"80050c8c",
  2194 => x"08ff8805",
  2195 => x"088c08ff",
  2196 => x"a8050805",
  2197 => x"8c08ff88",
  2198 => x"050c8c08",
  2199 => x"ffa80508",
  2200 => x"8c08ff88",
  2201 => x"050826b1",
  2202 => x"388c08ff",
  2203 => x"8805088c",
  2204 => x"08fee805",
  2205 => x"0827a238",
  2206 => x"8c08ff80",
  2207 => x"0508ff05",
  2208 => x"8c08ff80",
  2209 => x"050c8c08",
  2210 => x"ff880508",
  2211 => x"8c08ffa8",
  2212 => x"0508058c",
  2213 => x"08ff8805",
  2214 => x"0c8c08ff",
  2215 => x"8805088c",
  2216 => x"08fee805",
  2217 => x"08318c08",
  2218 => x"ff88050c",
  2219 => x"8c08ff88",
  2220 => x"05088c08",
  2221 => x"fef80508",
  2222 => x"53705254",
  2223 => x"88d33f80",
  2224 => x"08708c08",
  2225 => x"feec050c",
  2226 => x"8c08fef8",
  2227 => x"0508538c",
  2228 => x"08ff8805",
  2229 => x"08525488",
  2230 => x"933f8008",
  2231 => x"708c08ff",
  2232 => x"84050c8c",
  2233 => x"08ff8405",
  2234 => x"088c08fe",
  2235 => x"fc050829",
  2236 => x"708c08fe",
  2237 => x"e8050c8c",
  2238 => x"08feec05",
  2239 => x"0870902b",
  2240 => x"8c08ffa0",
  2241 => x"050883ff",
  2242 => x"ff067072",
  2243 => x"078c08fe",
  2244 => x"ec050c52",
  2245 => x"58515154",
  2246 => x"8c08feec",
  2247 => x"05088c08",
  2248 => x"fee80508",
  2249 => x"2780e138",
  2250 => x"8c08ff84",
  2251 => x"0508ff05",
  2252 => x"8c08ff84",
  2253 => x"050c8c08",
  2254 => x"feec0508",
  2255 => x"8c08ffa8",
  2256 => x"0508058c",
  2257 => x"08feec05",
  2258 => x"0c8c08ff",
  2259 => x"a805088c",
  2260 => x"08feec05",
  2261 => x"0826b138",
  2262 => x"8c08feec",
  2263 => x"05088c08",
  2264 => x"fee80508",
  2265 => x"27a2388c",
  2266 => x"08ff8405",
  2267 => x"08ff058c",
  2268 => x"08ff8405",
  2269 => x"0c8c08fe",
  2270 => x"ec05088c",
  2271 => x"08ffa805",
  2272 => x"08058c08",
  2273 => x"feec050c",
  2274 => x"8c08feec",
  2275 => x"05088c08",
  2276 => x"fee80508",
  2277 => x"318c08fe",
  2278 => x"ec050c8c",
  2279 => x"08ff8005",
  2280 => x"0870902b",
  2281 => x"708c08ff",
  2282 => x"84050807",
  2283 => x"8c08ff98",
  2284 => x"050c8c08",
  2285 => x"feec0508",
  2286 => x"8c08ffa0",
  2287 => x"050c8c08",
  2288 => x"ff980508",
  2289 => x"83ffff06",
  2290 => x"8c08ff80",
  2291 => x"050c8c08",
  2292 => x"ff980508",
  2293 => x"902a8c08",
  2294 => x"ff88050c",
  2295 => x"8c08ffac",
  2296 => x"050883ff",
  2297 => x"ff068c08",
  2298 => x"ff84050c",
  2299 => x"8c08ffac",
  2300 => x"0508902a",
  2301 => x"8c08fee4",
  2302 => x"050c8c08",
  2303 => x"ff800508",
  2304 => x"8c08ff84",
  2305 => x"05082970",
  2306 => x"8c08fee8",
  2307 => x"050c8c08",
  2308 => x"ff800508",
  2309 => x"8c08fee4",
  2310 => x"05082970",
  2311 => x"8c08feec",
  2312 => x"050c8c08",
  2313 => x"ff880508",
  2314 => x"8c08ff84",
  2315 => x"05082970",
  2316 => x"8c08fef8",
  2317 => x"050c8c08",
  2318 => x"ff880508",
  2319 => x"8c08fee4",
  2320 => x"05082970",
  2321 => x"8c08fefc",
  2322 => x"050c8c08",
  2323 => x"fee80508",
  2324 => x"902a8c08",
  2325 => x"feec0508",
  2326 => x"118c08fe",
  2327 => x"ec050c8c",
  2328 => x"08feec05",
  2329 => x"088c08fe",
  2330 => x"f8050805",
  2331 => x"8c08feec",
  2332 => x"050c5151",
  2333 => x"51515151",
  2334 => x"548c08fe",
  2335 => x"ec05088c",
  2336 => x"08fef805",
  2337 => x"08279138",
  2338 => x"8c08fefc",
  2339 => x"05088480",
  2340 => x"80058c08",
  2341 => x"fefc050c",
  2342 => x"8c08feec",
  2343 => x"0508902a",
  2344 => x"8c08fefc",
  2345 => x"0508118c",
  2346 => x"08fef005",
  2347 => x"0c8c08fe",
  2348 => x"ec050883",
  2349 => x"ffff0670",
  2350 => x"902b8c08",
  2351 => x"fee80508",
  2352 => x"83ffff06",
  2353 => x"70128c08",
  2354 => x"fef4050c",
  2355 => x"52575154",
  2356 => x"8c08fef0",
  2357 => x"05088c08",
  2358 => x"ffa00508",
  2359 => x"26a6388c",
  2360 => x"08fef005",
  2361 => x"088c08ff",
  2362 => x"a005082e",
  2363 => x"09810680",
  2364 => x"fe388c08",
  2365 => x"fef40508",
  2366 => x"8c08ffa4",
  2367 => x"05082684",
  2368 => x"3880ec39",
  2369 => x"8c08ff98",
  2370 => x"0508ff05",
  2371 => x"8c08ff98",
  2372 => x"050c8c08",
  2373 => x"fef40508",
  2374 => x"8c08ffac",
  2375 => x"0508318c",
  2376 => x"08fee405",
  2377 => x"0c8c08fe",
  2378 => x"f005088c",
  2379 => x"08ffa805",
  2380 => x"0831708c",
  2381 => x"08fec805",
  2382 => x"0c548c08",
  2383 => x"fef40508",
  2384 => x"8c08fee4",
  2385 => x"0508278f",
  2386 => x"388c08fe",
  2387 => x"c80508ff",
  2388 => x"058c08fe",
  2389 => x"c8050c8c",
  2390 => x"08fec805",
  2391 => x"088c08fe",
  2392 => x"f0050c8c",
  2393 => x"08fee405",
  2394 => x"088c08fe",
  2395 => x"f4050c80",
  2396 => x"0b8c08ff",
  2397 => x"94050c8c",
  2398 => x"08c80508",
  2399 => x"802e81b1",
  2400 => x"388c08ff",
  2401 => x"a405088c",
  2402 => x"08fef405",
  2403 => x"08318c08",
  2404 => x"fee4050c",
  2405 => x"8c08ffa0",
  2406 => x"05088c08",
  2407 => x"fef00508",
  2408 => x"31708c08",
  2409 => x"fec4050c",
  2410 => x"548c08ff",
  2411 => x"a405088c",
  2412 => x"08fee405",
  2413 => x"08278f38",
  2414 => x"8c08fec4",
  2415 => x"0508ff05",
  2416 => x"8c08fec4",
  2417 => x"050c8c08",
  2418 => x"fec40508",
  2419 => x"8c08ffa0",
  2420 => x"050c8c08",
  2421 => x"fee40508",
  2422 => x"8c08ffa4",
  2423 => x"050c8c08",
  2424 => x"ffa00508",
  2425 => x"8c08ff90",
  2426 => x"05082b8c",
  2427 => x"08ffa405",
  2428 => x"088c08ff",
  2429 => x"8c05082a",
  2430 => x"7072078c",
  2431 => x"08ffb405",
  2432 => x"0c8c08ff",
  2433 => x"a005088c",
  2434 => x"08ff8c05",
  2435 => x"082a8c08",
  2436 => x"ffb0050c",
  2437 => x"8c08c805",
  2438 => x"08585555",
  2439 => x"8c08ffb0",
  2440 => x"05088c08",
  2441 => x"ffb40508",
  2442 => x"56547376",
  2443 => x"0c748417",
  2444 => x"0c800b8c",
  2445 => x"08fedc05",
  2446 => x"0c800b8c",
  2447 => x"08fee005",
  2448 => x"0c8c08ff",
  2449 => x"9405088c",
  2450 => x"08fedc05",
  2451 => x"0c8c08ff",
  2452 => x"9805088c",
  2453 => x"08fee005",
  2454 => x"0c8c08fe",
  2455 => x"dc05088c",
  2456 => x"08fee005",
  2457 => x"08565473",
  2458 => x"8c08c005",
  2459 => x"0c748c08",
  2460 => x"c4050c8c",
  2461 => x"08c00508",
  2462 => x"8c08c405",
  2463 => x"08565473",
  2464 => x"8c08dc05",
  2465 => x"0c748c08",
  2466 => x"e0050c8c",
  2467 => x"08fc0508",
  2468 => x"802eb338",
  2469 => x"8c08c005",
  2470 => x"548c08dc",
  2471 => x"05088c08",
  2472 => x"e0050857",
  2473 => x"55745275",
  2474 => x"537351d8",
  2475 => x"d73f8c08",
  2476 => x"c005088c",
  2477 => x"08c40508",
  2478 => x"5654738c",
  2479 => x"08dc050c",
  2480 => x"748c08e0",
  2481 => x"050c8c08",
  2482 => x"dc05088c",
  2483 => x"08e00508",
  2484 => x"8c088805",
  2485 => x"08585654",
  2486 => x"73760c74",
  2487 => x"84170c8c",
  2488 => x"08880508",
  2489 => x"800cb63d",
  2490 => x"0d8c0c04",
  2491 => x"8c08028c",
  2492 => x"0cfd3d0d",
  2493 => x"80538c08",
  2494 => x"8c050852",
  2495 => x"8c088805",
  2496 => x"085182de",
  2497 => x"3f800870",
  2498 => x"800c5485",
  2499 => x"3d0d8c0c",
  2500 => x"048c0802",
  2501 => x"8c0cfd3d",
  2502 => x"0d81538c",
  2503 => x"088c0508",
  2504 => x"528c0888",
  2505 => x"05085182",
  2506 => x"b93f8008",
  2507 => x"70800c54",
  2508 => x"853d0d8c",
  2509 => x"0c048c08",
  2510 => x"028c0cf9",
  2511 => x"3d0d800b",
  2512 => x"8c08fc05",
  2513 => x"0c8c0888",
  2514 => x"05088025",
  2515 => x"ab388c08",
  2516 => x"88050830",
  2517 => x"8c088805",
  2518 => x"0c800b8c",
  2519 => x"08f4050c",
  2520 => x"8c08fc05",
  2521 => x"08883881",
  2522 => x"0b8c08f4",
  2523 => x"050c8c08",
  2524 => x"f405088c",
  2525 => x"08fc050c",
  2526 => x"8c088c05",
  2527 => x"088025ab",
  2528 => x"388c088c",
  2529 => x"0508308c",
  2530 => x"088c050c",
  2531 => x"800b8c08",
  2532 => x"f0050c8c",
  2533 => x"08fc0508",
  2534 => x"8838810b",
  2535 => x"8c08f005",
  2536 => x"0c8c08f0",
  2537 => x"05088c08",
  2538 => x"fc050c80",
  2539 => x"538c088c",
  2540 => x"0508528c",
  2541 => x"08880508",
  2542 => x"5181a73f",
  2543 => x"8008708c",
  2544 => x"08f8050c",
  2545 => x"548c08fc",
  2546 => x"0508802e",
  2547 => x"8c388c08",
  2548 => x"f8050830",
  2549 => x"8c08f805",
  2550 => x"0c8c08f8",
  2551 => x"05087080",
  2552 => x"0c54893d",
  2553 => x"0d8c0c04",
  2554 => x"8c08028c",
  2555 => x"0cfb3d0d",
  2556 => x"800b8c08",
  2557 => x"fc050c8c",
  2558 => x"08880508",
  2559 => x"80259338",
  2560 => x"8c088805",
  2561 => x"08308c08",
  2562 => x"88050c81",
  2563 => x"0b8c08fc",
  2564 => x"050c8c08",
  2565 => x"8c050880",
  2566 => x"258c388c",
  2567 => x"088c0508",
  2568 => x"308c088c",
  2569 => x"050c8153",
  2570 => x"8c088c05",
  2571 => x"08528c08",
  2572 => x"88050851",
  2573 => x"ad3f8008",
  2574 => x"708c08f8",
  2575 => x"050c548c",
  2576 => x"08fc0508",
  2577 => x"802e8c38",
  2578 => x"8c08f805",
  2579 => x"08308c08",
  2580 => x"f8050c8c",
  2581 => x"08f80508",
  2582 => x"70800c54",
  2583 => x"873d0d8c",
  2584 => x"0c048c08",
  2585 => x"028c0cfd",
  2586 => x"3d0d810b",
  2587 => x"8c08fc05",
  2588 => x"0c800b8c",
  2589 => x"08f8050c",
  2590 => x"8c088c05",
  2591 => x"088c0888",
  2592 => x"050827ac",
  2593 => x"388c08fc",
  2594 => x"0508802e",
  2595 => x"a338800b",
  2596 => x"8c088c05",
  2597 => x"08249938",
  2598 => x"8c088c05",
  2599 => x"08108c08",
  2600 => x"8c050c8c",
  2601 => x"08fc0508",
  2602 => x"108c08fc",
  2603 => x"050cc939",
  2604 => x"8c08fc05",
  2605 => x"08802e80",
  2606 => x"c9388c08",
  2607 => x"8c05088c",
  2608 => x"08880508",
  2609 => x"26a1388c",
  2610 => x"08880508",
  2611 => x"8c088c05",
  2612 => x"08318c08",
  2613 => x"88050c8c",
  2614 => x"08f80508",
  2615 => x"8c08fc05",
  2616 => x"08078c08",
  2617 => x"f8050c8c",
  2618 => x"08fc0508",
  2619 => x"812a8c08",
  2620 => x"fc050c8c",
  2621 => x"088c0508",
  2622 => x"812a8c08",
  2623 => x"8c050cff",
  2624 => x"af398c08",
  2625 => x"90050880",
  2626 => x"2e8f388c",
  2627 => x"08880508",
  2628 => x"708c08f4",
  2629 => x"050c518d",
  2630 => x"398c08f8",
  2631 => x"0508708c",
  2632 => x"08f4050c",
  2633 => x"518c08f4",
  2634 => x"0508800c",
  2635 => x"853d0d8c",
  2636 => x"0c04ff3d",
  2637 => x"0d735281",
  2638 => x"81c80851",
  2639 => x"963f833d",
  2640 => x"0d04ff3d",
  2641 => x"0d735281",
  2642 => x"81c80851",
  2643 => x"90953f83",
  2644 => x"3d0d04f3",
  2645 => x"3d0d7f61",
  2646 => x"8b1170f8",
  2647 => x"065c5555",
  2648 => x"5e729626",
  2649 => x"83389059",
  2650 => x"80792474",
  2651 => x"7a260753",
  2652 => x"80547274",
  2653 => x"2e098106",
  2654 => x"80cb387d",
  2655 => x"518ce33f",
  2656 => x"7883f726",
  2657 => x"80c63878",
  2658 => x"832a7010",
  2659 => x"101080f9",
  2660 => x"c0058c11",
  2661 => x"0859595a",
  2662 => x"76782e83",
  2663 => x"b0388417",
  2664 => x"08fc0656",
  2665 => x"8c170888",
  2666 => x"1808718c",
  2667 => x"120c8812",
  2668 => x"0c587517",
  2669 => x"84110881",
  2670 => x"0784120c",
  2671 => x"537d518c",
  2672 => x"a23f8817",
  2673 => x"5473800c",
  2674 => x"8f3d0d04",
  2675 => x"78892a79",
  2676 => x"832a5b53",
  2677 => x"72802ebf",
  2678 => x"3878862a",
  2679 => x"b8055a84",
  2680 => x"7327b438",
  2681 => x"80db135a",
  2682 => x"947327ab",
  2683 => x"38788c2a",
  2684 => x"80ee055a",
  2685 => x"80d47327",
  2686 => x"9e38788f",
  2687 => x"2a80f705",
  2688 => x"5a82d473",
  2689 => x"27913878",
  2690 => x"922a80fc",
  2691 => x"055a8ad4",
  2692 => x"73278438",
  2693 => x"80fe5a79",
  2694 => x"10101080",
  2695 => x"f9c0058c",
  2696 => x"11085855",
  2697 => x"76752ea3",
  2698 => x"38841708",
  2699 => x"fc06707a",
  2700 => x"31555673",
  2701 => x"8f2488d5",
  2702 => x"38738025",
  2703 => x"fee6388c",
  2704 => x"17085776",
  2705 => x"752e0981",
  2706 => x"06df3881",
  2707 => x"1a5a80f9",
  2708 => x"d0085776",
  2709 => x"80f9c82e",
  2710 => x"82c03884",
  2711 => x"1708fc06",
  2712 => x"707a3155",
  2713 => x"56738f24",
  2714 => x"81f93880",
  2715 => x"f9c80b80",
  2716 => x"f9d40c80",
  2717 => x"f9c80b80",
  2718 => x"f9d00c73",
  2719 => x"8025feb2",
  2720 => x"3883ff76",
  2721 => x"2783df38",
  2722 => x"75892a76",
  2723 => x"832a5553",
  2724 => x"72802ebf",
  2725 => x"3875862a",
  2726 => x"b8055484",
  2727 => x"7327b438",
  2728 => x"80db1354",
  2729 => x"947327ab",
  2730 => x"38758c2a",
  2731 => x"80ee0554",
  2732 => x"80d47327",
  2733 => x"9e38758f",
  2734 => x"2a80f705",
  2735 => x"5482d473",
  2736 => x"27913875",
  2737 => x"922a80fc",
  2738 => x"05548ad4",
  2739 => x"73278438",
  2740 => x"80fe5473",
  2741 => x"10101080",
  2742 => x"f9c00588",
  2743 => x"11085658",
  2744 => x"74782e86",
  2745 => x"cf388415",
  2746 => x"08fc0653",
  2747 => x"7573278d",
  2748 => x"38881508",
  2749 => x"5574782e",
  2750 => x"098106ea",
  2751 => x"388c1508",
  2752 => x"80f9c00b",
  2753 => x"84050871",
  2754 => x"8c1a0c76",
  2755 => x"881a0c78",
  2756 => x"88130c78",
  2757 => x"8c180c5d",
  2758 => x"58795380",
  2759 => x"7a2483e6",
  2760 => x"3872822c",
  2761 => x"81712b5c",
  2762 => x"537a7c26",
  2763 => x"8198387b",
  2764 => x"7b065372",
  2765 => x"82f13879",
  2766 => x"fc068405",
  2767 => x"5a7a1070",
  2768 => x"7d06545b",
  2769 => x"7282e038",
  2770 => x"841a5af1",
  2771 => x"3988178c",
  2772 => x"11085858",
  2773 => x"76782e09",
  2774 => x"8106fcc2",
  2775 => x"38821a5a",
  2776 => x"fdec3978",
  2777 => x"17798107",
  2778 => x"84190c70",
  2779 => x"80f9d40c",
  2780 => x"7080f9d0",
  2781 => x"0c80f9c8",
  2782 => x"0b8c120c",
  2783 => x"8c110888",
  2784 => x"120c7481",
  2785 => x"0784120c",
  2786 => x"74117571",
  2787 => x"0c51537d",
  2788 => x"5188d03f",
  2789 => x"881754fc",
  2790 => x"ac3980f9",
  2791 => x"c00b8405",
  2792 => x"087a545c",
  2793 => x"798025fe",
  2794 => x"f83882da",
  2795 => x"397a097c",
  2796 => x"067080f9",
  2797 => x"c00b8405",
  2798 => x"0c5c7a10",
  2799 => x"5b7a7c26",
  2800 => x"85387a85",
  2801 => x"b83880f9",
  2802 => x"c00b8805",
  2803 => x"08708412",
  2804 => x"08fc0670",
  2805 => x"7c317c72",
  2806 => x"268f7225",
  2807 => x"0757575c",
  2808 => x"5d557280",
  2809 => x"2e80db38",
  2810 => x"797a1680",
  2811 => x"f9b8081b",
  2812 => x"90115a55",
  2813 => x"575b80f9",
  2814 => x"b408ff2e",
  2815 => x"8838a08f",
  2816 => x"13e08006",
  2817 => x"5776527d",
  2818 => x"5187d93f",
  2819 => x"80085480",
  2820 => x"08ff2e90",
  2821 => x"38800876",
  2822 => x"27829938",
  2823 => x"7480f9c0",
  2824 => x"2e829138",
  2825 => x"80f9c00b",
  2826 => x"88050855",
  2827 => x"841508fc",
  2828 => x"06707a31",
  2829 => x"7a72268f",
  2830 => x"72250752",
  2831 => x"55537283",
  2832 => x"e6387479",
  2833 => x"81078417",
  2834 => x"0c791670",
  2835 => x"80f9c00b",
  2836 => x"88050c75",
  2837 => x"81078412",
  2838 => x"0c547e52",
  2839 => x"5787843f",
  2840 => x"881754fa",
  2841 => x"e0397583",
  2842 => x"2a705454",
  2843 => x"80742481",
  2844 => x"9b387282",
  2845 => x"2c81712b",
  2846 => x"80f9c408",
  2847 => x"077080f9",
  2848 => x"c00b8405",
  2849 => x"0c751010",
  2850 => x"1080f9c0",
  2851 => x"05881108",
  2852 => x"585a5d53",
  2853 => x"778c180c",
  2854 => x"7488180c",
  2855 => x"7688190c",
  2856 => x"768c160c",
  2857 => x"fcf33979",
  2858 => x"7a101010",
  2859 => x"80f9c005",
  2860 => x"7057595d",
  2861 => x"8c150857",
  2862 => x"76752ea3",
  2863 => x"38841708",
  2864 => x"fc06707a",
  2865 => x"31555673",
  2866 => x"8f2483ca",
  2867 => x"38738025",
  2868 => x"8481388c",
  2869 => x"17085776",
  2870 => x"752e0981",
  2871 => x"06df3888",
  2872 => x"15811b70",
  2873 => x"8306555b",
  2874 => x"5572c938",
  2875 => x"7c830653",
  2876 => x"72802efd",
  2877 => x"b838ff1d",
  2878 => x"f819595d",
  2879 => x"88180878",
  2880 => x"2eea38fd",
  2881 => x"b539831a",
  2882 => x"53fc9639",
  2883 => x"83147082",
  2884 => x"2c81712b",
  2885 => x"80f9c408",
  2886 => x"077080f9",
  2887 => x"c00b8405",
  2888 => x"0c761010",
  2889 => x"1080f9c0",
  2890 => x"05881108",
  2891 => x"595b5e51",
  2892 => x"53fee139",
  2893 => x"80f98408",
  2894 => x"17588008",
  2895 => x"762e818d",
  2896 => x"3880f9b4",
  2897 => x"08ff2e83",
  2898 => x"ec387376",
  2899 => x"311880f9",
  2900 => x"840c7387",
  2901 => x"06705753",
  2902 => x"72802e88",
  2903 => x"38887331",
  2904 => x"70155556",
  2905 => x"76149fff",
  2906 => x"06a08071",
  2907 => x"31177054",
  2908 => x"7f535753",
  2909 => x"84ee3f80",
  2910 => x"08538008",
  2911 => x"ff2e81a0",
  2912 => x"3880f984",
  2913 => x"08167080",
  2914 => x"f9840c74",
  2915 => x"7580f9c0",
  2916 => x"0b88050c",
  2917 => x"74763118",
  2918 => x"70810751",
  2919 => x"5556587b",
  2920 => x"80f9c02e",
  2921 => x"839c3879",
  2922 => x"8f2682cb",
  2923 => x"38810b84",
  2924 => x"150c8415",
  2925 => x"08fc0670",
  2926 => x"7a317a72",
  2927 => x"268f7225",
  2928 => x"07525553",
  2929 => x"72802efc",
  2930 => x"f93880db",
  2931 => x"3980089f",
  2932 => x"ff065372",
  2933 => x"feeb3877",
  2934 => x"80f9840c",
  2935 => x"80f9c00b",
  2936 => x"8805087b",
  2937 => x"18810784",
  2938 => x"120c5580",
  2939 => x"f9b00878",
  2940 => x"27863877",
  2941 => x"80f9b00c",
  2942 => x"80f9ac08",
  2943 => x"7827fcac",
  2944 => x"387780f9",
  2945 => x"ac0c8415",
  2946 => x"08fc0670",
  2947 => x"7a317a72",
  2948 => x"268f7225",
  2949 => x"07525553",
  2950 => x"72802efc",
  2951 => x"a5388839",
  2952 => x"80745456",
  2953 => x"fedb397d",
  2954 => x"5183b83f",
  2955 => x"800b800c",
  2956 => x"8f3d0d04",
  2957 => x"73538074",
  2958 => x"24a93872",
  2959 => x"822c8171",
  2960 => x"2b80f9c4",
  2961 => x"08077080",
  2962 => x"f9c00b84",
  2963 => x"050c5d53",
  2964 => x"778c180c",
  2965 => x"7488180c",
  2966 => x"7688190c",
  2967 => x"768c160c",
  2968 => x"f9b73983",
  2969 => x"1470822c",
  2970 => x"81712b80",
  2971 => x"f9c40807",
  2972 => x"7080f9c0",
  2973 => x"0b84050c",
  2974 => x"5e5153d4",
  2975 => x"397b7b06",
  2976 => x"5372fca3",
  2977 => x"38841a7b",
  2978 => x"105c5af1",
  2979 => x"39ff1a81",
  2980 => x"11515af7",
  2981 => x"b9397817",
  2982 => x"79810784",
  2983 => x"190c8c18",
  2984 => x"08881908",
  2985 => x"718c120c",
  2986 => x"88120c59",
  2987 => x"7080f9d4",
  2988 => x"0c7080f9",
  2989 => x"d00c80f9",
  2990 => x"c80b8c12",
  2991 => x"0c8c1108",
  2992 => x"88120c74",
  2993 => x"81078412",
  2994 => x"0c741175",
  2995 => x"710c5153",
  2996 => x"f9bd3975",
  2997 => x"17841108",
  2998 => x"81078412",
  2999 => x"0c538c17",
  3000 => x"08881808",
  3001 => x"718c120c",
  3002 => x"88120c58",
  3003 => x"7d5181f3",
  3004 => x"3f881754",
  3005 => x"f5cf3972",
  3006 => x"84150cf4",
  3007 => x"1af80670",
  3008 => x"841e0881",
  3009 => x"0607841e",
  3010 => x"0c701d54",
  3011 => x"5b850b84",
  3012 => x"140c850b",
  3013 => x"88140c8f",
  3014 => x"7b27fdcf",
  3015 => x"38881c52",
  3016 => x"7d5184bf",
  3017 => x"3f80f9c0",
  3018 => x"0b880508",
  3019 => x"80f98408",
  3020 => x"5955fdb7",
  3021 => x"397780f9",
  3022 => x"840c7380",
  3023 => x"f9b40cfc",
  3024 => x"91397284",
  3025 => x"150cfda3",
  3026 => x"39fc3d0d",
  3027 => x"7670797b",
  3028 => x"55555555",
  3029 => x"8f72278c",
  3030 => x"38727507",
  3031 => x"83065170",
  3032 => x"802ea738",
  3033 => x"ff125271",
  3034 => x"ff2e9838",
  3035 => x"72708105",
  3036 => x"54337470",
  3037 => x"81055634",
  3038 => x"ff125271",
  3039 => x"ff2e0981",
  3040 => x"06ea3874",
  3041 => x"800c863d",
  3042 => x"0d047451",
  3043 => x"72708405",
  3044 => x"54087170",
  3045 => x"8405530c",
  3046 => x"72708405",
  3047 => x"54087170",
  3048 => x"8405530c",
  3049 => x"72708405",
  3050 => x"54087170",
  3051 => x"8405530c",
  3052 => x"72708405",
  3053 => x"54087170",
  3054 => x"8405530c",
  3055 => x"f0125271",
  3056 => x"8f26c938",
  3057 => x"83722795",
  3058 => x"38727084",
  3059 => x"05540871",
  3060 => x"70840553",
  3061 => x"0cfc1252",
  3062 => x"718326ed",
  3063 => x"387054ff",
  3064 => x"83390404",
  3065 => x"fd3d0d80",
  3066 => x"0b81d998",
  3067 => x"0c765187",
  3068 => x"c83f8008",
  3069 => x"538008ff",
  3070 => x"2e883872",
  3071 => x"800c853d",
  3072 => x"0d0481d9",
  3073 => x"98085473",
  3074 => x"802ef038",
  3075 => x"7574710c",
  3076 => x"5272800c",
  3077 => x"853d0d04",
  3078 => x"fb3d0d77",
  3079 => x"79707207",
  3080 => x"83065354",
  3081 => x"52709338",
  3082 => x"71737308",
  3083 => x"54565471",
  3084 => x"73082e80",
  3085 => x"c4387375",
  3086 => x"54527133",
  3087 => x"7081ff06",
  3088 => x"52547080",
  3089 => x"2e9d3872",
  3090 => x"33557075",
  3091 => x"2e098106",
  3092 => x"95388112",
  3093 => x"81147133",
  3094 => x"7081ff06",
  3095 => x"54565452",
  3096 => x"70e53872",
  3097 => x"33557381",
  3098 => x"ff067581",
  3099 => x"ff067171",
  3100 => x"31800c52",
  3101 => x"52873d0d",
  3102 => x"04710970",
  3103 => x"f7fbfdff",
  3104 => x"140670f8",
  3105 => x"84828180",
  3106 => x"06515151",
  3107 => x"70973884",
  3108 => x"14841671",
  3109 => x"08545654",
  3110 => x"7175082e",
  3111 => x"dc387375",
  3112 => x"5452ff96",
  3113 => x"39800b80",
  3114 => x"0c873d0d",
  3115 => x"04fb3d0d",
  3116 => x"77705256",
  3117 => x"feac3f80",
  3118 => x"f9c00b88",
  3119 => x"05088411",
  3120 => x"08fc0670",
  3121 => x"7b319fef",
  3122 => x"05e08006",
  3123 => x"e0800556",
  3124 => x"5653a080",
  3125 => x"74249438",
  3126 => x"80527551",
  3127 => x"fe863f80",
  3128 => x"f9c80815",
  3129 => x"53728008",
  3130 => x"2e8f3875",
  3131 => x"51fdf43f",
  3132 => x"80537280",
  3133 => x"0c873d0d",
  3134 => x"04733052",
  3135 => x"7551fde4",
  3136 => x"3f8008ff",
  3137 => x"2ea83880",
  3138 => x"f9c00b88",
  3139 => x"05087575",
  3140 => x"31810784",
  3141 => x"120c5380",
  3142 => x"f9840874",
  3143 => x"3180f984",
  3144 => x"0c7551fd",
  3145 => x"be3f810b",
  3146 => x"800c873d",
  3147 => x"0d048052",
  3148 => x"7551fdb0",
  3149 => x"3f80f9c0",
  3150 => x"0b880508",
  3151 => x"80087131",
  3152 => x"56538f75",
  3153 => x"25ffa438",
  3154 => x"800880f9",
  3155 => x"b4083180",
  3156 => x"f9840c74",
  3157 => x"81078414",
  3158 => x"0c7551fd",
  3159 => x"863f8053",
  3160 => x"ff9039f6",
  3161 => x"3d0d7c7e",
  3162 => x"545b7280",
  3163 => x"2e828338",
  3164 => x"7a51fcee",
  3165 => x"3ff81384",
  3166 => x"110870fe",
  3167 => x"06701384",
  3168 => x"1108fc06",
  3169 => x"5d585954",
  3170 => x"5880f9c8",
  3171 => x"08752e82",
  3172 => x"de387884",
  3173 => x"160c8073",
  3174 => x"8106545a",
  3175 => x"727a2e81",
  3176 => x"d5387815",
  3177 => x"84110881",
  3178 => x"06515372",
  3179 => x"a0387817",
  3180 => x"577981e6",
  3181 => x"38881508",
  3182 => x"537280f9",
  3183 => x"c82e82f9",
  3184 => x"388c1508",
  3185 => x"708c150c",
  3186 => x"7388120c",
  3187 => x"56768107",
  3188 => x"84190c76",
  3189 => x"1877710c",
  3190 => x"53798191",
  3191 => x"3883ff77",
  3192 => x"2781c838",
  3193 => x"76892a77",
  3194 => x"832a5653",
  3195 => x"72802ebf",
  3196 => x"3876862a",
  3197 => x"b8055584",
  3198 => x"7327b438",
  3199 => x"80db1355",
  3200 => x"947327ab",
  3201 => x"38768c2a",
  3202 => x"80ee0555",
  3203 => x"80d47327",
  3204 => x"9e38768f",
  3205 => x"2a80f705",
  3206 => x"5582d473",
  3207 => x"27913876",
  3208 => x"922a80fc",
  3209 => x"05558ad4",
  3210 => x"73278438",
  3211 => x"80fe5574",
  3212 => x"10101080",
  3213 => x"f9c00588",
  3214 => x"11085556",
  3215 => x"73762e82",
  3216 => x"b3388414",
  3217 => x"08fc0653",
  3218 => x"7673278d",
  3219 => x"38881408",
  3220 => x"5473762e",
  3221 => x"098106ea",
  3222 => x"388c1408",
  3223 => x"708c1a0c",
  3224 => x"74881a0c",
  3225 => x"7888120c",
  3226 => x"56778c15",
  3227 => x"0c7a51fa",
  3228 => x"f23f8c3d",
  3229 => x"0d047708",
  3230 => x"78713159",
  3231 => x"77058819",
  3232 => x"08545772",
  3233 => x"80f9c82e",
  3234 => x"80e0388c",
  3235 => x"1808708c",
  3236 => x"150c7388",
  3237 => x"120c56fe",
  3238 => x"89398815",
  3239 => x"088c1608",
  3240 => x"708c130c",
  3241 => x"5788170c",
  3242 => x"fea33976",
  3243 => x"832a7054",
  3244 => x"55807524",
  3245 => x"81983872",
  3246 => x"822c8171",
  3247 => x"2b80f9c4",
  3248 => x"080780f9",
  3249 => x"c00b8405",
  3250 => x"0c537410",
  3251 => x"101080f9",
  3252 => x"c0058811",
  3253 => x"08555675",
  3254 => x"8c190c73",
  3255 => x"88190c77",
  3256 => x"88170c77",
  3257 => x"8c150cff",
  3258 => x"8439815a",
  3259 => x"fdb43978",
  3260 => x"17738106",
  3261 => x"54577298",
  3262 => x"38770878",
  3263 => x"71315977",
  3264 => x"058c1908",
  3265 => x"881a0871",
  3266 => x"8c120c88",
  3267 => x"120c5757",
  3268 => x"76810784",
  3269 => x"190c7780",
  3270 => x"f9c00b88",
  3271 => x"050c80f9",
  3272 => x"bc087726",
  3273 => x"fec73880",
  3274 => x"f9b80852",
  3275 => x"7a51fafd",
  3276 => x"3f7a51f9",
  3277 => x"ae3ffeba",
  3278 => x"3981788c",
  3279 => x"150c7888",
  3280 => x"150c738c",
  3281 => x"1a0c7388",
  3282 => x"1a0c5afd",
  3283 => x"80398315",
  3284 => x"70822c81",
  3285 => x"712b80f9",
  3286 => x"c4080780",
  3287 => x"f9c00b84",
  3288 => x"050c5153",
  3289 => x"74101010",
  3290 => x"80f9c005",
  3291 => x"88110855",
  3292 => x"56fee439",
  3293 => x"74538075",
  3294 => x"24a73872",
  3295 => x"822c8171",
  3296 => x"2b80f9c4",
  3297 => x"080780f9",
  3298 => x"c00b8405",
  3299 => x"0c53758c",
  3300 => x"190c7388",
  3301 => x"190c7788",
  3302 => x"170c778c",
  3303 => x"150cfdcd",
  3304 => x"39831570",
  3305 => x"822c8171",
  3306 => x"2b80f9c4",
  3307 => x"080780f9",
  3308 => x"c00b8405",
  3309 => x"0c5153d6",
  3310 => x"39fe3d0d",
  3311 => x"8188f008",
  3312 => x"51708a38",
  3313 => x"81d99c70",
  3314 => x"8188f00c",
  3315 => x"51707512",
  3316 => x"5252ff53",
  3317 => x"7087fb80",
  3318 => x"80268838",
  3319 => x"708188f0",
  3320 => x"0c715372",
  3321 => x"800c843d",
  3322 => x"0d04fd3d",
  3323 => x"0d800b80",
  3324 => x"f8ec0854",
  3325 => x"5472812e",
  3326 => x"9e387381",
  3327 => x"88f40cff",
  3328 => x"a0ff3fff",
  3329 => x"9ffa3f81",
  3330 => x"88c85281",
  3331 => x"51ffa9ae",
  3332 => x"3f800851",
  3333 => x"80e13f72",
  3334 => x"8188f40c",
  3335 => x"ffa0e23f",
  3336 => x"ff9fdd3f",
  3337 => x"8188c852",
  3338 => x"8151ffa9",
  3339 => x"913f8008",
  3340 => x"5180c43f",
  3341 => x"00ff3900",
  3342 => x"ff39f43d",
  3343 => x"0d7e8188",
  3344 => x"e8087008",
  3345 => x"7081ff06",
  3346 => x"923df805",
  3347 => x"55515a57",
  3348 => x"59ffa19a",
  3349 => x"3f805477",
  3350 => x"557b7d58",
  3351 => x"5276538e",
  3352 => x"3df00551",
  3353 => x"c0c03f79",
  3354 => x"7b58790c",
  3355 => x"76841a0c",
  3356 => x"78800c8e",
  3357 => x"3d0d04f7",
  3358 => x"3d0d7b81",
  3359 => x"81c80882",
  3360 => x"c811085a",
  3361 => x"545a7780",
  3362 => x"2e80da38",
  3363 => x"81881884",
  3364 => x"1908ff05",
  3365 => x"81712b59",
  3366 => x"55598074",
  3367 => x"2480ea38",
  3368 => x"807424b5",
  3369 => x"3873822b",
  3370 => x"78118805",
  3371 => x"56568180",
  3372 => x"19087706",
  3373 => x"5372802e",
  3374 => x"b6387816",
  3375 => x"70085353",
  3376 => x"79517408",
  3377 => x"53722dff",
  3378 => x"14fc17fc",
  3379 => x"1779812c",
  3380 => x"5a575754",
  3381 => x"738025d6",
  3382 => x"38770858",
  3383 => x"77ffad38",
  3384 => x"8181c808",
  3385 => x"53bc1308",
  3386 => x"a5387951",
  3387 => x"fec63f74",
  3388 => x"0853722d",
  3389 => x"ff14fc17",
  3390 => x"fc177981",
  3391 => x"2c5a5757",
  3392 => x"54738025",
  3393 => x"ffa838d1",
  3394 => x"398057ff",
  3395 => x"93397251",
  3396 => x"bc130853",
  3397 => x"722d7951",
  3398 => x"fe9a3fff",
  3399 => x"3d0d8188",
  3400 => x"d00bfc05",
  3401 => x"70085252",
  3402 => x"70ff2e91",
  3403 => x"38702dfc",
  3404 => x"12700852",
  3405 => x"5270ff2e",
  3406 => x"098106f1",
  3407 => x"38833d0d",
  3408 => x"0404ffa0",
  3409 => x"873f0400",
  3410 => x"00000040",
  3411 => x"30313233",
  3412 => x"34353637",
  3413 => x"38390000",
  3414 => x"44485259",
  3415 => x"53544f4e",
  3416 => x"45205052",
  3417 => x"4f475241",
  3418 => x"4d2c2053",
  3419 => x"4f4d4520",
  3420 => x"53545249",
  3421 => x"4e470000",
  3422 => x"44485259",
  3423 => x"53544f4e",
  3424 => x"45205052",
  3425 => x"4f475241",
  3426 => x"4d2c2031",
  3427 => x"27535420",
  3428 => x"53545249",
  3429 => x"4e470000",
  3430 => x"44687279",
  3431 => x"73746f6e",
  3432 => x"65204265",
  3433 => x"6e63686d",
  3434 => x"61726b2c",
  3435 => x"20566572",
  3436 => x"73696f6e",
  3437 => x"20322e31",
  3438 => x"20284c61",
  3439 => x"6e677561",
  3440 => x"67653a20",
  3441 => x"43290a00",
  3442 => x"50726f67",
  3443 => x"72616d20",
  3444 => x"636f6d70",
  3445 => x"696c6564",
  3446 => x"20776974",
  3447 => x"68202772",
  3448 => x"65676973",
  3449 => x"74657227",
  3450 => x"20617474",
  3451 => x"72696275",
  3452 => x"74650a00",
  3453 => x"45786563",
  3454 => x"7574696f",
  3455 => x"6e207374",
  3456 => x"61727473",
  3457 => x"2c202564",
  3458 => x"2072756e",
  3459 => x"73207468",
  3460 => x"726f7567",
  3461 => x"68204468",
  3462 => x"72797374",
  3463 => x"6f6e650a",
  3464 => x"00000000",
  3465 => x"44485259",
  3466 => x"53544f4e",
  3467 => x"45205052",
  3468 => x"4f475241",
  3469 => x"4d2c2032",
  3470 => x"274e4420",
  3471 => x"53545249",
  3472 => x"4e470000",
  3473 => x"45786563",
  3474 => x"7574696f",
  3475 => x"6e20656e",
  3476 => x"64730a00",
  3477 => x"46696e61",
  3478 => x"6c207661",
  3479 => x"6c756573",
  3480 => x"206f6620",
  3481 => x"74686520",
  3482 => x"76617269",
  3483 => x"61626c65",
  3484 => x"73207573",
  3485 => x"65642069",
  3486 => x"6e207468",
  3487 => x"65206265",
  3488 => x"6e63686d",
  3489 => x"61726b3a",
  3490 => x"0a000000",
  3491 => x"496e745f",
  3492 => x"476c6f62",
  3493 => x"3a202020",
  3494 => x"20202020",
  3495 => x"20202020",
  3496 => x"2025640a",
  3497 => x"00000000",
  3498 => x"20202020",
  3499 => x"20202020",
  3500 => x"73686f75",
  3501 => x"6c642062",
  3502 => x"653a2020",
  3503 => x"2025640a",
  3504 => x"00000000",
  3505 => x"426f6f6c",
  3506 => x"5f476c6f",
  3507 => x"623a2020",
  3508 => x"20202020",
  3509 => x"20202020",
  3510 => x"2025640a",
  3511 => x"00000000",
  3512 => x"43685f31",
  3513 => x"5f476c6f",
  3514 => x"623a2020",
  3515 => x"20202020",
  3516 => x"20202020",
  3517 => x"2025630a",
  3518 => x"00000000",
  3519 => x"20202020",
  3520 => x"20202020",
  3521 => x"73686f75",
  3522 => x"6c642062",
  3523 => x"653a2020",
  3524 => x"2025630a",
  3525 => x"00000000",
  3526 => x"43685f32",
  3527 => x"5f476c6f",
  3528 => x"623a2020",
  3529 => x"20202020",
  3530 => x"20202020",
  3531 => x"2025630a",
  3532 => x"00000000",
  3533 => x"4172725f",
  3534 => x"315f476c",
  3535 => x"6f625b38",
  3536 => x"5d3a2020",
  3537 => x"20202020",
  3538 => x"2025640a",
  3539 => x"00000000",
  3540 => x"4172725f",
  3541 => x"325f476c",
  3542 => x"6f625b38",
  3543 => x"5d5b375d",
  3544 => x"3a202020",
  3545 => x"2025640a",
  3546 => x"00000000",
  3547 => x"20202020",
  3548 => x"20202020",
  3549 => x"73686f75",
  3550 => x"6c642062",
  3551 => x"653a2020",
  3552 => x"204e756d",
  3553 => x"6265725f",
  3554 => x"4f665f52",
  3555 => x"756e7320",
  3556 => x"2b203130",
  3557 => x"0a000000",
  3558 => x"5074725f",
  3559 => x"476c6f62",
  3560 => x"2d3e0a00",
  3561 => x"20205074",
  3562 => x"725f436f",
  3563 => x"6d703a20",
  3564 => x"20202020",
  3565 => x"20202020",
  3566 => x"2025640a",
  3567 => x"00000000",
  3568 => x"20202020",
  3569 => x"20202020",
  3570 => x"73686f75",
  3571 => x"6c642062",
  3572 => x"653a2020",
  3573 => x"2028696d",
  3574 => x"706c656d",
  3575 => x"656e7461",
  3576 => x"74696f6e",
  3577 => x"2d646570",
  3578 => x"656e6465",
  3579 => x"6e74290a",
  3580 => x"00000000",
  3581 => x"20204469",
  3582 => x"7363723a",
  3583 => x"20202020",
  3584 => x"20202020",
  3585 => x"20202020",
  3586 => x"2025640a",
  3587 => x"00000000",
  3588 => x"2020456e",
  3589 => x"756d5f43",
  3590 => x"6f6d703a",
  3591 => x"20202020",
  3592 => x"20202020",
  3593 => x"2025640a",
  3594 => x"00000000",
  3595 => x"2020496e",
  3596 => x"745f436f",
  3597 => x"6d703a20",
  3598 => x"20202020",
  3599 => x"20202020",
  3600 => x"2025640a",
  3601 => x"00000000",
  3602 => x"20205374",
  3603 => x"725f436f",
  3604 => x"6d703a20",
  3605 => x"20202020",
  3606 => x"20202020",
  3607 => x"2025730a",
  3608 => x"00000000",
  3609 => x"20202020",
  3610 => x"20202020",
  3611 => x"73686f75",
  3612 => x"6c642062",
  3613 => x"653a2020",
  3614 => x"20444852",
  3615 => x"5953544f",
  3616 => x"4e452050",
  3617 => x"524f4752",
  3618 => x"414d2c20",
  3619 => x"534f4d45",
  3620 => x"20535452",
  3621 => x"494e470a",
  3622 => x"00000000",
  3623 => x"4e657874",
  3624 => x"5f507472",
  3625 => x"5f476c6f",
  3626 => x"622d3e0a",
  3627 => x"00000000",
  3628 => x"20202020",
  3629 => x"20202020",
  3630 => x"73686f75",
  3631 => x"6c642062",
  3632 => x"653a2020",
  3633 => x"2028696d",
  3634 => x"706c656d",
  3635 => x"656e7461",
  3636 => x"74696f6e",
  3637 => x"2d646570",
  3638 => x"656e6465",
  3639 => x"6e74292c",
  3640 => x"2073616d",
  3641 => x"65206173",
  3642 => x"2061626f",
  3643 => x"76650a00",
  3644 => x"496e745f",
  3645 => x"315f4c6f",
  3646 => x"633a2020",
  3647 => x"20202020",
  3648 => x"20202020",
  3649 => x"2025640a",
  3650 => x"00000000",
  3651 => x"496e745f",
  3652 => x"325f4c6f",
  3653 => x"633a2020",
  3654 => x"20202020",
  3655 => x"20202020",
  3656 => x"2025640a",
  3657 => x"00000000",
  3658 => x"496e745f",
  3659 => x"335f4c6f",
  3660 => x"633a2020",
  3661 => x"20202020",
  3662 => x"20202020",
  3663 => x"2025640a",
  3664 => x"00000000",
  3665 => x"456e756d",
  3666 => x"5f4c6f63",
  3667 => x"3a202020",
  3668 => x"20202020",
  3669 => x"20202020",
  3670 => x"2025640a",
  3671 => x"00000000",
  3672 => x"5374725f",
  3673 => x"315f4c6f",
  3674 => x"633a2020",
  3675 => x"20202020",
  3676 => x"20202020",
  3677 => x"2025730a",
  3678 => x"00000000",
  3679 => x"20202020",
  3680 => x"20202020",
  3681 => x"73686f75",
  3682 => x"6c642062",
  3683 => x"653a2020",
  3684 => x"20444852",
  3685 => x"5953544f",
  3686 => x"4e452050",
  3687 => x"524f4752",
  3688 => x"414d2c20",
  3689 => x"31275354",
  3690 => x"20535452",
  3691 => x"494e470a",
  3692 => x"00000000",
  3693 => x"5374725f",
  3694 => x"325f4c6f",
  3695 => x"633a2020",
  3696 => x"20202020",
  3697 => x"20202020",
  3698 => x"2025730a",
  3699 => x"00000000",
  3700 => x"20202020",
  3701 => x"20202020",
  3702 => x"73686f75",
  3703 => x"6c642062",
  3704 => x"653a2020",
  3705 => x"20444852",
  3706 => x"5953544f",
  3707 => x"4e452050",
  3708 => x"524f4752",
  3709 => x"414d2c20",
  3710 => x"32274e44",
  3711 => x"20535452",
  3712 => x"494e470a",
  3713 => x"00000000",
  3714 => x"55736572",
  3715 => x"2074696d",
  3716 => x"653a2025",
  3717 => x"640a0000",
  3718 => x"4d696372",
  3719 => x"6f736563",
  3720 => x"6f6e6473",
  3721 => x"20666f72",
  3722 => x"206f6e65",
  3723 => x"2072756e",
  3724 => x"20746872",
  3725 => x"6f756768",
  3726 => x"20446872",
  3727 => x"7973746f",
  3728 => x"6e653a20",
  3729 => x"00000000",
  3730 => x"2564200a",
  3731 => x"00000000",
  3732 => x"44687279",
  3733 => x"73746f6e",
  3734 => x"65732070",
  3735 => x"65722053",
  3736 => x"65636f6e",
  3737 => x"643a2020",
  3738 => x"20202020",
  3739 => x"20202020",
  3740 => x"20202020",
  3741 => x"20202020",
  3742 => x"20202020",
  3743 => x"00000000",
  3744 => x"56415820",
  3745 => x"4d495053",
  3746 => x"20726174",
  3747 => x"696e6720",
  3748 => x"2a203130",
  3749 => x"3030203d",
  3750 => x"20256420",
  3751 => x"0a000000",
  3752 => x"50726f67",
  3753 => x"72616d20",
  3754 => x"636f6d70",
  3755 => x"696c6564",
  3756 => x"20776974",
  3757 => x"686f7574",
  3758 => x"20277265",
  3759 => x"67697374",
  3760 => x"65722720",
  3761 => x"61747472",
  3762 => x"69627574",
  3763 => x"650a0000",
  3764 => x"4d656173",
  3765 => x"75726564",
  3766 => x"2074696d",
  3767 => x"6520746f",
  3768 => x"6f20736d",
  3769 => x"616c6c20",
  3770 => x"746f206f",
  3771 => x"62746169",
  3772 => x"6e206d65",
  3773 => x"616e696e",
  3774 => x"6766756c",
  3775 => x"20726573",
  3776 => x"756c7473",
  3777 => x"0a000000",
  3778 => x"506c6561",
  3779 => x"73652069",
  3780 => x"6e637265",
  3781 => x"61736520",
  3782 => x"6e756d62",
  3783 => x"6572206f",
  3784 => x"66207275",
  3785 => x"6e730a00",
  3786 => x"44485259",
  3787 => x"53544f4e",
  3788 => x"45205052",
  3789 => x"4f475241",
  3790 => x"4d2c2033",
  3791 => x"27524420",
  3792 => x"53545249",
  3793 => x"4e470000",
  3794 => x"00010202",
  3795 => x"03030303",
  3796 => x"04040404",
  3797 => x"04040404",
  3798 => x"05050505",
  3799 => x"05050505",
  3800 => x"05050505",
  3801 => x"05050505",
  3802 => x"06060606",
  3803 => x"06060606",
  3804 => x"06060606",
  3805 => x"06060606",
  3806 => x"06060606",
  3807 => x"06060606",
  3808 => x"06060606",
  3809 => x"06060606",
  3810 => x"07070707",
  3811 => x"07070707",
  3812 => x"07070707",
  3813 => x"07070707",
  3814 => x"07070707",
  3815 => x"07070707",
  3816 => x"07070707",
  3817 => x"07070707",
  3818 => x"07070707",
  3819 => x"07070707",
  3820 => x"07070707",
  3821 => x"07070707",
  3822 => x"07070707",
  3823 => x"07070707",
  3824 => x"07070707",
  3825 => x"07070707",
  3826 => x"08080808",
  3827 => x"08080808",
  3828 => x"08080808",
  3829 => x"08080808",
  3830 => x"08080808",
  3831 => x"08080808",
  3832 => x"08080808",
  3833 => x"08080808",
  3834 => x"08080808",
  3835 => x"08080808",
  3836 => x"08080808",
  3837 => x"08080808",
  3838 => x"08080808",
  3839 => x"08080808",
  3840 => x"08080808",
  3841 => x"08080808",
  3842 => x"08080808",
  3843 => x"08080808",
  3844 => x"08080808",
  3845 => x"08080808",
  3846 => x"08080808",
  3847 => x"08080808",
  3848 => x"08080808",
  3849 => x"08080808",
  3850 => x"08080808",
  3851 => x"08080808",
  3852 => x"08080808",
  3853 => x"08080808",
  3854 => x"08080808",
  3855 => x"08080808",
  3856 => x"08080808",
  3857 => x"08080808",
  3858 => x"43000000",
  3859 => x"64756d6d",
  3860 => x"792e6578",
  3861 => x"65000000",
  3862 => x"00ffffff",
  3863 => x"ff00ffff",
  3864 => x"ffff00ff",
  3865 => x"ffffff00",
  3866 => x"00000000",
  3867 => x"00000000",
  3868 => x"00000000",
  3869 => x"00004458",
  3870 => x"0000000a",
  3871 => x"00000000",
  3872 => x"00000032",
  3873 => x"00000000",
  3874 => x"00000000",
  3875 => x"00000000",
  3876 => x"00000000",
  3877 => x"00000000",
  3878 => x"00000000",
  3879 => x"00000000",
  3880 => x"00000000",
  3881 => x"00000000",
  3882 => x"00000000",
  3883 => x"00000000",
  3884 => x"00000000",
  3885 => x"ffffffff",
  3886 => x"00000000",
  3887 => x"00020000",
  3888 => x"00000000",
  3889 => x"00000000",
  3890 => x"00003cc0",
  3891 => x"00003cc0",
  3892 => x"00003cc8",
  3893 => x"00003cc8",
  3894 => x"00003cd0",
  3895 => x"00003cd0",
  3896 => x"00003cd8",
  3897 => x"00003cd8",
  3898 => x"00003ce0",
  3899 => x"00003ce0",
  3900 => x"00003ce8",
  3901 => x"00003ce8",
  3902 => x"00003cf0",
  3903 => x"00003cf0",
  3904 => x"00003cf8",
  3905 => x"00003cf8",
  3906 => x"00003d00",
  3907 => x"00003d00",
  3908 => x"00003d08",
  3909 => x"00003d08",
  3910 => x"00003d10",
  3911 => x"00003d10",
  3912 => x"00003d18",
  3913 => x"00003d18",
  3914 => x"00003d20",
  3915 => x"00003d20",
  3916 => x"00003d28",
  3917 => x"00003d28",
  3918 => x"00003d30",
  3919 => x"00003d30",
  3920 => x"00003d38",
  3921 => x"00003d38",
  3922 => x"00003d40",
  3923 => x"00003d40",
  3924 => x"00003d48",
  3925 => x"00003d48",
  3926 => x"00003d50",
  3927 => x"00003d50",
  3928 => x"00003d58",
  3929 => x"00003d58",
  3930 => x"00003d60",
  3931 => x"00003d60",
  3932 => x"00003d68",
  3933 => x"00003d68",
  3934 => x"00003d70",
  3935 => x"00003d70",
  3936 => x"00003d78",
  3937 => x"00003d78",
  3938 => x"00003d80",
  3939 => x"00003d80",
  3940 => x"00003d88",
  3941 => x"00003d88",
  3942 => x"00003d90",
  3943 => x"00003d90",
  3944 => x"00003d98",
  3945 => x"00003d98",
  3946 => x"00003da0",
  3947 => x"00003da0",
  3948 => x"00003da8",
  3949 => x"00003da8",
  3950 => x"00003db0",
  3951 => x"00003db0",
  3952 => x"00003db8",
  3953 => x"00003db8",
  3954 => x"00003dc0",
  3955 => x"00003dc0",
  3956 => x"00003dc8",
  3957 => x"00003dc8",
  3958 => x"00003dd0",
  3959 => x"00003dd0",
  3960 => x"00003dd8",
  3961 => x"00003dd8",
  3962 => x"00003de0",
  3963 => x"00003de0",
  3964 => x"00003de8",
  3965 => x"00003de8",
  3966 => x"00003df0",
  3967 => x"00003df0",
  3968 => x"00003df8",
  3969 => x"00003df8",
  3970 => x"00003e00",
  3971 => x"00003e00",
  3972 => x"00003e08",
  3973 => x"00003e08",
  3974 => x"00003e10",
  3975 => x"00003e10",
  3976 => x"00003e18",
  3977 => x"00003e18",
  3978 => x"00003e20",
  3979 => x"00003e20",
  3980 => x"00003e28",
  3981 => x"00003e28",
  3982 => x"00003e30",
  3983 => x"00003e30",
  3984 => x"00003e38",
  3985 => x"00003e38",
  3986 => x"00003e40",
  3987 => x"00003e40",
  3988 => x"00003e48",
  3989 => x"00003e48",
  3990 => x"00003e50",
  3991 => x"00003e50",
  3992 => x"00003e58",
  3993 => x"00003e58",
  3994 => x"00003e60",
  3995 => x"00003e60",
  3996 => x"00003e68",
  3997 => x"00003e68",
  3998 => x"00003e70",
  3999 => x"00003e70",
  4000 => x"00003e78",
  4001 => x"00003e78",
  4002 => x"00003e80",
  4003 => x"00003e80",
  4004 => x"00003e88",
  4005 => x"00003e88",
  4006 => x"00003e90",
  4007 => x"00003e90",
  4008 => x"00003e98",
  4009 => x"00003e98",
  4010 => x"00003ea0",
  4011 => x"00003ea0",
  4012 => x"00003ea8",
  4013 => x"00003ea8",
  4014 => x"00003eb0",
  4015 => x"00003eb0",
  4016 => x"00003eb8",
  4017 => x"00003eb8",
  4018 => x"00003ec0",
  4019 => x"00003ec0",
  4020 => x"00003ec8",
  4021 => x"00003ec8",
  4022 => x"00003ed0",
  4023 => x"00003ed0",
  4024 => x"00003ed8",
  4025 => x"00003ed8",
  4026 => x"00003ee0",
  4027 => x"00003ee0",
  4028 => x"00003ee8",
  4029 => x"00003ee8",
  4030 => x"00003ef0",
  4031 => x"00003ef0",
  4032 => x"00003ef8",
  4033 => x"00003ef8",
  4034 => x"00003f00",
  4035 => x"00003f00",
  4036 => x"00003f08",
  4037 => x"00003f08",
  4038 => x"00003f10",
  4039 => x"00003f10",
  4040 => x"00003f18",
  4041 => x"00003f18",
  4042 => x"00003f20",
  4043 => x"00003f20",
  4044 => x"00003f28",
  4045 => x"00003f28",
  4046 => x"00003f30",
  4047 => x"00003f30",
  4048 => x"00003f38",
  4049 => x"00003f38",
  4050 => x"00003f40",
  4051 => x"00003f40",
  4052 => x"00003f48",
  4053 => x"00003f48",
  4054 => x"00003f50",
  4055 => x"00003f50",
  4056 => x"00003f58",
  4057 => x"00003f58",
  4058 => x"00003f60",
  4059 => x"00003f60",
  4060 => x"00003f68",
  4061 => x"00003f68",
  4062 => x"00003f70",
  4063 => x"00003f70",
  4064 => x"00003f78",
  4065 => x"00003f78",
  4066 => x"00003f80",
  4067 => x"00003f80",
  4068 => x"00003f88",
  4069 => x"00003f88",
  4070 => x"00003f90",
  4071 => x"00003f90",
  4072 => x"00003f98",
  4073 => x"00003f98",
  4074 => x"00003fa0",
  4075 => x"00003fa0",
  4076 => x"00003fa8",
  4077 => x"00003fa8",
  4078 => x"00003fb0",
  4079 => x"00003fb0",
  4080 => x"00003fb8",
  4081 => x"00003fb8",
  4082 => x"00003fc0",
  4083 => x"00003fc0",
  4084 => x"00003fc8",
  4085 => x"00003fc8",
  4086 => x"00003fd0",
  4087 => x"00003fd0",
  4088 => x"00003fd8",
  4089 => x"00003fd8",
  4090 => x"00003fe0",
  4091 => x"00003fe0",
  4092 => x"00003fe8",
  4093 => x"00003fe8",
  4094 => x"00003ff0",
  4095 => x"00003ff0",
  4096 => x"00003ff8",
  4097 => x"00003ff8",
  4098 => x"00004000",
  4099 => x"00004000",
  4100 => x"00004008",
  4101 => x"00004008",
  4102 => x"00004010",
  4103 => x"00004010",
  4104 => x"00004018",
  4105 => x"00004018",
  4106 => x"00004020",
  4107 => x"00004020",
  4108 => x"00004028",
  4109 => x"00004028",
  4110 => x"00004030",
  4111 => x"00004030",
  4112 => x"00004038",
  4113 => x"00004038",
  4114 => x"00004040",
  4115 => x"00004040",
  4116 => x"00004048",
  4117 => x"00004048",
  4118 => x"00004050",
  4119 => x"00004050",
  4120 => x"00004058",
  4121 => x"00004058",
  4122 => x"00004060",
  4123 => x"00004060",
  4124 => x"00004068",
  4125 => x"00004068",
  4126 => x"00004070",
  4127 => x"00004070",
  4128 => x"00004078",
  4129 => x"00004078",
  4130 => x"00004080",
  4131 => x"00004080",
  4132 => x"00004088",
  4133 => x"00004088",
  4134 => x"00004090",
  4135 => x"00004090",
  4136 => x"00004098",
  4137 => x"00004098",
  4138 => x"000040a0",
  4139 => x"000040a0",
  4140 => x"000040a8",
  4141 => x"000040a8",
  4142 => x"000040b0",
  4143 => x"000040b0",
  4144 => x"000040b8",
  4145 => x"000040b8",
  4146 => x"000040cc",
  4147 => x"00000000",
  4148 => x"00004334",
  4149 => x"00004390",
  4150 => x"000043ec",
  4151 => x"00000000",
  4152 => x"00000000",
  4153 => x"00000000",
  4154 => x"00000000",
  4155 => x"00000000",
  4156 => x"00000000",
  4157 => x"00000000",
  4158 => x"00000000",
  4159 => x"00000000",
  4160 => x"00003c48",
  4161 => x"00000000",
  4162 => x"00000000",
  4163 => x"00000000",
  4164 => x"00000000",
  4165 => x"00000000",
  4166 => x"00000000",
  4167 => x"00000000",
  4168 => x"00000000",
  4169 => x"00000000",
  4170 => x"00000000",
  4171 => x"00000000",
  4172 => x"00000000",
  4173 => x"00000000",
  4174 => x"00000000",
  4175 => x"00000000",
  4176 => x"00000000",
  4177 => x"00000000",
  4178 => x"00000000",
  4179 => x"00000000",
  4180 => x"00000000",
  4181 => x"00000000",
  4182 => x"00000000",
  4183 => x"00000000",
  4184 => x"00000000",
  4185 => x"00000000",
  4186 => x"00000000",
  4187 => x"00000000",
  4188 => x"00000000",
  4189 => x"00000001",
  4190 => x"330eabcd",
  4191 => x"1234e66d",
  4192 => x"deec0005",
  4193 => x"000b0000",
  4194 => x"00000000",
  4195 => x"00000000",
  4196 => x"00000000",
  4197 => x"00000000",
  4198 => x"00000000",
  4199 => x"00000000",
  4200 => x"00000000",
  4201 => x"00000000",
  4202 => x"00000000",
  4203 => x"00000000",
  4204 => x"00000000",
  4205 => x"00000000",
  4206 => x"00000000",
  4207 => x"00000000",
  4208 => x"00000000",
  4209 => x"00000000",
  4210 => x"00000000",
  4211 => x"00000000",
  4212 => x"00000000",
  4213 => x"00000000",
  4214 => x"00000000",
  4215 => x"00000000",
  4216 => x"00000000",
  4217 => x"00000000",
  4218 => x"00000000",
  4219 => x"00000000",
  4220 => x"00000000",
  4221 => x"00000000",
  4222 => x"00000000",
  4223 => x"00000000",
  4224 => x"00000000",
  4225 => x"00000000",
  4226 => x"00000000",
  4227 => x"00000000",
  4228 => x"00000000",
  4229 => x"00000000",
  4230 => x"00000000",
  4231 => x"00000000",
  4232 => x"00000000",
  4233 => x"00000000",
  4234 => x"00000000",
  4235 => x"00000000",
  4236 => x"00000000",
  4237 => x"00000000",
  4238 => x"00000000",
  4239 => x"00000000",
  4240 => x"00000000",
  4241 => x"00000000",
  4242 => x"00000000",
  4243 => x"00000000",
  4244 => x"00000000",
  4245 => x"00000000",
  4246 => x"00000000",
  4247 => x"00000000",
  4248 => x"00000000",
  4249 => x"00000000",
  4250 => x"00000000",
  4251 => x"00000000",
  4252 => x"00000000",
  4253 => x"00000000",
  4254 => x"00000000",
  4255 => x"00000000",
  4256 => x"00000000",
  4257 => x"00000000",
  4258 => x"00000000",
  4259 => x"00000000",
  4260 => x"00000000",
  4261 => x"00000000",
  4262 => x"00000000",
  4263 => x"00000000",
  4264 => x"00000000",
  4265 => x"00000000",
  4266 => x"00000000",
  4267 => x"00000000",
  4268 => x"00000000",
  4269 => x"00000000",
  4270 => x"00000000",
  4271 => x"00000000",
  4272 => x"00000000",
  4273 => x"00000000",
  4274 => x"00000000",
  4275 => x"00000000",
  4276 => x"00000000",
  4277 => x"00000000",
  4278 => x"00000000",
  4279 => x"00000000",
  4280 => x"00000000",
  4281 => x"00000000",
  4282 => x"00000000",
  4283 => x"00000000",
  4284 => x"00000000",
  4285 => x"00000000",
  4286 => x"00000000",
  4287 => x"00000000",
  4288 => x"00000000",
  4289 => x"00000000",
  4290 => x"00000000",
  4291 => x"00000000",
  4292 => x"00000000",
  4293 => x"00000000",
  4294 => x"00000000",
  4295 => x"00000000",
  4296 => x"00000000",
  4297 => x"00000000",
  4298 => x"00000000",
  4299 => x"00000000",
  4300 => x"00000000",
  4301 => x"00000000",
  4302 => x"00000000",
  4303 => x"00000000",
  4304 => x"00000000",
  4305 => x"00000000",
  4306 => x"00000000",
  4307 => x"00000000",
  4308 => x"00000000",
  4309 => x"00000000",
  4310 => x"00000000",
  4311 => x"00000000",
  4312 => x"00000000",
  4313 => x"00000000",
  4314 => x"00000000",
  4315 => x"00000000",
  4316 => x"00000000",
  4317 => x"00000000",
  4318 => x"00000000",
  4319 => x"00000000",
  4320 => x"00000000",
  4321 => x"00000000",
  4322 => x"00000000",
  4323 => x"00000000",
  4324 => x"00000000",
  4325 => x"00000000",
  4326 => x"00000000",
  4327 => x"00000000",
  4328 => x"00000000",
  4329 => x"00000000",
  4330 => x"00000000",
  4331 => x"00000000",
  4332 => x"00000000",
  4333 => x"00000000",
  4334 => x"00000000",
  4335 => x"00000000",
  4336 => x"00000000",
  4337 => x"00000000",
  4338 => x"00000000",
  4339 => x"00000000",
  4340 => x"00000000",
  4341 => x"00000000",
  4342 => x"00000000",
  4343 => x"00000000",
  4344 => x"00000000",
  4345 => x"00000000",
  4346 => x"00000000",
  4347 => x"00000000",
  4348 => x"00000000",
  4349 => x"00000000",
  4350 => x"00000000",
  4351 => x"00000000",
  4352 => x"00000000",
  4353 => x"00000000",
  4354 => x"00000000",
  4355 => x"00000000",
  4356 => x"00000000",
  4357 => x"00000000",
  4358 => x"00000000",
  4359 => x"00000000",
  4360 => x"00000000",
  4361 => x"00000000",
  4362 => x"00000000",
  4363 => x"00000000",
  4364 => x"00000000",
  4365 => x"00000000",
  4366 => x"00000000",
  4367 => x"00000000",
  4368 => x"00000000",
  4369 => x"00000000",
  4370 => x"00003c4c",
  4371 => x"ffffffff",
  4372 => x"00000000",
  4373 => x"ffffffff",
  4374 => x"00000000",
  4375 => x"00000000",

others => x"00000000"
);
begin
   busy_o <= re_i; -- we're done on the cycle after we serve the read request

   do_ram:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if we_i='1' then
            ram(to_integer(addr_i)) <= write_i;
         end if;
         addr_r <= addr_i;
      end if;
   end process do_ram;
   read_o <= ram(to_integer(addr_r));
end architecture Xilinx; -- Entity: SinglePortRAM

