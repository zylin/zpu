-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80e3e40c",
     3 => x"3a0b0b80",
     4 => x"dd980400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80dde12d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80e3",
   162 => x"d0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80c0",
   171 => x"ff2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80c2",
   179 => x"b12d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80e3e00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"d7823f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80e3e008",
   281 => x"802ea438",
   282 => x"80e3e408",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80f3",
   286 => x"e40c82a0",
   287 => x"800b80f3",
   288 => x"e80c8290",
   289 => x"800b80f3",
   290 => x"ec0c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"f3e40cf8",
   294 => x"80808280",
   295 => x"0b80f3e8",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"f3ec0c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80f3e40c",
   302 => x"80c0a880",
   303 => x"940b80f3",
   304 => x"e80c0b0b",
   305 => x"80dfb40b",
   306 => x"80f3ec0c",
   307 => x"04ff3d0d",
   308 => x"80f3f033",
   309 => x"5170a738",
   310 => x"80e3ec08",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"e3ec0c70",
   315 => x"2d80e3ec",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80f3",
   319 => x"f034833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80f3e008",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"f3e0510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404fd3d",
   333 => x"0d80e3fc",
   334 => x"0876b0ea",
   335 => x"2994120c",
   336 => x"54850b98",
   337 => x"150c9814",
   338 => x"08708106",
   339 => x"515372f6",
   340 => x"38853d0d",
   341 => x"04ff3d0d",
   342 => x"80e3fc08",
   343 => x"74101075",
   344 => x"10059412",
   345 => x"0c52850b",
   346 => x"98130c98",
   347 => x"12087081",
   348 => x"06515170",
   349 => x"f638833d",
   350 => x"0d04803d",
   351 => x"0d725180",
   352 => x"71278738",
   353 => x"ff115170",
   354 => x"fb38823d",
   355 => x"0d04803d",
   356 => x"0d80e3fc",
   357 => x"0851870b",
   358 => x"84120c82",
   359 => x"3d0d0480",
   360 => x"3d0d80e4",
   361 => x"800851b6",
   362 => x"0b8c120c",
   363 => x"830b8812",
   364 => x"0c823d0d",
   365 => x"04ff3d0d",
   366 => x"80e48008",
   367 => x"52841208",
   368 => x"70810651",
   369 => x"5170802e",
   370 => x"f4387108",
   371 => x"7081ff06",
   372 => x"800c5183",
   373 => x"3d0d04fe",
   374 => x"3d0d0293",
   375 => x"053380e4",
   376 => x"80085353",
   377 => x"84120870",
   378 => x"822a7081",
   379 => x"06515151",
   380 => x"70802ef0",
   381 => x"3872720c",
   382 => x"843d0d04",
   383 => x"fe3d0d02",
   384 => x"93053353",
   385 => x"728a2e9e",
   386 => x"3880e480",
   387 => x"08528412",
   388 => x"0870822a",
   389 => x"70810651",
   390 => x"51517080",
   391 => x"2ef03872",
   392 => x"720c843d",
   393 => x"0d0480e4",
   394 => x"80085284",
   395 => x"12087082",
   396 => x"2a708106",
   397 => x"51515170",
   398 => x"802ef038",
   399 => x"8d720c84",
   400 => x"12087082",
   401 => x"2a708106",
   402 => x"51515170",
   403 => x"802effbe",
   404 => x"38cd39fd",
   405 => x"3d0d7570",
   406 => x"33525470",
   407 => x"802eaa38",
   408 => x"7080e480",
   409 => x"08535381",
   410 => x"1454728a",
   411 => x"2e9f3884",
   412 => x"12087082",
   413 => x"2a708106",
   414 => x"51515170",
   415 => x"802ef038",
   416 => x"72720c73",
   417 => x"335372df",
   418 => x"38853d0d",
   419 => x"04841208",
   420 => x"70822a70",
   421 => x"81065151",
   422 => x"5170802e",
   423 => x"f0388d72",
   424 => x"0c841208",
   425 => x"70822a70",
   426 => x"81065151",
   427 => x"5170802e",
   428 => x"ffbd38cc",
   429 => x"39f53d0d",
   430 => x"7e028405",
   431 => x"b705338c",
   432 => x"3d5b5557",
   433 => x"8b5380df",
   434 => x"b8527851",
   435 => x"b7ba3f82",
   436 => x"5673882e",
   437 => x"96388456",
   438 => x"73902e8f",
   439 => x"38885673",
   440 => x"a02e8838",
   441 => x"74567480",
   442 => x"2ea73802",
   443 => x"a5055876",
   444 => x"8f065473",
   445 => x"892680ce",
   446 => x"387518b0",
   447 => x"15555573",
   448 => x"75347684",
   449 => x"2aff1770",
   450 => x"81ff0658",
   451 => x"555775df",
   452 => x"38787933",
   453 => x"55577380",
   454 => x"2ea83873",
   455 => x"80e48008",
   456 => x"56568117",
   457 => x"57758a2e",
   458 => x"b9388415",
   459 => x"0870822a",
   460 => x"81065954",
   461 => x"77802ef2",
   462 => x"3875750c",
   463 => x"76335675",
   464 => x"e1388d3d",
   465 => x"0d047518",
   466 => x"b7155555",
   467 => x"73753476",
   468 => x"842aff17",
   469 => x"7081ff06",
   470 => x"58555775",
   471 => x"ff9138ff",
   472 => x"b0398415",
   473 => x"0870822a",
   474 => x"81065954",
   475 => x"77802ef2",
   476 => x"388d750c",
   477 => x"84150870",
   478 => x"822a8106",
   479 => x"59547780",
   480 => x"2effa738",
   481 => x"ffb339f8",
   482 => x"3d0d7a7c",
   483 => x"59538073",
   484 => x"56577673",
   485 => x"2480dc38",
   486 => x"7717548a",
   487 => x"527451b1",
   488 => x"b93f8008",
   489 => x"b0055372",
   490 => x"74348117",
   491 => x"578a5274",
   492 => x"51b1823f",
   493 => x"80085580",
   494 => x"08de3880",
   495 => x"08779f2a",
   496 => x"1870812c",
   497 => x"5b565680",
   498 => x"79259e38",
   499 => x"7717ff05",
   500 => x"55751870",
   501 => x"33555374",
   502 => x"33733473",
   503 => x"75348116",
   504 => x"ff165656",
   505 => x"787624e9",
   506 => x"38761856",
   507 => x"8076348a",
   508 => x"3d0d04ad",
   509 => x"78708105",
   510 => x"5a347230",
   511 => x"78185555",
   512 => x"8a527451",
   513 => x"b0d43f80",
   514 => x"08b00553",
   515 => x"72743481",
   516 => x"17578a52",
   517 => x"7451b09d",
   518 => x"3f800855",
   519 => x"8008fef8",
   520 => x"38ff9839",
   521 => x"803d0d80",
   522 => x"e3f80851",
   523 => x"800b8412",
   524 => x"0cfe800a",
   525 => x"0b88120c",
   526 => x"800b80f4",
   527 => x"8034800b",
   528 => x"80f3fc34",
   529 => x"823d0d04",
   530 => x"fd3d0d02",
   531 => x"97053352",
   532 => x"718a2eb0",
   533 => x"3880f480",
   534 => x"33701010",
   535 => x"1180f3fc",
   536 => x"33719029",
   537 => x"0570882b",
   538 => x"750780e3",
   539 => x"f8085271",
   540 => x"0c525253",
   541 => x"80f3fc33",
   542 => x"81055473",
   543 => x"80f3fc34",
   544 => x"853d0d04",
   545 => x"80f48033",
   546 => x"7081ff06",
   547 => x"525270a3",
   548 => x"26933881",
   549 => x"12537280",
   550 => x"f4803480",
   551 => x"0b80f3fc",
   552 => x"34853d0d",
   553 => x"04800b80",
   554 => x"f4803480",
   555 => x"0b80f3fc",
   556 => x"34ef39fb",
   557 => x"3d0d7770",
   558 => x"33525370",
   559 => x"802ebc38",
   560 => x"7080e3f8",
   561 => x"08555281",
   562 => x"1353718a",
   563 => x"2eb13880",
   564 => x"f4803370",
   565 => x"10101180",
   566 => x"f3fc3371",
   567 => x"90290570",
   568 => x"882b7507",
   569 => x"770c80f3",
   570 => x"fc338105",
   571 => x"59525255",
   572 => x"7580f3fc",
   573 => x"34723352",
   574 => x"71cd3887",
   575 => x"3d0d0480",
   576 => x"f4803370",
   577 => x"81ff0652",
   578 => x"5270a326",
   579 => x"98388112",
   580 => x"557480f4",
   581 => x"8034800b",
   582 => x"80f3fc34",
   583 => x"72335271",
   584 => x"ffa538d7",
   585 => x"39800b80",
   586 => x"f4803480",
   587 => x"0b80f3fc",
   588 => x"34ea39fb",
   589 => x"3d0d7770",
   590 => x"71337081",
   591 => x"ff065455",
   592 => x"55557080",
   593 => x"2eb13880",
   594 => x"e4800852",
   595 => x"7281ff06",
   596 => x"81155553",
   597 => x"728a2e80",
   598 => x"e8388412",
   599 => x"0870822a",
   600 => x"81065151",
   601 => x"70802ef2",
   602 => x"3872720c",
   603 => x"73337081",
   604 => x"ff065753",
   605 => x"75d63874",
   606 => x"75335253",
   607 => x"70802ebd",
   608 => x"387080e3",
   609 => x"f8085552",
   610 => x"81135371",
   611 => x"8a2e80d6",
   612 => x"3880f480",
   613 => x"33701010",
   614 => x"1180f3fc",
   615 => x"33719029",
   616 => x"0570882b",
   617 => x"7507770c",
   618 => x"80f3fc33",
   619 => x"81055951",
   620 => x"52557580",
   621 => x"f3fc3472",
   622 => x"335271cc",
   623 => x"38873d0d",
   624 => x"04841208",
   625 => x"70822a81",
   626 => x"06515675",
   627 => x"802ef238",
   628 => x"8d720c84",
   629 => x"12087082",
   630 => x"2a810651",
   631 => x"5170802e",
   632 => x"fef838ff",
   633 => x"843980f4",
   634 => x"80337081",
   635 => x"ff065652",
   636 => x"74a32699",
   637 => x"38811251",
   638 => x"7080f480",
   639 => x"34800b80",
   640 => x"f3fc3472",
   641 => x"335271fe",
   642 => x"ff38ffb1",
   643 => x"39800b80",
   644 => x"f4803480",
   645 => x"0b80f3fc",
   646 => x"34e939f5",
   647 => x"3d0d7e02",
   648 => x"8405b705",
   649 => x"338c3d5b",
   650 => x"55578b53",
   651 => x"80dfb852",
   652 => x"7851b0d4",
   653 => x"3f825673",
   654 => x"882e9638",
   655 => x"84567390",
   656 => x"2e8f3888",
   657 => x"5673a02e",
   658 => x"88387456",
   659 => x"74802ea7",
   660 => x"3802a505",
   661 => x"58768f06",
   662 => x"54738926",
   663 => x"81953875",
   664 => x"18b01555",
   665 => x"55737534",
   666 => x"76842aff",
   667 => x"177081ff",
   668 => x"06585557",
   669 => x"75df3878",
   670 => x"79335557",
   671 => x"73802ea9",
   672 => x"387380e4",
   673 => x"80085656",
   674 => x"81175775",
   675 => x"8a2e80ff",
   676 => x"38841508",
   677 => x"70822a81",
   678 => x"06515473",
   679 => x"802ef238",
   680 => x"75750c76",
   681 => x"335675e0",
   682 => x"38787933",
   683 => x"55567380",
   684 => x"2ebd3873",
   685 => x"80e3f808",
   686 => x"58558116",
   687 => x"56748a2e",
   688 => x"80f23880",
   689 => x"f4803370",
   690 => x"10101180",
   691 => x"f3fc3371",
   692 => x"90290570",
   693 => x"882b7807",
   694 => x"7a0c80f3",
   695 => x"fc338105",
   696 => x"52525558",
   697 => x"7380f3fc",
   698 => x"34753355",
   699 => x"74cc388d",
   700 => x"3d0d0475",
   701 => x"18b71555",
   702 => x"55737534",
   703 => x"76842aff",
   704 => x"177081ff",
   705 => x"06585557",
   706 => x"75feca38",
   707 => x"fee93984",
   708 => x"15087082",
   709 => x"2a810651",
   710 => x"5877802e",
   711 => x"f2388d75",
   712 => x"0c841508",
   713 => x"70822a81",
   714 => x"06515473",
   715 => x"802efee1",
   716 => x"38feed39",
   717 => x"80f48033",
   718 => x"7081ff06",
   719 => x"5a5578a3",
   720 => x"26993881",
   721 => x"15587780",
   722 => x"f4803480",
   723 => x"0b80f3fc",
   724 => x"34753355",
   725 => x"74fee338",
   726 => x"ff953980",
   727 => x"0b80f480",
   728 => x"34800b80",
   729 => x"f3fc34e9",
   730 => x"39803d0d",
   731 => x"80e3f408",
   732 => x"5181ff0b",
   733 => x"88120c82",
   734 => x"3d0d04f8",
   735 => x"3d0d7a59",
   736 => x"f881c08e",
   737 => x"8055a00b",
   738 => x"80e3f408",
   739 => x"80e3fc08",
   740 => x"5a585674",
   741 => x"84180c74",
   742 => x"9f2a7510",
   743 => x"07557880",
   744 => x"2e973875",
   745 => x"802ebb38",
   746 => x"ff167584",
   747 => x"190c759f",
   748 => x"2a761007",
   749 => x"565678eb",
   750 => x"387754af",
   751 => x"d7c20b94",
   752 => x"190c850b",
   753 => x"98190c98",
   754 => x"14087081",
   755 => x"06515372",
   756 => x"802ec038",
   757 => x"98140870",
   758 => x"81065153",
   759 => x"72e938ff",
   760 => x"b2398a3d",
   761 => x"0d04fd3d",
   762 => x"0d80e3f4",
   763 => x"085480d5",
   764 => x"0b84150c",
   765 => x"80e48008",
   766 => x"52841208",
   767 => x"81065170",
   768 => x"802ef638",
   769 => x"71087081",
   770 => x"ff06f611",
   771 => x"52545170",
   772 => x"ae268c38",
   773 => x"70101080",
   774 => x"e2840551",
   775 => x"70080484",
   776 => x"12087082",
   777 => x"2a708106",
   778 => x"51515170",
   779 => x"802ef038",
   780 => x"ab720c72",
   781 => x"8a2eaa38",
   782 => x"84120870",
   783 => x"822a7081",
   784 => x"06515151",
   785 => x"70802ef0",
   786 => x"3872720c",
   787 => x"84120870",
   788 => x"822a8106",
   789 => x"51537280",
   790 => x"2ef238ad",
   791 => x"720cff99",
   792 => x"39841208",
   793 => x"70822a70",
   794 => x"81065151",
   795 => x"5170802e",
   796 => x"f0388d72",
   797 => x"0c841208",
   798 => x"70822a70",
   799 => x"81065151",
   800 => x"5170802e",
   801 => x"ffb238c1",
   802 => x"3981ff0b",
   803 => x"84150cfe",
   804 => x"e83980ff",
   805 => x"0b84150c",
   806 => x"fedf39bf",
   807 => x"0b84150c",
   808 => x"fed7399f",
   809 => x"0b84150c",
   810 => x"fecf398f",
   811 => x"0b84150c",
   812 => x"fec73987",
   813 => x"0b84150c",
   814 => x"febf3983",
   815 => x"0b84150c",
   816 => x"feb73981",
   817 => x"0b84150c",
   818 => x"feaf3980",
   819 => x"0b84150c",
   820 => x"fea739ff",
   821 => x"3d0d80e3",
   822 => x"f4085271",
   823 => x"08708f06",
   824 => x"7071842b",
   825 => x"0784150c",
   826 => x"51517108",
   827 => x"708f0670",
   828 => x"71842b07",
   829 => x"84150c51",
   830 => x"51e139fc",
   831 => x"3d0d029a",
   832 => x"05220284",
   833 => x"059e0522",
   834 => x"028805a2",
   835 => x"052280e3",
   836 => x"f0085556",
   837 => x"54559012",
   838 => x"0870832a",
   839 => x"70810651",
   840 => x"515170f2",
   841 => x"3874902b",
   842 => x"738b2b07",
   843 => x"74862b07",
   844 => x"81079013",
   845 => x"0c863d0d",
   846 => x"04fd3d0d",
   847 => x"02960522",
   848 => x"0284059a",
   849 => x"052280e3",
   850 => x"f0085454",
   851 => x"54901208",
   852 => x"70832a70",
   853 => x"81065151",
   854 => x"5170f238",
   855 => x"738b2b73",
   856 => x"862b0782",
   857 => x"0790130c",
   858 => x"90120870",
   859 => x"832a8106",
   860 => x"555173f4",
   861 => x"38901208",
   862 => x"70902a80",
   863 => x"0c54853d",
   864 => x"0d04ff3d",
   865 => x"0d80e3f0",
   866 => x"0852ff0b",
   867 => x"84130cfc",
   868 => x"94800b88",
   869 => x"130c82d0",
   870 => x"affdfb0b",
   871 => x"8c130c80",
   872 => x"c0720c71",
   873 => x"0870862a",
   874 => x"70810651",
   875 => x"515170f3",
   876 => x"38901208",
   877 => x"70832a70",
   878 => x"81065151",
   879 => x"5170f238",
   880 => x"81fc8081",
   881 => x"0b90130c",
   882 => x"90120870",
   883 => x"832a7081",
   884 => x"06515151",
   885 => x"70f23880",
   886 => x"fdc0810b",
   887 => x"90130c83",
   888 => x"3d0d04f5",
   889 => x"3d0d80e3",
   890 => x"f00857ff",
   891 => x"0b84180c",
   892 => x"fc809b0b",
   893 => x"88180c82",
   894 => x"8ba1968a",
   895 => x"0b8c180c",
   896 => x"a4b40b94",
   897 => x"180c8186",
   898 => x"a10b9818",
   899 => x"0c80dfc4",
   900 => x"0b80dfc4",
   901 => x"33545672",
   902 => x"802eab38",
   903 => x"7280e480",
   904 => x"08555581",
   905 => x"1656748a",
   906 => x"2e85f638",
   907 => x"84140870",
   908 => x"822a7081",
   909 => x"06515153",
   910 => x"72802ef0",
   911 => x"3874740c",
   912 => x"75335574",
   913 => x"de3880df",
   914 => x"d80b80df",
   915 => x"d8335456",
   916 => x"72802eab",
   917 => x"3880e480",
   918 => x"08735654",
   919 => x"81165674",
   920 => x"8a2e85e6",
   921 => x"38841408",
   922 => x"70822a70",
   923 => x"81065151",
   924 => x"5372802e",
   925 => x"f0387474",
   926 => x"0c753355",
   927 => x"74de3876",
   928 => x"0852a051",
   929 => x"f0af3f80",
   930 => x"dfe80b80",
   931 => x"dfe83354",
   932 => x"5672802e",
   933 => x"a93880e4",
   934 => x"80087356",
   935 => x"54811656",
   936 => x"748a2e85",
   937 => x"ce388414",
   938 => x"0870822a",
   939 => x"81065153",
   940 => x"72802ef2",
   941 => x"3874740c",
   942 => x"75335574",
   943 => x"e03880e3",
   944 => x"f0088411",
   945 => x"085354a0",
   946 => x"51efea3f",
   947 => x"80dff80b",
   948 => x"80dff833",
   949 => x"54567280",
   950 => x"2ea93880",
   951 => x"e4800873",
   952 => x"56548116",
   953 => x"56748a2e",
   954 => x"85ae3884",
   955 => x"14087082",
   956 => x"2a810651",
   957 => x"5372802e",
   958 => x"f2387474",
   959 => x"0c753355",
   960 => x"74e03880",
   961 => x"e3f00888",
   962 => x"11085355",
   963 => x"a051efa5",
   964 => x"3f80e088",
   965 => x"0b80e088",
   966 => x"33545672",
   967 => x"802ea938",
   968 => x"80e48008",
   969 => x"73565481",
   970 => x"1656748a",
   971 => x"2e858e38",
   972 => x"84140870",
   973 => x"822a8106",
   974 => x"51537280",
   975 => x"2ef23874",
   976 => x"740c7533",
   977 => x"5574e038",
   978 => x"80e3f008",
   979 => x"8c110853",
   980 => x"56a051ee",
   981 => x"e03f80e0",
   982 => x"980b80e0",
   983 => x"98335456",
   984 => x"72802ea9",
   985 => x"3880e480",
   986 => x"08735654",
   987 => x"81165674",
   988 => x"8a2e84ee",
   989 => x"38841408",
   990 => x"70822a81",
   991 => x"06515372",
   992 => x"802ef238",
   993 => x"74740c75",
   994 => x"335574e0",
   995 => x"3880e3f0",
   996 => x"08901108",
   997 => x"5354a051",
   998 => x"ee9b3f80",
   999 => x"e0a80b80",
  1000 => x"e0a83354",
  1001 => x"5672802e",
  1002 => x"a93880e4",
  1003 => x"80087356",
  1004 => x"54811656",
  1005 => x"748a2e84",
  1006 => x"ce388414",
  1007 => x"0870822a",
  1008 => x"81065153",
  1009 => x"72802ef2",
  1010 => x"3874740c",
  1011 => x"75335574",
  1012 => x"e03880e3",
  1013 => x"f0089411",
  1014 => x"085355a0",
  1015 => x"51edd63f",
  1016 => x"80e0b80b",
  1017 => x"80e0b833",
  1018 => x"54567280",
  1019 => x"2ea93880",
  1020 => x"e4800873",
  1021 => x"56548116",
  1022 => x"56748a2e",
  1023 => x"84ae3884",
  1024 => x"14087082",
  1025 => x"2a810651",
  1026 => x"5372802e",
  1027 => x"f2387474",
  1028 => x"0c753355",
  1029 => x"74e03880",
  1030 => x"e3f00898",
  1031 => x"11085356",
  1032 => x"a051ed91",
  1033 => x"3f80e0c8",
  1034 => x"0b80e0c8",
  1035 => x"33545672",
  1036 => x"802ea938",
  1037 => x"80e48008",
  1038 => x"73565481",
  1039 => x"1656748a",
  1040 => x"2e848e38",
  1041 => x"84140870",
  1042 => x"822a8106",
  1043 => x"51537280",
  1044 => x"2ef23874",
  1045 => x"740c7533",
  1046 => x"5574e038",
  1047 => x"80e3f008",
  1048 => x"9c110853",
  1049 => x"54a051ec",
  1050 => x"cc3f80e0",
  1051 => x"d80b80e0",
  1052 => x"d8335456",
  1053 => x"72802ea9",
  1054 => x"3880e480",
  1055 => x"08735654",
  1056 => x"81165674",
  1057 => x"8a2e83ee",
  1058 => x"38841408",
  1059 => x"70822a81",
  1060 => x"06515372",
  1061 => x"802ef238",
  1062 => x"74740c75",
  1063 => x"335574e0",
  1064 => x"3880e3f0",
  1065 => x"08a01108",
  1066 => x"5355a051",
  1067 => x"ec873f80",
  1068 => x"e0e80b80",
  1069 => x"e0e83354",
  1070 => x"5672802e",
  1071 => x"a93880e4",
  1072 => x"80087356",
  1073 => x"54811656",
  1074 => x"748a2e83",
  1075 => x"ce388414",
  1076 => x"0870822a",
  1077 => x"81065153",
  1078 => x"72802ef2",
  1079 => x"3874740c",
  1080 => x"75335574",
  1081 => x"e03880e3",
  1082 => x"f008a411",
  1083 => x"085356a0",
  1084 => x"51ebc23f",
  1085 => x"80e48008",
  1086 => x"54841408",
  1087 => x"70822a81",
  1088 => x"06565374",
  1089 => x"802ef238",
  1090 => x"8d740c84",
  1091 => x"14087082",
  1092 => x"2a810657",
  1093 => x"5775802e",
  1094 => x"f2388a74",
  1095 => x"0c8d3d0d",
  1096 => x"04841408",
  1097 => x"70822a70",
  1098 => x"81065151",
  1099 => x"5372802e",
  1100 => x"f0388d74",
  1101 => x"0c841408",
  1102 => x"70822a70",
  1103 => x"81065151",
  1104 => x"5372802e",
  1105 => x"f9e638f9",
  1106 => x"f4398414",
  1107 => x"0870822a",
  1108 => x"70810651",
  1109 => x"51537280",
  1110 => x"2ef0388d",
  1111 => x"740c8414",
  1112 => x"0870822a",
  1113 => x"70810651",
  1114 => x"51537280",
  1115 => x"2ef9f638",
  1116 => x"fa843984",
  1117 => x"14087082",
  1118 => x"2a810651",
  1119 => x"5776802e",
  1120 => x"f2388d74",
  1121 => x"0c841408",
  1122 => x"70822a81",
  1123 => x"06515372",
  1124 => x"802efa92",
  1125 => x"38fa9e39",
  1126 => x"84140870",
  1127 => x"822a8106",
  1128 => x"51577680",
  1129 => x"2ef2388d",
  1130 => x"740c8414",
  1131 => x"0870822a",
  1132 => x"81065153",
  1133 => x"72802efa",
  1134 => x"b238fabe",
  1135 => x"39841408",
  1136 => x"70822a81",
  1137 => x"06515776",
  1138 => x"802ef238",
  1139 => x"8d740c84",
  1140 => x"14087082",
  1141 => x"2a810651",
  1142 => x"5372802e",
  1143 => x"fad238fa",
  1144 => x"de398414",
  1145 => x"0870822a",
  1146 => x"81065157",
  1147 => x"76802ef2",
  1148 => x"388d740c",
  1149 => x"84140870",
  1150 => x"822a8106",
  1151 => x"51537280",
  1152 => x"2efaf238",
  1153 => x"fafe3984",
  1154 => x"14087082",
  1155 => x"2a810651",
  1156 => x"5776802e",
  1157 => x"f2388d74",
  1158 => x"0c841408",
  1159 => x"70822a81",
  1160 => x"06515372",
  1161 => x"802efb92",
  1162 => x"38fb9e39",
  1163 => x"84140870",
  1164 => x"822a8106",
  1165 => x"51577680",
  1166 => x"2ef2388d",
  1167 => x"740c8414",
  1168 => x"0870822a",
  1169 => x"81065153",
  1170 => x"72802efb",
  1171 => x"b238fbbe",
  1172 => x"39841408",
  1173 => x"70822a81",
  1174 => x"06515776",
  1175 => x"802ef238",
  1176 => x"8d740c84",
  1177 => x"14087082",
  1178 => x"2a810651",
  1179 => x"5372802e",
  1180 => x"fbd238fb",
  1181 => x"de398414",
  1182 => x"0870822a",
  1183 => x"81065157",
  1184 => x"76802ef2",
  1185 => x"388d740c",
  1186 => x"84140870",
  1187 => x"822a8106",
  1188 => x"51537280",
  1189 => x"2efbf238",
  1190 => x"fbfe3984",
  1191 => x"14087082",
  1192 => x"2a810651",
  1193 => x"5776802e",
  1194 => x"f2388d74",
  1195 => x"0c841408",
  1196 => x"70822a81",
  1197 => x"06515372",
  1198 => x"802efc92",
  1199 => x"38fc9e39",
  1200 => x"ee3d0d80",
  1201 => x"0b80e484",
  1202 => x"08575574",
  1203 => x"76279a38",
  1204 => x"75753154",
  1205 => x"73fa8080",
  1206 => x"82aa1634",
  1207 => x"811580e4",
  1208 => x"84085755",
  1209 => x"757526e8",
  1210 => x"38800bfa",
  1211 => x"80808280",
  1212 => x"349b0bfa",
  1213 => x"80808281",
  1214 => x"34a10bfa",
  1215 => x"80808282",
  1216 => x"3480e80b",
  1217 => x"fa808082",
  1218 => x"833480cb",
  1219 => x"0bfa8080",
  1220 => x"8284348a",
  1221 => x"0bfa8080",
  1222 => x"828534de",
  1223 => x"0bfa8080",
  1224 => x"828634ff",
  1225 => x"ad0bfa80",
  1226 => x"80828734",
  1227 => x"ffbe0bfa",
  1228 => x"80808288",
  1229 => x"34ef0bfa",
  1230 => x"80808289",
  1231 => x"34800bfa",
  1232 => x"8080828a",
  1233 => x"34a00bfa",
  1234 => x"8080828b",
  1235 => x"34880bfa",
  1236 => x"8080828c",
  1237 => x"34800bfa",
  1238 => x"8080828d",
  1239 => x"3480c50b",
  1240 => x"fa808082",
  1241 => x"8e34800b",
  1242 => x"fa808082",
  1243 => x"8f349d16",
  1244 => x"7083ffff",
  1245 => x"0670882a",
  1246 => x"575b5474",
  1247 => x"fa808082",
  1248 => x"903479fa",
  1249 => x"80808291",
  1250 => x"34800bfa",
  1251 => x"80808292",
  1252 => x"34800bfa",
  1253 => x"80808293",
  1254 => x"3480c00b",
  1255 => x"fa808082",
  1256 => x"9434800b",
  1257 => x"fa808082",
  1258 => x"9534ff0b",
  1259 => x"fa808082",
  1260 => x"9634910b",
  1261 => x"fa808082",
  1262 => x"973480e7",
  1263 => x"0bfa8080",
  1264 => x"829834ff",
  1265 => x"8d0bfa80",
  1266 => x"80829934",
  1267 => x"8a0bfa80",
  1268 => x"80829a34",
  1269 => x"800bfa80",
  1270 => x"80829b34",
  1271 => x"800bfa80",
  1272 => x"80829c34",
  1273 => x"820bfa80",
  1274 => x"80829d34",
  1275 => x"8a0bfa80",
  1276 => x"80829e34",
  1277 => x"800bfa80",
  1278 => x"80829f34",
  1279 => x"800bfa80",
  1280 => x"8082a034",
  1281 => x"810bfa80",
  1282 => x"8082a134",
  1283 => x"930bfa80",
  1284 => x"8082a234",
  1285 => x"ffba0bfa",
  1286 => x"808082a3",
  1287 => x"34930bfa",
  1288 => x"808082a4",
  1289 => x"34ffba0b",
  1290 => x"fa808082",
  1291 => x"a5348816",
  1292 => x"7083ffff",
  1293 => x"0670882a",
  1294 => x"5a585977",
  1295 => x"fa808082",
  1296 => x"a63476fa",
  1297 => x"808082a7",
  1298 => x"34ff9f0b",
  1299 => x"fa808082",
  1300 => x"a834e30b",
  1301 => x"fa808082",
  1302 => x"a934fa80",
  1303 => x"8082800b",
  1304 => x"fa808080",
  1305 => x"840caa16",
  1306 => x"b0800785",
  1307 => x"0a0c80e3",
  1308 => x"f0085885",
  1309 => x"0a0b9419",
  1310 => x"0c91780c",
  1311 => x"850a0870",
  1312 => x"8b2a8106",
  1313 => x"575975f4",
  1314 => x"3880e0f8",
  1315 => x"0b80e0f8",
  1316 => x"337081ff",
  1317 => x"065c5657",
  1318 => x"79802eb8",
  1319 => x"387480e4",
  1320 => x"80085656",
  1321 => x"7581ff06",
  1322 => x"81185856",
  1323 => x"758a2e87",
  1324 => x"b8388415",
  1325 => x"0870822a",
  1326 => x"8106555a",
  1327 => x"73802ef2",
  1328 => x"3875750c",
  1329 => x"76337081",
  1330 => x"ff065556",
  1331 => x"73d63880",
  1332 => x"e0f83355",
  1333 => x"80e0f875",
  1334 => x"81ff0655",
  1335 => x"5673802e",
  1336 => x"bd387380",
  1337 => x"e3f80858",
  1338 => x"55811656",
  1339 => x"748a2e89",
  1340 => x"993880f4",
  1341 => x"80337010",
  1342 => x"101180f3",
  1343 => x"fc337190",
  1344 => x"29057088",
  1345 => x"2b78077a",
  1346 => x"0c80f3fc",
  1347 => x"33810551",
  1348 => x"51555973",
  1349 => x"80f3fc34",
  1350 => x"75335574",
  1351 => x"cc387708",
  1352 => x"923d5a56",
  1353 => x"8b5380df",
  1354 => x"b8527851",
  1355 => x"9ada3f88",
  1356 => x"02840580",
  1357 => x"c1055957",
  1358 => x"758f0654",
  1359 => x"73892688",
  1360 => x"98387618",
  1361 => x"b0155555",
  1362 => x"73753475",
  1363 => x"842aff18",
  1364 => x"7081ff06",
  1365 => x"59565676",
  1366 => x"df387879",
  1367 => x"33555773",
  1368 => x"802ea938",
  1369 => x"80e48008",
  1370 => x"74575581",
  1371 => x"1757758a",
  1372 => x"2e869b38",
  1373 => x"84150870",
  1374 => x"822a8106",
  1375 => x"595a7780",
  1376 => x"2ef23875",
  1377 => x"750c7633",
  1378 => x"5675e038",
  1379 => x"78793355",
  1380 => x"5673802e",
  1381 => x"bd387380",
  1382 => x"e3f80858",
  1383 => x"55811656",
  1384 => x"748a2e87",
  1385 => x"bd3880f4",
  1386 => x"80337010",
  1387 => x"101180f3",
  1388 => x"fc337190",
  1389 => x"29057088",
  1390 => x"2b78077a",
  1391 => x"0c80f3fc",
  1392 => x"33810558",
  1393 => x"5a555a74",
  1394 => x"80f3fc34",
  1395 => x"75335574",
  1396 => x"cc3880e1",
  1397 => x"8c0b80e1",
  1398 => x"8c337081",
  1399 => x"ff065757",
  1400 => x"5774802e",
  1401 => x"b63880e4",
  1402 => x"80085575",
  1403 => x"81ff0681",
  1404 => x"18585675",
  1405 => x"8a2e85bb",
  1406 => x"38841508",
  1407 => x"70822a81",
  1408 => x"065b5479",
  1409 => x"802ef238",
  1410 => x"75750c76",
  1411 => x"337081ff",
  1412 => x"065a5678",
  1413 => x"d63880e1",
  1414 => x"8c335680",
  1415 => x"e18c7681",
  1416 => x"ff065557",
  1417 => x"73802ebd",
  1418 => x"387380e3",
  1419 => x"f8085755",
  1420 => x"81175774",
  1421 => x"8a2e87f2",
  1422 => x"3880f480",
  1423 => x"33701010",
  1424 => x"1180f3fc",
  1425 => x"33719029",
  1426 => x"0570882b",
  1427 => x"7807790c",
  1428 => x"80f3fc33",
  1429 => x"8105585c",
  1430 => x"55597480",
  1431 => x"f3fc3476",
  1432 => x"335574cc",
  1433 => x"3880e3f0",
  1434 => x"08841108",
  1435 => x"903d5b57",
  1436 => x"578b5380",
  1437 => x"dfb85278",
  1438 => x"51988d3f",
  1439 => x"88028405",
  1440 => x"b5055957",
  1441 => x"758f0654",
  1442 => x"73892685",
  1443 => x"c3387618",
  1444 => x"b0155555",
  1445 => x"73753475",
  1446 => x"842aff18",
  1447 => x"7081ff06",
  1448 => x"59565676",
  1449 => x"df387879",
  1450 => x"33555773",
  1451 => x"802ea938",
  1452 => x"80e48008",
  1453 => x"74575581",
  1454 => x"1757758a",
  1455 => x"2e849938",
  1456 => x"84150870",
  1457 => x"822a8106",
  1458 => x"5b587980",
  1459 => x"2ef23875",
  1460 => x"750c7633",
  1461 => x"5675e038",
  1462 => x"78793355",
  1463 => x"5673802e",
  1464 => x"bd387380",
  1465 => x"e3f80858",
  1466 => x"55811656",
  1467 => x"748a2e86",
  1468 => x"913880f4",
  1469 => x"80337010",
  1470 => x"101180f3",
  1471 => x"fc337190",
  1472 => x"29057088",
  1473 => x"2b78077a",
  1474 => x"0c80f3fc",
  1475 => x"33810558",
  1476 => x"5c555874",
  1477 => x"80f3fc34",
  1478 => x"75335574",
  1479 => x"cc3880e1",
  1480 => x"a00b80e1",
  1481 => x"a0337081",
  1482 => x"ff065757",
  1483 => x"5774802e",
  1484 => x"b63880e4",
  1485 => x"80085575",
  1486 => x"81ff0681",
  1487 => x"18585675",
  1488 => x"8a2e83b9",
  1489 => x"38841508",
  1490 => x"70822a81",
  1491 => x"06595477",
  1492 => x"802ef238",
  1493 => x"75750c76",
  1494 => x"337081ff",
  1495 => x"065a5678",
  1496 => x"d63880e1",
  1497 => x"a0335680",
  1498 => x"e1a07681",
  1499 => x"ff065557",
  1500 => x"73802ebd",
  1501 => x"387380e3",
  1502 => x"f8085755",
  1503 => x"81175774",
  1504 => x"8a2e84d6",
  1505 => x"3880f480",
  1506 => x"33701010",
  1507 => x"1180f3fc",
  1508 => x"33719029",
  1509 => x"0570882b",
  1510 => x"7807790c",
  1511 => x"80f3fc33",
  1512 => x"8105585a",
  1513 => x"5b597480",
  1514 => x"f3fc3476",
  1515 => x"335574cc",
  1516 => x"38850a08",
  1517 => x"8c3d5a56",
  1518 => x"8b5380df",
  1519 => x"b8527851",
  1520 => x"95c63f88",
  1521 => x"028405a9",
  1522 => x"05595775",
  1523 => x"8f065473",
  1524 => x"892682f3",
  1525 => x"387618b0",
  1526 => x"15555573",
  1527 => x"75347584",
  1528 => x"2aff1870",
  1529 => x"81ff0659",
  1530 => x"565676df",
  1531 => x"38787933",
  1532 => x"55577380",
  1533 => x"2ea93880",
  1534 => x"e4800874",
  1535 => x"57558117",
  1536 => x"57758a2e",
  1537 => x"829c3884",
  1538 => x"15087082",
  1539 => x"2a810659",
  1540 => x"5477802e",
  1541 => x"f2387575",
  1542 => x"0c763356",
  1543 => x"75e03878",
  1544 => x"79335556",
  1545 => x"73802ebd",
  1546 => x"387380e3",
  1547 => x"f8085855",
  1548 => x"81165674",
  1549 => x"8a2e82fa",
  1550 => x"3880f480",
  1551 => x"33701010",
  1552 => x"1180f3fc",
  1553 => x"33719029",
  1554 => x"0570882b",
  1555 => x"78077a0c",
  1556 => x"80f3fc33",
  1557 => x"8105585a",
  1558 => x"5b547480",
  1559 => x"f3fc3475",
  1560 => x"335574cc",
  1561 => x"38943d0d",
  1562 => x"04841508",
  1563 => x"70822a81",
  1564 => x"06555a73",
  1565 => x"802ef238",
  1566 => x"8d750c84",
  1567 => x"15087082",
  1568 => x"2a810655",
  1569 => x"5a73802e",
  1570 => x"f8a838f8",
  1571 => x"b4398415",
  1572 => x"0870822a",
  1573 => x"8106595a",
  1574 => x"77802ef2",
  1575 => x"388d750c",
  1576 => x"84150870",
  1577 => x"822a8106",
  1578 => x"595a7780",
  1579 => x"2ef9c538",
  1580 => x"f9d13984",
  1581 => x"15087082",
  1582 => x"2a810659",
  1583 => x"5977802e",
  1584 => x"f2388d75",
  1585 => x"0c841508",
  1586 => x"70822a81",
  1587 => x"065b5479",
  1588 => x"802efaa5",
  1589 => x"38fab139",
  1590 => x"84150870",
  1591 => x"822a8106",
  1592 => x"5b587980",
  1593 => x"2ef2388d",
  1594 => x"750c8415",
  1595 => x"0870822a",
  1596 => x"81065b58",
  1597 => x"79802efb",
  1598 => x"c738fbd3",
  1599 => x"39841508",
  1600 => x"70822a81",
  1601 => x"065b5979",
  1602 => x"802ef238",
  1603 => x"8d750c84",
  1604 => x"15087082",
  1605 => x"2a810659",
  1606 => x"5477802e",
  1607 => x"fca738fc",
  1608 => x"b3398415",
  1609 => x"0870822a",
  1610 => x"81065954",
  1611 => x"77802ef2",
  1612 => x"388d750c",
  1613 => x"84150870",
  1614 => x"822a8106",
  1615 => x"59547780",
  1616 => x"2efdc438",
  1617 => x"fdd03976",
  1618 => x"18b71555",
  1619 => x"55fd8c39",
  1620 => x"7618b715",
  1621 => x"5555fabc",
  1622 => x"397618b7",
  1623 => x"155555f7",
  1624 => x"e73980f4",
  1625 => x"80337081",
  1626 => x"ff065a55",
  1627 => x"78a32681",
  1628 => x"ef388115",
  1629 => x"587780f4",
  1630 => x"8034800b",
  1631 => x"80f3fc34",
  1632 => x"75335574",
  1633 => x"f89738f8",
  1634 => x"c93980f4",
  1635 => x"80337081",
  1636 => x"ff065a55",
  1637 => x"78a32681",
  1638 => x"b8388115",
  1639 => x"5a7980f4",
  1640 => x"8034800b",
  1641 => x"80f3fc34",
  1642 => x"75335574",
  1643 => x"f6bb38f6",
  1644 => x"ed3980f4",
  1645 => x"80337081",
  1646 => x"ff065a55",
  1647 => x"78a32681",
  1648 => x"da388115",
  1649 => x"587780f4",
  1650 => x"8034800b",
  1651 => x"80f3fc34",
  1652 => x"75335574",
  1653 => x"fcda38fd",
  1654 => x"8c3980f4",
  1655 => x"80337081",
  1656 => x"ff065955",
  1657 => x"77a32681",
  1658 => x"a3388115",
  1659 => x"5a7980f4",
  1660 => x"8034800b",
  1661 => x"80f3fc34",
  1662 => x"76335574",
  1663 => x"fafe38fb",
  1664 => x"b03980f4",
  1665 => x"80337081",
  1666 => x"ff065a55",
  1667 => x"78a32680",
  1668 => x"ec388115",
  1669 => x"5a7980f4",
  1670 => x"8034800b",
  1671 => x"80f3fc34",
  1672 => x"75335574",
  1673 => x"f9c338f9",
  1674 => x"f53980f4",
  1675 => x"80337081",
  1676 => x"ff065b55",
  1677 => x"79a326b7",
  1678 => x"38811558",
  1679 => x"7780f480",
  1680 => x"34800b80",
  1681 => x"f3fc3476",
  1682 => x"335574f7",
  1683 => x"e338f895",
  1684 => x"39800b80",
  1685 => x"f4803480",
  1686 => x"0b80f3fc",
  1687 => x"34fec939",
  1688 => x"800b80f4",
  1689 => x"8034800b",
  1690 => x"80f3fc34",
  1691 => x"fe923980",
  1692 => x"0b80f480",
  1693 => x"34800b80",
  1694 => x"f3fc34cb",
  1695 => x"39800b80",
  1696 => x"f4803480",
  1697 => x"0b80f3fc",
  1698 => x"34ff9539",
  1699 => x"800b80f4",
  1700 => x"8034800b",
  1701 => x"80f3fc34",
  1702 => x"fede3980",
  1703 => x"0b80f480",
  1704 => x"34800b80",
  1705 => x"f3fc34fe",
  1706 => x"a739f73d",
  1707 => x"0d80e3f4",
  1708 => x"08700881",
  1709 => x"0a0680e3",
  1710 => x"fc08565a",
  1711 => x"53870b84",
  1712 => x"150c80e3",
  1713 => x"f8085780",
  1714 => x"0b84180c",
  1715 => x"fe800a0b",
  1716 => x"88180c80",
  1717 => x"0b80f480",
  1718 => x"34800b80",
  1719 => x"f3fc3480",
  1720 => x"e4800855",
  1721 => x"b60b8c16",
  1722 => x"0c830b88",
  1723 => x"160c81ff",
  1724 => x"0b88140c",
  1725 => x"80e3f008",
  1726 => x"54ff0b84",
  1727 => x"150cfc94",
  1728 => x"800b8815",
  1729 => x"0c82d0af",
  1730 => x"fdfb0b8c",
  1731 => x"150c80c0",
  1732 => x"740c7308",
  1733 => x"70862a81",
  1734 => x"06575a75",
  1735 => x"f5389014",
  1736 => x"0870832a",
  1737 => x"81065458",
  1738 => x"72f43881",
  1739 => x"fc80810b",
  1740 => x"90150c90",
  1741 => x"14087083",
  1742 => x"2a81065b",
  1743 => x"5679f438",
  1744 => x"80fdc081",
  1745 => x"0b90150c",
  1746 => x"80e1b40b",
  1747 => x"80e1b433",
  1748 => x"7081ff06",
  1749 => x"5a555677",
  1750 => x"802eb138",
  1751 => x"7381ff06",
  1752 => x"81175754",
  1753 => x"738a2e84",
  1754 => x"eb388415",
  1755 => x"0870822a",
  1756 => x"81065b58",
  1757 => x"79802ef2",
  1758 => x"3873750c",
  1759 => x"75337081",
  1760 => x"ff065b54",
  1761 => x"79d63880",
  1762 => x"e1b43354",
  1763 => x"80e1b474",
  1764 => x"81ff0654",
  1765 => x"5672802e",
  1766 => x"b8387254",
  1767 => x"81165673",
  1768 => x"8a2e85ec",
  1769 => x"3880f480",
  1770 => x"33701010",
  1771 => x"1180f3fc",
  1772 => x"33719029",
  1773 => x"0570882b",
  1774 => x"77077a0c",
  1775 => x"80f3fc33",
  1776 => x"81055d52",
  1777 => x"54587980",
  1778 => x"f3fc3475",
  1779 => x"335473cc",
  1780 => x"3880e1b8",
  1781 => x"0b80e1b8",
  1782 => x"337081ff",
  1783 => x"06555556",
  1784 => x"72802eb1",
  1785 => x"387381ff",
  1786 => x"06811757",
  1787 => x"54738a2e",
  1788 => x"84873884",
  1789 => x"15087082",
  1790 => x"2a81065b",
  1791 => x"5379802e",
  1792 => x"f2387375",
  1793 => x"0c753370",
  1794 => x"81ff065b",
  1795 => x"5479d638",
  1796 => x"80e1b833",
  1797 => x"5480e1b8",
  1798 => x"7481ff06",
  1799 => x"54567280",
  1800 => x"2eb83872",
  1801 => x"54811656",
  1802 => x"738a2e85",
  1803 => x"8b3880f4",
  1804 => x"80337010",
  1805 => x"101180f3",
  1806 => x"fc337190",
  1807 => x"29057088",
  1808 => x"2b77077a",
  1809 => x"0c80f3fc",
  1810 => x"3381055d",
  1811 => x"51545879",
  1812 => x"80f3fc34",
  1813 => x"75335473",
  1814 => x"cc387880",
  1815 => x"2e85d738",
  1816 => x"80e1c00b",
  1817 => x"80e1c033",
  1818 => x"7081ff06",
  1819 => x"55555672",
  1820 => x"802eb138",
  1821 => x"7381ff06",
  1822 => x"81175754",
  1823 => x"738a2e83",
  1824 => x"9d388415",
  1825 => x"0870822a",
  1826 => x"81065b53",
  1827 => x"79802ef2",
  1828 => x"3873750c",
  1829 => x"75337081",
  1830 => x"ff065b54",
  1831 => x"79d63880",
  1832 => x"e1c03354",
  1833 => x"80e1c074",
  1834 => x"81ff0654",
  1835 => x"5672802e",
  1836 => x"b8387254",
  1837 => x"81165673",
  1838 => x"8a2e84d2",
  1839 => x"3880f480",
  1840 => x"33701010",
  1841 => x"1180f3fc",
  1842 => x"33719029",
  1843 => x"0570882b",
  1844 => x"77077a0c",
  1845 => x"80f3fc33",
  1846 => x"81055d51",
  1847 => x"54587980",
  1848 => x"f3fc3475",
  1849 => x"335473cc",
  1850 => x"3880e1d0",
  1851 => x"0b80e1d0",
  1852 => x"337081ff",
  1853 => x"06555556",
  1854 => x"72802eb1",
  1855 => x"387381ff",
  1856 => x"06811757",
  1857 => x"54738a2e",
  1858 => x"82b93884",
  1859 => x"15087082",
  1860 => x"2a81065b",
  1861 => x"5379802e",
  1862 => x"f2387375",
  1863 => x"0c753370",
  1864 => x"81ff065b",
  1865 => x"5479d638",
  1866 => x"80e1d033",
  1867 => x"5480e1d0",
  1868 => x"7481ff06",
  1869 => x"54557280",
  1870 => x"2eb83872",
  1871 => x"54811555",
  1872 => x"738a2e82",
  1873 => x"a33880f4",
  1874 => x"80337010",
  1875 => x"101180f3",
  1876 => x"fc337190",
  1877 => x"29057088",
  1878 => x"2b77077a",
  1879 => x"0c80f3fc",
  1880 => x"33810557",
  1881 => x"58545a73",
  1882 => x"80f3fc34",
  1883 => x"74335473",
  1884 => x"cc38eacc",
  1885 => x"3ff881c0",
  1886 => x"8e8055a0",
  1887 => x"0b80e3f4",
  1888 => x"0880e3fc",
  1889 => x"085a5856",
  1890 => x"7484180c",
  1891 => x"749f2a75",
  1892 => x"10075578",
  1893 => x"802e9838",
  1894 => x"75802e82",
  1895 => x"c238ff16",
  1896 => x"7584190c",
  1897 => x"759f2a76",
  1898 => x"10075656",
  1899 => x"78ea3877",
  1900 => x"54afd7c2",
  1901 => x"0b94190c",
  1902 => x"850b9819",
  1903 => x"0c981408",
  1904 => x"81065372",
  1905 => x"802ec138",
  1906 => x"98140881",
  1907 => x"065372ed",
  1908 => x"38ffb539",
  1909 => x"84150870",
  1910 => x"822a8106",
  1911 => x"5b587980",
  1912 => x"2ef2388d",
  1913 => x"750c8415",
  1914 => x"0870822a",
  1915 => x"81065b58",
  1916 => x"79802efa",
  1917 => x"f538fb81",
  1918 => x"39841508",
  1919 => x"70822a81",
  1920 => x"065b5379",
  1921 => x"802ef238",
  1922 => x"8d750c84",
  1923 => x"15087082",
  1924 => x"2a81065b",
  1925 => x"5379802e",
  1926 => x"fbd938fb",
  1927 => x"e5398415",
  1928 => x"0870822a",
  1929 => x"81065b53",
  1930 => x"79802ef2",
  1931 => x"388d750c",
  1932 => x"84150870",
  1933 => x"822a8106",
  1934 => x"5b537980",
  1935 => x"2efcc338",
  1936 => x"fccf3984",
  1937 => x"15087082",
  1938 => x"2a81065b",
  1939 => x"5379802e",
  1940 => x"f2388d75",
  1941 => x"0c841508",
  1942 => x"70822a81",
  1943 => x"065b5379",
  1944 => x"802efda7",
  1945 => x"38fdb339",
  1946 => x"80f48033",
  1947 => x"7081ff06",
  1948 => x"575475a3",
  1949 => x"2680eb38",
  1950 => x"81145877",
  1951 => x"80f48034",
  1952 => x"800b80f3",
  1953 => x"fc347433",
  1954 => x"5473fdb1",
  1955 => x"38fde339",
  1956 => x"80f48033",
  1957 => x"7081ff06",
  1958 => x"545472a3",
  1959 => x"2680e038",
  1960 => x"81145877",
  1961 => x"80f48034",
  1962 => x"800b80f3",
  1963 => x"fc347533",
  1964 => x"5473f9e8",
  1965 => x"38fa9a39",
  1966 => x"80f48033",
  1967 => x"7081ff06",
  1968 => x"595477a3",
  1969 => x"26ab3881",
  1970 => x"14537280",
  1971 => x"f4803480",
  1972 => x"0b80f3fc",
  1973 => x"34753354",
  1974 => x"73faca38",
  1975 => x"fafc3987",
  1976 => x"9a3f800b",
  1977 => x"80f48034",
  1978 => x"800b80f3",
  1979 => x"fc34ff96",
  1980 => x"39800b80",
  1981 => x"f4803480",
  1982 => x"0b80f3fc",
  1983 => x"34d73980",
  1984 => x"0b80f480",
  1985 => x"34800b80",
  1986 => x"f3fc34ff",
  1987 => x"a13980f4",
  1988 => x"80337081",
  1989 => x"ff065954",
  1990 => x"77a32682",
  1991 => x"89388114",
  1992 => x"537280f4",
  1993 => x"8034800b",
  1994 => x"80f3fc34",
  1995 => x"75335473",
  1996 => x"fb8238fb",
  1997 => x"b43980e1",
  1998 => x"f40b80e1",
  1999 => x"f4337081",
  2000 => x"ff065555",
  2001 => x"5672802e",
  2002 => x"b1387381",
  2003 => x"ff068117",
  2004 => x"5754738a",
  2005 => x"2e819c38",
  2006 => x"84150870",
  2007 => x"822a8106",
  2008 => x"5b537980",
  2009 => x"2ef23873",
  2010 => x"750c7533",
  2011 => x"7081ff06",
  2012 => x"5b5479d6",
  2013 => x"3880e1f4",
  2014 => x"335480e1",
  2015 => x"f47481ff",
  2016 => x"06545672",
  2017 => x"802efae1",
  2018 => x"38728117",
  2019 => x"5754738a",
  2020 => x"2ebb3880",
  2021 => x"f4803370",
  2022 => x"10101180",
  2023 => x"f3fc3371",
  2024 => x"90290570",
  2025 => x"882b7707",
  2026 => x"7a0c80f3",
  2027 => x"fc338105",
  2028 => x"5d515458",
  2029 => x"7980f3fc",
  2030 => x"34753354",
  2031 => x"73802efa",
  2032 => x"a8388116",
  2033 => x"56738a2e",
  2034 => x"098106c7",
  2035 => x"3880f480",
  2036 => x"337081ff",
  2037 => x"06595477",
  2038 => x"a326bd38",
  2039 => x"81145372",
  2040 => x"80f48034",
  2041 => x"800b80f3",
  2042 => x"fc347533",
  2043 => x"5473d338",
  2044 => x"f9f73984",
  2045 => x"15087082",
  2046 => x"2a81065b",
  2047 => x"5379802e",
  2048 => x"f2388d75",
  2049 => x"0c841508",
  2050 => x"70822a81",
  2051 => x"065b5379",
  2052 => x"802efec4",
  2053 => x"38fed039",
  2054 => x"800b80f4",
  2055 => x"8034800b",
  2056 => x"80f3fc34",
  2057 => x"c539800b",
  2058 => x"80f48034",
  2059 => x"800b80f3",
  2060 => x"fc34fdf8",
  2061 => x"398c0802",
  2062 => x"8c0cfd3d",
  2063 => x"0d80538c",
  2064 => x"088c0508",
  2065 => x"528c0888",
  2066 => x"05085182",
  2067 => x"de3f8008",
  2068 => x"70800c54",
  2069 => x"853d0d8c",
  2070 => x"0c048c08",
  2071 => x"028c0cfd",
  2072 => x"3d0d8153",
  2073 => x"8c088c05",
  2074 => x"08528c08",
  2075 => x"88050851",
  2076 => x"82b93f80",
  2077 => x"0870800c",
  2078 => x"54853d0d",
  2079 => x"8c0c048c",
  2080 => x"08028c0c",
  2081 => x"f93d0d80",
  2082 => x"0b8c08fc",
  2083 => x"050c8c08",
  2084 => x"88050880",
  2085 => x"25ab388c",
  2086 => x"08880508",
  2087 => x"308c0888",
  2088 => x"050c800b",
  2089 => x"8c08f405",
  2090 => x"0c8c08fc",
  2091 => x"05088838",
  2092 => x"810b8c08",
  2093 => x"f4050c8c",
  2094 => x"08f40508",
  2095 => x"8c08fc05",
  2096 => x"0c8c088c",
  2097 => x"05088025",
  2098 => x"ab388c08",
  2099 => x"8c050830",
  2100 => x"8c088c05",
  2101 => x"0c800b8c",
  2102 => x"08f0050c",
  2103 => x"8c08fc05",
  2104 => x"08883881",
  2105 => x"0b8c08f0",
  2106 => x"050c8c08",
  2107 => x"f005088c",
  2108 => x"08fc050c",
  2109 => x"80538c08",
  2110 => x"8c050852",
  2111 => x"8c088805",
  2112 => x"085181a7",
  2113 => x"3f800870",
  2114 => x"8c08f805",
  2115 => x"0c548c08",
  2116 => x"fc050880",
  2117 => x"2e8c388c",
  2118 => x"08f80508",
  2119 => x"308c08f8",
  2120 => x"050c8c08",
  2121 => x"f8050870",
  2122 => x"800c5489",
  2123 => x"3d0d8c0c",
  2124 => x"048c0802",
  2125 => x"8c0cfb3d",
  2126 => x"0d800b8c",
  2127 => x"08fc050c",
  2128 => x"8c088805",
  2129 => x"08802593",
  2130 => x"388c0888",
  2131 => x"0508308c",
  2132 => x"0888050c",
  2133 => x"810b8c08",
  2134 => x"fc050c8c",
  2135 => x"088c0508",
  2136 => x"80258c38",
  2137 => x"8c088c05",
  2138 => x"08308c08",
  2139 => x"8c050c81",
  2140 => x"538c088c",
  2141 => x"0508528c",
  2142 => x"08880508",
  2143 => x"51ad3f80",
  2144 => x"08708c08",
  2145 => x"f8050c54",
  2146 => x"8c08fc05",
  2147 => x"08802e8c",
  2148 => x"388c08f8",
  2149 => x"0508308c",
  2150 => x"08f8050c",
  2151 => x"8c08f805",
  2152 => x"0870800c",
  2153 => x"54873d0d",
  2154 => x"8c0c048c",
  2155 => x"08028c0c",
  2156 => x"fd3d0d81",
  2157 => x"0b8c08fc",
  2158 => x"050c800b",
  2159 => x"8c08f805",
  2160 => x"0c8c088c",
  2161 => x"05088c08",
  2162 => x"88050827",
  2163 => x"ac388c08",
  2164 => x"fc050880",
  2165 => x"2ea33880",
  2166 => x"0b8c088c",
  2167 => x"05082499",
  2168 => x"388c088c",
  2169 => x"0508108c",
  2170 => x"088c050c",
  2171 => x"8c08fc05",
  2172 => x"08108c08",
  2173 => x"fc050cc9",
  2174 => x"398c08fc",
  2175 => x"0508802e",
  2176 => x"80c9388c",
  2177 => x"088c0508",
  2178 => x"8c088805",
  2179 => x"0826a138",
  2180 => x"8c088805",
  2181 => x"088c088c",
  2182 => x"0508318c",
  2183 => x"0888050c",
  2184 => x"8c08f805",
  2185 => x"088c08fc",
  2186 => x"0508078c",
  2187 => x"08f8050c",
  2188 => x"8c08fc05",
  2189 => x"08812a8c",
  2190 => x"08fc050c",
  2191 => x"8c088c05",
  2192 => x"08812a8c",
  2193 => x"088c050c",
  2194 => x"ffaf398c",
  2195 => x"08900508",
  2196 => x"802e8f38",
  2197 => x"8c088805",
  2198 => x"08708c08",
  2199 => x"f4050c51",
  2200 => x"8d398c08",
  2201 => x"f8050870",
  2202 => x"8c08f405",
  2203 => x"0c518c08",
  2204 => x"f4050880",
  2205 => x"0c853d0d",
  2206 => x"8c0c0480",
  2207 => x"3d0d8651",
  2208 => x"84963f81",
  2209 => x"5198d73f",
  2210 => x"fc3d0d76",
  2211 => x"70797b55",
  2212 => x"5555558f",
  2213 => x"72278c38",
  2214 => x"72750783",
  2215 => x"06517080",
  2216 => x"2ea738ff",
  2217 => x"125271ff",
  2218 => x"2e983872",
  2219 => x"70810554",
  2220 => x"33747081",
  2221 => x"055634ff",
  2222 => x"125271ff",
  2223 => x"2e098106",
  2224 => x"ea387480",
  2225 => x"0c863d0d",
  2226 => x"04745172",
  2227 => x"70840554",
  2228 => x"08717084",
  2229 => x"05530c72",
  2230 => x"70840554",
  2231 => x"08717084",
  2232 => x"05530c72",
  2233 => x"70840554",
  2234 => x"08717084",
  2235 => x"05530c72",
  2236 => x"70840554",
  2237 => x"08717084",
  2238 => x"05530cf0",
  2239 => x"1252718f",
  2240 => x"26c93883",
  2241 => x"72279538",
  2242 => x"72708405",
  2243 => x"54087170",
  2244 => x"8405530c",
  2245 => x"fc125271",
  2246 => x"8326ed38",
  2247 => x"7054ff83",
  2248 => x"39fd3d0d",
  2249 => x"755384d8",
  2250 => x"1308802e",
  2251 => x"8a388053",
  2252 => x"72800c85",
  2253 => x"3d0d0481",
  2254 => x"80527251",
  2255 => x"83d83f80",
  2256 => x"0884d814",
  2257 => x"0cff5380",
  2258 => x"08802ee4",
  2259 => x"38800854",
  2260 => x"9f538074",
  2261 => x"70840556",
  2262 => x"0cff1353",
  2263 => x"807324ce",
  2264 => x"38807470",
  2265 => x"8405560c",
  2266 => x"ff135372",
  2267 => x"8025e338",
  2268 => x"ffbc39fd",
  2269 => x"3d0d7577",
  2270 => x"55539f74",
  2271 => x"278d3896",
  2272 => x"730cff52",
  2273 => x"71800c85",
  2274 => x"3d0d0484",
  2275 => x"d8130852",
  2276 => x"71802e93",
  2277 => x"38731010",
  2278 => x"12700879",
  2279 => x"720c5152",
  2280 => x"71800c85",
  2281 => x"3d0d0472",
  2282 => x"51fef63f",
  2283 => x"ff528008",
  2284 => x"d33884d8",
  2285 => x"13087410",
  2286 => x"10117008",
  2287 => x"7a720c51",
  2288 => x"5152dd39",
  2289 => x"f93d0d79",
  2290 => x"7b585676",
  2291 => x"9f2680e8",
  2292 => x"3884d816",
  2293 => x"08547380",
  2294 => x"2eaa3876",
  2295 => x"10101470",
  2296 => x"08555573",
  2297 => x"802eba38",
  2298 => x"80587381",
  2299 => x"2e8f3873",
  2300 => x"ff2ea338",
  2301 => x"80750c76",
  2302 => x"51732d80",
  2303 => x"5877800c",
  2304 => x"893d0d04",
  2305 => x"7551fe99",
  2306 => x"3fff5880",
  2307 => x"08ef3884",
  2308 => x"d8160854",
  2309 => x"c6399676",
  2310 => x"0c810b80",
  2311 => x"0c893d0d",
  2312 => x"04755181",
  2313 => x"ed3f7653",
  2314 => x"80085275",
  2315 => x"5181ad3f",
  2316 => x"8008800c",
  2317 => x"893d0d04",
  2318 => x"96760cff",
  2319 => x"0b800c89",
  2320 => x"3d0d04fc",
  2321 => x"3d0d7678",
  2322 => x"5653ff54",
  2323 => x"749f26b1",
  2324 => x"3884d813",
  2325 => x"08527180",
  2326 => x"2eae3874",
  2327 => x"10101270",
  2328 => x"08535381",
  2329 => x"5471802e",
  2330 => x"98388254",
  2331 => x"71ff2e91",
  2332 => x"38835471",
  2333 => x"812e8a38",
  2334 => x"80730c74",
  2335 => x"51712d80",
  2336 => x"5473800c",
  2337 => x"863d0d04",
  2338 => x"7251fd95",
  2339 => x"3f8008f1",
  2340 => x"3884d813",
  2341 => x"0852c439",
  2342 => x"ff3d0d73",
  2343 => x"5280e488",
  2344 => x"0851fea0",
  2345 => x"3f833d0d",
  2346 => x"04fe3d0d",
  2347 => x"75537452",
  2348 => x"80e48808",
  2349 => x"51fdbc3f",
  2350 => x"843d0d04",
  2351 => x"803d0d80",
  2352 => x"e4880851",
  2353 => x"fcdb3f82",
  2354 => x"3d0d04ff",
  2355 => x"3d0d7352",
  2356 => x"80e48808",
  2357 => x"51feec3f",
  2358 => x"833d0d04",
  2359 => x"fc3d0d80",
  2360 => x"0b80f484",
  2361 => x"0c785277",
  2362 => x"5192e73f",
  2363 => x"80085480",
  2364 => x"08ff2e88",
  2365 => x"3873800c",
  2366 => x"863d0d04",
  2367 => x"80f48408",
  2368 => x"5574802e",
  2369 => x"f0387675",
  2370 => x"710c5373",
  2371 => x"800c863d",
  2372 => x"0d0492b9",
  2373 => x"3f04f33d",
  2374 => x"0d7f618b",
  2375 => x"1170f806",
  2376 => x"5c55555e",
  2377 => x"72962683",
  2378 => x"38905980",
  2379 => x"7924747a",
  2380 => x"26075380",
  2381 => x"5472742e",
  2382 => x"09810680",
  2383 => x"cb387d51",
  2384 => x"8bca3f78",
  2385 => x"83f72680",
  2386 => x"c6387883",
  2387 => x"2a701010",
  2388 => x"1080ebc4",
  2389 => x"058c1108",
  2390 => x"59595a76",
  2391 => x"782e83b0",
  2392 => x"38841708",
  2393 => x"fc06568c",
  2394 => x"17088818",
  2395 => x"08718c12",
  2396 => x"0c88120c",
  2397 => x"58751784",
  2398 => x"11088107",
  2399 => x"84120c53",
  2400 => x"7d518b89",
  2401 => x"3f881754",
  2402 => x"73800c8f",
  2403 => x"3d0d0478",
  2404 => x"892a7983",
  2405 => x"2a5b5372",
  2406 => x"802ebf38",
  2407 => x"78862ab8",
  2408 => x"055a8473",
  2409 => x"27b43880",
  2410 => x"db135a94",
  2411 => x"7327ab38",
  2412 => x"788c2a80",
  2413 => x"ee055a80",
  2414 => x"d473279e",
  2415 => x"38788f2a",
  2416 => x"80f7055a",
  2417 => x"82d47327",
  2418 => x"91387892",
  2419 => x"2a80fc05",
  2420 => x"5a8ad473",
  2421 => x"27843880",
  2422 => x"fe5a7910",
  2423 => x"101080eb",
  2424 => x"c4058c11",
  2425 => x"08585576",
  2426 => x"752ea338",
  2427 => x"841708fc",
  2428 => x"06707a31",
  2429 => x"5556738f",
  2430 => x"2488d538",
  2431 => x"738025fe",
  2432 => x"e6388c17",
  2433 => x"08577675",
  2434 => x"2e098106",
  2435 => x"df38811a",
  2436 => x"5a80ebd4",
  2437 => x"08577680",
  2438 => x"ebcc2e82",
  2439 => x"c0388417",
  2440 => x"08fc0670",
  2441 => x"7a315556",
  2442 => x"738f2481",
  2443 => x"f93880eb",
  2444 => x"cc0b80eb",
  2445 => x"d80c80eb",
  2446 => x"cc0b80eb",
  2447 => x"d40c7380",
  2448 => x"25feb238",
  2449 => x"83ff7627",
  2450 => x"83df3875",
  2451 => x"892a7683",
  2452 => x"2a555372",
  2453 => x"802ebf38",
  2454 => x"75862ab8",
  2455 => x"05548473",
  2456 => x"27b43880",
  2457 => x"db135494",
  2458 => x"7327ab38",
  2459 => x"758c2a80",
  2460 => x"ee055480",
  2461 => x"d473279e",
  2462 => x"38758f2a",
  2463 => x"80f70554",
  2464 => x"82d47327",
  2465 => x"91387592",
  2466 => x"2a80fc05",
  2467 => x"548ad473",
  2468 => x"27843880",
  2469 => x"fe547310",
  2470 => x"101080eb",
  2471 => x"c4058811",
  2472 => x"08565874",
  2473 => x"782e86cf",
  2474 => x"38841508",
  2475 => x"fc065375",
  2476 => x"73278d38",
  2477 => x"88150855",
  2478 => x"74782e09",
  2479 => x"8106ea38",
  2480 => x"8c150880",
  2481 => x"ebc40b84",
  2482 => x"0508718c",
  2483 => x"1a0c7688",
  2484 => x"1a0c7888",
  2485 => x"130c788c",
  2486 => x"180c5d58",
  2487 => x"7953807a",
  2488 => x"2483e638",
  2489 => x"72822c81",
  2490 => x"712b5c53",
  2491 => x"7a7c2681",
  2492 => x"98387b7b",
  2493 => x"06537282",
  2494 => x"f13879fc",
  2495 => x"0684055a",
  2496 => x"7a10707d",
  2497 => x"06545b72",
  2498 => x"82e03884",
  2499 => x"1a5af139",
  2500 => x"88178c11",
  2501 => x"08585876",
  2502 => x"782e0981",
  2503 => x"06fcc238",
  2504 => x"821a5afd",
  2505 => x"ec397817",
  2506 => x"79810784",
  2507 => x"190c7080",
  2508 => x"ebd80c70",
  2509 => x"80ebd40c",
  2510 => x"80ebcc0b",
  2511 => x"8c120c8c",
  2512 => x"11088812",
  2513 => x"0c748107",
  2514 => x"84120c74",
  2515 => x"1175710c",
  2516 => x"51537d51",
  2517 => x"87b73f88",
  2518 => x"1754fcac",
  2519 => x"3980ebc4",
  2520 => x"0b840508",
  2521 => x"7a545c79",
  2522 => x"8025fef8",
  2523 => x"3882da39",
  2524 => x"7a097c06",
  2525 => x"7080ebc4",
  2526 => x"0b84050c",
  2527 => x"5c7a105b",
  2528 => x"7a7c2685",
  2529 => x"387a85b8",
  2530 => x"3880ebc4",
  2531 => x"0b880508",
  2532 => x"70841208",
  2533 => x"fc06707c",
  2534 => x"317c7226",
  2535 => x"8f722507",
  2536 => x"57575c5d",
  2537 => x"5572802e",
  2538 => x"80db3879",
  2539 => x"7a1680eb",
  2540 => x"bc081b90",
  2541 => x"115a5557",
  2542 => x"5b80ebb8",
  2543 => x"08ff2e88",
  2544 => x"38a08f13",
  2545 => x"e0800657",
  2546 => x"76527d51",
  2547 => x"86c03f80",
  2548 => x"08548008",
  2549 => x"ff2e9038",
  2550 => x"80087627",
  2551 => x"82993874",
  2552 => x"80ebc42e",
  2553 => x"82913880",
  2554 => x"ebc40b88",
  2555 => x"05085584",
  2556 => x"1508fc06",
  2557 => x"707a317a",
  2558 => x"72268f72",
  2559 => x"25075255",
  2560 => x"537283e6",
  2561 => x"38747981",
  2562 => x"0784170c",
  2563 => x"79167080",
  2564 => x"ebc40b88",
  2565 => x"050c7581",
  2566 => x"0784120c",
  2567 => x"547e5257",
  2568 => x"85eb3f88",
  2569 => x"1754fae0",
  2570 => x"3975832a",
  2571 => x"70545480",
  2572 => x"7424819b",
  2573 => x"3872822c",
  2574 => x"81712b80",
  2575 => x"ebc80807",
  2576 => x"7080ebc4",
  2577 => x"0b84050c",
  2578 => x"75101010",
  2579 => x"80ebc405",
  2580 => x"88110858",
  2581 => x"5a5d5377",
  2582 => x"8c180c74",
  2583 => x"88180c76",
  2584 => x"88190c76",
  2585 => x"8c160cfc",
  2586 => x"f339797a",
  2587 => x"10101080",
  2588 => x"ebc40570",
  2589 => x"57595d8c",
  2590 => x"15085776",
  2591 => x"752ea338",
  2592 => x"841708fc",
  2593 => x"06707a31",
  2594 => x"5556738f",
  2595 => x"2483ca38",
  2596 => x"73802584",
  2597 => x"81388c17",
  2598 => x"08577675",
  2599 => x"2e098106",
  2600 => x"df388815",
  2601 => x"811b7083",
  2602 => x"06555b55",
  2603 => x"72c9387c",
  2604 => x"83065372",
  2605 => x"802efdb8",
  2606 => x"38ff1df8",
  2607 => x"19595d88",
  2608 => x"1808782e",
  2609 => x"ea38fdb5",
  2610 => x"39831a53",
  2611 => x"fc963983",
  2612 => x"1470822c",
  2613 => x"81712b80",
  2614 => x"ebc80807",
  2615 => x"7080ebc4",
  2616 => x"0b84050c",
  2617 => x"76101010",
  2618 => x"80ebc405",
  2619 => x"88110859",
  2620 => x"5b5e5153",
  2621 => x"fee13980",
  2622 => x"eb880817",
  2623 => x"58800876",
  2624 => x"2e818d38",
  2625 => x"80ebb808",
  2626 => x"ff2e83ec",
  2627 => x"38737631",
  2628 => x"1880eb88",
  2629 => x"0c738706",
  2630 => x"70575372",
  2631 => x"802e8838",
  2632 => x"88733170",
  2633 => x"15555676",
  2634 => x"149fff06",
  2635 => x"a0807131",
  2636 => x"1770547f",
  2637 => x"53575383",
  2638 => x"d53f8008",
  2639 => x"538008ff",
  2640 => x"2e81a038",
  2641 => x"80eb8808",
  2642 => x"167080eb",
  2643 => x"880c7475",
  2644 => x"80ebc40b",
  2645 => x"88050c74",
  2646 => x"76311870",
  2647 => x"81075155",
  2648 => x"56587b80",
  2649 => x"ebc42e83",
  2650 => x"9c38798f",
  2651 => x"2682cb38",
  2652 => x"810b8415",
  2653 => x"0c841508",
  2654 => x"fc06707a",
  2655 => x"317a7226",
  2656 => x"8f722507",
  2657 => x"52555372",
  2658 => x"802efcf9",
  2659 => x"3880db39",
  2660 => x"80089fff",
  2661 => x"065372fe",
  2662 => x"eb387780",
  2663 => x"eb880c80",
  2664 => x"ebc40b88",
  2665 => x"05087b18",
  2666 => x"81078412",
  2667 => x"0c5580eb",
  2668 => x"b4087827",
  2669 => x"86387780",
  2670 => x"ebb40c80",
  2671 => x"ebb00878",
  2672 => x"27fcac38",
  2673 => x"7780ebb0",
  2674 => x"0c841508",
  2675 => x"fc06707a",
  2676 => x"317a7226",
  2677 => x"8f722507",
  2678 => x"52555372",
  2679 => x"802efca5",
  2680 => x"38883980",
  2681 => x"745456fe",
  2682 => x"db397d51",
  2683 => x"829f3f80",
  2684 => x"0b800c8f",
  2685 => x"3d0d0473",
  2686 => x"53807424",
  2687 => x"a9387282",
  2688 => x"2c81712b",
  2689 => x"80ebc808",
  2690 => x"077080eb",
  2691 => x"c40b8405",
  2692 => x"0c5d5377",
  2693 => x"8c180c74",
  2694 => x"88180c76",
  2695 => x"88190c76",
  2696 => x"8c160cf9",
  2697 => x"b7398314",
  2698 => x"70822c81",
  2699 => x"712b80eb",
  2700 => x"c8080770",
  2701 => x"80ebc40b",
  2702 => x"84050c5e",
  2703 => x"5153d439",
  2704 => x"7b7b0653",
  2705 => x"72fca338",
  2706 => x"841a7b10",
  2707 => x"5c5af139",
  2708 => x"ff1a8111",
  2709 => x"515af7b9",
  2710 => x"39781779",
  2711 => x"81078419",
  2712 => x"0c8c1808",
  2713 => x"88190871",
  2714 => x"8c120c88",
  2715 => x"120c5970",
  2716 => x"80ebd80c",
  2717 => x"7080ebd4",
  2718 => x"0c80ebcc",
  2719 => x"0b8c120c",
  2720 => x"8c110888",
  2721 => x"120c7481",
  2722 => x"0784120c",
  2723 => x"74117571",
  2724 => x"0c5153f9",
  2725 => x"bd397517",
  2726 => x"84110881",
  2727 => x"0784120c",
  2728 => x"538c1708",
  2729 => x"88180871",
  2730 => x"8c120c88",
  2731 => x"120c587d",
  2732 => x"5180da3f",
  2733 => x"881754f5",
  2734 => x"cf397284",
  2735 => x"150cf41a",
  2736 => x"f8067084",
  2737 => x"1e088106",
  2738 => x"07841e0c",
  2739 => x"701d545b",
  2740 => x"850b8414",
  2741 => x"0c850b88",
  2742 => x"140c8f7b",
  2743 => x"27fdcf38",
  2744 => x"881c527d",
  2745 => x"5182903f",
  2746 => x"80ebc40b",
  2747 => x"88050880",
  2748 => x"eb880859",
  2749 => x"55fdb739",
  2750 => x"7780eb88",
  2751 => x"0c7380eb",
  2752 => x"b80cfc91",
  2753 => x"39728415",
  2754 => x"0cfda339",
  2755 => x"0404fd3d",
  2756 => x"0d800b80",
  2757 => x"f4840c76",
  2758 => x"5186cc3f",
  2759 => x"80085380",
  2760 => x"08ff2e88",
  2761 => x"3872800c",
  2762 => x"853d0d04",
  2763 => x"80f48408",
  2764 => x"5473802e",
  2765 => x"f0387574",
  2766 => x"710c5272",
  2767 => x"800c853d",
  2768 => x"0d04fb3d",
  2769 => x"0d777052",
  2770 => x"56c23f80",
  2771 => x"ebc40b88",
  2772 => x"05088411",
  2773 => x"08fc0670",
  2774 => x"7b319fef",
  2775 => x"05e08006",
  2776 => x"e0800556",
  2777 => x"5653a080",
  2778 => x"74249438",
  2779 => x"80527551",
  2780 => x"ff9c3f80",
  2781 => x"ebcc0815",
  2782 => x"53728008",
  2783 => x"2e8f3875",
  2784 => x"51ff8a3f",
  2785 => x"80537280",
  2786 => x"0c873d0d",
  2787 => x"04733052",
  2788 => x"7551fefa",
  2789 => x"3f8008ff",
  2790 => x"2ea83880",
  2791 => x"ebc40b88",
  2792 => x"05087575",
  2793 => x"31810784",
  2794 => x"120c5380",
  2795 => x"eb880874",
  2796 => x"3180eb88",
  2797 => x"0c7551fe",
  2798 => x"d43f810b",
  2799 => x"800c873d",
  2800 => x"0d048052",
  2801 => x"7551fec6",
  2802 => x"3f80ebc4",
  2803 => x"0b880508",
  2804 => x"80087131",
  2805 => x"56538f75",
  2806 => x"25ffa438",
  2807 => x"800880eb",
  2808 => x"b8083180",
  2809 => x"eb880c74",
  2810 => x"81078414",
  2811 => x"0c7551fe",
  2812 => x"9c3f8053",
  2813 => x"ff9039f6",
  2814 => x"3d0d7c7e",
  2815 => x"545b7280",
  2816 => x"2e828338",
  2817 => x"7a51fe84",
  2818 => x"3ff81384",
  2819 => x"110870fe",
  2820 => x"06701384",
  2821 => x"1108fc06",
  2822 => x"5d585954",
  2823 => x"5880ebcc",
  2824 => x"08752e82",
  2825 => x"de387884",
  2826 => x"160c8073",
  2827 => x"8106545a",
  2828 => x"727a2e81",
  2829 => x"d5387815",
  2830 => x"84110881",
  2831 => x"06515372",
  2832 => x"a0387817",
  2833 => x"577981e6",
  2834 => x"38881508",
  2835 => x"537280eb",
  2836 => x"cc2e82f9",
  2837 => x"388c1508",
  2838 => x"708c150c",
  2839 => x"7388120c",
  2840 => x"56768107",
  2841 => x"84190c76",
  2842 => x"1877710c",
  2843 => x"53798191",
  2844 => x"3883ff77",
  2845 => x"2781c838",
  2846 => x"76892a77",
  2847 => x"832a5653",
  2848 => x"72802ebf",
  2849 => x"3876862a",
  2850 => x"b8055584",
  2851 => x"7327b438",
  2852 => x"80db1355",
  2853 => x"947327ab",
  2854 => x"38768c2a",
  2855 => x"80ee0555",
  2856 => x"80d47327",
  2857 => x"9e38768f",
  2858 => x"2a80f705",
  2859 => x"5582d473",
  2860 => x"27913876",
  2861 => x"922a80fc",
  2862 => x"05558ad4",
  2863 => x"73278438",
  2864 => x"80fe5574",
  2865 => x"10101080",
  2866 => x"ebc40588",
  2867 => x"11085556",
  2868 => x"73762e82",
  2869 => x"b3388414",
  2870 => x"08fc0653",
  2871 => x"7673278d",
  2872 => x"38881408",
  2873 => x"5473762e",
  2874 => x"098106ea",
  2875 => x"388c1408",
  2876 => x"708c1a0c",
  2877 => x"74881a0c",
  2878 => x"7888120c",
  2879 => x"56778c15",
  2880 => x"0c7a51fc",
  2881 => x"883f8c3d",
  2882 => x"0d047708",
  2883 => x"78713159",
  2884 => x"77058819",
  2885 => x"08545772",
  2886 => x"80ebcc2e",
  2887 => x"80e0388c",
  2888 => x"1808708c",
  2889 => x"150c7388",
  2890 => x"120c56fe",
  2891 => x"89398815",
  2892 => x"088c1608",
  2893 => x"708c130c",
  2894 => x"5788170c",
  2895 => x"fea33976",
  2896 => x"832a7054",
  2897 => x"55807524",
  2898 => x"81983872",
  2899 => x"822c8171",
  2900 => x"2b80ebc8",
  2901 => x"080780eb",
  2902 => x"c40b8405",
  2903 => x"0c537410",
  2904 => x"101080eb",
  2905 => x"c4058811",
  2906 => x"08555675",
  2907 => x"8c190c73",
  2908 => x"88190c77",
  2909 => x"88170c77",
  2910 => x"8c150cff",
  2911 => x"8439815a",
  2912 => x"fdb43978",
  2913 => x"17738106",
  2914 => x"54577298",
  2915 => x"38770878",
  2916 => x"71315977",
  2917 => x"058c1908",
  2918 => x"881a0871",
  2919 => x"8c120c88",
  2920 => x"120c5757",
  2921 => x"76810784",
  2922 => x"190c7780",
  2923 => x"ebc40b88",
  2924 => x"050c80eb",
  2925 => x"c0087726",
  2926 => x"fec73880",
  2927 => x"ebbc0852",
  2928 => x"7a51fafe",
  2929 => x"3f7a51fa",
  2930 => x"c43ffeba",
  2931 => x"3981788c",
  2932 => x"150c7888",
  2933 => x"150c738c",
  2934 => x"1a0c7388",
  2935 => x"1a0c5afd",
  2936 => x"80398315",
  2937 => x"70822c81",
  2938 => x"712b80eb",
  2939 => x"c8080780",
  2940 => x"ebc40b84",
  2941 => x"050c5153",
  2942 => x"74101010",
  2943 => x"80ebc405",
  2944 => x"88110855",
  2945 => x"56fee439",
  2946 => x"74538075",
  2947 => x"24a73872",
  2948 => x"822c8171",
  2949 => x"2b80ebc8",
  2950 => x"080780eb",
  2951 => x"c40b8405",
  2952 => x"0c53758c",
  2953 => x"190c7388",
  2954 => x"190c7788",
  2955 => x"170c778c",
  2956 => x"150cfdcd",
  2957 => x"39831570",
  2958 => x"822c8171",
  2959 => x"2b80ebc8",
  2960 => x"080780eb",
  2961 => x"c40b8405",
  2962 => x"0c5153d6",
  2963 => x"39810b80",
  2964 => x"0c04803d",
  2965 => x"0d72812e",
  2966 => x"8938800b",
  2967 => x"800c823d",
  2968 => x"0d047351",
  2969 => x"80f83ffe",
  2970 => x"3d0d80f3",
  2971 => x"f4085170",
  2972 => x"8a3880f4",
  2973 => x"887080f3",
  2974 => x"f40c5170",
  2975 => x"75125252",
  2976 => x"ff537087",
  2977 => x"fb808026",
  2978 => x"88387080",
  2979 => x"f3f40c71",
  2980 => x"5372800c",
  2981 => x"843d0d04",
  2982 => x"fd3d0d80",
  2983 => x"0b80e3e4",
  2984 => x"08545472",
  2985 => x"812e9c38",
  2986 => x"7380f3f8",
  2987 => x"0cffabb0",
  2988 => x"3fffaacc",
  2989 => x"3f80f3cc",
  2990 => x"528151d7",
  2991 => x"ed3f8008",
  2992 => x"51a23f72",
  2993 => x"80f3f80c",
  2994 => x"ffab953f",
  2995 => x"ffaab13f",
  2996 => x"80f3cc52",
  2997 => x"8151d7d2",
  2998 => x"3f800851",
  2999 => x"873f00ff",
  3000 => x"3900ff39",
  3001 => x"f73d0d7b",
  3002 => x"80e48808",
  3003 => x"82c81108",
  3004 => x"5a545a77",
  3005 => x"802e80da",
  3006 => x"38818818",
  3007 => x"841908ff",
  3008 => x"0581712b",
  3009 => x"59555980",
  3010 => x"742480ea",
  3011 => x"38807424",
  3012 => x"b5387382",
  3013 => x"2b781188",
  3014 => x"05565681",
  3015 => x"80190877",
  3016 => x"06537280",
  3017 => x"2eb63878",
  3018 => x"16700853",
  3019 => x"53795174",
  3020 => x"0853722d",
  3021 => x"ff14fc17",
  3022 => x"fc177981",
  3023 => x"2c5a5757",
  3024 => x"54738025",
  3025 => x"d6387708",
  3026 => x"5877ffad",
  3027 => x"3880e488",
  3028 => x"0853bc13",
  3029 => x"08a53879",
  3030 => x"51ff833f",
  3031 => x"74085372",
  3032 => x"2dff14fc",
  3033 => x"17fc1779",
  3034 => x"812c5a57",
  3035 => x"57547380",
  3036 => x"25ffa838",
  3037 => x"d1398057",
  3038 => x"ff933972",
  3039 => x"51bc1308",
  3040 => x"53722d79",
  3041 => x"51fed73f",
  3042 => x"ff3d0d80",
  3043 => x"f3d40bfc",
  3044 => x"05700852",
  3045 => x"5270ff2e",
  3046 => x"9138702d",
  3047 => x"fc127008",
  3048 => x"525270ff",
  3049 => x"2e098106",
  3050 => x"f138833d",
  3051 => x"0d0404ff",
  3052 => x"aa9b3f04",
  3053 => x"00000040",
  3054 => x"30782020",
  3055 => x"20202020",
  3056 => x"20200000",
  3057 => x"0a677265",
  3058 => x"74682072",
  3059 => x"65676973",
  3060 => x"74657273",
  3061 => x"3a000000",
  3062 => x"0a636f6e",
  3063 => x"74726f6c",
  3064 => x"3a202020",
  3065 => x"20202000",
  3066 => x"0a737461",
  3067 => x"7475733a",
  3068 => x"20202020",
  3069 => x"20202000",
  3070 => x"0a6d6163",
  3071 => x"5f6d7362",
  3072 => x"3a202020",
  3073 => x"20202000",
  3074 => x"0a6d6163",
  3075 => x"5f6c7362",
  3076 => x"3a202020",
  3077 => x"20202000",
  3078 => x"0a6d6469",
  3079 => x"6f5f636f",
  3080 => x"6e74726f",
  3081 => x"6c3a2000",
  3082 => x"0a74785f",
  3083 => x"706f696e",
  3084 => x"7465723a",
  3085 => x"20202000",
  3086 => x"0a72785f",
  3087 => x"706f696e",
  3088 => x"7465723a",
  3089 => x"20202000",
  3090 => x"0a656463",
  3091 => x"6c5f6970",
  3092 => x"3a202020",
  3093 => x"20202000",
  3094 => x"0a686173",
  3095 => x"685f6d73",
  3096 => x"623a2020",
  3097 => x"20202000",
  3098 => x"0a686173",
  3099 => x"685f6c73",
  3100 => x"623a2020",
  3101 => x"20202000",
  3102 => x"0a677265",
  3103 => x"74682d3e",
  3104 => x"636f6e74",
  3105 => x"726f6c20",
  3106 => x"3a000000",
  3107 => x"0a677265",
  3108 => x"74682d3e",
  3109 => x"73746174",
  3110 => x"75732020",
  3111 => x"3a000000",
  3112 => x"0a646573",
  3113 => x"63722d3e",
  3114 => x"636f6e74",
  3115 => x"726f6c20",
  3116 => x"3a000000",
  3117 => x"0a0a0000",
  3118 => x"74657374",
  3119 => x"2e632000",
  3120 => x"286f6e20",
  3121 => x"73696d75",
  3122 => x"6c61746f",
  3123 => x"72290a00",
  3124 => x"636f6d70",
  3125 => x"696c6564",
  3126 => x"3a204175",
  3127 => x"67203139",
  3128 => x"20323031",
  3129 => x"30202031",
  3130 => x"363a3337",
  3131 => x"3a34390a",
  3132 => x"00000000",
  3133 => x"286f6e20",
  3134 => x"68617264",
  3135 => x"77617265",
  3136 => x"290a0000",
  3137 => x"00000bf9",
  3138 => x"00000c1f",
  3139 => x"00000c1f",
  3140 => x"00000bf9",
  3141 => x"00000c1f",
  3142 => x"00000c1f",
  3143 => x"00000c1f",
  3144 => x"00000c1f",
  3145 => x"00000c1f",
  3146 => x"00000c1f",
  3147 => x"00000c1f",
  3148 => x"00000c1f",
  3149 => x"00000c1f",
  3150 => x"00000c1f",
  3151 => x"00000c1f",
  3152 => x"00000c1f",
  3153 => x"00000c1f",
  3154 => x"00000c1f",
  3155 => x"00000c1f",
  3156 => x"00000c1f",
  3157 => x"00000c1f",
  3158 => x"00000c1f",
  3159 => x"00000c1f",
  3160 => x"00000c1f",
  3161 => x"00000c1f",
  3162 => x"00000c1f",
  3163 => x"00000c1f",
  3164 => x"00000c1f",
  3165 => x"00000c1f",
  3166 => x"00000c1f",
  3167 => x"00000c1f",
  3168 => x"00000c1f",
  3169 => x"00000c1f",
  3170 => x"00000c1f",
  3171 => x"00000c1f",
  3172 => x"00000c1f",
  3173 => x"00000c1f",
  3174 => x"00000c1f",
  3175 => x"00000ccb",
  3176 => x"00000cc3",
  3177 => x"00000cbb",
  3178 => x"00000cb3",
  3179 => x"00000cab",
  3180 => x"00000ca3",
  3181 => x"00000c9b",
  3182 => x"00000c92",
  3183 => x"00000c89",
  3184 => x"43000000",
  3185 => x"64756d6d",
  3186 => x"792e6578",
  3187 => x"65000000",
  3188 => x"00ffffff",
  3189 => x"ff00ffff",
  3190 => x"ffff00ff",
  3191 => x"ffffff00",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00000000",
  3195 => x"000039dc",
  3196 => x"80000c00",
  3197 => x"80000800",
  3198 => x"80000600",
  3199 => x"80000200",
  3200 => x"80000100",
  3201 => x"00000040",
  3202 => x"0000320c",
  3203 => x"00000000",
  3204 => x"00003474",
  3205 => x"000034d0",
  3206 => x"0000352c",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"000031c0",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"00000000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000001",
  3246 => x"330eabcd",
  3247 => x"1234e66d",
  3248 => x"deec0005",
  3249 => x"000b0000",
  3250 => x"00000000",
  3251 => x"00000000",
  3252 => x"00000000",
  3253 => x"00000000",
  3254 => x"00000000",
  3255 => x"00000000",
  3256 => x"00000000",
  3257 => x"00000000",
  3258 => x"00000000",
  3259 => x"00000000",
  3260 => x"00000000",
  3261 => x"00000000",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00000000",
  3265 => x"00000000",
  3266 => x"00000000",
  3267 => x"00000000",
  3268 => x"00000000",
  3269 => x"00000000",
  3270 => x"00000000",
  3271 => x"00000000",
  3272 => x"00000000",
  3273 => x"00000000",
  3274 => x"00000000",
  3275 => x"00000000",
  3276 => x"00000000",
  3277 => x"00000000",
  3278 => x"00000000",
  3279 => x"00000000",
  3280 => x"00000000",
  3281 => x"00000000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"00000000",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00000000",
  3288 => x"00000000",
  3289 => x"00000000",
  3290 => x"00000000",
  3291 => x"00000000",
  3292 => x"00000000",
  3293 => x"00000000",
  3294 => x"00000000",
  3295 => x"00000000",
  3296 => x"00000000",
  3297 => x"00000000",
  3298 => x"00000000",
  3299 => x"00000000",
  3300 => x"00000000",
  3301 => x"00000000",
  3302 => x"00000000",
  3303 => x"00000000",
  3304 => x"00000000",
  3305 => x"00000000",
  3306 => x"00000000",
  3307 => x"00000000",
  3308 => x"00000000",
  3309 => x"00000000",
  3310 => x"00000000",
  3311 => x"00000000",
  3312 => x"00000000",
  3313 => x"00000000",
  3314 => x"00000000",
  3315 => x"00000000",
  3316 => x"00000000",
  3317 => x"00000000",
  3318 => x"00000000",
  3319 => x"00000000",
  3320 => x"00000000",
  3321 => x"00000000",
  3322 => x"00000000",
  3323 => x"00000000",
  3324 => x"00000000",
  3325 => x"00000000",
  3326 => x"00000000",
  3327 => x"00000000",
  3328 => x"00000000",
  3329 => x"00000000",
  3330 => x"00000000",
  3331 => x"00000000",
  3332 => x"00000000",
  3333 => x"00000000",
  3334 => x"00000000",
  3335 => x"00000000",
  3336 => x"00000000",
  3337 => x"00000000",
  3338 => x"00000000",
  3339 => x"00000000",
  3340 => x"00000000",
  3341 => x"00000000",
  3342 => x"00000000",
  3343 => x"00000000",
  3344 => x"00000000",
  3345 => x"00000000",
  3346 => x"00000000",
  3347 => x"00000000",
  3348 => x"00000000",
  3349 => x"00000000",
  3350 => x"00000000",
  3351 => x"00000000",
  3352 => x"00000000",
  3353 => x"00000000",
  3354 => x"00000000",
  3355 => x"00000000",
  3356 => x"00000000",
  3357 => x"00000000",
  3358 => x"00000000",
  3359 => x"00000000",
  3360 => x"00000000",
  3361 => x"00000000",
  3362 => x"00000000",
  3363 => x"00000000",
  3364 => x"00000000",
  3365 => x"00000000",
  3366 => x"00000000",
  3367 => x"00000000",
  3368 => x"00000000",
  3369 => x"00000000",
  3370 => x"00000000",
  3371 => x"00000000",
  3372 => x"00000000",
  3373 => x"00000000",
  3374 => x"00000000",
  3375 => x"00000000",
  3376 => x"00000000",
  3377 => x"00000000",
  3378 => x"00000000",
  3379 => x"00000000",
  3380 => x"00000000",
  3381 => x"00000000",
  3382 => x"00000000",
  3383 => x"00000000",
  3384 => x"00000000",
  3385 => x"00000000",
  3386 => x"00000000",
  3387 => x"00000000",
  3388 => x"00000000",
  3389 => x"00000000",
  3390 => x"00000000",
  3391 => x"00000000",
  3392 => x"00000000",
  3393 => x"00000000",
  3394 => x"00000000",
  3395 => x"00000000",
  3396 => x"00000000",
  3397 => x"00000000",
  3398 => x"00000000",
  3399 => x"00000000",
  3400 => x"00000000",
  3401 => x"00000000",
  3402 => x"00000000",
  3403 => x"00000000",
  3404 => x"00000000",
  3405 => x"00000000",
  3406 => x"00000000",
  3407 => x"00000000",
  3408 => x"00000000",
  3409 => x"00000000",
  3410 => x"00000000",
  3411 => x"00000000",
  3412 => x"00000000",
  3413 => x"00000000",
  3414 => x"00000000",
  3415 => x"00000000",
  3416 => x"00000000",
  3417 => x"00000000",
  3418 => x"00000000",
  3419 => x"00000000",
  3420 => x"00000000",
  3421 => x"00000000",
  3422 => x"00000000",
  3423 => x"00000000",
  3424 => x"00000000",
  3425 => x"00000000",
  3426 => x"00000000",
  3427 => x"00000000",
  3428 => x"00000000",
  3429 => x"00000000",
  3430 => x"00000000",
  3431 => x"00000000",
  3432 => x"00000000",
  3433 => x"00000000",
  3434 => x"00000000",
  3435 => x"00000000",
  3436 => x"00000000",
  3437 => x"00000000",
  3438 => x"ffffffff",
  3439 => x"00000000",
  3440 => x"00020000",
  3441 => x"00000000",
  3442 => x"00000000",
  3443 => x"000035c4",
  3444 => x"000035c4",
  3445 => x"000035cc",
  3446 => x"000035cc",
  3447 => x"000035d4",
  3448 => x"000035d4",
  3449 => x"000035dc",
  3450 => x"000035dc",
  3451 => x"000035e4",
  3452 => x"000035e4",
  3453 => x"000035ec",
  3454 => x"000035ec",
  3455 => x"000035f4",
  3456 => x"000035f4",
  3457 => x"000035fc",
  3458 => x"000035fc",
  3459 => x"00003604",
  3460 => x"00003604",
  3461 => x"0000360c",
  3462 => x"0000360c",
  3463 => x"00003614",
  3464 => x"00003614",
  3465 => x"0000361c",
  3466 => x"0000361c",
  3467 => x"00003624",
  3468 => x"00003624",
  3469 => x"0000362c",
  3470 => x"0000362c",
  3471 => x"00003634",
  3472 => x"00003634",
  3473 => x"0000363c",
  3474 => x"0000363c",
  3475 => x"00003644",
  3476 => x"00003644",
  3477 => x"0000364c",
  3478 => x"0000364c",
  3479 => x"00003654",
  3480 => x"00003654",
  3481 => x"0000365c",
  3482 => x"0000365c",
  3483 => x"00003664",
  3484 => x"00003664",
  3485 => x"0000366c",
  3486 => x"0000366c",
  3487 => x"00003674",
  3488 => x"00003674",
  3489 => x"0000367c",
  3490 => x"0000367c",
  3491 => x"00003684",
  3492 => x"00003684",
  3493 => x"0000368c",
  3494 => x"0000368c",
  3495 => x"00003694",
  3496 => x"00003694",
  3497 => x"0000369c",
  3498 => x"0000369c",
  3499 => x"000036a4",
  3500 => x"000036a4",
  3501 => x"000036ac",
  3502 => x"000036ac",
  3503 => x"000036b4",
  3504 => x"000036b4",
  3505 => x"000036bc",
  3506 => x"000036bc",
  3507 => x"000036c4",
  3508 => x"000036c4",
  3509 => x"000036cc",
  3510 => x"000036cc",
  3511 => x"000036d4",
  3512 => x"000036d4",
  3513 => x"000036dc",
  3514 => x"000036dc",
  3515 => x"000036e4",
  3516 => x"000036e4",
  3517 => x"000036ec",
  3518 => x"000036ec",
  3519 => x"000036f4",
  3520 => x"000036f4",
  3521 => x"000036fc",
  3522 => x"000036fc",
  3523 => x"00003704",
  3524 => x"00003704",
  3525 => x"0000370c",
  3526 => x"0000370c",
  3527 => x"00003714",
  3528 => x"00003714",
  3529 => x"0000371c",
  3530 => x"0000371c",
  3531 => x"00003724",
  3532 => x"00003724",
  3533 => x"0000372c",
  3534 => x"0000372c",
  3535 => x"00003734",
  3536 => x"00003734",
  3537 => x"0000373c",
  3538 => x"0000373c",
  3539 => x"00003744",
  3540 => x"00003744",
  3541 => x"0000374c",
  3542 => x"0000374c",
  3543 => x"00003754",
  3544 => x"00003754",
  3545 => x"0000375c",
  3546 => x"0000375c",
  3547 => x"00003764",
  3548 => x"00003764",
  3549 => x"0000376c",
  3550 => x"0000376c",
  3551 => x"00003774",
  3552 => x"00003774",
  3553 => x"0000377c",
  3554 => x"0000377c",
  3555 => x"00003784",
  3556 => x"00003784",
  3557 => x"0000378c",
  3558 => x"0000378c",
  3559 => x"00003794",
  3560 => x"00003794",
  3561 => x"0000379c",
  3562 => x"0000379c",
  3563 => x"000037a4",
  3564 => x"000037a4",
  3565 => x"000037ac",
  3566 => x"000037ac",
  3567 => x"000037b4",
  3568 => x"000037b4",
  3569 => x"000037bc",
  3570 => x"000037bc",
  3571 => x"000037c4",
  3572 => x"000037c4",
  3573 => x"000037cc",
  3574 => x"000037cc",
  3575 => x"000037d4",
  3576 => x"000037d4",
  3577 => x"000037dc",
  3578 => x"000037dc",
  3579 => x"000037e4",
  3580 => x"000037e4",
  3581 => x"000037ec",
  3582 => x"000037ec",
  3583 => x"000037f4",
  3584 => x"000037f4",
  3585 => x"000037fc",
  3586 => x"000037fc",
  3587 => x"00003804",
  3588 => x"00003804",
  3589 => x"0000380c",
  3590 => x"0000380c",
  3591 => x"00003814",
  3592 => x"00003814",
  3593 => x"0000381c",
  3594 => x"0000381c",
  3595 => x"00003824",
  3596 => x"00003824",
  3597 => x"0000382c",
  3598 => x"0000382c",
  3599 => x"00003834",
  3600 => x"00003834",
  3601 => x"0000383c",
  3602 => x"0000383c",
  3603 => x"00003844",
  3604 => x"00003844",
  3605 => x"0000384c",
  3606 => x"0000384c",
  3607 => x"00003854",
  3608 => x"00003854",
  3609 => x"0000385c",
  3610 => x"0000385c",
  3611 => x"00003864",
  3612 => x"00003864",
  3613 => x"0000386c",
  3614 => x"0000386c",
  3615 => x"00003874",
  3616 => x"00003874",
  3617 => x"0000387c",
  3618 => x"0000387c",
  3619 => x"00003884",
  3620 => x"00003884",
  3621 => x"0000388c",
  3622 => x"0000388c",
  3623 => x"00003894",
  3624 => x"00003894",
  3625 => x"0000389c",
  3626 => x"0000389c",
  3627 => x"000038a4",
  3628 => x"000038a4",
  3629 => x"000038ac",
  3630 => x"000038ac",
  3631 => x"000038b4",
  3632 => x"000038b4",
  3633 => x"000038bc",
  3634 => x"000038bc",
  3635 => x"000038c4",
  3636 => x"000038c4",
  3637 => x"000038cc",
  3638 => x"000038cc",
  3639 => x"000038d4",
  3640 => x"000038d4",
  3641 => x"000038dc",
  3642 => x"000038dc",
  3643 => x"000038e4",
  3644 => x"000038e4",
  3645 => x"000038ec",
  3646 => x"000038ec",
  3647 => x"000038f4",
  3648 => x"000038f4",
  3649 => x"000038fc",
  3650 => x"000038fc",
  3651 => x"00003904",
  3652 => x"00003904",
  3653 => x"0000390c",
  3654 => x"0000390c",
  3655 => x"00003914",
  3656 => x"00003914",
  3657 => x"0000391c",
  3658 => x"0000391c",
  3659 => x"00003924",
  3660 => x"00003924",
  3661 => x"0000392c",
  3662 => x"0000392c",
  3663 => x"00003934",
  3664 => x"00003934",
  3665 => x"0000393c",
  3666 => x"0000393c",
  3667 => x"00003944",
  3668 => x"00003944",
  3669 => x"0000394c",
  3670 => x"0000394c",
  3671 => x"00003954",
  3672 => x"00003954",
  3673 => x"0000395c",
  3674 => x"0000395c",
  3675 => x"00003964",
  3676 => x"00003964",
  3677 => x"0000396c",
  3678 => x"0000396c",
  3679 => x"00003974",
  3680 => x"00003974",
  3681 => x"0000397c",
  3682 => x"0000397c",
  3683 => x"00003984",
  3684 => x"00003984",
  3685 => x"0000398c",
  3686 => x"0000398c",
  3687 => x"00003994",
  3688 => x"00003994",
  3689 => x"0000399c",
  3690 => x"0000399c",
  3691 => x"000039a4",
  3692 => x"000039a4",
  3693 => x"000039ac",
  3694 => x"000039ac",
  3695 => x"000039b4",
  3696 => x"000039b4",
  3697 => x"000039bc",
  3698 => x"000039bc",
  3699 => x"000031c4",
  3700 => x"ffffffff",
  3701 => x"00000000",
  3702 => x"ffffffff",
  3703 => x"00000000",
  3704 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
