library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


library zylin;
use zylin.zpu_config.all;
use zylin.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"800b0b0b",
1 => x"0b0b8070",
2 => x"0b0b818a",
3 => x"880c3a0b",
4 => x"0b80fae8",
5 => x"04000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"80fbba2d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"530b0b51",
38 => x"04000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"0b0b5104",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"530b0b51",
55 => x"04000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"0b0b5104",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"72728072",
73 => x"8106ff05",
74 => x"09720605",
75 => x"71105272",
76 => x"0a100a53",
77 => x"0b0b72eb",
78 => x"38515153",
79 => x"0b0b5104",
80 => x"720a722b",
81 => x"0a530b0b",
82 => x"51040000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"0607530b",
101 => x"0b510400",
102 => x"00000000",
103 => x"00000000",
104 => x"7171530b",
105 => x"0b510406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"0b0b5104",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"530b0b51",
125 => x"04000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"0505530b",
138 => x"0b510400",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07530b0b",
147 => x"51040000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b8189",
162 => x"f4738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88ac0400",
166 => x"00000000",
167 => x"00000000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0b8f",
171 => x"e42d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0b91",
179 => x"9c2d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70540b0b",
188 => x"71067309",
189 => x"727405ff",
190 => x"05060751",
191 => x"51510400",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"0570540b",
196 => x"0b710673",
197 => x"09727405",
198 => x"ff050607",
199 => x"51515104",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"818a840c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"0571530b",
250 => x"0b510400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83cd3f80",
257 => x"fd803f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"0b0b5104",
267 => x"7381ff06",
268 => x"73830609",
269 => x"81058305",
270 => x"1010102b",
271 => x"0772fc06",
272 => x"0c515104",
273 => x"3c047070",
274 => x"0b0b819a",
275 => x"90085284",
276 => x"0b720508",
277 => x"70810651",
278 => x"510b0b70",
279 => x"f2387108",
280 => x"81ff0680",
281 => x"0c505004",
282 => x"70700b0b",
283 => x"819a9008",
284 => x"52840b72",
285 => x"0508700a",
286 => x"100a7081",
287 => x"06515151",
288 => x"0b0b70ed",
289 => x"3873720c",
290 => x"50500481",
291 => x"8a840880",
292 => x"2ea83883",
293 => x"80800b0b",
294 => x"0b819a90",
295 => x"0c82a080",
296 => x"0b0b0b81",
297 => x"9a940c82",
298 => x"90800b81",
299 => x"9aa40c0b",
300 => x"0b819a98",
301 => x"0b819aa8",
302 => x"0c04f880",
303 => x"8080a40b",
304 => x"0b0b819a",
305 => x"900cf880",
306 => x"8082800b",
307 => x"0b0b819a",
308 => x"940cf880",
309 => x"8084800b",
310 => x"819aa40c",
311 => x"f8808080",
312 => x"940b819a",
313 => x"a80cf880",
314 => x"80809c0b",
315 => x"819aa00c",
316 => x"f8808080",
317 => x"a00b819a",
318 => x"ac0c04f2",
319 => x"3d0d600b",
320 => x"0b819a94",
321 => x"08565d82",
322 => x"750c8059",
323 => x"805a800b",
324 => x"8f3d7110",
325 => x"10177008",
326 => x"5a575d5b",
327 => x"807781ff",
328 => x"067c832b",
329 => x"5658520b",
330 => x"76530b0b",
331 => x"7b5183ae",
332 => x"3f7d7f7a",
333 => x"72077c72",
334 => x"07717160",
335 => x"8105415f",
336 => x"5d5b5957",
337 => x"557a8724",
338 => x"bf380b0b",
339 => x"819a9408",
340 => x"7b101071",
341 => x"05700859",
342 => x"51558077",
343 => x"81ff067c",
344 => x"832b5658",
345 => x"520b7653",
346 => x"0b0b7b51",
347 => x"82f03f7d",
348 => x"7f7a7207",
349 => x"7c720771",
350 => x"71608105",
351 => x"415f5d5b",
352 => x"59575587",
353 => x"7b25c338",
354 => x"767d0c77",
355 => x"841e0c7c",
356 => x"800c903d",
357 => x"0d047070",
358 => x"819a9c33",
359 => x"510b0b70",
360 => x"aa38818a",
361 => x"90087008",
362 => x"52520b70",
363 => x"802e9638",
364 => x"84720581",
365 => x"8a900c70",
366 => x"2d818a90",
367 => x"08700852",
368 => x"520b70ec",
369 => x"38810b81",
370 => x"9a9c3450",
371 => x"50040470",
372 => x"0b0b819a",
373 => x"8c08802e",
374 => x"8e380b0b",
375 => x"0b0b800b",
376 => x"802e0981",
377 => x"06833850",
378 => x"040b0b81",
379 => x"9a8c510b",
380 => x"0b0bf48c",
381 => x"3f500404",
382 => x"8c08028c",
383 => x"0cfa3d0d",
384 => x"800b8c08",
385 => x"fc050c8c",
386 => x"08fc0508",
387 => x"892481b9",
388 => x"388c08f0",
389 => x"05705253",
390 => x"0b0bfddf",
391 => x"3f8c08f4",
392 => x"05088c08",
393 => x"f8050c8c",
394 => x"08f80508",
395 => x"520b0b81",
396 => x"85b45187",
397 => x"c53f0b0b",
398 => x"8185c051",
399 => x"8a8b3f0b",
400 => x"0b8185d0",
401 => x"518a823f",
402 => x"fc0b819a",
403 => x"b00c819a",
404 => x"b008812c",
405 => x"530b0b72",
406 => x"fe2e8438",
407 => x"87903f8a",
408 => x"0b819ab4",
409 => x"0c819ab4",
410 => x"08819ab0",
411 => x"0829530b",
412 => x"0b72d82e",
413 => x"843886f6",
414 => x"3f8a0b81",
415 => x"9ab00c84",
416 => x"e2ad800b",
417 => x"819ab40c",
418 => x"819ab408",
419 => x"819ab008",
420 => x"29530b0b",
421 => x"72afd7c2",
422 => x"802e8438",
423 => x"86d03f81",
424 => x"0a0b819a",
425 => x"b00cff0b",
426 => x"819ab40c",
427 => x"819ab408",
428 => x"819ab008",
429 => x"25843886",
430 => x"b53f8c08",
431 => x"fc050881",
432 => x"058c08fc",
433 => x"050cfebf",
434 => x"398c08fc",
435 => x"05088a2e",
436 => x"8438869a",
437 => x"3f72800c",
438 => x"883d0d8c",
439 => x"0c048c08",
440 => x"028c0cf5",
441 => x"3d0d8c08",
442 => x"9405089f",
443 => x"388c088c",
444 => x"05088c08",
445 => x"9005088c",
446 => x"08880508",
447 => x"5856540b",
448 => x"0b73760c",
449 => x"7484170c",
450 => x"81cd3980",
451 => x"0b8c08f0",
452 => x"050c800b",
453 => x"8c08f405",
454 => x"0c8c088c",
455 => x"05088c08",
456 => x"90050856",
457 => x"540b0b73",
458 => x"8c08f005",
459 => x"0c748c08",
460 => x"f4050c8c",
461 => x"08f8058c",
462 => x"08f00556",
463 => x"56887054",
464 => x"0b0b7553",
465 => x"0b0b7652",
466 => x"540b0b85",
467 => x"ef3fa00b",
468 => x"8c089405",
469 => x"08318c08",
470 => x"ec050c8c",
471 => x"08ec0508",
472 => x"80249f38",
473 => x"800b8c08",
474 => x"f4050c8c",
475 => x"08ec0508",
476 => x"308c08fc",
477 => x"0508712b",
478 => x"8c08f005",
479 => x"0c540b0b",
480 => x"bb398c08",
481 => x"fc05088c",
482 => x"08ec0508",
483 => x"2a8c08e8",
484 => x"050c8c08",
485 => x"fc05088c",
486 => x"08940508",
487 => x"2b8c08f4",
488 => x"050c8c08",
489 => x"f805088c",
490 => x"08940508",
491 => x"2b708c08",
492 => x"e8050807",
493 => x"8c08f005",
494 => x"0c540b0b",
495 => x"8c08f005",
496 => x"088c08f4",
497 => x"05088c08",
498 => x"88050858",
499 => x"56540b0b",
500 => x"73760c74",
501 => x"84170c8c",
502 => x"08880508",
503 => x"800c8d3d",
504 => x"0d8c0c04",
505 => x"8c08028c",
506 => x"0cf93d0d",
507 => x"800b8c08",
508 => x"fc050c8c",
509 => x"08880508",
510 => x"8025ab38",
511 => x"8c088805",
512 => x"08308c08",
513 => x"88050c80",
514 => x"0b8c08f4",
515 => x"050c8c08",
516 => x"fc050888",
517 => x"38810b8c",
518 => x"08f4050c",
519 => x"8c08f405",
520 => x"088c08fc",
521 => x"050c8c08",
522 => x"8c050880",
523 => x"25ab388c",
524 => x"088c0508",
525 => x"308c088c",
526 => x"050c800b",
527 => x"8c08f005",
528 => x"0c8c08fc",
529 => x"05088838",
530 => x"810b8c08",
531 => x"f0050c8c",
532 => x"08f00508",
533 => x"8c08fc05",
534 => x"0c80530b",
535 => x"0b8c088c",
536 => x"0508528c",
537 => x"08880508",
538 => x"5181b13f",
539 => x"8008708c",
540 => x"08f8050c",
541 => x"540b0b8c",
542 => x"08fc0508",
543 => x"802e8c38",
544 => x"8c08f805",
545 => x"08308c08",
546 => x"f8050c8c",
547 => x"08f80508",
548 => x"70800c54",
549 => x"0b0b893d",
550 => x"0d8c0c04",
551 => x"8c08028c",
552 => x"0cfb3d0d",
553 => x"800b8c08",
554 => x"fc050c8c",
555 => x"08880508",
556 => x"80259338",
557 => x"8c088805",
558 => x"08308c08",
559 => x"88050c81",
560 => x"0b8c08fc",
561 => x"050c8c08",
562 => x"8c050880",
563 => x"258c388c",
564 => x"088c0508",
565 => x"308c088c",
566 => x"050c8153",
567 => x"0b0b8c08",
568 => x"8c050852",
569 => x"8c088805",
570 => x"0851b13f",
571 => x"8008708c",
572 => x"08f8050c",
573 => x"540b0b8c",
574 => x"08fc0508",
575 => x"802e8c38",
576 => x"8c08f805",
577 => x"08308c08",
578 => x"f8050c8c",
579 => x"08f80508",
580 => x"70800c54",
581 => x"0b0b873d",
582 => x"0d8c0c04",
583 => x"8c08028c",
584 => x"0c707070",
585 => x"70810b8c",
586 => x"08fc050c",
587 => x"800b8c08",
588 => x"f8050c8c",
589 => x"088c0508",
590 => x"8c088805",
591 => x"0827ac38",
592 => x"8c08fc05",
593 => x"08802ea3",
594 => x"38800b8c",
595 => x"088c0508",
596 => x"2499388c",
597 => x"088c0508",
598 => x"108c088c",
599 => x"050c8c08",
600 => x"fc050810",
601 => x"8c08fc05",
602 => x"0cc9398c",
603 => x"08fc0508",
604 => x"802e80c9",
605 => x"388c088c",
606 => x"05088c08",
607 => x"88050826",
608 => x"a1388c08",
609 => x"8805088c",
610 => x"088c0508",
611 => x"318c0888",
612 => x"050c8c08",
613 => x"f805088c",
614 => x"08fc0508",
615 => x"078c08f8",
616 => x"050c8c08",
617 => x"fc050881",
618 => x"2a8c08fc",
619 => x"050c8c08",
620 => x"8c050881",
621 => x"2a8c088c",
622 => x"050cffaf",
623 => x"398c0890",
624 => x"0508802e",
625 => x"8f388c08",
626 => x"88050870",
627 => x"8c08f405",
628 => x"0c518d39",
629 => x"8c08f805",
630 => x"08708c08",
631 => x"f4050c51",
632 => x"8c08f405",
633 => x"08800c50",
634 => x"5050508c",
635 => x"0c047086",
636 => x"5186a03f",
637 => x"815180e7",
638 => x"be3ffc3d",
639 => x"0d873d70",
640 => x"70840552",
641 => x"0856530b",
642 => x"0b745281",
643 => x"8a940888",
644 => x"71050852",
645 => x"540b0b9f",
646 => x"e73f863d",
647 => x"0d047070",
648 => x"7070863d",
649 => x"8805530b",
650 => x"0b765275",
651 => x"88710508",
652 => x"52540b0b",
653 => x"9fca3f50",
654 => x"50505004",
655 => x"fc3d0d76",
656 => x"70797b55",
657 => x"5555558f",
658 => x"72278e38",
659 => x"72750783",
660 => x"06510b0b",
661 => x"70802eaf",
662 => x"38ff7205",
663 => x"520b0b71",
664 => x"ff2e9d38",
665 => x"72708105",
666 => x"540b0b33",
667 => x"74708105",
668 => x"5634ff72",
669 => x"05520b0b",
670 => x"71ff2e09",
671 => x"8106e538",
672 => x"74800c86",
673 => x"3d0d0474",
674 => x"51727084",
675 => x"05540b0b",
676 => x"08717084",
677 => x"05530b0b",
678 => x"0c727084",
679 => x"05540b0b",
680 => x"08717084",
681 => x"05530b0b",
682 => x"0c727084",
683 => x"05540b0b",
684 => x"08717084",
685 => x"05530b0b",
686 => x"0c727084",
687 => x"05540b0b",
688 => x"08717084",
689 => x"05530b0b",
690 => x"0cf07205",
691 => x"520b0b71",
692 => x"8f26ffb5",
693 => x"38837227",
694 => x"9c387270",
695 => x"8405540b",
696 => x"0b087170",
697 => x"8405530b",
698 => x"0b0cfc72",
699 => x"05520b0b",
700 => x"718326e6",
701 => x"3870540b",
702 => x"0bfede39",
703 => x"f73d0d7c",
704 => x"7052530b",
705 => x"0b858c3f",
706 => x"72540b0b",
707 => x"80085581",
708 => x"85e05681",
709 => x"57800881",
710 => x"055a8b3d",
711 => x"e4710559",
712 => x"530b0b82",
713 => x"59f47305",
714 => x"527b8871",
715 => x"05085253",
716 => x"0b0bb7ce",
717 => x"3f800830",
718 => x"70800807",
719 => x"9f2c8a07",
720 => x"800c530b",
721 => x"0b8b3d0d",
722 => x"04707073",
723 => x"52818a94",
724 => x"0851ffa8",
725 => x"3f505004",
726 => x"70707070",
727 => x"75530b0b",
728 => x"84d87305",
729 => x"08802e8d",
730 => x"3880530b",
731 => x"0b72800c",
732 => x"50505050",
733 => x"04818052",
734 => x"725180c1",
735 => x"cc3f8008",
736 => x"84d8140c",
737 => x"ff530b0b",
738 => x"8008802e",
739 => x"e0388008",
740 => x"540b0b9f",
741 => x"530b0b80",
742 => x"74708405",
743 => x"560cff73",
744 => x"05530b0b",
745 => x"807324c1",
746 => x"38807470",
747 => x"8405560c",
748 => x"ff730553",
749 => x"0b0b7280",
750 => x"25dd38ff",
751 => x"ac397070",
752 => x"70707577",
753 => x"55530b0b",
754 => x"9f742790",
755 => x"3896730c",
756 => x"ff520b0b",
757 => x"71800c50",
758 => x"50505004",
759 => x"84d87305",
760 => x"08520b0b",
761 => x"71802e97",
762 => x"38731010",
763 => x"72057008",
764 => x"79720c51",
765 => x"520b0b71",
766 => x"800c5050",
767 => x"50500472",
768 => x"51fed53f",
769 => x"ff528008",
770 => x"c93884d8",
771 => x"73050874",
772 => x"10107105",
773 => x"70087a72",
774 => x"0c515152",
775 => x"d839f93d",
776 => x"0d797b58",
777 => x"560b769f",
778 => x"2680f138",
779 => x"84d81608",
780 => x"540b0b73",
781 => x"802ead38",
782 => x"76101014",
783 => x"70085555",
784 => x"0b73802e",
785 => x"be388058",
786 => x"73812e8f",
787 => x"3873ff2e",
788 => x"a7388075",
789 => x"0c765173",
790 => x"2d80580b",
791 => x"0b77800c",
792 => x"893d0d04",
793 => x"7551fdf0",
794 => x"3fff5880",
795 => x"08ed3884",
796 => x"d8160854",
797 => x"0b0bc139",
798 => x"96760c81",
799 => x"0b800c89",
800 => x"3d0d0475",
801 => x"5182873f",
802 => x"76530b0b",
803 => x"80085275",
804 => x"5181be3f",
805 => x"8008800c",
806 => x"893d0d04",
807 => x"96760cff",
808 => x"0b800c89",
809 => x"3d0d04fc",
810 => x"3d0d7678",
811 => x"56530b0b",
812 => x"ff540b0b",
813 => x"749f2680",
814 => x"c13884d8",
815 => x"73050852",
816 => x"0b0b7180",
817 => x"2ebb3874",
818 => x"10107205",
819 => x"7008530b",
820 => x"0b530b0b",
821 => x"81540b0b",
822 => x"71802e9e",
823 => x"3882540b",
824 => x"0b71ff2e",
825 => x"95388354",
826 => x"0b0b7181",
827 => x"2e8c3880",
828 => x"730c7451",
829 => x"712d8054",
830 => x"0b0b7380",
831 => x"0c863d0d",
832 => x"047251fc",
833 => x"d33f8008",
834 => x"f13884d8",
835 => x"73050852",
836 => x"ffb53970",
837 => x"70735281",
838 => x"8a940851",
839 => x"fe803f50",
840 => x"50047070",
841 => x"7075530b",
842 => x"0b745281",
843 => x"8a940851",
844 => x"fd8c3f50",
845 => x"50500470",
846 => x"818a9408",
847 => x"51fc993f",
848 => x"50047070",
849 => x"7352818a",
850 => x"940851fe",
851 => x"da3f5050",
852 => x"04fc3d0d",
853 => x"800b819a",
854 => x"b80c7852",
855 => x"775180df",
856 => x"bc3f8008",
857 => x"540b0b80",
858 => x"08ff2e88",
859 => x"3873800c",
860 => x"863d0d04",
861 => x"819ab808",
862 => x"550b0b74",
863 => x"802eee38",
864 => x"7675710c",
865 => x"530b0b73",
866 => x"800c863d",
867 => x"0d0480df",
868 => x"873f0470",
869 => x"70707075",
870 => x"70718306",
871 => x"530b0b55",
872 => x"5270bf38",
873 => x"71700870",
874 => x"09f7fbfd",
875 => x"ff720506",
876 => x"70f88482",
877 => x"81800651",
878 => x"5152530b",
879 => x"0b70a138",
880 => x"84730570",
881 => x"087009f7",
882 => x"fbfdff72",
883 => x"050670f8",
884 => x"84828180",
885 => x"06515152",
886 => x"530b0b70",
887 => x"802ee138",
888 => x"72520b0b",
889 => x"7133510b",
890 => x"0b70802e",
891 => x"8c388172",
892 => x"05703352",
893 => x"520b70f6",
894 => x"38717431",
895 => x"800c5050",
896 => x"50500470",
897 => x"70707076",
898 => x"88710508",
899 => x"540b0b54",
900 => x"0b0b728d",
901 => x"38728415",
902 => x"0c72800c",
903 => x"50505050",
904 => x"04735275",
905 => x"51b1db3f",
906 => x"800b8815",
907 => x"0c800b84",
908 => x"150c8008",
909 => x"800c5050",
910 => x"505004fd",
911 => x"ad3d0d82",
912 => x"d63d0882",
913 => x"d83d0882",
914 => x"da3d0882",
915 => x"dc3d0844",
916 => x"5b454980",
917 => x"70658c05",
918 => x"2270832a",
919 => x"81327081",
920 => x"06515959",
921 => x"4947750b",
922 => x"672e0981",
923 => x"068c3863",
924 => x"90050867",
925 => x"2e098106",
926 => x"92386351",
927 => x"a2e03fff",
928 => x"56800881",
929 => x"ec38638c",
930 => x"0522570b",
931 => x"0b769a06",
932 => x"560b0b75",
933 => x"8a2ebf38",
934 => x"82c13d70",
935 => x"7182d43d",
936 => x"0c5b4380",
937 => x"0b82d43d",
938 => x"0c800b82",
939 => x"d33d0c80",
940 => x"46785b80",
941 => x"79337081",
942 => x"ff065959",
943 => x"56760b76",
944 => x"2e833881",
945 => x"5676a52e",
946 => x"81b13875",
947 => x"802e81ab",
948 => x"38811959",
949 => x"de39638e",
950 => x"05227090",
951 => x"2b575880",
952 => x"7624ffb4",
953 => x"3876fd06",
954 => x"560b0b75",
955 => x"82a33d23",
956 => x"77028405",
957 => x"89860523",
958 => x"639c0508",
959 => x"82a73d0c",
960 => x"63a40508",
961 => x"82a93d0c",
962 => x"9f3d7082",
963 => x"a13d0c82",
964 => x"a43d0c88",
965 => x"800b82a2",
966 => x"3d0c8880",
967 => x"0b82a53d",
968 => x"0c800b82",
969 => x"a63d0c60",
970 => x"530b0b78",
971 => x"52829f3d",
972 => x"70525695",
973 => x"cb3f8008",
974 => x"57800b80",
975 => x"08248e38",
976 => x"7551a39b",
977 => x"3f800880",
978 => x"2e8338ff",
979 => x"5782a23d",
980 => x"2270862a",
981 => x"70810651",
982 => x"57580b75",
983 => x"802e9038",
984 => x"638c0522",
985 => x"80c00756",
986 => x"0b0b7564",
987 => x"8c052376",
988 => x"560b0b75",
989 => x"800c82d5",
990 => x"3d0d0478",
991 => x"7b31570b",
992 => x"0b76802e",
993 => x"b1387a7a",
994 => x"0c76841b",
995 => x"0c82d33d",
996 => x"081782d4",
997 => x"3d0c881a",
998 => x"82d33d08",
999 => x"81710582",
1000 => x"d53d0c81",
1001 => x"71055157",
1002 => x"5a0b7587",
1003 => x"2480cb38",
1004 => x"65177933",
1005 => x"59460b77",
1006 => x"81ff0656",
1007 => x"0b0b7580",
1008 => x"2e93fe38",
1009 => x"81195980",
1010 => x"70714743",
1011 => x"5fff5e7e",
1012 => x"82d53d34",
1013 => x"7833580b",
1014 => x"0b7781ff",
1015 => x"06811a5a",
1016 => x"5de01d56",
1017 => x"0b0b7580",
1018 => x"d82687a1",
1019 => x"38751010",
1020 => x"81868405",
1021 => x"560b0b75",
1022 => x"080482d5",
1023 => x"3df00552",
1024 => x"6351fbff",
1025 => x"3f80088a",
1026 => x"a5386266",
1027 => x"187a335a",
1028 => x"475affa2",
1029 => x"397e9007",
1030 => x"5f0b0b7e",
1031 => x"842a7081",
1032 => x"0651560b",
1033 => x"0b7592ba",
1034 => x"387e862a",
1035 => x"70810651",
1036 => x"560b0b75",
1037 => x"802e92aa",
1038 => x"38606184",
1039 => x"05827205",
1040 => x"225a4256",
1041 => x"815c800b",
1042 => x"82d53d34",
1043 => x"7d42807e",
1044 => x"2486387e",
1045 => x"feff065f",
1046 => x"62783070",
1047 => x"7a079f2a",
1048 => x"64307066",
1049 => x"079f2a72",
1050 => x"07525951",
1051 => x"585b0b76",
1052 => x"802e918d",
1053 => x"387b812e",
1054 => x"8b9d3881",
1055 => x"7c259281",
1056 => x"387b822e",
1057 => x"8bd63881",
1058 => x"88e85b0b",
1059 => x"0b7a51fa",
1060 => x"823f8008",
1061 => x"5c0b0b7b",
1062 => x"5e7b6225",
1063 => x"8338615e",
1064 => x"82d43d33",
1065 => x"7081ff06",
1066 => x"57580b75",
1067 => x"802e90ba",
1068 => x"38811e5e",
1069 => x"7e818406",
1070 => x"400b0b7f",
1071 => x"80fa3864",
1072 => x"7e315780",
1073 => x"0b772580",
1074 => x"ef389077",
1075 => x"25b93881",
1076 => x"85e47a0c",
1077 => x"900b841b",
1078 => x"0c82d33d",
1079 => x"08900582",
1080 => x"d43d0c88",
1081 => x"1a82d33d",
1082 => x"08817105",
1083 => x"82d53d0c",
1084 => x"81710551",
1085 => x"575a0b75",
1086 => x"872485aa",
1087 => x"38f01757",
1088 => x"0b0b7690",
1089 => x"24c93881",
1090 => x"85e47a0c",
1091 => x"76841b0c",
1092 => x"82d33d08",
1093 => x"1782d43d",
1094 => x"0c881a82",
1095 => x"d33d0881",
1096 => x"710582d5",
1097 => x"3d0c8171",
1098 => x"0551575a",
1099 => x"0b758724",
1100 => x"8ff63882",
1101 => x"d43d3358",
1102 => x"0b0b7781",
1103 => x"ff06560b",
1104 => x"0b75802e",
1105 => x"86e83882",
1106 => x"d53dfc71",
1107 => x"057b0c58",
1108 => x"810b841b",
1109 => x"0c82d33d",
1110 => x"08810582",
1111 => x"d43d0c88",
1112 => x"1a82d33d",
1113 => x"08817105",
1114 => x"82d53d0c",
1115 => x"81710551",
1116 => x"575a0b75",
1117 => x"87248789",
1118 => x"387f8180",
1119 => x"2e84d738",
1120 => x"617c3157",
1121 => x"800b7725",
1122 => x"80fa3890",
1123 => x"7725b938",
1124 => x"8185f47a",
1125 => x"0c900b84",
1126 => x"1b0c82d3",
1127 => x"3d089005",
1128 => x"82d43d0c",
1129 => x"881a82d3",
1130 => x"3d088171",
1131 => x"0582d53d",
1132 => x"0c817105",
1133 => x"51575a0b",
1134 => x"75872484",
1135 => x"8138f017",
1136 => x"570b0b76",
1137 => x"9024c938",
1138 => x"8185f47a",
1139 => x"0c76841b",
1140 => x"0c82d33d",
1141 => x"081782d4",
1142 => x"3d0c881a",
1143 => x"82d33d08",
1144 => x"81710582",
1145 => x"d53d0c81",
1146 => x"71055157",
1147 => x"5a877625",
1148 => x"933882d5",
1149 => x"3df00552",
1150 => x"6351f887",
1151 => x"3f800886",
1152 => x"ad38625a",
1153 => x"7a0b7a0c",
1154 => x"7b841b0c",
1155 => x"82d33d08",
1156 => x"1c82d43d",
1157 => x"0c881a82",
1158 => x"d33d0881",
1159 => x"710582d5",
1160 => x"3d0c8171",
1161 => x"0551575a",
1162 => x"0b758724",
1163 => x"84eb387e",
1164 => x"822a7081",
1165 => x"0651560b",
1166 => x"0b75802e",
1167 => x"81813864",
1168 => x"7e315780",
1169 => x"0b772580",
1170 => x"f6389077",
1171 => x"25b93881",
1172 => x"85e47a0c",
1173 => x"900b841b",
1174 => x"0c82d33d",
1175 => x"08900582",
1176 => x"d43d0c88",
1177 => x"1a82d33d",
1178 => x"08817105",
1179 => x"82d53d0c",
1180 => x"81710551",
1181 => x"575a0b75",
1182 => x"87248485",
1183 => x"38f01757",
1184 => x"0b0b7690",
1185 => x"24c93881",
1186 => x"85e47a0c",
1187 => x"76841b0c",
1188 => x"82d33d08",
1189 => x"1782d43d",
1190 => x"0c82d23d",
1191 => x"08817105",
1192 => x"82d43d0c",
1193 => x"81710551",
1194 => x"56870b76",
1195 => x"25913882",
1196 => x"d53df005",
1197 => x"526351f6",
1198 => x"ca3f8008",
1199 => x"84f0387d",
1200 => x"567d6525",
1201 => x"83386456",
1202 => x"65164682",
1203 => x"d33d0884",
1204 => x"cb38800b",
1205 => x"82d33d0c",
1206 => x"625a6680",
1207 => x"2ef7d238",
1208 => x"6651b2d6",
1209 => x"3f80795c",
1210 => x"47f7c839",
1211 => x"7e90075f",
1212 => x"0b0b7e84",
1213 => x"2a708106",
1214 => x"51560b0b",
1215 => x"758cd538",
1216 => x"7e862a70",
1217 => x"81065156",
1218 => x"0b0b7580",
1219 => x"2e8cc538",
1220 => x"60618405",
1221 => x"82720522",
1222 => x"5a425680",
1223 => x"5c800b82",
1224 => x"d53d34fa",
1225 => x"a7397e90",
1226 => x"075f0b0b",
1227 => x"7e842a70",
1228 => x"81065156",
1229 => x"0b0b758c",
1230 => x"89387e86",
1231 => x"2a708106",
1232 => x"51560b0b",
1233 => x"75802e8b",
1234 => x"f9386061",
1235 => x"84057108",
1236 => x"902b7090",
1237 => x"2c515a42",
1238 => x"56807824",
1239 => x"89ac3881",
1240 => x"5cf9e939",
1241 => x"60618405",
1242 => x"71084742",
1243 => x"56648025",
1244 => x"f8e23864",
1245 => x"30457e84",
1246 => x"07793359",
1247 => x"5ff8d839",
1248 => x"8119597e",
1249 => x"90077933",
1250 => x"595ff8cb",
1251 => x"397c802e",
1252 => x"8caf3882",
1253 => x"b73d5b7c",
1254 => x"0b7b3481",
1255 => x"5c800b82",
1256 => x"d53d34f9",
1257 => x"f03982d5",
1258 => x"3df00552",
1259 => x"6351f4d3",
1260 => x"3f800882",
1261 => x"f93862f0",
1262 => x"18585afa",
1263 => x"c33982d5",
1264 => x"3df00552",
1265 => x"6351f4bb",
1266 => x"3f800882",
1267 => x"e13862f0",
1268 => x"18585afb",
1269 => x"ec39647e",
1270 => x"3157800b",
1271 => x"7725fba0",
1272 => x"38907725",
1273 => x"b9388185",
1274 => x"f47a0c90",
1275 => x"0b841b0c",
1276 => x"82d33d08",
1277 => x"900582d4",
1278 => x"3d0c881a",
1279 => x"82d33d08",
1280 => x"81710582",
1281 => x"d53d0c81",
1282 => x"71055157",
1283 => x"5a0b7587",
1284 => x"2480d638",
1285 => x"f017570b",
1286 => x"0b769024",
1287 => x"c9388185",
1288 => x"f47a0c76",
1289 => x"841b0c82",
1290 => x"d33d0817",
1291 => x"82d43d0c",
1292 => x"881a82d3",
1293 => x"3d088171",
1294 => x"0582d53d",
1295 => x"0c817105",
1296 => x"51575a87",
1297 => x"7625fab8",
1298 => x"3882d53d",
1299 => x"f0055263",
1300 => x"51f3b03f",
1301 => x"800881d6",
1302 => x"3862627d",
1303 => x"31585a0b",
1304 => x"768024fa",
1305 => x"a638fb9c",
1306 => x"3982d53d",
1307 => x"f0055263",
1308 => x"51f3903f",
1309 => x"800881b6",
1310 => x"3862f018",
1311 => x"585aff97",
1312 => x"3982d53d",
1313 => x"f0055263",
1314 => x"51f2f83f",
1315 => x"8008819e",
1316 => x"3862f018",
1317 => x"585afbe8",
1318 => x"3982d53d",
1319 => x"f0055263",
1320 => x"51f2e03f",
1321 => x"80088186",
1322 => x"38625afb",
1323 => x"82397e0a",
1324 => x"100a7081",
1325 => x"0651560b",
1326 => x"0b75802e",
1327 => x"f9bb38b0",
1328 => x"0b82b73d",
1329 => x"347c0284",
1330 => x"0589d505",
1331 => x"3482d53d",
1332 => x"ff84057a",
1333 => x"0c820b84",
1334 => x"1b0c82d3",
1335 => x"3d088205",
1336 => x"82d43d0c",
1337 => x"881a82d3",
1338 => x"3d088171",
1339 => x"0582d53d",
1340 => x"0c817105",
1341 => x"51575a87",
1342 => x"7625f8fd",
1343 => x"3882d53d",
1344 => x"58f01852",
1345 => x"6351f1fb",
1346 => x"3f8008a2",
1347 => x"38625a7f",
1348 => x"81802e09",
1349 => x"8106f8e8",
1350 => x"38fdbb39",
1351 => x"82d53df0",
1352 => x"05526351",
1353 => x"f1dd3f80",
1354 => x"08802efb",
1355 => x"a5386680",
1356 => x"2e863866",
1357 => x"51ae833f",
1358 => x"638c0522",
1359 => x"70862a70",
1360 => x"8106685a",
1361 => x"5157440b",
1362 => x"75802ef4",
1363 => x"a238ff56",
1364 => x"f49f3980",
1365 => x"0b82d53d",
1366 => x"34606184",
1367 => x"0571085d",
1368 => x"42567a80",
1369 => x"2e88d138",
1370 => x"7c80d32e",
1371 => x"85aa387e",
1372 => x"842a7081",
1373 => x"0651560b",
1374 => x"0b75859c",
1375 => x"38807e24",
1376 => x"f689387d",
1377 => x"530b0b75",
1378 => x"527a51ba",
1379 => x"d03f7d5c",
1380 => x"8008802e",
1381 => x"f5ff3880",
1382 => x"087b315c",
1383 => x"7d0b7c25",
1384 => x"f5f3387d",
1385 => x"5cf5ee39",
1386 => x"7e842a70",
1387 => x"81065156",
1388 => x"0b0b7587",
1389 => x"bb387e86",
1390 => x"2a708106",
1391 => x"51560b0b",
1392 => x"75802e87",
1393 => x"ab386061",
1394 => x"84057108",
1395 => x"52425665",
1396 => x"0b762378",
1397 => x"5bf1dc39",
1398 => x"78337081",
1399 => x"ff065758",
1400 => x"0b7580ec",
1401 => x"2efb9938",
1402 => x"7e900778",
1403 => x"81ff0681",
1404 => x"1b5b5e5f",
1405 => x"f3eb3960",
1406 => x"61840571",
1407 => x"085a4256",
1408 => x"820b8189",
1409 => x"84607207",
1410 => x"41495c80",
1411 => x"f85d800b",
1412 => x"82d53d34",
1413 => x"f4b63989",
1414 => x"7827a838",
1415 => x"ff1b5b8a",
1416 => x"52775180",
1417 => x"d8b43f80",
1418 => x"08b00556",
1419 => x"0b0b757b",
1420 => x"348a5277",
1421 => x"5180d7f6",
1422 => x"3f800858",
1423 => x"0b0b7789",
1424 => x"26da38ff",
1425 => x"1bb01957",
1426 => x"5b0b750b",
1427 => x"7b3482d5",
1428 => x"3d707c31",
1429 => x"ffb0055d",
1430 => x"56f4ba39",
1431 => x"ff1b788f",
1432 => x"06690557",
1433 => x"5b0b7533",
1434 => x"7b347784",
1435 => x"2a580b0b",
1436 => x"77802eda",
1437 => x"38ff1b78",
1438 => x"8f066905",
1439 => x"575b0b75",
1440 => x"337b3477",
1441 => x"842a580b",
1442 => x"0b77d138",
1443 => x"c1397e80",
1444 => x"c0077933",
1445 => x"595ff2bf",
1446 => x"3982b73d",
1447 => x"5b7c80c3",
1448 => x"2e91387e",
1449 => x"842a7081",
1450 => x"0651560b",
1451 => x"0b75802e",
1452 => x"82c83888",
1453 => x"530b0b80",
1454 => x"529d3d70",
1455 => x"5256bbcf",
1456 => x"3f75540b",
1457 => x"0b606184",
1458 => x"05710855",
1459 => x"7c540b0b",
1460 => x"6a530b0b",
1461 => x"425686e8",
1462 => x"3f80085c",
1463 => x"8008ff2e",
1464 => x"fccc3880",
1465 => x"0b82d53d",
1466 => x"34f3aa39",
1467 => x"78708105",
1468 => x"5a335d0b",
1469 => x"0b7caa2e",
1470 => x"85ef3880",
1471 => x"0bd01e71",
1472 => x"4057570b",
1473 => x"758926f1",
1474 => x"d8387610",
1475 => x"10107710",
1476 => x"057d05d0",
1477 => x"05797081",
1478 => x"055b33d0",
1479 => x"7105585e",
1480 => x"57897627",
1481 => x"e538765e",
1482 => x"76ff25f1",
1483 => x"b438ff5e",
1484 => x"f1af3981",
1485 => x"89987f84",
1486 => x"2a708106",
1487 => x"5157480b",
1488 => x"75818a38",
1489 => x"7e862a70",
1490 => x"81065156",
1491 => x"0b0b7580",
1492 => x"2e80fa38",
1493 => x"60618405",
1494 => x"82720522",
1495 => x"5a425682",
1496 => x"7f810657",
1497 => x"5c77802e",
1498 => x"f1dc3875",
1499 => x"802ef1d6",
1500 => x"387e7c07",
1501 => x"5f800b82",
1502 => x"d53d34f1",
1503 => x"cf39ab0b",
1504 => x"82d53d34",
1505 => x"783358f0",
1506 => x"ce398057",
1507 => x"0b0b7610",
1508 => x"10107710",
1509 => x"057d05d0",
1510 => x"05797081",
1511 => x"055b33d0",
1512 => x"7105585e",
1513 => x"57897627",
1514 => x"e3387645",
1515 => x"f0b3397e",
1516 => x"81800779",
1517 => x"33595ff0",
1518 => x"9e398189",
1519 => x"847f842a",
1520 => x"70810651",
1521 => x"57480b75",
1522 => x"802efef8",
1523 => x"38606184",
1524 => x"0571085a",
1525 => x"4256ff87",
1526 => x"397e8107",
1527 => x"7933595f",
1528 => x"eff53982",
1529 => x"d43d3356",
1530 => x"0b0b75ef",
1531 => x"e738a00b",
1532 => x"82d53d34",
1533 => x"783358ef",
1534 => x"de396061",
1535 => x"84054256",
1536 => x"8316337b",
1537 => x"34815cf7",
1538 => x"94397730",
1539 => x"58ad0b82",
1540 => x"d53d3481",
1541 => x"5cf0b539",
1542 => x"7a4a8070",
1543 => x"585c8853",
1544 => x"0b0b7b52",
1545 => x"9b3d7052",
1546 => x"58b8e43f",
1547 => x"7b7e2481",
1548 => x"94387610",
1549 => x"106a0556",
1550 => x"0b0b7508",
1551 => x"802eb638",
1552 => x"77540b0b",
1553 => x"7508530b",
1554 => x"0b82d53d",
1555 => x"ff880552",
1556 => x"685183ec",
1557 => x"3f8008ff",
1558 => x"2ef9d338",
1559 => x"80081c56",
1560 => x"0b0b757e",
1561 => x"248f3881",
1562 => x"17765d57",
1563 => x"757e2e09",
1564 => x"8106ffbe",
1565 => x"387b802e",
1566 => x"f09b3881",
1567 => x"1c526851",
1568 => x"a7c73f80",
1569 => x"08478008",
1570 => x"802ef9ac",
1571 => x"3888530b",
1572 => x"0b805277",
1573 => x"51b7f83f",
1574 => x"77557b54",
1575 => x"0b0b82d5",
1576 => x"3df69405",
1577 => x"530b0b66",
1578 => x"52685184",
1579 => x"8a3f8008",
1580 => x"7c2e0981",
1581 => x"06f8f738",
1582 => x"66678008",
1583 => x"05575b80",
1584 => x"7634efd1",
1585 => x"3977557b",
1586 => x"540b0b82",
1587 => x"d53df694",
1588 => x"05530b0b",
1589 => x"7b526851",
1590 => x"83dd3f80",
1591 => x"085c8008",
1592 => x"ff2ef8ca",
1593 => x"387a4aff",
1594 => x"8c397e0a",
1595 => x"100a7081",
1596 => x"0651560b",
1597 => x"0b75802e",
1598 => x"efba3882",
1599 => x"1e5eefb4",
1600 => x"397bfaca",
1601 => x"387e8106",
1602 => x"560b0b75",
1603 => x"802efabe",
1604 => x"380289ff",
1605 => x"055bb00b",
1606 => x"7b3482d5",
1607 => x"3d707c31",
1608 => x"ffb0055d",
1609 => x"56eeee39",
1610 => x"82d53df0",
1611 => x"05526351",
1612 => x"e9d13f80",
1613 => x"08f7f738",
1614 => x"6282d53d",
1615 => x"33595aef",
1616 => x"f7396061",
1617 => x"84057108",
1618 => x"5a425677",
1619 => x"8025f48f",
1620 => x"38fdb739",
1621 => x"60618405",
1622 => x"71085a42",
1623 => x"56805cf3",
1624 => x"bc396061",
1625 => x"84057108",
1626 => x"5a425681",
1627 => x"5cedd739",
1628 => x"60618405",
1629 => x"71086871",
1630 => x"0c527a5d",
1631 => x"4256eab3",
1632 => x"397bee83",
1633 => x"38ff1b78",
1634 => x"b706b007",
1635 => x"585b0b76",
1636 => x"0b7b3477",
1637 => x"832a580b",
1638 => x"0b77ea38",
1639 => x"7e810656",
1640 => x"0b0b7580",
1641 => x"2ef9a738",
1642 => x"76b02ef9",
1643 => x"a138ff1b",
1644 => x"5bb00b7b",
1645 => x"34fee339",
1646 => x"8189ac5b",
1647 => x"865cedd5",
1648 => x"3982d33d",
1649 => x"088a3880",
1650 => x"0b82d33d",
1651 => x"0cf6df39",
1652 => x"82d53df0",
1653 => x"05526351",
1654 => x"e8a93f80",
1655 => x"08f6cf38",
1656 => x"800b82d3",
1657 => x"3d0cf6c6",
1658 => x"39606184",
1659 => x"05710840",
1660 => x"42567d80",
1661 => x"25ebdd38",
1662 => x"ff793359",
1663 => x"5eebd839",
1664 => x"fc3d0d81",
1665 => x"8a940855",
1666 => x"b8150880",
1667 => x"2e973878",
1668 => x"540b0b77",
1669 => x"530b0b76",
1670 => x"52818a94",
1671 => x"0851e89b",
1672 => x"3f863d0d",
1673 => x"04745190",
1674 => x"c13f7854",
1675 => x"0b0b7753",
1676 => x"0b0b7652",
1677 => x"818a9408",
1678 => x"51e8803f",
1679 => x"863d0d04",
1680 => x"f63d0d7c",
1681 => x"7e615956",
1682 => x"58805674",
1683 => x"0b762ea0",
1684 => x"3876540b",
1685 => x"0b7e530b",
1686 => x"0b745277",
1687 => x"5182d53f",
1688 => x"80085580",
1689 => x"08ff2ea6",
1690 => x"3874800c",
1691 => x"8c3d0d04",
1692 => x"76540b0b",
1693 => x"75530b0b",
1694 => x"8c3df405",
1695 => x"52775182",
1696 => x"b33f8008",
1697 => x"558008ff",
1698 => x"2e098106",
1699 => x"dc388077",
1700 => x"0c818a78",
1701 => x"0c74800c",
1702 => x"8c3d0d04",
1703 => x"70707070",
1704 => x"77540b0b",
1705 => x"76530b0b",
1706 => x"7552818a",
1707 => x"940851ff",
1708 => x"8f3f5050",
1709 => x"505004ec",
1710 => x"3d0d6668",
1711 => x"6a6c6e73",
1712 => x"5c405d42",
1713 => x"42420b60",
1714 => x"802e819b",
1715 => x"38806008",
1716 => x"5a5d0b0b",
1717 => x"7c7a2781",
1718 => x"8338933d",
1719 => x"5b7b0884",
1720 => x"1d087d56",
1721 => x"7a08557c",
1722 => x"540b0b63",
1723 => x"530b0b40",
1724 => x"5efecd3f",
1725 => x"80085880",
1726 => x"08ff2e80",
1727 => x"fa38807a",
1728 => x"80083156",
1729 => x"567c7526",
1730 => x"83388156",
1731 => x"80087a27",
1732 => x"80da3875",
1733 => x"802e80d4",
1734 => x"3880081d",
1735 => x"5d60802e",
1736 => x"a7388056",
1737 => x"0b0b7580",
1738 => x"08259738",
1739 => x"751b550b",
1740 => x"0b743377",
1741 => x"70810559",
1742 => x"34811656",
1743 => x"770b7624",
1744 => x"eb387f08",
1745 => x"8405600c",
1746 => x"78708405",
1747 => x"5a08550b",
1748 => x"0b74802e",
1749 => x"b138797d",
1750 => x"26ff8238",
1751 => x"7c550b0b",
1752 => x"74800c96",
1753 => x"3d0d04ff",
1754 => x"5afee239",
1755 => x"7d7c0c7e",
1756 => x"841d0c7c",
1757 => x"55e83981",
1758 => x"8a620c80",
1759 => x"7c0c8008",
1760 => x"800c963d",
1761 => x"0d046080",
1762 => x"2e843874",
1763 => x"600c747c",
1764 => x"0cff1d80",
1765 => x"0c963d0d",
1766 => x"04fc3d0d",
1767 => x"79557854",
1768 => x"0b0b7753",
1769 => x"0b0b7652",
1770 => x"818a9408",
1771 => x"51fe883f",
1772 => x"863d0d04",
1773 => x"f83d0d7b",
1774 => x"7d7f8191",
1775 => x"94540b0b",
1776 => x"595755e3",
1777 => x"ce3f8008",
1778 => x"81269838",
1779 => x"74540b0b",
1780 => x"74802e88",
1781 => x"38757534",
1782 => x"81540b0b",
1783 => x"73800c8a",
1784 => x"3d0d0481",
1785 => x"89b45281",
1786 => x"919451be",
1787 => x"c93f8008",
1788 => x"81d93880",
1789 => x"08540b0b",
1790 => x"74802ee0",
1791 => x"3880ff76",
1792 => x"25d338ff",
1793 => x"8016530b",
1794 => x"0b8eff73",
1795 => x"2785b838",
1796 => x"f0801653",
1797 => x"0b0b83ef",
1798 => x"ff732782",
1799 => x"d038fc80",
1800 => x"8016530b",
1801 => x"0b80fbff",
1802 => x"ff732785",
1803 => x"c2388fff",
1804 => x"0a16530b",
1805 => x"0bf7c00a",
1806 => x"73278689",
1807 => x"38ff540b",
1808 => x"0bc00a76",
1809 => x"25ff9538",
1810 => x"75820a06",
1811 => x"709e2c70",
1812 => x"fc075151",
1813 => x"530b0b72",
1814 => x"75708105",
1815 => x"57347581",
1816 => x"fc0a0670",
1817 => x"982aff80",
1818 => x"0751530b",
1819 => x"0b727570",
1820 => x"81055734",
1821 => x"7587f080",
1822 => x"80067092",
1823 => x"2aff8007",
1824 => x"51530b0b",
1825 => x"72757081",
1826 => x"05573475",
1827 => x"8fe08006",
1828 => x"708c2aff",
1829 => x"80075153",
1830 => x"0b0b7275",
1831 => x"70810557",
1832 => x"34759fc0",
1833 => x"0670862a",
1834 => x"ff800751",
1835 => x"530b0b72",
1836 => x"75708105",
1837 => x"573475ff",
1838 => x"bf06ff80",
1839 => x"07530b0b",
1840 => x"72753486",
1841 => x"0b800c8a",
1842 => x"3d0d0481",
1843 => x"89bc5281",
1844 => x"919451bc",
1845 => x"e13f8008",
1846 => x"81f93875",
1847 => x"81ff0676",
1848 => x"882c7081",
1849 => x"ff068008",
1850 => x"5759540b",
1851 => x"0b587480",
1852 => x"2efde938",
1853 => x"76802efd",
1854 => x"d3388008",
1855 => x"80ff1870",
1856 => x"81ff0651",
1857 => x"540b0b56",
1858 => x"729e2683",
1859 => x"38815680",
1860 => x"08a01870",
1861 => x"81ff0651",
1862 => x"540b0b54",
1863 => x"0b0b728f",
1864 => x"26853881",
1865 => x"540b0b75",
1866 => x"7407530b",
1867 => x"0b72802e",
1868 => x"b4388008",
1869 => x"c019540b",
1870 => x"0b5672be",
1871 => x"26833881",
1872 => x"568008ff",
1873 => x"80197081",
1874 => x"ff065154",
1875 => x"0b0b540b",
1876 => x"0b7280fc",
1877 => x"26853881",
1878 => x"540b0b75",
1879 => x"7407530b",
1880 => x"0b7280da",
1881 => x"38ff0b80",
1882 => x"0c8a3d0d",
1883 => x"04fcd080",
1884 => x"16530b0b",
1885 => x"ff540b0b",
1886 => x"8fff7327",
1887 => x"fcde3875",
1888 => x"83e08006",
1889 => x"708c2ae0",
1890 => x"0751530b",
1891 => x"0b727570",
1892 => x"81055734",
1893 => x"759fc006",
1894 => x"70862aff",
1895 => x"80075153",
1896 => x"0b0b7275",
1897 => x"70810557",
1898 => x"3475ffbf",
1899 => x"06ff8007",
1900 => x"530b0b72",
1901 => x"7534830b",
1902 => x"800c8a3d",
1903 => x"0d047675",
1904 => x"70810557",
1905 => x"34777534",
1906 => x"82540b0b",
1907 => x"73800c8a",
1908 => x"3d0d0481",
1909 => x"89c45281",
1910 => x"919451ba",
1911 => x"d93f8008",
1912 => x"80eb3875",
1913 => x"81ff0676",
1914 => x"882c7081",
1915 => x"ff068008",
1916 => x"5759540b",
1917 => x"0b587480",
1918 => x"2efbe138",
1919 => x"76802efb",
1920 => x"cb388008",
1921 => x"530b0b81",
1922 => x"a0772785",
1923 => x"3881530b",
1924 => x"0b7681ff",
1925 => x"2efece38",
1926 => x"81707406",
1927 => x"540b0b54",
1928 => x"0b0b7280",
1929 => x"2efebe38",
1930 => x"8008530b",
1931 => x"0b81a078",
1932 => x"27853873",
1933 => x"530b0b77",
1934 => x"81ff2efe",
1935 => x"a8387274",
1936 => x"06530b0b",
1937 => x"72802efe",
1938 => x"9c38fef2",
1939 => x"398189cc",
1940 => x"52819194",
1941 => x"51b9df3f",
1942 => x"8008faf0",
1943 => x"38800876",
1944 => x"81ff0677",
1945 => x"882c7081",
1946 => x"ff065955",
1947 => x"59598154",
1948 => x"0b0b7480",
1949 => x"2efae538",
1950 => x"75802e82",
1951 => x"b438df16",
1952 => x"530b0b72",
1953 => x"80dd26fd",
1954 => x"dc38df18",
1955 => x"530b0b72",
1956 => x"80dd26fd",
1957 => x"d0387608",
1958 => x"9c387377",
1959 => x"0c9b7570",
1960 => x"81055734",
1961 => x"a4757081",
1962 => x"05573480",
1963 => x"c2757081",
1964 => x"05573483",
1965 => x"59757570",
1966 => x"81055734",
1967 => x"77753482",
1968 => x"19800c8a",
1969 => x"3d0d0475",
1970 => x"8fc00670",
1971 => x"862ac007",
1972 => x"51530b0b",
1973 => x"72757081",
1974 => x"05573475",
1975 => x"ffbf06ff",
1976 => x"8007530b",
1977 => x"0b727534",
1978 => x"82540b0b",
1979 => x"fdde3975",
1980 => x"80f08080",
1981 => x"0670922a",
1982 => x"f0075153",
1983 => x"0b0b7275",
1984 => x"70810557",
1985 => x"34758fe0",
1986 => x"8006708c",
1987 => x"2aff8007",
1988 => x"51530b0b",
1989 => x"72757081",
1990 => x"05573475",
1991 => x"9fc00670",
1992 => x"862aff80",
1993 => x"0751530b",
1994 => x"0b727570",
1995 => x"81055734",
1996 => x"75ffbf06",
1997 => x"ff800753",
1998 => x"0b0b7275",
1999 => x"34840b80",
2000 => x"0c8a3d0d",
2001 => x"047581c0",
2002 => x"0a067098",
2003 => x"2af80751",
2004 => x"530b0b72",
2005 => x"75708105",
2006 => x"57347587",
2007 => x"f0808006",
2008 => x"70922aff",
2009 => x"80075153",
2010 => x"0b0b7275",
2011 => x"70810557",
2012 => x"34758fe0",
2013 => x"8006708c",
2014 => x"2aff8007",
2015 => x"51530b0b",
2016 => x"72757081",
2017 => x"05573475",
2018 => x"9fc00670",
2019 => x"862aff80",
2020 => x"0751530b",
2021 => x"0b727570",
2022 => x"81055734",
2023 => x"75ffbf06",
2024 => x"ff800753",
2025 => x"0b0b7275",
2026 => x"34850b80",
2027 => x"0c8a3d0d",
2028 => x"04760880",
2029 => x"2e9d3880",
2030 => x"08770c9b",
2031 => x"75708105",
2032 => x"5734a875",
2033 => x"70810557",
2034 => x"3480c275",
2035 => x"70810557",
2036 => x"34835977",
2037 => x"75348119",
2038 => x"800c8a3d",
2039 => x"0d04fa3d",
2040 => x"0d78818a",
2041 => x"9408540b",
2042 => x"0b55b873",
2043 => x"0508802e",
2044 => x"81ce388c",
2045 => x"15227083",
2046 => x"ffff0670",
2047 => x"832a8132",
2048 => x"70810651",
2049 => x"55555672",
2050 => x"802e80ea",
2051 => x"3873842a",
2052 => x"81328106",
2053 => x"57ff530b",
2054 => x"0b76818b",
2055 => x"3873822a",
2056 => x"70810651",
2057 => x"530b0b72",
2058 => x"802ebf38",
2059 => x"b0150854",
2060 => x"0b0b7380",
2061 => x"2e9e3880",
2062 => x"c015530b",
2063 => x"0b73732e",
2064 => x"8f387352",
2065 => x"818a9408",
2066 => x"5188a53f",
2067 => x"8c152256",
2068 => x"76b0160c",
2069 => x"75db0653",
2070 => x"0b0b728c",
2071 => x"1623800b",
2072 => x"84160c90",
2073 => x"1508750c",
2074 => x"72560b0b",
2075 => x"75880753",
2076 => x"0b0b728c",
2077 => x"16239015",
2078 => x"08802e80",
2079 => x"cb388c15",
2080 => x"22708106",
2081 => x"55530b0b",
2082 => x"73a43872",
2083 => x"0a100a70",
2084 => x"81065153",
2085 => x"0b0b7287",
2086 => x"38941508",
2087 => x"540b0b73",
2088 => x"88160c80",
2089 => x"530b0b72",
2090 => x"800c883d",
2091 => x"0d04800b",
2092 => x"88160c94",
2093 => x"15083098",
2094 => x"160c8053",
2095 => x"0b0be839",
2096 => x"725183a6",
2097 => x"3ffeac39",
2098 => x"745194c6",
2099 => x"3f8c1522",
2100 => x"70810655",
2101 => x"530b0b73",
2102 => x"802effaf",
2103 => x"38d039f8",
2104 => x"3d0d7a58",
2105 => x"0b0b7780",
2106 => x"2e81a938",
2107 => x"818a9408",
2108 => x"540b0bb8",
2109 => x"1408802e",
2110 => x"80f9388c",
2111 => x"18227090",
2112 => x"2b70902c",
2113 => x"70832a81",
2114 => x"3281065c",
2115 => x"5157540b",
2116 => x"0b7880d7",
2117 => x"38901808",
2118 => x"570b0b76",
2119 => x"802e80cb",
2120 => x"38770877",
2121 => x"3177790c",
2122 => x"7683067a",
2123 => x"5855550b",
2124 => x"73853894",
2125 => x"1808560b",
2126 => x"0b758819",
2127 => x"0c807525",
2128 => x"aa387453",
2129 => x"0b0b7652",
2130 => x"9c180851",
2131 => x"a4180854",
2132 => x"0b0b732d",
2133 => x"800b8008",
2134 => x"2580cd38",
2135 => x"80081775",
2136 => x"80083156",
2137 => x"570b7480",
2138 => x"24d83880",
2139 => x"0b800c8a",
2140 => x"3d0d0473",
2141 => x"5181f33f",
2142 => x"8c182270",
2143 => x"902b7090",
2144 => x"2c70832a",
2145 => x"81328106",
2146 => x"5c515754",
2147 => x"0b0b78db",
2148 => x"38ff8239",
2149 => x"80c1df52",
2150 => x"818a9408",
2151 => x"5191973f",
2152 => x"8008800c",
2153 => x"8a3d0d04",
2154 => x"8c182280",
2155 => x"c007540b",
2156 => x"0b738c19",
2157 => x"23ff0b80",
2158 => x"0c8a3d0d",
2159 => x"04707251",
2160 => x"800b710c",
2161 => x"800b8472",
2162 => x"050c800b",
2163 => x"8872050c",
2164 => x"028e0522",
2165 => x"8c720523",
2166 => x"02920522",
2167 => x"8e720523",
2168 => x"800b9072",
2169 => x"050c800b",
2170 => x"9472050c",
2171 => x"800b9872",
2172 => x"050c709c",
2173 => x"72050c80",
2174 => x"f3d60ba0",
2175 => x"72050c80",
2176 => x"f4a90ba4",
2177 => x"72050c80",
2178 => x"f5bc0ba8",
2179 => x"72050c80",
2180 => x"f6960bac",
2181 => x"72050c50",
2182 => x"04fa3d0d",
2183 => x"797080dc",
2184 => x"298c7105",
2185 => x"540b0b7a",
2186 => x"530b0b56",
2187 => x"57949a3f",
2188 => x"80088008",
2189 => x"55568008",
2190 => x"802ea838",
2191 => x"80088c05",
2192 => x"540b0b80",
2193 => x"0b80080c",
2194 => x"76800884",
2195 => x"050c7380",
2196 => x"0888050c",
2197 => x"74530b0b",
2198 => x"80527351",
2199 => x"a4b13f75",
2200 => x"540b0b73",
2201 => x"800c883d",
2202 => x"0d04fc3d",
2203 => x"0d7680c7",
2204 => x"940bbc72",
2205 => x"050c5581",
2206 => x"0bb8160c",
2207 => x"800b84dc",
2208 => x"160c830b",
2209 => x"84e0160c",
2210 => x"84e81584",
2211 => x"e4160c74",
2212 => x"540b0b80",
2213 => x"530b0b84",
2214 => x"52841508",
2215 => x"51fe9e3f",
2216 => x"74540b0b",
2217 => x"81530b0b",
2218 => x"89528815",
2219 => x"0851fe8d",
2220 => x"3f74540b",
2221 => x"0b82530b",
2222 => x"0b8a528c",
2223 => x"150851fd",
2224 => x"fc3f863d",
2225 => x"0d04f93d",
2226 => x"0d79818a",
2227 => x"9408540b",
2228 => x"0b57b873",
2229 => x"0508802e",
2230 => x"80ce3884",
2231 => x"dc730556",
2232 => x"88160884",
2233 => x"1708ff05",
2234 => x"55558074",
2235 => x"24a2388c",
2236 => x"15227090",
2237 => x"2b70902c",
2238 => x"51540b0b",
2239 => x"5872802e",
2240 => x"80cd3880",
2241 => x"dc15ff15",
2242 => x"55550b73",
2243 => x"8025e038",
2244 => x"7508530b",
2245 => x"0b72802e",
2246 => x"9f387256",
2247 => x"88160884",
2248 => x"1708ff05",
2249 => x"5555c339",
2250 => x"7251febe",
2251 => x"3f818a94",
2252 => x"0884dc05",
2253 => x"56ffa939",
2254 => x"84527651",
2255 => x"fddb3f80",
2256 => x"08760c80",
2257 => x"08802e80",
2258 => x"c0388008",
2259 => x"56ce3981",
2260 => x"0b8c1623",
2261 => x"72750c72",
2262 => x"88160c72",
2263 => x"84160c72",
2264 => x"90160c72",
2265 => x"94160c72",
2266 => x"98160cff",
2267 => x"0b8e1623",
2268 => x"72b0160c",
2269 => x"72b4160c",
2270 => x"7280c416",
2271 => x"0c7280c8",
2272 => x"160c7480",
2273 => x"0c893d0d",
2274 => x"048c770c",
2275 => x"800b800c",
2276 => x"893d0d04",
2277 => x"707080c1",
2278 => x"df527351",
2279 => x"8d983f50",
2280 => x"50047081",
2281 => x"8a940851",
2282 => x"eb3f5004",
2283 => x"fb3d0d77",
2284 => x"705256a3",
2285 => x"873f8191",
2286 => x"f00b8805",
2287 => x"08847105",
2288 => x"08fc0670",
2289 => x"7b319fef",
2290 => x"05e08006",
2291 => x"e0800556",
2292 => x"56530b0b",
2293 => x"a0807424",
2294 => x"96388052",
2295 => x"7551abbb",
2296 => x"3f8191f8",
2297 => x"0815530b",
2298 => x"0b728008",
2299 => x"2e913875",
2300 => x"51a2ca3f",
2301 => x"80530b0b",
2302 => x"72800c87",
2303 => x"3d0d0473",
2304 => x"30527551",
2305 => x"ab953f80",
2306 => x"08ff2eab",
2307 => x"388191f0",
2308 => x"0b880508",
2309 => x"75753181",
2310 => x"07847205",
2311 => x"0c530b0b",
2312 => x"8191b408",
2313 => x"74318191",
2314 => x"b40c7551",
2315 => x"a28f3f81",
2316 => x"0b800c87",
2317 => x"3d0d0480",
2318 => x"527551aa",
2319 => x"de3f8191",
2320 => x"f00b8805",
2321 => x"08800871",
2322 => x"3156530b",
2323 => x"0b8f7525",
2324 => x"ff9d3880",
2325 => x"088191e4",
2326 => x"08318191",
2327 => x"b40c7481",
2328 => x"0784140c",
2329 => x"7551a1d5",
2330 => x"3f80530b",
2331 => x"0bff8939",
2332 => x"f63d0d7c",
2333 => x"7e540b0b",
2334 => x"5b72802e",
2335 => x"82a2387a",
2336 => x"51a1b93f",
2337 => x"f8730584",
2338 => x"71050870",
2339 => x"fe067073",
2340 => x"05847105",
2341 => x"08fc065d",
2342 => x"5859540b",
2343 => x"0b588191",
2344 => x"f808752e",
2345 => x"83833878",
2346 => x"84160c80",
2347 => x"73810654",
2348 => x"0b0b5a72",
2349 => x"0b7a2e81",
2350 => x"eb387815",
2351 => x"84710508",
2352 => x"81065153",
2353 => x"0b0b72a3",
2354 => x"38781757",
2355 => x"7981fc38",
2356 => x"88150853",
2357 => x"0b0b7281",
2358 => x"91f82e83",
2359 => x"9c388c15",
2360 => x"08708c15",
2361 => x"0c738872",
2362 => x"050c5676",
2363 => x"81078419",
2364 => x"0c761877",
2365 => x"710c530b",
2366 => x"0b79819f",
2367 => x"3883ff77",
2368 => x"2781da38",
2369 => x"76892a77",
2370 => x"832a5653",
2371 => x"0b0b7280",
2372 => x"2e80c038",
2373 => x"76862ab8",
2374 => x"05558473",
2375 => x"27b53880",
2376 => x"db730555",
2377 => x"947327ab",
2378 => x"38768c2a",
2379 => x"80ee0555",
2380 => x"80d47327",
2381 => x"9e38768f",
2382 => x"2a80f705",
2383 => x"5582d473",
2384 => x"27913876",
2385 => x"922a80fc",
2386 => x"05558ad4",
2387 => x"73278438",
2388 => x"80fe550b",
2389 => x"0b741010",
2390 => x"108191f0",
2391 => x"05887105",
2392 => x"0855560b",
2393 => x"730b762e",
2394 => x"82cd3884",
2395 => x"1408fc06",
2396 => x"530b0b76",
2397 => x"73278f38",
2398 => x"88140854",
2399 => x"0b0b7376",
2400 => x"2e098106",
2401 => x"e6388c14",
2402 => x"08708c1a",
2403 => x"0c74881a",
2404 => x"0c788872",
2405 => x"050c5677",
2406 => x"8c150c7a",
2407 => x"519f9e3f",
2408 => x"8c3d0d04",
2409 => x"77087871",
2410 => x"31597705",
2411 => x"88190854",
2412 => x"0b0b5772",
2413 => x"8191f82e",
2414 => x"80ea388c",
2415 => x"1808708c",
2416 => x"150c7388",
2417 => x"72050c56",
2418 => x"fdf03988",
2419 => x"15088c16",
2420 => x"08708c73",
2421 => x"050c5788",
2422 => x"170cfe8f",
2423 => x"3976832a",
2424 => x"70540b0b",
2425 => x"55800b75",
2426 => x"2481a338",
2427 => x"72822c81",
2428 => x"712b8191",
2429 => x"f4080781",
2430 => x"91f00b84",
2431 => x"050c530b",
2432 => x"0b741010",
2433 => x"108191f0",
2434 => x"05887105",
2435 => x"0855560b",
2436 => x"0b758c19",
2437 => x"0c738819",
2438 => x"0c778817",
2439 => x"0c778c15",
2440 => x"0cfef839",
2441 => x"815afd92",
2442 => x"39781773",
2443 => x"8106540b",
2444 => x"0b57729a",
2445 => x"38770878",
2446 => x"71315977",
2447 => x"058c1908",
2448 => x"881a0871",
2449 => x"8c72050c",
2450 => x"8872050c",
2451 => x"57570b0b",
2452 => x"76810784",
2453 => x"190c7781",
2454 => x"91f00b88",
2455 => x"050c8191",
2456 => x"ec087726",
2457 => x"feb53881",
2458 => x"91e80852",
2459 => x"7a51fabc",
2460 => x"3f7a519d",
2461 => x"c83ffea8",
2462 => x"3981788c",
2463 => x"150c7888",
2464 => x"150c738c",
2465 => x"1a0c7388",
2466 => x"1a0c5afc",
2467 => x"de398315",
2468 => x"70822c81",
2469 => x"712b8191",
2470 => x"f4080781",
2471 => x"91f00b84",
2472 => x"050c5153",
2473 => x"0b0b7410",
2474 => x"10108191",
2475 => x"f0058871",
2476 => x"05085556",
2477 => x"fed93974",
2478 => x"530b0b80",
2479 => x"7524a938",
2480 => x"72822c81",
2481 => x"712b8191",
2482 => x"f4080781",
2483 => x"91f00b84",
2484 => x"050c530b",
2485 => x"0b758c19",
2486 => x"0c738819",
2487 => x"0c778817",
2488 => x"0c778c15",
2489 => x"0cfdb439",
2490 => x"83157082",
2491 => x"2c81712b",
2492 => x"8191f408",
2493 => x"078191f0",
2494 => x"0b84050c",
2495 => x"51530b0b",
2496 => x"d439f23d",
2497 => x"0d606288",
2498 => x"71050870",
2499 => x"57575f5a",
2500 => x"74802e81",
2501 => x"9f388c1a",
2502 => x"2270832a",
2503 => x"81327081",
2504 => x"06515558",
2505 => x"0b738638",
2506 => x"901a0893",
2507 => x"387951f1",
2508 => x"ad3fff54",
2509 => x"0b0b8008",
2510 => x"80fa388c",
2511 => x"1a22587d",
2512 => x"08578078",
2513 => x"83ffff06",
2514 => x"700a100a",
2515 => x"70810651",
2516 => x"56575573",
2517 => x"0b752e80",
2518 => x"e2387491",
2519 => x"38760884",
2520 => x"18088819",
2521 => x"5956590b",
2522 => x"74802ef1",
2523 => x"3874540b",
2524 => x"0b888075",
2525 => x"27863888",
2526 => x"80540b0b",
2527 => x"73530b0b",
2528 => x"78529c1a",
2529 => x"0851a41a",
2530 => x"08540b0b",
2531 => x"732d800b",
2532 => x"80082583",
2533 => x"86388008",
2534 => x"19758008",
2535 => x"317f8805",
2536 => x"08800831",
2537 => x"70618805",
2538 => x"0c565659",
2539 => x"73ffab38",
2540 => x"80540b0b",
2541 => x"73800c90",
2542 => x"3d0d0475",
2543 => x"81327081",
2544 => x"06764151",
2545 => x"540b0b73",
2546 => x"802e81d0",
2547 => x"38749138",
2548 => x"76088418",
2549 => x"08881959",
2550 => x"56590b74",
2551 => x"802ef138",
2552 => x"881a0878",
2553 => x"83ffff06",
2554 => x"70892a70",
2555 => x"81065156",
2556 => x"59567380",
2557 => x"2e839e38",
2558 => x"7575278f",
2559 => x"3877872a",
2560 => x"70810651",
2561 => x"540b0b73",
2562 => x"82d63874",
2563 => x"76278338",
2564 => x"74560b0b",
2565 => x"75530b0b",
2566 => x"78527908",
2567 => x"5196f93f",
2568 => x"881a0876",
2569 => x"31881b0c",
2570 => x"7908167a",
2571 => x"0c74560b",
2572 => x"0b751975",
2573 => x"77317f88",
2574 => x"05087831",
2575 => x"70618805",
2576 => x"0c565659",
2577 => x"73802efe",
2578 => x"e7388c1a",
2579 => x"2258fefd",
2580 => x"39777854",
2581 => x"0b0b7953",
2582 => x"0b0b7b52",
2583 => x"5696b93f",
2584 => x"881a0878",
2585 => x"31881b0c",
2586 => x"7908187a",
2587 => x"0c7c7631",
2588 => x"5d0b0b7c",
2589 => x"8e387951",
2590 => x"f0e53f80",
2591 => x"08819c38",
2592 => x"80085f75",
2593 => x"19757731",
2594 => x"7f880508",
2595 => x"78317061",
2596 => x"88050c56",
2597 => x"56597380",
2598 => x"2efe9538",
2599 => x"74819438",
2600 => x"76088418",
2601 => x"08881959",
2602 => x"56590b74",
2603 => x"802ef138",
2604 => x"74530b0b",
2605 => x"8a527851",
2606 => x"94a33f80",
2607 => x"08793181",
2608 => x"055d8008",
2609 => x"84388115",
2610 => x"5d815f7c",
2611 => x"58747d27",
2612 => x"83387458",
2613 => x"941a0888",
2614 => x"1b087105",
2615 => x"575c807a",
2616 => x"085c540b",
2617 => x"0b901a08",
2618 => x"7b278538",
2619 => x"81540b0b",
2620 => x"75782585",
2621 => x"387380c2",
2622 => x"387b7824",
2623 => x"fed3387b",
2624 => x"530b0b78",
2625 => x"529c1a08",
2626 => x"51a41a08",
2627 => x"540b0b73",
2628 => x"2d800856",
2629 => x"80088024",
2630 => x"fed3388c",
2631 => x"1a2280c0",
2632 => x"07540b0b",
2633 => x"738c1b23",
2634 => x"ff540b0b",
2635 => x"73800c90",
2636 => x"3d0d047e",
2637 => x"ff9538fe",
2638 => x"f7397553",
2639 => x"0b0b7852",
2640 => x"7a5194d4",
2641 => x"3f790816",
2642 => x"7a0c7951",
2643 => x"ef913f80",
2644 => x"08c9387c",
2645 => x"76315d0b",
2646 => x"0b7cfea7",
2647 => x"38fe9739",
2648 => x"901a087a",
2649 => x"08713176",
2650 => x"71057056",
2651 => x"5a575281",
2652 => x"8a940851",
2653 => x"97c83f80",
2654 => x"08802eff",
2655 => x"9e388008",
2656 => x"901b0c80",
2657 => x"08167a0c",
2658 => x"77941b0c",
2659 => x"74881b0c",
2660 => x"7456fcf7",
2661 => x"39790858",
2662 => x"901a0878",
2663 => x"27853881",
2664 => x"540b0b75",
2665 => x"75278438",
2666 => x"73bd3894",
2667 => x"1a08560b",
2668 => x"0b757526",
2669 => x"80e13875",
2670 => x"530b0b78",
2671 => x"529c1a08",
2672 => x"51a41a08",
2673 => x"540b0b73",
2674 => x"2d800856",
2675 => x"80088024",
2676 => x"fcdd388c",
2677 => x"1a2280c0",
2678 => x"07540b0b",
2679 => x"738c1b23",
2680 => x"ff540b0b",
2681 => x"fec63975",
2682 => x"530b0b78",
2683 => x"52775193",
2684 => x"a73f7908",
2685 => x"167a0c79",
2686 => x"51ede43f",
2687 => x"8008802e",
2688 => x"fcad388c",
2689 => x"1a2280c0",
2690 => x"07540b0b",
2691 => x"738c1b23",
2692 => x"ff540b0b",
2693 => x"fe963974",
2694 => x"75540b0b",
2695 => x"79530b0b",
2696 => x"78525692",
2697 => x"f33f881a",
2698 => x"08753188",
2699 => x"1b0c7908",
2700 => x"157a0cfb",
2701 => x"fa39f93d",
2702 => x"0d797b58",
2703 => x"530b0b80",
2704 => x"0b818a94",
2705 => x"08530b0b",
2706 => x"5672722e",
2707 => x"80d03884",
2708 => x"dc730555",
2709 => x"0b0b7476",
2710 => x"2e80c338",
2711 => x"88150884",
2712 => x"1608ff05",
2713 => x"540b0b54",
2714 => x"0b0b8073",
2715 => x"24a3388c",
2716 => x"14227090",
2717 => x"2b70902c",
2718 => x"51530b0b",
2719 => x"587180ed",
2720 => x"3880dc14",
2721 => x"ff14540b",
2722 => x"0b540b0b",
2723 => x"728025df",
2724 => x"38740855",
2725 => x"0b0b74c4",
2726 => x"38818a94",
2727 => x"085284dc",
2728 => x"7205550b",
2729 => x"0b74802e",
2730 => x"bd388815",
2731 => x"08841608",
2732 => x"ff05540b",
2733 => x"0b540b0b",
2734 => x"807324a2",
2735 => x"388c1422",
2736 => x"70902b70",
2737 => x"902c5153",
2738 => x"0b0b5871",
2739 => x"b33880dc",
2740 => x"14ff1454",
2741 => x"0b0b540b",
2742 => x"0b728025",
2743 => x"e0387408",
2744 => x"550b0b74",
2745 => x"c5387580",
2746 => x"0c893d0d",
2747 => x"04735176",
2748 => x"2d758008",
2749 => x"0780dc15",
2750 => x"ff155555",
2751 => x"56ff8d39",
2752 => x"7351762d",
2753 => x"75800807",
2754 => x"80dc15ff",
2755 => x"15555556",
2756 => x"c839ea3d",
2757 => x"0d688c71",
2758 => x"0522700a",
2759 => x"100a8106",
2760 => x"57585674",
2761 => x"80ee388e",
2762 => x"16227090",
2763 => x"2b70902c",
2764 => x"51555880",
2765 => x"7424b538",
2766 => x"983dc405",
2767 => x"530b0b73",
2768 => x"52818a94",
2769 => x"0851a298",
2770 => x"3f800b80",
2771 => x"08249938",
2772 => x"7983e080",
2773 => x"06540b0b",
2774 => x"7380c080",
2775 => x"2e819f38",
2776 => x"73828080",
2777 => x"2e81a138",
2778 => x"8c162257",
2779 => x"0b0b7690",
2780 => x"8007540b",
2781 => x"0b738c17",
2782 => x"23888052",
2783 => x"818a9408",
2784 => x"5181c63f",
2785 => x"80089f38",
2786 => x"8c162282",
2787 => x"07540b0b",
2788 => x"738c1723",
2789 => x"80c31670",
2790 => x"770c9017",
2791 => x"0c810b94",
2792 => x"170c983d",
2793 => x"0d04818a",
2794 => x"940880c7",
2795 => x"940bbc72",
2796 => x"050c540b",
2797 => x"0b8c1622",
2798 => x"81800754",
2799 => x"0b0b738c",
2800 => x"17238008",
2801 => x"760c8008",
2802 => x"90170c88",
2803 => x"800b9417",
2804 => x"0c74802e",
2805 => x"cd388e16",
2806 => x"2270902b",
2807 => x"70902c53",
2808 => x"0b0b5558",
2809 => x"aacb3f80",
2810 => x"08802eff",
2811 => x"b5388c16",
2812 => x"22810754",
2813 => x"0b0b738c",
2814 => x"1723983d",
2815 => x"0d04810b",
2816 => x"8c172258",
2817 => x"55fee539",
2818 => x"a8160880",
2819 => x"f5bc2e09",
2820 => x"8106fed4",
2821 => x"388c1622",
2822 => x"88800754",
2823 => x"0b0b738c",
2824 => x"17238880",
2825 => x"0b80cc17",
2826 => x"0cfece39",
2827 => x"70707352",
2828 => x"818a9408",
2829 => x"51933f50",
2830 => x"50047070",
2831 => x"7352818a",
2832 => x"940851f0",
2833 => x"ab3f5050",
2834 => x"04f33d0d",
2835 => x"7f618b71",
2836 => x"0570f806",
2837 => x"5c55555e",
2838 => x"72962683",
2839 => x"38905980",
2840 => x"0b792474",
2841 => x"7a260753",
2842 => x"0b0b8054",
2843 => x"0b0b7274",
2844 => x"2e098106",
2845 => x"80d4387d",
2846 => x"5191c13f",
2847 => x"7883f726",
2848 => x"80cf3878",
2849 => x"832a7010",
2850 => x"10108191",
2851 => x"f0058c71",
2852 => x"05085959",
2853 => x"5a76782e",
2854 => x"83e73884",
2855 => x"1708fc06",
2856 => x"568c1708",
2857 => x"88180871",
2858 => x"8c72050c",
2859 => x"8872050c",
2860 => x"58751784",
2861 => x"71050881",
2862 => x"07847205",
2863 => x"0c530b0b",
2864 => x"7d5190f9",
2865 => x"3f881754",
2866 => x"0b0b7380",
2867 => x"0c8f3d0d",
2868 => x"0478892a",
2869 => x"79832a5b",
2870 => x"530b0b72",
2871 => x"802e80c0",
2872 => x"3878862a",
2873 => x"b8055a84",
2874 => x"7327b538",
2875 => x"80db7305",
2876 => x"5a947327",
2877 => x"ab38788c",
2878 => x"2a80ee05",
2879 => x"5a80d473",
2880 => x"279e3878",
2881 => x"8f2a80f7",
2882 => x"055a82d4",
2883 => x"73279138",
2884 => x"78922a80",
2885 => x"fc055a8a",
2886 => x"d4732784",
2887 => x"3880fe5a",
2888 => x"0b0b7910",
2889 => x"10108191",
2890 => x"f0058c71",
2891 => x"05085855",
2892 => x"0b760b75",
2893 => x"2ea63884",
2894 => x"1708fc06",
2895 => x"707a3155",
2896 => x"560b738f",
2897 => x"2489c638",
2898 => x"738025fe",
2899 => x"d4388c17",
2900 => x"08570b0b",
2901 => x"76752e09",
2902 => x"8106dc38",
2903 => x"811a5a81",
2904 => x"92800857",
2905 => x"0b0b7681",
2906 => x"91f82e82",
2907 => x"ed388417",
2908 => x"08fc0670",
2909 => x"7a315556",
2910 => x"0b738f24",
2911 => x"829c3881",
2912 => x"91f80b81",
2913 => x"92840c81",
2914 => x"91f80b81",
2915 => x"92800c73",
2916 => x"8025fe9d",
2917 => x"3883ff76",
2918 => x"27849d38",
2919 => x"75892a76",
2920 => x"832a5553",
2921 => x"0b0b7280",
2922 => x"2e80cc38",
2923 => x"75862ab8",
2924 => x"05540b0b",
2925 => x"847327bf",
2926 => x"3880db73",
2927 => x"05540b0b",
2928 => x"947327b3",
2929 => x"38758c2a",
2930 => x"80ee0554",
2931 => x"0b0b80d4",
2932 => x"7327a438",
2933 => x"758f2a80",
2934 => x"f705540b",
2935 => x"0b82d473",
2936 => x"27953875",
2937 => x"922a80fc",
2938 => x"05540b0b",
2939 => x"8ad47327",
2940 => x"863880fe",
2941 => x"540b0b73",
2942 => x"10101081",
2943 => x"91f00588",
2944 => x"71050856",
2945 => x"580b740b",
2946 => x"782e87a0",
2947 => x"38841508",
2948 => x"fc06530b",
2949 => x"0b757327",
2950 => x"8f388815",
2951 => x"08550b0b",
2952 => x"74782e09",
2953 => x"8106e638",
2954 => x"8c150881",
2955 => x"91f00b84",
2956 => x"0508718c",
2957 => x"1a0c7688",
2958 => x"1a0c7888",
2959 => x"73050c78",
2960 => x"8c180c5d",
2961 => x"5879530b",
2962 => x"0b807a24",
2963 => x"84983872",
2964 => x"822c8171",
2965 => x"2b5c530b",
2966 => x"0b7a7c26",
2967 => x"81ac387b",
2968 => x"7b06530b",
2969 => x"0b728398",
2970 => x"3879fc06",
2971 => x"84055a7a",
2972 => x"10707d06",
2973 => x"540b0b5b",
2974 => x"72838538",
2975 => x"841a5aef",
2976 => x"3988178c",
2977 => x"71050858",
2978 => x"580b760b",
2979 => x"782e0981",
2980 => x"06fc8838",
2981 => x"821a5afd",
2982 => x"c6397817",
2983 => x"79810784",
2984 => x"190c7081",
2985 => x"92840c70",
2986 => x"8192800c",
2987 => x"8191f80b",
2988 => x"8c72050c",
2989 => x"8c710508",
2990 => x"8872050c",
2991 => x"74810784",
2992 => x"72050c74",
2993 => x"71057571",
2994 => x"0c51530b",
2995 => x"0b7d518c",
2996 => x"ec3f8817",
2997 => x"540b0bfb",
2998 => x"f1398191",
2999 => x"f00b8405",
3000 => x"087a540b",
3001 => x"0b5c7980",
3002 => x"25fee438",
3003 => x"82f8397a",
3004 => x"097c0670",
3005 => x"8191f00b",
3006 => x"84050c5c",
3007 => x"7a105b0b",
3008 => x"0b7a7c26",
3009 => x"85387a85",
3010 => x"f2388191",
3011 => x"f00b8805",
3012 => x"08708472",
3013 => x"0508fc06",
3014 => x"707c317c",
3015 => x"72268f72",
3016 => x"25075757",
3017 => x"5c5d5572",
3018 => x"802e80e3",
3019 => x"38797a16",
3020 => x"8191e808",
3021 => x"1b907105",
3022 => x"5a55575b",
3023 => x"8191e408",
3024 => x"ff2e8938",
3025 => x"a08f7305",
3026 => x"e0800657",
3027 => x"0b0b7652",
3028 => x"7d5194c7",
3029 => x"3f800854",
3030 => x"0b0b8008",
3031 => x"ff2e9038",
3032 => x"80087627",
3033 => x"82b33874",
3034 => x"8191f02e",
3035 => x"82ab3881",
3036 => x"91f00b88",
3037 => x"05085584",
3038 => x"1508fc06",
3039 => x"707a317a",
3040 => x"72268f72",
3041 => x"25075255",
3042 => x"530b0b72",
3043 => x"84913874",
3044 => x"79810784",
3045 => x"170c7916",
3046 => x"708191f0",
3047 => x"0b88050c",
3048 => x"75810784",
3049 => x"72050c54",
3050 => x"0b0b7e52",
3051 => x"578b8e3f",
3052 => x"8817540b",
3053 => x"0bfa9339",
3054 => x"75832a70",
3055 => x"540b0b54",
3056 => x"0b0b8074",
3057 => x"2481a738",
3058 => x"72822c81",
3059 => x"712b8191",
3060 => x"f4080770",
3061 => x"8191f00b",
3062 => x"84050c75",
3063 => x"10101081",
3064 => x"91f00588",
3065 => x"71050858",
3066 => x"5a5d530b",
3067 => x"0b778c18",
3068 => x"0c748818",
3069 => x"0c768819",
3070 => x"0c768c16",
3071 => x"0cfcc639",
3072 => x"797a1010",
3073 => x"108191f0",
3074 => x"05705759",
3075 => x"5d8c1508",
3076 => x"570b0b76",
3077 => x"752ea638",
3078 => x"841708fc",
3079 => x"06707a31",
3080 => x"55560b73",
3081 => x"8f2483ef",
3082 => x"38738025",
3083 => x"84af388c",
3084 => x"1708570b",
3085 => x"0b76752e",
3086 => x"098106dc",
3087 => x"38881581",
3088 => x"1b708306",
3089 => x"555b5572",
3090 => x"c4387c83",
3091 => x"06530b0b",
3092 => x"72802efd",
3093 => x"9a38ff1d",
3094 => x"f819595d",
3095 => x"88180878",
3096 => x"2ee838fd",
3097 => x"9739831a",
3098 => x"530b0bfb",
3099 => x"e2398314",
3100 => x"70822c81",
3101 => x"712b8191",
3102 => x"f4080770",
3103 => x"8191f00b",
3104 => x"84050c76",
3105 => x"10101081",
3106 => x"91f00588",
3107 => x"71050859",
3108 => x"5b5e5153",
3109 => x"0b0bfed5",
3110 => x"398191b4",
3111 => x"08175880",
3112 => x"08762e81",
3113 => x"99388191",
3114 => x"e408ff2e",
3115 => x"849b3873",
3116 => x"76311881",
3117 => x"91b40c73",
3118 => x"87067057",
3119 => x"530b0b72",
3120 => x"802e8838",
3121 => x"88733170",
3122 => x"15555676",
3123 => x"149fff06",
3124 => x"a0807131",
3125 => x"1770540b",
3126 => x"0b7f530b",
3127 => x"0b57530b",
3128 => x"0b91b83f",
3129 => x"8008530b",
3130 => x"0b8008ff",
3131 => x"2e81a738",
3132 => x"8191b408",
3133 => x"16708191",
3134 => x"b40c7475",
3135 => x"8191f00b",
3136 => x"88050c74",
3137 => x"76311870",
3138 => x"81075155",
3139 => x"56587b81",
3140 => x"91f02e83",
3141 => x"c138798f",
3142 => x"2682ee38",
3143 => x"810b8415",
3144 => x"0c841508",
3145 => x"fc06707a",
3146 => x"317a7226",
3147 => x"8f722507",
3148 => x"5255530b",
3149 => x"0b72802e",
3150 => x"fcd53880",
3151 => x"e2398008",
3152 => x"9fff0653",
3153 => x"0b0b72fe",
3154 => x"dd387781",
3155 => x"91b40c81",
3156 => x"91f00b88",
3157 => x"05087b18",
3158 => x"81078472",
3159 => x"050c5581",
3160 => x"91e00878",
3161 => x"27863877",
3162 => x"8191e00c",
3163 => x"8191dc08",
3164 => x"7827fc83",
3165 => x"38778191",
3166 => x"dc0c8415",
3167 => x"08fc0670",
3168 => x"7a317a72",
3169 => x"268f7225",
3170 => x"07525553",
3171 => x"0b0b7280",
3172 => x"2efbfc38",
3173 => x"8a398074",
3174 => x"540b0b56",
3175 => x"fed2397d",
3176 => x"51879a3f",
3177 => x"800b800c",
3178 => x"8f3d0d04",
3179 => x"73530b0b",
3180 => x"807424ab",
3181 => x"3872822c",
3182 => x"81712b81",
3183 => x"91f40807",
3184 => x"708191f0",
3185 => x"0b84050c",
3186 => x"5d530b0b",
3187 => x"778c180c",
3188 => x"7488180c",
3189 => x"7688190c",
3190 => x"768c160c",
3191 => x"f8e73983",
3192 => x"1470822c",
3193 => x"81712b81",
3194 => x"91f40807",
3195 => x"708191f0",
3196 => x"0b84050c",
3197 => x"5e51530b",
3198 => x"0bd2397b",
3199 => x"7b06530b",
3200 => x"0b72fbfc",
3201 => x"38841a7b",
3202 => x"105c5aef",
3203 => x"39ff1a81",
3204 => x"7105515a",
3205 => x"f6c93978",
3206 => x"17798107",
3207 => x"84190c8c",
3208 => x"18088819",
3209 => x"08718c72",
3210 => x"050c8872",
3211 => x"050c5970",
3212 => x"8192840c",
3213 => x"70819280",
3214 => x"0c8191f8",
3215 => x"0b8c7205",
3216 => x"0c8c7105",
3217 => x"08887205",
3218 => x"0c748107",
3219 => x"8472050c",
3220 => x"74710575",
3221 => x"710c5153",
3222 => x"0b0bf8f1",
3223 => x"39751784",
3224 => x"71050881",
3225 => x"07847205",
3226 => x"0c530b0b",
3227 => x"8c170888",
3228 => x"1808718c",
3229 => x"72050c88",
3230 => x"72050c58",
3231 => x"7d5185bd",
3232 => x"3f881754",
3233 => x"0b0bf4c2",
3234 => x"39728415",
3235 => x"0cf41af8",
3236 => x"0670841e",
3237 => x"08810607",
3238 => x"841e0c70",
3239 => x"1d540b0b",
3240 => x"5b850b84",
3241 => x"140c850b",
3242 => x"88140c8f",
3243 => x"7b27fdaf",
3244 => x"38881c52",
3245 => x"7d51e3b8",
3246 => x"3f8191f0",
3247 => x"0b880508",
3248 => x"8191b408",
3249 => x"5955fd97",
3250 => x"39778191",
3251 => x"b40c7381",
3252 => x"91e40cfb",
3253 => x"e2397284",
3254 => x"150cfd83",
3255 => x"39fa3d0d",
3256 => x"7a790288",
3257 => x"05a70533",
3258 => x"5652530b",
3259 => x"0b837327",
3260 => x"8c387083",
3261 => x"06520b0b",
3262 => x"71802eb1",
3263 => x"38ff7305",
3264 => x"530b0b72",
3265 => x"ff2e9b38",
3266 => x"70335273",
3267 => x"0b722e94",
3268 => x"38817105",
3269 => x"ff14540b",
3270 => x"0b5172ff",
3271 => x"2e098106",
3272 => x"e7388051",
3273 => x"0b0b7080",
3274 => x"0c883d0d",
3275 => x"04707257",
3276 => x"55835175",
3277 => x"82802914",
3278 => x"ff720552",
3279 => x"560b7080",
3280 => x"25f13883",
3281 => x"732780cb",
3282 => x"38740876",
3283 => x"327009f7",
3284 => x"fbfdff72",
3285 => x"050670f8",
3286 => x"84828180",
3287 => x"06515151",
3288 => x"0b0b7080",
3289 => x"2e9e3874",
3290 => x"51805270",
3291 => x"3357730b",
3292 => x"772effb0",
3293 => x"38817105",
3294 => x"81730553",
3295 => x"0b0b5183",
3296 => x"7227e838",
3297 => x"fc730584",
3298 => x"1656530b",
3299 => x"0b728326",
3300 => x"ffb73874",
3301 => x"51fee639",
3302 => x"fa3d0d78",
3303 => x"7a7c7272",
3304 => x"72575757",
3305 => x"5956560b",
3306 => x"740b7627",
3307 => x"be387615",
3308 => x"51750b71",
3309 => x"27b53870",
3310 => x"7717ff14",
3311 => x"540b0b55",
3312 => x"530b0b71",
3313 => x"ff2e9d38",
3314 => x"ff14ff14",
3315 => x"540b0b54",
3316 => x"0b0b7233",
3317 => x"7434ff72",
3318 => x"05520b0b",
3319 => x"71ff2e09",
3320 => x"8106e538",
3321 => x"75800c88",
3322 => x"3d0d0476",
3323 => x"8f269c38",
3324 => x"ff720552",
3325 => x"0b0b71ff",
3326 => x"2eea3872",
3327 => x"70810554",
3328 => x"0b0b3374",
3329 => x"70810556",
3330 => x"34e63974",
3331 => x"76078306",
3332 => x"510b0b70",
3333 => x"db387575",
3334 => x"540b0b51",
3335 => x"72708405",
3336 => x"540b0b08",
3337 => x"71708405",
3338 => x"530b0b0c",
3339 => x"72708405",
3340 => x"540b0b08",
3341 => x"71708405",
3342 => x"530b0b0c",
3343 => x"72708405",
3344 => x"540b0b08",
3345 => x"71708405",
3346 => x"530b0b0c",
3347 => x"72708405",
3348 => x"540b0b08",
3349 => x"71708405",
3350 => x"530b0b0c",
3351 => x"f0720552",
3352 => x"0b0b718f",
3353 => x"26ffb538",
3354 => x"8372279c",
3355 => x"38727084",
3356 => x"05540b0b",
3357 => x"08717084",
3358 => x"05530b0b",
3359 => x"0cfc7205",
3360 => x"520b0b71",
3361 => x"8326e638",
3362 => x"70540b0b",
3363 => x"fee239fc",
3364 => x"3d0d7679",
3365 => x"71028c05",
3366 => x"9f053357",
3367 => x"55530b0b",
3368 => x"55837227",
3369 => x"8c387483",
3370 => x"06510b0b",
3371 => x"70802ea8",
3372 => x"38ff7205",
3373 => x"520b0b71",
3374 => x"ff2e9638",
3375 => x"73737081",
3376 => x"055534ff",
3377 => x"7205520b",
3378 => x"0b71ff2e",
3379 => x"098106ec",
3380 => x"3874800c",
3381 => x"863d0d04",
3382 => x"7474882b",
3383 => x"75077071",
3384 => x"902b0751",
3385 => x"540b0b51",
3386 => x"8f7227b0",
3387 => x"38727170",
3388 => x"8405530b",
3389 => x"0b0c7271",
3390 => x"70840553",
3391 => x"0b0b0c72",
3392 => x"71708405",
3393 => x"530b0b0c",
3394 => x"72717084",
3395 => x"05530b0b",
3396 => x"0cf07205",
3397 => x"520b0b71",
3398 => x"8f26d238",
3399 => x"83722795",
3400 => x"38727170",
3401 => x"8405530b",
3402 => x"0b0cfc72",
3403 => x"05520b0b",
3404 => x"718326ed",
3405 => x"3870530b",
3406 => x"0bfef639",
3407 => x"0404ef3d",
3408 => x"0d636567",
3409 => x"405d420b",
3410 => x"7b802e85",
3411 => x"ab386151",
3412 => x"eb3ff81c",
3413 => x"70847205",
3414 => x"0870fc06",
3415 => x"70628b05",
3416 => x"70f80641",
3417 => x"59455b5c",
3418 => x"41579674",
3419 => x"2782e238",
3420 => x"807b247e",
3421 => x"7c260759",
3422 => x"80540b0b",
3423 => x"78742e09",
3424 => x"810682c6",
3425 => x"38777b25",
3426 => x"82913877",
3427 => x"178191f0",
3428 => x"0b880508",
3429 => x"5e560b7c",
3430 => x"0b762e84",
3431 => x"ea388416",
3432 => x"0870fe06",
3433 => x"17847105",
3434 => x"08810651",
3435 => x"55550b73",
3436 => x"82a43874",
3437 => x"fc06597c",
3438 => x"762e858f",
3439 => x"3877195f",
3440 => x"0b0b7e7b",
3441 => x"25829438",
3442 => x"79810654",
3443 => x"0b0b7382",
3444 => x"dc387677",
3445 => x"08318471",
3446 => x"0508fc06",
3447 => x"565a7580",
3448 => x"2e93387c",
3449 => x"762e859c",
3450 => x"38741918",
3451 => x"590b0b78",
3452 => x"7b2584b0",
3453 => x"3879802e",
3454 => x"82b33877",
3455 => x"15567a0b",
3456 => x"762482a9",
3457 => x"388c1a08",
3458 => x"881b0871",
3459 => x"8c72050c",
3460 => x"8872050c",
3461 => x"55797659",
3462 => x"57881761",
3463 => x"fc055759",
3464 => x"0b75a426",
3465 => x"86ab387b",
3466 => x"79555593",
3467 => x"762780cf",
3468 => x"387b7084",
3469 => x"055d087c",
3470 => x"56790c74",
3471 => x"70840556",
3472 => x"088c180c",
3473 => x"9017540b",
3474 => x"0b9b7627",
3475 => x"b2387470",
3476 => x"84055608",
3477 => x"740c7470",
3478 => x"84055608",
3479 => x"94180c98",
3480 => x"17540b0b",
3481 => x"a3762797",
3482 => x"38747084",
3483 => x"05560874",
3484 => x"0c747084",
3485 => x"0556089c",
3486 => x"180ca017",
3487 => x"540b0b74",
3488 => x"70840556",
3489 => x"08747084",
3490 => x"05560c74",
3491 => x"70840556",
3492 => x"08747084",
3493 => x"05560c74",
3494 => x"08740c77",
3495 => x"7b31560b",
3496 => x"0b758f26",
3497 => x"80d13884",
3498 => x"17088106",
3499 => x"78078418",
3500 => x"0c771784",
3501 => x"71050881",
3502 => x"07847205",
3503 => x"0c540b0b",
3504 => x"6151fcf9",
3505 => x"3f881754",
3506 => x"0b0b7380",
3507 => x"0c933d0d",
3508 => x"04905bfd",
3509 => x"9b397856",
3510 => x"fdee398c",
3511 => x"16088817",
3512 => x"08718c72",
3513 => x"050c8872",
3514 => x"050c557e",
3515 => x"707c3157",
3516 => x"588f7627",
3517 => x"ffb1387a",
3518 => x"17841808",
3519 => x"81067c07",
3520 => x"84190c76",
3521 => x"81078472",
3522 => x"050c7671",
3523 => x"05847105",
3524 => x"08810784",
3525 => x"72050c55",
3526 => x"88055261",
3527 => x"51dad13f",
3528 => x"6151fc99",
3529 => x"3f881754",
3530 => x"0b0bff9e",
3531 => x"397d5261",
3532 => x"51ea963f",
3533 => x"80085980",
3534 => x"08802e81",
3535 => x"ab388008",
3536 => x"f8056084",
3537 => x"0508fe06",
3538 => x"61055557",
3539 => x"0b0b7674",
3540 => x"2e848d38",
3541 => x"fc18560b",
3542 => x"0b75a426",
3543 => x"81b0387b",
3544 => x"80085555",
3545 => x"93762780",
3546 => x"dc387470",
3547 => x"84055608",
3548 => x"80087084",
3549 => x"05800c0c",
3550 => x"80087570",
3551 => x"84055708",
3552 => x"71708405",
3553 => x"530b0b0c",
3554 => x"540b0b9b",
3555 => x"7627b638",
3556 => x"74708405",
3557 => x"56087470",
3558 => x"8405560c",
3559 => x"74708405",
3560 => x"56087470",
3561 => x"8405560c",
3562 => x"a3762799",
3563 => x"38747084",
3564 => x"05560874",
3565 => x"70840556",
3566 => x"0c747084",
3567 => x"05560874",
3568 => x"70840556",
3569 => x"0c747084",
3570 => x"05560874",
3571 => x"70840556",
3572 => x"0c747084",
3573 => x"05560874",
3574 => x"70840556",
3575 => x"0c740874",
3576 => x"0c7b5261",
3577 => x"51d9893f",
3578 => x"6151fad1",
3579 => x"3f78540b",
3580 => x"0b73800c",
3581 => x"933d0d04",
3582 => x"7d526151",
3583 => x"e8cb3f80",
3584 => x"08800c93",
3585 => x"3d0d0484",
3586 => x"160855fb",
3587 => x"a6397553",
3588 => x"0b0b7b52",
3589 => x"800851ff",
3590 => x"a4a23f7b",
3591 => x"526151d8",
3592 => x"cf3fc539",
3593 => x"8c160888",
3594 => x"1708718c",
3595 => x"72050c88",
3596 => x"72050c55",
3597 => x"8c1a0888",
3598 => x"1b08718c",
3599 => x"72050c88",
3600 => x"72050c55",
3601 => x"79795957",
3602 => x"fbcf3977",
3603 => x"19901c55",
3604 => x"550b730b",
3605 => x"7524faf0",
3606 => x"387a1770",
3607 => x"8191f00b",
3608 => x"88050c75",
3609 => x"7c318107",
3610 => x"8472050c",
3611 => x"5d841708",
3612 => x"81067b07",
3613 => x"84180c61",
3614 => x"51f9c23f",
3615 => x"8817540b",
3616 => x"0bfcc739",
3617 => x"74191890",
3618 => x"1c555d0b",
3619 => x"730b7d24",
3620 => x"fae3388c",
3621 => x"1a08881b",
3622 => x"08718c72",
3623 => x"050c8872",
3624 => x"050c5588",
3625 => x"1a61fc05",
3626 => x"57590b75",
3627 => x"a42681bc",
3628 => x"387b7955",
3629 => x"55937627",
3630 => x"80cf387b",
3631 => x"7084055d",
3632 => x"087c5679",
3633 => x"0c747084",
3634 => x"0556088c",
3635 => x"1b0c901a",
3636 => x"540b0b9b",
3637 => x"7627b238",
3638 => x"74708405",
3639 => x"5608740c",
3640 => x"74708405",
3641 => x"5608941b",
3642 => x"0c981a54",
3643 => x"0b0ba376",
3644 => x"27973874",
3645 => x"70840556",
3646 => x"08740c74",
3647 => x"70840556",
3648 => x"089c1b0c",
3649 => x"a01a540b",
3650 => x"0b747084",
3651 => x"05560874",
3652 => x"70840556",
3653 => x"0c747084",
3654 => x"05560874",
3655 => x"70840556",
3656 => x"0c740874",
3657 => x"0c7a1a70",
3658 => x"8191f00b",
3659 => x"88050c7d",
3660 => x"7c318107",
3661 => x"8472050c",
3662 => x"540b0b84",
3663 => x"1a088106",
3664 => x"7b07841b",
3665 => x"0c6151f7",
3666 => x"f43f7854",
3667 => x"0b0bfda1",
3668 => x"3975530b",
3669 => x"0b7b5278",
3670 => x"51ffa1e0",
3671 => x"3ffabc39",
3672 => x"841708fc",
3673 => x"06186058",
3674 => x"58fab039",
3675 => x"75530b0b",
3676 => x"7b527851",
3677 => x"ffa1c53f",
3678 => x"7a1a7081",
3679 => x"91f00b88",
3680 => x"050c7d7c",
3681 => x"31810784",
3682 => x"72050c54",
3683 => x"0b0b841a",
3684 => x"0881067b",
3685 => x"07841b0c",
3686 => x"ffab3970",
3687 => x"70707080",
3688 => x"0b819ab8",
3689 => x"0c765187",
3690 => x"853f8008",
3691 => x"530b0b80",
3692 => x"08ff2e89",
3693 => x"3872800c",
3694 => x"50505050",
3695 => x"04819ab8",
3696 => x"08540b0b",
3697 => x"73802eed",
3698 => x"38757471",
3699 => x"0c527280",
3700 => x"0c505050",
3701 => x"5004f93d",
3702 => x"0d797c55",
3703 => x"7b540b0b",
3704 => x"8e710522",
3705 => x"70902b70",
3706 => x"902c5557",
3707 => x"818a9408",
3708 => x"530b0b58",
3709 => x"5685e33f",
3710 => x"80085780",
3711 => x"0b800824",
3712 => x"933880d0",
3713 => x"16088008",
3714 => x"0580d017",
3715 => x"0c76800c",
3716 => x"893d0d04",
3717 => x"8c162283",
3718 => x"dfff0655",
3719 => x"0b0b748c",
3720 => x"17237680",
3721 => x"0c893d0d",
3722 => x"04fa3d0d",
3723 => x"788c7105",
3724 => x"2270882a",
3725 => x"70810651",
3726 => x"57585674",
3727 => x"b1388c16",
3728 => x"2283dfff",
3729 => x"06550b0b",
3730 => x"748c1723",
3731 => x"7a540b0b",
3732 => x"79530b0b",
3733 => x"8e162270",
3734 => x"902b7090",
3735 => x"2c540b0b",
3736 => x"56818a94",
3737 => x"08525682",
3738 => x"fe3f883d",
3739 => x"0d048254",
3740 => x"0b0b8053",
3741 => x"0b0b8e16",
3742 => x"2270902b",
3743 => x"70902c54",
3744 => x"0b0b5681",
3745 => x"8a940852",
3746 => x"5784913f",
3747 => x"8c162283",
3748 => x"dfff0655",
3749 => x"0b0b748c",
3750 => x"17237a54",
3751 => x"0b0b7953",
3752 => x"0b0b8e16",
3753 => x"2270902b",
3754 => x"70902c54",
3755 => x"0b0b5681",
3756 => x"8a940852",
3757 => x"5682b03f",
3758 => x"883d0d04",
3759 => x"f93d0d79",
3760 => x"7c557b54",
3761 => x"0b0b8e71",
3762 => x"05227090",
3763 => x"2b70902c",
3764 => x"5557818a",
3765 => x"9408530b",
3766 => x"0b585683",
3767 => x"bf3f8008",
3768 => x"578008ff",
3769 => x"2e9b388c",
3770 => x"1622a080",
3771 => x"07550b0b",
3772 => x"748c1723",
3773 => x"800880d0",
3774 => x"170c7680",
3775 => x"0c893d0d",
3776 => x"048c1622",
3777 => x"83dfff06",
3778 => x"550b0b74",
3779 => x"8c172376",
3780 => x"800c893d",
3781 => x"0d047070",
3782 => x"70748e71",
3783 => x"05227090",
3784 => x"2b70902c",
3785 => x"55515153",
3786 => x"0b0b818a",
3787 => x"94085181",
3788 => x"f43f5050",
3789 => x"5004fb3d",
3790 => x"0d777970",
3791 => x"72078306",
3792 => x"530b0b54",
3793 => x"0b0b5270",
3794 => x"99387173",
3795 => x"7308540b",
3796 => x"0b56540b",
3797 => x"0b717308",
3798 => x"2e80d038",
3799 => x"7375540b",
3800 => x"0b520b0b",
3801 => x"71337081",
3802 => x"ff065254",
3803 => x"0b0b7080",
3804 => x"2ea33872",
3805 => x"3355700b",
3806 => x"752e0981",
3807 => x"069a3881",
3808 => x"72058114",
3809 => x"71337081",
3810 => x"ff06540b",
3811 => x"0b56540b",
3812 => x"0b5270df",
3813 => x"38723355",
3814 => x"7381ff06",
3815 => x"7581ff06",
3816 => x"71713180",
3817 => x"0c525287",
3818 => x"3d0d0471",
3819 => x"0970f7fb",
3820 => x"fdff1406",
3821 => x"70f88482",
3822 => x"81800651",
3823 => x"51510b0b",
3824 => x"709d3884",
3825 => x"14841671",
3826 => x"08540b0b",
3827 => x"56540b0b",
3828 => x"7175082e",
3829 => x"d6387375",
3830 => x"540b0b52",
3831 => x"ff843980",
3832 => x"0b800c87",
3833 => x"3d0d04fb",
3834 => x"3d0d800b",
3835 => x"819ab80c",
3836 => x"7a530b0b",
3837 => x"79527851",
3838 => x"83c33f80",
3839 => x"08558008",
3840 => x"ff2e8838",
3841 => x"74800c87",
3842 => x"3d0d0481",
3843 => x"9ab80856",
3844 => x"0b0b7580",
3845 => x"2eee3877",
3846 => x"76710c54",
3847 => x"0b0b7480",
3848 => x"0c873d0d",
3849 => x"04707070",
3850 => x"70800b81",
3851 => x"9ab80c76",
3852 => x"5185db3f",
3853 => x"8008530b",
3854 => x"0b8008ff",
3855 => x"2e893872",
3856 => x"800c5050",
3857 => x"50500481",
3858 => x"9ab80854",
3859 => x"0b0b7380",
3860 => x"2eed3875",
3861 => x"74710c52",
3862 => x"72800c50",
3863 => x"50505004",
3864 => x"fc3d0d80",
3865 => x"0b819ab8",
3866 => x"0c785277",
3867 => x"51889c3f",
3868 => x"8008540b",
3869 => x"0b8008ff",
3870 => x"2e883873",
3871 => x"800c863d",
3872 => x"0d04819a",
3873 => x"b808550b",
3874 => x"0b74802e",
3875 => x"ee387675",
3876 => x"710c530b",
3877 => x"0b73800c",
3878 => x"863d0d04",
3879 => x"fb3d0d80",
3880 => x"0b819ab8",
3881 => x"0c7a530b",
3882 => x"0b795278",
3883 => x"5185e63f",
3884 => x"80085580",
3885 => x"08ff2e88",
3886 => x"3874800c",
3887 => x"873d0d04",
3888 => x"819ab808",
3889 => x"560b0b75",
3890 => x"802eee38",
3891 => x"7776710c",
3892 => x"540b0b74",
3893 => x"800c873d",
3894 => x"0d04fb3d",
3895 => x"0d800b81",
3896 => x"9ab80c7a",
3897 => x"530b0b79",
3898 => x"52785182",
3899 => x"cd3f8008",
3900 => x"558008ff",
3901 => x"2e883874",
3902 => x"800c873d",
3903 => x"0d04819a",
3904 => x"b808560b",
3905 => x"0b75802e",
3906 => x"ee387776",
3907 => x"710c540b",
3908 => x"0b74800c",
3909 => x"873d0d04",
3910 => x"810b800c",
3911 => x"04707281",
3912 => x"2e873880",
3913 => x"0b800c50",
3914 => x"04735181",
3915 => x"8a3f7070",
3916 => x"70819abc",
3917 => x"08510b0b",
3918 => x"708a3881",
3919 => x"9ac47081",
3920 => x"9abc0c51",
3921 => x"0b0b7075",
3922 => x"72055252",
3923 => x"ff530b0b",
3924 => x"7087fb80",
3925 => x"80268a38",
3926 => x"70819abc",
3927 => x"0c71530b",
3928 => x"0b72800c",
3929 => x"50505004",
3930 => x"70707070",
3931 => x"800b818a",
3932 => x"8808540b",
3933 => x"0b540b0b",
3934 => x"72812e9e",
3935 => x"3873819a",
3936 => x"c00cff8e",
3937 => x"863fff8c",
3938 => x"f73f8199",
3939 => x"f8528151",
3940 => x"ff90e53f",
3941 => x"80085187",
3942 => x"d53f7281",
3943 => x"9ac00cff",
3944 => x"8de93fff",
3945 => x"8cda3f81",
3946 => x"99f85281",
3947 => x"51ff90c8",
3948 => x"3f800851",
3949 => x"87b83f00",
3950 => x"ff3900ff",
3951 => x"39f53d0d",
3952 => x"7e60819a",
3953 => x"c008705b",
3954 => x"585b5b75",
3955 => x"80c63877",
3956 => x"7a25a338",
3957 => x"771b7033",
3958 => x"7081ff06",
3959 => x"58585975",
3960 => x"8a2e9a38",
3961 => x"7681ff06",
3962 => x"51ff8cfc",
3963 => x"3f811858",
3964 => x"790b7824",
3965 => x"df387980",
3966 => x"0c8d3d0d",
3967 => x"048d51ff",
3968 => x"8ce63f78",
3969 => x"337081ff",
3970 => x"065257ff",
3971 => x"8cda3f81",
3972 => x"1858dd39",
3973 => x"79557a54",
3974 => x"0b0b7d53",
3975 => x"0b0b8552",
3976 => x"8d3dfc05",
3977 => x"51ff8c9c",
3978 => x"3f800856",
3979 => x"86b93f7b",
3980 => x"80080c75",
3981 => x"800c8d3d",
3982 => x"0d04f63d",
3983 => x"0d7d7f81",
3984 => x"9ac00870",
3985 => x"5a585a5a",
3986 => x"7580ca38",
3987 => x"767925b6",
3988 => x"38761a56",
3989 => x"ff8bef3f",
3990 => x"80087634",
3991 => x"800b8008",
3992 => x"81ff0657",
3993 => x"580b758a",
3994 => x"2ea73875",
3995 => x"8d327030",
3996 => x"7080257a",
3997 => x"07515156",
3998 => x"0b0b75bf",
3999 => x"38811757",
4000 => x"780b7724",
4001 => x"cc387656",
4002 => x"0b0b7580",
4003 => x"0c8c3d0d",
4004 => x"048158d7",
4005 => x"39785579",
4006 => x"540b0b7c",
4007 => x"530b0b84",
4008 => x"528c3dfc",
4009 => x"0551ff8b",
4010 => x"9b3f8008",
4011 => x"5685b83f",
4012 => x"7a80080c",
4013 => x"75800c8c",
4014 => x"3d0d0481",
4015 => x"1756c939",
4016 => x"f93d0d79",
4017 => x"57819ac0",
4018 => x"08802eb2",
4019 => x"387651ff",
4020 => x"9dc13f7b",
4021 => x"567a5580",
4022 => x"08810554",
4023 => x"0b0b7653",
4024 => x"0b0b8252",
4025 => x"893dfc05",
4026 => x"51ff8ad8",
4027 => x"3f800857",
4028 => x"84f53f77",
4029 => x"80080c76",
4030 => x"800c893d",
4031 => x"0d0484e7",
4032 => x"3f850b80",
4033 => x"080cff0b",
4034 => x"800c893d",
4035 => x"0d04fb3d",
4036 => x"0d819ac0",
4037 => x"08705654",
4038 => x"0b0b7388",
4039 => x"3874800c",
4040 => x"873d0d04",
4041 => x"77530b0b",
4042 => x"8352873d",
4043 => x"fc0551ff",
4044 => x"8a923f80",
4045 => x"08540b0b",
4046 => x"84ad3f75",
4047 => x"80080c73",
4048 => x"800c873d",
4049 => x"0d04ff0b",
4050 => x"800c04fb",
4051 => x"3d0d7755",
4052 => x"819ac008",
4053 => x"802eae38",
4054 => x"7451ff9c",
4055 => x"b63f8008",
4056 => x"8105540b",
4057 => x"0b74530b",
4058 => x"0b875287",
4059 => x"3dfc0551",
4060 => x"ff89d13f",
4061 => x"80085583",
4062 => x"ee3f7580",
4063 => x"080c7480",
4064 => x"0c873d0d",
4065 => x"0483e03f",
4066 => x"850b8008",
4067 => x"0cff0b80",
4068 => x"0c873d0d",
4069 => x"04fa3d0d",
4070 => x"819ac008",
4071 => x"802ea738",
4072 => x"7a557954",
4073 => x"0b0b7853",
4074 => x"0b0b8652",
4075 => x"883dfc05",
4076 => x"51ff8990",
4077 => x"3f800856",
4078 => x"83ad3f76",
4079 => x"80080c75",
4080 => x"800c883d",
4081 => x"0d04839f",
4082 => x"3f9d0b80",
4083 => x"080cff0b",
4084 => x"800c883d",
4085 => x"0d04fb3d",
4086 => x"0d777956",
4087 => x"56807054",
4088 => x"0b0b540b",
4089 => x"0b737525",
4090 => x"9f387410",
4091 => x"1010f805",
4092 => x"52721670",
4093 => x"3370742b",
4094 => x"76078116",
4095 => x"f8165656",
4096 => x"56515174",
4097 => x"7324ea38",
4098 => x"73800c87",
4099 => x"3d0d04fc",
4100 => x"3d0d7678",
4101 => x"5555bc53",
4102 => x"0b0b8052",
4103 => x"7351e8ef",
4104 => x"3f845274",
4105 => x"51ffaf3f",
4106 => x"80087423",
4107 => x"84528415",
4108 => x"51ffa33f",
4109 => x"80088215",
4110 => x"23845288",
4111 => x"1551ff96",
4112 => x"3f800884",
4113 => x"150c8452",
4114 => x"8c1551ff",
4115 => x"893f8008",
4116 => x"88152384",
4117 => x"52901551",
4118 => x"fefc3f80",
4119 => x"088a1523",
4120 => x"84529415",
4121 => x"51feef3f",
4122 => x"80088c15",
4123 => x"23845298",
4124 => x"1551fee2",
4125 => x"3f80088e",
4126 => x"15238852",
4127 => x"9c1551fe",
4128 => x"d53f8008",
4129 => x"90150c86",
4130 => x"3d0d04e9",
4131 => x"3d0d6a81",
4132 => x"9ac00857",
4133 => x"570b7593",
4134 => x"3880c080",
4135 => x"0b84180c",
4136 => x"75ac180c",
4137 => x"75800c99",
4138 => x"3d0d0489",
4139 => x"3d70556a",
4140 => x"540b0b55",
4141 => x"8a52993d",
4142 => x"ffbc0551",
4143 => x"ff87853f",
4144 => x"80087753",
4145 => x"0b0b7552",
4146 => x"56fec43f",
4147 => x"81993f77",
4148 => x"80080c75",
4149 => x"800c993d",
4150 => x"0d04e93d",
4151 => x"0d695781",
4152 => x"9ac00880",
4153 => x"2ebb3876",
4154 => x"51ff99a7",
4155 => x"3f893d70",
4156 => x"56800881",
4157 => x"05557754",
4158 => x"0b0b568f",
4159 => x"52993dff",
4160 => x"bc0551ff",
4161 => x"86be3f80",
4162 => x"086b530b",
4163 => x"0b765257",
4164 => x"fdfd3f80",
4165 => x"d23f7780",
4166 => x"080c7680",
4167 => x"0c993d0d",
4168 => x"0480c43f",
4169 => x"850b8008",
4170 => x"0cff0b80",
4171 => x"0c993d0d",
4172 => x"04fc3d0d",
4173 => x"81540b0b",
4174 => x"819ac008",
4175 => x"88387380",
4176 => x"0c863d0d",
4177 => x"0476530b",
4178 => x"0b97b952",
4179 => x"863dfc05",
4180 => x"51ff85f0",
4181 => x"3f800854",
4182 => x"0b0b8c3f",
4183 => x"7480080c",
4184 => x"73800c86",
4185 => x"3d0d0481",
4186 => x"8a940880",
4187 => x"0c04f73d",
4188 => x"0d7b818a",
4189 => x"940882c8",
4190 => x"7105085a",
4191 => x"540b0b5a",
4192 => x"77802e80",
4193 => x"eb388188",
4194 => x"18841908",
4195 => x"ff058171",
4196 => x"2b595559",
4197 => x"80742481",
4198 => x"80388074",
4199 => x"2480c138",
4200 => x"73822b78",
4201 => x"71058805",
4202 => x"56568180",
4203 => x"19087706",
4204 => x"530b0b72",
4205 => x"802e80c3",
4206 => x"38781670",
4207 => x"08530b0b",
4208 => x"530b0b79",
4209 => x"51740853",
4210 => x"0b0b722d",
4211 => x"ff14fc17",
4212 => x"fc177981",
4213 => x"2c5a5757",
4214 => x"540b0b73",
4215 => x"8025cb38",
4216 => x"7708580b",
4217 => x"0b77ff9e",
4218 => x"38818a94",
4219 => x"08530b0b",
4220 => x"bc730508",
4221 => x"a9387951",
4222 => x"f7bd3f74",
4223 => x"08530b0b",
4224 => x"722dff14",
4225 => x"fc17fc17",
4226 => x"79812c5a",
4227 => x"5757540b",
4228 => x"0b738025",
4229 => x"ff9438c8",
4230 => x"398057fe",
4231 => x"fd397251",
4232 => x"bc730508",
4233 => x"530b0b72",
4234 => x"2d7951f7",
4235 => x"8a3f8c08",
4236 => x"028c0c70",
4237 => x"70707080",
4238 => x"530b0b8c",
4239 => x"088c0508",
4240 => x"528c0888",
4241 => x"050851ff",
4242 => x"8dd23f80",
4243 => x"0870800c",
4244 => x"540b0b50",
4245 => x"5050508c",
4246 => x"0c048c08",
4247 => x"028c0c70",
4248 => x"70707081",
4249 => x"530b0b8c",
4250 => x"088c0508",
4251 => x"528c0888",
4252 => x"050851ff",
4253 => x"8da63f80",
4254 => x"0870800c",
4255 => x"540b0b50",
4256 => x"5050508c",
4257 => x"0c047070",
4258 => x"819a800b",
4259 => x"fc057008",
4260 => x"52520b70",
4261 => x"ff2e9338",
4262 => x"702dfc72",
4263 => x"05700852",
4264 => x"520b70ff",
4265 => x"2e098106",
4266 => x"ef385050",
4267 => x"0404ff85",
4268 => x"e53f0400",
4269 => x"4379636c",
4270 => x"65732025",
4271 => x"640a0000",
4272 => x"48656c6c",
4273 => x"6f20776f",
4274 => x"726c6420",
4275 => x"310a0000",
4276 => x"48656c6c",
4277 => x"6f20776f",
4278 => x"726c6420",
4279 => x"320a0000",
4280 => x"0a000000",
4281 => x"20202020",
4282 => x"20202020",
4283 => x"20202020",
4284 => x"20202020",
4285 => x"30303030",
4286 => x"30303030",
4287 => x"30303030",
4288 => x"30303030",
4289 => x"000017e3",
4290 => x"0000138d",
4291 => x"0000138d",
4292 => x"000017d9",
4293 => x"0000138d",
4294 => x"0000138d",
4295 => x"0000138d",
4296 => x"0000138d",
4297 => x"0000138d",
4298 => x"0000138d",
4299 => x"00001364",
4300 => x"0000177e",
4301 => x"0000138d",
4302 => x"00001376",
4303 => x"000016ec",
4304 => x"0000138d",
4305 => x"000017af",
4306 => x"0000178a",
4307 => x"0000178a",
4308 => x"0000178a",
4309 => x"0000178a",
4310 => x"0000178a",
4311 => x"0000178a",
4312 => x"0000178a",
4313 => x"0000178a",
4314 => x"0000178a",
4315 => x"0000138d",
4316 => x"0000138d",
4317 => x"0000138d",
4318 => x"0000138d",
4319 => x"0000138d",
4320 => x"0000138d",
4321 => x"0000138d",
4322 => x"0000138d",
4323 => x"0000138d",
4324 => x"00001699",
4325 => x"00001326",
4326 => x"0000138d",
4327 => x"0000138d",
4328 => x"0000138d",
4329 => x"0000138d",
4330 => x"0000138d",
4331 => x"0000138d",
4332 => x"0000138d",
4333 => x"0000138d",
4334 => x"0000138d",
4335 => x"0000138d",
4336 => x"000012ec",
4337 => x"0000138d",
4338 => x"0000138d",
4339 => x"0000138d",
4340 => x"00001553",
4341 => x"0000138d",
4342 => x"00001015",
4343 => x"0000138d",
4344 => x"0000138d",
4345 => x"00001733",
4346 => x"0000138d",
4347 => x"0000138d",
4348 => x"0000138d",
4349 => x"0000138d",
4350 => x"0000138d",
4351 => x"0000138d",
4352 => x"0000138d",
4353 => x"0000138d",
4354 => x"0000138d",
4355 => x"0000138d",
4356 => x"00001699",
4357 => x"0000132a",
4358 => x"0000138d",
4359 => x"0000138d",
4360 => x"0000138d",
4361 => x"0000168e",
4362 => x"0000132a",
4363 => x"0000138d",
4364 => x"0000138d",
4365 => x"000015d8",
4366 => x"0000138d",
4367 => x"000015a8",
4368 => x"000012f0",
4369 => x"000015f7",
4370 => x"00001383",
4371 => x"0000138d",
4372 => x"00001553",
4373 => x"0000138d",
4374 => x"00001019",
4375 => x"0000138d",
4376 => x"0000138d",
4377 => x"000017ba",
4378 => x"62756720",
4379 => x"696e2076",
4380 => x"66707269",
4381 => x"6e74663a",
4382 => x"20626164",
4383 => x"20626173",
4384 => x"65000000",
4385 => x"30313233",
4386 => x"34353637",
4387 => x"38396162",
4388 => x"63646566",
4389 => x"00000000",
4390 => x"30313233",
4391 => x"34353637",
4392 => x"38394142",
4393 => x"43444546",
4394 => x"00000000",
4395 => x"286e756c",
4396 => x"6c290000",
4397 => x"432d5554",
4398 => x"462d3800",
4399 => x"432d534a",
4400 => x"49530000",
4401 => x"432d4555",
4402 => x"434a5000",
4403 => x"432d4a49",
4404 => x"53000000",
4405 => x"43000000",
4406 => x"2e000000",
4407 => x"49534f2d",
4408 => x"38383539",
4409 => x"2d310000",
4410 => x"64756d6d",
4411 => x"792e6578",
4412 => x"65000000",
4413 => x"00ffffff",
4414 => x"ff00ffff",
4415 => x"ffff00ff",
4416 => x"ffffff00",
4417 => x"00000000",
4418 => x"00000000",
4419 => x"00000000",
4420 => x"00004d08",
4421 => x"00004518",
4422 => x"00000000",
4423 => x"00004780",
4424 => x"000047dc",
4425 => x"00004838",
4426 => x"00000000",
4427 => x"00000000",
4428 => x"00000000",
4429 => x"00000000",
4430 => x"00000000",
4431 => x"00000000",
4432 => x"00000000",
4433 => x"00000000",
4434 => x"00000000",
4435 => x"000044d4",
4436 => x"00000000",
4437 => x"00000000",
4438 => x"00000000",
4439 => x"00000000",
4440 => x"00000000",
4441 => x"00000000",
4442 => x"00000000",
4443 => x"00000000",
4444 => x"00000000",
4445 => x"00000000",
4446 => x"00000000",
4447 => x"00000000",
4448 => x"00000000",
4449 => x"00000000",
4450 => x"00000000",
4451 => x"00000000",
4452 => x"00000000",
4453 => x"00000000",
4454 => x"00000000",
4455 => x"00000000",
4456 => x"00000000",
4457 => x"00000000",
4458 => x"00000000",
4459 => x"00000000",
4460 => x"00000000",
4461 => x"00000000",
4462 => x"00000000",
4463 => x"00000000",
4464 => x"00000001",
4465 => x"330eabcd",
4466 => x"1234e66d",
4467 => x"deec0005",
4468 => x"000b0000",
4469 => x"00000000",
4470 => x"00000000",
4471 => x"00000000",
4472 => x"00000000",
4473 => x"00000000",
4474 => x"00000000",
4475 => x"00000000",
4476 => x"00000000",
4477 => x"00000000",
4478 => x"00000000",
4479 => x"00000000",
4480 => x"00000000",
4481 => x"00000000",
4482 => x"00000000",
4483 => x"00000000",
4484 => x"00000000",
4485 => x"00000000",
4486 => x"00000000",
4487 => x"00000000",
4488 => x"00000000",
4489 => x"00000000",
4490 => x"00000000",
4491 => x"00000000",
4492 => x"00000000",
4493 => x"00000000",
4494 => x"00000000",
4495 => x"00000000",
4496 => x"00000000",
4497 => x"00000000",
4498 => x"00000000",
4499 => x"00000000",
4500 => x"00000000",
4501 => x"00000000",
4502 => x"00000000",
4503 => x"00000000",
4504 => x"00000000",
4505 => x"00000000",
4506 => x"00000000",
4507 => x"00000000",
4508 => x"00000000",
4509 => x"00000000",
4510 => x"00000000",
4511 => x"00000000",
4512 => x"00000000",
4513 => x"00000000",
4514 => x"00000000",
4515 => x"00000000",
4516 => x"00000000",
4517 => x"00000000",
4518 => x"00000000",
4519 => x"00000000",
4520 => x"00000000",
4521 => x"00000000",
4522 => x"00000000",
4523 => x"00000000",
4524 => x"00000000",
4525 => x"00000000",
4526 => x"00000000",
4527 => x"00000000",
4528 => x"00000000",
4529 => x"00000000",
4530 => x"00000000",
4531 => x"00000000",
4532 => x"00000000",
4533 => x"00000000",
4534 => x"00000000",
4535 => x"00000000",
4536 => x"00000000",
4537 => x"00000000",
4538 => x"00000000",
4539 => x"00000000",
4540 => x"00000000",
4541 => x"00000000",
4542 => x"00000000",
4543 => x"00000000",
4544 => x"00000000",
4545 => x"00000000",
4546 => x"00000000",
4547 => x"00000000",
4548 => x"00000000",
4549 => x"00000000",
4550 => x"00000000",
4551 => x"00000000",
4552 => x"00000000",
4553 => x"00000000",
4554 => x"00000000",
4555 => x"00000000",
4556 => x"00000000",
4557 => x"00000000",
4558 => x"00000000",
4559 => x"00000000",
4560 => x"00000000",
4561 => x"00000000",
4562 => x"00000000",
4563 => x"00000000",
4564 => x"00000000",
4565 => x"00000000",
4566 => x"00000000",
4567 => x"00000000",
4568 => x"00000000",
4569 => x"00000000",
4570 => x"00000000",
4571 => x"00000000",
4572 => x"00000000",
4573 => x"00000000",
4574 => x"00000000",
4575 => x"00000000",
4576 => x"00000000",
4577 => x"00000000",
4578 => x"00000000",
4579 => x"00000000",
4580 => x"00000000",
4581 => x"00000000",
4582 => x"00000000",
4583 => x"00000000",
4584 => x"00000000",
4585 => x"00000000",
4586 => x"00000000",
4587 => x"00000000",
4588 => x"00000000",
4589 => x"00000000",
4590 => x"00000000",
4591 => x"00000000",
4592 => x"00000000",
4593 => x"00000000",
4594 => x"00000000",
4595 => x"00000000",
4596 => x"00000000",
4597 => x"00000000",
4598 => x"00000000",
4599 => x"00000000",
4600 => x"00000000",
4601 => x"00000000",
4602 => x"00000000",
4603 => x"00000000",
4604 => x"00000000",
4605 => x"00000000",
4606 => x"00000000",
4607 => x"00000000",
4608 => x"00000000",
4609 => x"00000000",
4610 => x"00000000",
4611 => x"00000000",
4612 => x"00000000",
4613 => x"00000000",
4614 => x"00000000",
4615 => x"00000000",
4616 => x"00000000",
4617 => x"00000000",
4618 => x"00000000",
4619 => x"00000000",
4620 => x"00000000",
4621 => x"00000000",
4622 => x"00000000",
4623 => x"00000000",
4624 => x"00000000",
4625 => x"00000000",
4626 => x"00000000",
4627 => x"00000000",
4628 => x"00000000",
4629 => x"00000000",
4630 => x"00000000",
4631 => x"00000000",
4632 => x"00000000",
4633 => x"00000000",
4634 => x"00000000",
4635 => x"00000000",
4636 => x"00000000",
4637 => x"00000000",
4638 => x"00000000",
4639 => x"00000000",
4640 => x"00000000",
4641 => x"00000000",
4642 => x"00000000",
4643 => x"00000000",
4644 => x"00000000",
4645 => x"43000000",
4646 => x"00000000",
4647 => x"00000000",
4648 => x"00000000",
4649 => x"00000000",
4650 => x"00000000",
4651 => x"00000001",
4652 => x"000044dc",
4653 => x"00000000",
4654 => x"00000000",
4655 => x"00000000",
4656 => x"00000000",
4657 => x"00000000",
4658 => x"00000000",
4659 => x"00000000",
4660 => x"00000000",
4661 => x"00000000",
4662 => x"00000000",
4663 => x"00000000",
4664 => x"00000000",
4665 => x"ffffffff",
4666 => x"00000000",
4667 => x"00020000",
4668 => x"00000000",
4669 => x"00000000",
4670 => x"000048f0",
4671 => x"000048f0",
4672 => x"000048f8",
4673 => x"000048f8",
4674 => x"00004900",
4675 => x"00004900",
4676 => x"00004908",
4677 => x"00004908",
4678 => x"00004910",
4679 => x"00004910",
4680 => x"00004918",
4681 => x"00004918",
4682 => x"00004920",
4683 => x"00004920",
4684 => x"00004928",
4685 => x"00004928",
4686 => x"00004930",
4687 => x"00004930",
4688 => x"00004938",
4689 => x"00004938",
4690 => x"00004940",
4691 => x"00004940",
4692 => x"00004948",
4693 => x"00004948",
4694 => x"00004950",
4695 => x"00004950",
4696 => x"00004958",
4697 => x"00004958",
4698 => x"00004960",
4699 => x"00004960",
4700 => x"00004968",
4701 => x"00004968",
4702 => x"00004970",
4703 => x"00004970",
4704 => x"00004978",
4705 => x"00004978",
4706 => x"00004980",
4707 => x"00004980",
4708 => x"00004988",
4709 => x"00004988",
4710 => x"00004990",
4711 => x"00004990",
4712 => x"00004998",
4713 => x"00004998",
4714 => x"000049a0",
4715 => x"000049a0",
4716 => x"000049a8",
4717 => x"000049a8",
4718 => x"000049b0",
4719 => x"000049b0",
4720 => x"000049b8",
4721 => x"000049b8",
4722 => x"000049c0",
4723 => x"000049c0",
4724 => x"000049c8",
4725 => x"000049c8",
4726 => x"000049d0",
4727 => x"000049d0",
4728 => x"000049d8",
4729 => x"000049d8",
4730 => x"000049e0",
4731 => x"000049e0",
4732 => x"000049e8",
4733 => x"000049e8",
4734 => x"000049f0",
4735 => x"000049f0",
4736 => x"000049f8",
4737 => x"000049f8",
4738 => x"00004a00",
4739 => x"00004a00",
4740 => x"00004a08",
4741 => x"00004a08",
4742 => x"00004a10",
4743 => x"00004a10",
4744 => x"00004a18",
4745 => x"00004a18",
4746 => x"00004a20",
4747 => x"00004a20",
4748 => x"00004a28",
4749 => x"00004a28",
4750 => x"00004a30",
4751 => x"00004a30",
4752 => x"00004a38",
4753 => x"00004a38",
4754 => x"00004a40",
4755 => x"00004a40",
4756 => x"00004a48",
4757 => x"00004a48",
4758 => x"00004a50",
4759 => x"00004a50",
4760 => x"00004a58",
4761 => x"00004a58",
4762 => x"00004a60",
4763 => x"00004a60",
4764 => x"00004a68",
4765 => x"00004a68",
4766 => x"00004a70",
4767 => x"00004a70",
4768 => x"00004a78",
4769 => x"00004a78",
4770 => x"00004a80",
4771 => x"00004a80",
4772 => x"00004a88",
4773 => x"00004a88",
4774 => x"00004a90",
4775 => x"00004a90",
4776 => x"00004a98",
4777 => x"00004a98",
4778 => x"00004aa0",
4779 => x"00004aa0",
4780 => x"00004aa8",
4781 => x"00004aa8",
4782 => x"00004ab0",
4783 => x"00004ab0",
4784 => x"00004ab8",
4785 => x"00004ab8",
4786 => x"00004ac0",
4787 => x"00004ac0",
4788 => x"00004ac8",
4789 => x"00004ac8",
4790 => x"00004ad0",
4791 => x"00004ad0",
4792 => x"00004ad8",
4793 => x"00004ad8",
4794 => x"00004ae0",
4795 => x"00004ae0",
4796 => x"00004ae8",
4797 => x"00004ae8",
4798 => x"00004af0",
4799 => x"00004af0",
4800 => x"00004af8",
4801 => x"00004af8",
4802 => x"00004b00",
4803 => x"00004b00",
4804 => x"00004b08",
4805 => x"00004b08",
4806 => x"00004b10",
4807 => x"00004b10",
4808 => x"00004b18",
4809 => x"00004b18",
4810 => x"00004b20",
4811 => x"00004b20",
4812 => x"00004b28",
4813 => x"00004b28",
4814 => x"00004b30",
4815 => x"00004b30",
4816 => x"00004b38",
4817 => x"00004b38",
4818 => x"00004b40",
4819 => x"00004b40",
4820 => x"00004b48",
4821 => x"00004b48",
4822 => x"00004b50",
4823 => x"00004b50",
4824 => x"00004b58",
4825 => x"00004b58",
4826 => x"00004b60",
4827 => x"00004b60",
4828 => x"00004b68",
4829 => x"00004b68",
4830 => x"00004b70",
4831 => x"00004b70",
4832 => x"00004b78",
4833 => x"00004b78",
4834 => x"00004b80",
4835 => x"00004b80",
4836 => x"00004b88",
4837 => x"00004b88",
4838 => x"00004b90",
4839 => x"00004b90",
4840 => x"00004b98",
4841 => x"00004b98",
4842 => x"00004ba0",
4843 => x"00004ba0",
4844 => x"00004ba8",
4845 => x"00004ba8",
4846 => x"00004bb0",
4847 => x"00004bb0",
4848 => x"00004bb8",
4849 => x"00004bb8",
4850 => x"00004bc0",
4851 => x"00004bc0",
4852 => x"00004bc8",
4853 => x"00004bc8",
4854 => x"00004bd0",
4855 => x"00004bd0",
4856 => x"00004bd8",
4857 => x"00004bd8",
4858 => x"00004be0",
4859 => x"00004be0",
4860 => x"00004be8",
4861 => x"00004be8",
4862 => x"00004bf0",
4863 => x"00004bf0",
4864 => x"00004bf8",
4865 => x"00004bf8",
4866 => x"00004c00",
4867 => x"00004c00",
4868 => x"00004c08",
4869 => x"00004c08",
4870 => x"00004c10",
4871 => x"00004c10",
4872 => x"00004c18",
4873 => x"00004c18",
4874 => x"00004c20",
4875 => x"00004c20",
4876 => x"00004c28",
4877 => x"00004c28",
4878 => x"00004c30",
4879 => x"00004c30",
4880 => x"00004c38",
4881 => x"00004c38",
4882 => x"00004c40",
4883 => x"00004c40",
4884 => x"00004c48",
4885 => x"00004c48",
4886 => x"00004c50",
4887 => x"00004c50",
4888 => x"00004c58",
4889 => x"00004c58",
4890 => x"00004c60",
4891 => x"00004c60",
4892 => x"00004c68",
4893 => x"00004c68",
4894 => x"00004c70",
4895 => x"00004c70",
4896 => x"00004c78",
4897 => x"00004c78",
4898 => x"00004c80",
4899 => x"00004c80",
4900 => x"00004c88",
4901 => x"00004c88",
4902 => x"00004c90",
4903 => x"00004c90",
4904 => x"00004c98",
4905 => x"00004c98",
4906 => x"00004ca0",
4907 => x"00004ca0",
4908 => x"00004ca8",
4909 => x"00004ca8",
4910 => x"00004cb0",
4911 => x"00004cb0",
4912 => x"00004cb8",
4913 => x"00004cb8",
4914 => x"00004cc0",
4915 => x"00004cc0",
4916 => x"00004cc8",
4917 => x"00004cc8",
4918 => x"00004cd0",
4919 => x"00004cd0",
4920 => x"00004cd8",
4921 => x"00004cd8",
4922 => x"00004ce0",
4923 => x"00004ce0",
4924 => x"00004ce8",
4925 => x"00004ce8",
4926 => x"000044e8",
4927 => x"ffffffff",
4928 => x"00000000",
4929 => x"ffffffff",
4930 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(conv_integer(memAAddr)) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(conv_integer(memAAddr));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(conv_integer(memBAddr)) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(conv_integer(memBAddr));
		end if;
	end if;
end process;




end dualport_ram_arch;
