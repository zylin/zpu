-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"0b0b0b0b",
1 => x"80700b0b",
2 => x"80e2a40c",
3 => x"3a0b0b80",
4 => x"c6fc0400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"80c7c32d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80e2",
162 => x"90738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0baf",
171 => x"ac2d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0baf",
179 => x"f02d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80e2a00c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83d93f80",
257 => x"cbcf3f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"ff3d0d0b",
281 => x"0b80f294",
282 => x"08528412",
283 => x"08708106",
284 => x"515170f6",
285 => x"38710881",
286 => x"ff06800c",
287 => x"833d0d04",
288 => x"ff3d0d0b",
289 => x"0b80f294",
290 => x"08528412",
291 => x"08700a10",
292 => x"0a708106",
293 => x"51515170",
294 => x"f1387372",
295 => x"0c833d0d",
296 => x"0480e2a0",
297 => x"08802ea8",
298 => x"38838080",
299 => x"0b0b0b80",
300 => x"f2940c82",
301 => x"a0800b0b",
302 => x"0b80f298",
303 => x"0c829080",
304 => x"0b80f2a8",
305 => x"0c0b0b80",
306 => x"f29c0b80",
307 => x"f2ac0c04",
308 => x"f8808080",
309 => x"a40b0b0b",
310 => x"80f2940c",
311 => x"f8808082",
312 => x"800b0b0b",
313 => x"80f2980c",
314 => x"f8808084",
315 => x"800b80f2",
316 => x"a80cf880",
317 => x"8080940b",
318 => x"80f2ac0c",
319 => x"f8808080",
320 => x"9c0b80f2",
321 => x"a40cf880",
322 => x"8080a00b",
323 => x"80f2b00c",
324 => x"04f23d0d",
325 => x"600b0b80",
326 => x"f2980856",
327 => x"5d82750c",
328 => x"8059805a",
329 => x"800b8f3d",
330 => x"71101017",
331 => x"70085957",
332 => x"5d5b8076",
333 => x"81ff067c",
334 => x"832b5658",
335 => x"5276537b",
336 => x"519af33f",
337 => x"7d7f7a72",
338 => x"077c7207",
339 => x"71716081",
340 => x"05415f5d",
341 => x"5b595755",
342 => x"7a8724bb",
343 => x"380b0b80",
344 => x"f298087b",
345 => x"10101170",
346 => x"08585155",
347 => x"807681ff",
348 => x"067c832b",
349 => x"56585276",
350 => x"537b519a",
351 => x"b93f7d7f",
352 => x"7a72077c",
353 => x"72077171",
354 => x"60810541",
355 => x"5f5d5b59",
356 => x"5755877b",
357 => x"25c73876",
358 => x"7d0c7784",
359 => x"1e0c7c80",
360 => x"0c903d0d",
361 => x"04ff3d0d",
362 => x"80f2a033",
363 => x"5170a738",
364 => x"80e2ac08",
365 => x"70085252",
366 => x"70802e94",
367 => x"38841280",
368 => x"e2ac0c70",
369 => x"2d80e2ac",
370 => x"08700852",
371 => x"5270ee38",
372 => x"810b80f2",
373 => x"a034833d",
374 => x"0d040480",
375 => x"3d0d0b0b",
376 => x"80f29008",
377 => x"802e8e38",
378 => x"0b0b0b0b",
379 => x"800b802e",
380 => x"09810685",
381 => x"38823d0d",
382 => x"040b0b80",
383 => x"f290510b",
384 => x"0b0bf3fc",
385 => x"3f823d0d",
386 => x"0404ff3d",
387 => x"0d028f05",
388 => x"3352718a",
389 => x"2e8a3871",
390 => x"51fce53f",
391 => x"833d0d04",
392 => x"8d51fcdc",
393 => x"3f7151fc",
394 => x"d73f833d",
395 => x"0d04ce3d",
396 => x"0db53d70",
397 => x"70840552",
398 => x"088c8a5c",
399 => x"56a53d5e",
400 => x"5c807570",
401 => x"81055733",
402 => x"765b5558",
403 => x"73782e80",
404 => x"c1388e3d",
405 => x"5b73a52e",
406 => x"09810680",
407 => x"c5387870",
408 => x"81055a33",
409 => x"547380e4",
410 => x"2e81b638",
411 => x"7380e424",
412 => x"80c63873",
413 => x"80e32ea1",
414 => x"388052a5",
415 => x"51792d80",
416 => x"52735179",
417 => x"2d821858",
418 => x"78708105",
419 => x"5a335473",
420 => x"c4387780",
421 => x"0cb43d0d",
422 => x"047b841d",
423 => x"83123356",
424 => x"5d578052",
425 => x"7351792d",
426 => x"81187970",
427 => x"81055b33",
428 => x"555873ff",
429 => x"a038db39",
430 => x"7380f32e",
431 => x"098106ff",
432 => x"b8387b84",
433 => x"1d710859",
434 => x"5d568077",
435 => x"33555673",
436 => x"762e8d38",
437 => x"81167018",
438 => x"70335755",
439 => x"5674f538",
440 => x"ff165580",
441 => x"7625ffa0",
442 => x"38767081",
443 => x"05583354",
444 => x"80527351",
445 => x"792d8118",
446 => x"75ff1757",
447 => x"57588076",
448 => x"25ff8538",
449 => x"76708105",
450 => x"58335480",
451 => x"52735179",
452 => x"2d811875",
453 => x"ff175757",
454 => x"58758024",
455 => x"cc38fee8",
456 => x"397b841d",
457 => x"71087071",
458 => x"9f2c5953",
459 => x"595d5680",
460 => x"75248195",
461 => x"38757d7c",
462 => x"58565480",
463 => x"5773772e",
464 => x"098106b6",
465 => x"38b07b34",
466 => x"02b50556",
467 => x"7a762e97",
468 => x"38ff1656",
469 => x"75337570",
470 => x"81055734",
471 => x"8117577a",
472 => x"762e0981",
473 => x"06eb3880",
474 => x"7534767d",
475 => x"ff125758",
476 => x"56758024",
477 => x"fef338fe",
478 => x"8f398a52",
479 => x"7351a0f0",
480 => x"3f80080b",
481 => x"0b80d484",
482 => x"05337670",
483 => x"81055834",
484 => x"8a527351",
485 => x"a0963f80",
486 => x"08548008",
487 => x"802effac",
488 => x"388a5273",
489 => x"51a0c93f",
490 => x"80080b0b",
491 => x"80d48405",
492 => x"33767081",
493 => x"0558348a",
494 => x"5273519f",
495 => x"ef3f8008",
496 => x"548008ff",
497 => x"b538ff84",
498 => x"39745276",
499 => x"53b43dff",
500 => x"b8055195",
501 => x"b63fa33d",
502 => x"0856fed9",
503 => x"39803d0d",
504 => x"80c10b81",
505 => x"c0f43480",
506 => x"0b81c2d0",
507 => x"0c70800c",
508 => x"823d0d04",
509 => x"ff3d0d80",
510 => x"0b81c0f4",
511 => x"33525270",
512 => x"80c12e99",
513 => x"387181c2",
514 => x"d0080781",
515 => x"c2d00c80",
516 => x"c20b81c0",
517 => x"f8347080",
518 => x"0c833d0d",
519 => x"04810b81",
520 => x"c2d00807",
521 => x"81c2d00c",
522 => x"80c20b81",
523 => x"c0f83470",
524 => x"800c833d",
525 => x"0d04fd3d",
526 => x"0d757008",
527 => x"8a055353",
528 => x"81c0f433",
529 => x"517080c1",
530 => x"2e8b3873",
531 => x"f3387080",
532 => x"0c853d0d",
533 => x"04ff1270",
534 => x"81c0f008",
535 => x"31740c80",
536 => x"0c853d0d",
537 => x"04fc3d0d",
538 => x"81c0fc08",
539 => x"5574802e",
540 => x"8c387675",
541 => x"08710c81",
542 => x"c0fc0856",
543 => x"548c1553",
544 => x"81c0f008",
545 => x"528a5190",
546 => x"f03f7380",
547 => x"0c863d0d",
548 => x"04fb3d0d",
549 => x"77700856",
550 => x"56b05381",
551 => x"c0fc0852",
552 => x"7451acb4",
553 => x"3f850b8c",
554 => x"170c850b",
555 => x"8c160c75",
556 => x"08750c81",
557 => x"c0fc0854",
558 => x"73802e8a",
559 => x"38730875",
560 => x"0c81c0fc",
561 => x"08548c14",
562 => x"5381c0f0",
563 => x"08528a51",
564 => x"90a73f84",
565 => x"1508ad38",
566 => x"860b8c16",
567 => x"0c881552",
568 => x"88160851",
569 => x"8fb33f81",
570 => x"c0fc0870",
571 => x"08760c54",
572 => x"8c157054",
573 => x"548a5273",
574 => x"08518ffd",
575 => x"3f73800c",
576 => x"873d0d04",
577 => x"750854b0",
578 => x"53735275",
579 => x"51abc93f",
580 => x"73800c87",
581 => x"3d0d04d9",
582 => x"3d0db051",
583 => x"9eeb3f80",
584 => x"0881c0ec",
585 => x"0cb0519e",
586 => x"e03f8008",
587 => x"81c0fc0c",
588 => x"81c0ec08",
589 => x"80080c80",
590 => x"0b800884",
591 => x"050c820b",
592 => x"80088805",
593 => x"0ca80b80",
594 => x"088c050c",
595 => x"9f530b0b",
596 => x"80d49052",
597 => x"80089005",
598 => x"51aafd3f",
599 => x"a13d5e9f",
600 => x"530b0b80",
601 => x"d4b0527d",
602 => x"51aaed3f",
603 => x"8a0b80ff",
604 => x"b00c0b0b",
605 => x"80ded451",
606 => x"f9b43f0b",
607 => x"0b80d4d0",
608 => x"51f9ab3f",
609 => x"0b0b80de",
610 => x"d451f9a2",
611 => x"3f80e2b4",
612 => x"08802e8a",
613 => x"cf380b0b",
614 => x"80d58051",
615 => x"f9903f0b",
616 => x"0b80ded4",
617 => x"51f9873f",
618 => x"80e2b008",
619 => x"520b0b80",
620 => x"d5ac51f8",
621 => x"f93f80f2",
622 => x"cc51bbf8",
623 => x"3f810b9a",
624 => x"3d5e5b80",
625 => x"0b80e2b0",
626 => x"082582d6",
627 => x"38903d5f",
628 => x"80c10b81",
629 => x"c0f43481",
630 => x"0b81c2d0",
631 => x"0c80c20b",
632 => x"81c0f834",
633 => x"8240835a",
634 => x"9f530b0b",
635 => x"80d5dc52",
636 => x"7c51a9e4",
637 => x"3f814180",
638 => x"7d537e52",
639 => x"568f9e3f",
640 => x"8008762e",
641 => x"09810683",
642 => x"38815675",
643 => x"81c2d00c",
644 => x"7f705856",
645 => x"758325a2",
646 => x"38751010",
647 => x"16fd0542",
648 => x"a93dffa4",
649 => x"05538352",
650 => x"76518dcd",
651 => x"3f7f8105",
652 => x"70417058",
653 => x"56837624",
654 => x"e0386154",
655 => x"755380f2",
656 => x"d45281c1",
657 => x"88518dc1",
658 => x"3f81c0fc",
659 => x"08700858",
660 => x"58b05377",
661 => x"527651a8",
662 => x"ff3f850b",
663 => x"8c190c85",
664 => x"0b8c180c",
665 => x"7708770c",
666 => x"81c0fc08",
667 => x"5675802e",
668 => x"8a387508",
669 => x"770c81c0",
670 => x"fc08568c",
671 => x"165381c0",
672 => x"f008528a",
673 => x"518cf23f",
674 => x"84170888",
675 => x"e038860b",
676 => x"8c180c88",
677 => x"17528818",
678 => x"08518bfd",
679 => x"3f81c0fc",
680 => x"08700878",
681 => x"0c568c17",
682 => x"7054598a",
683 => x"52780851",
684 => x"8cc73f80",
685 => x"c10b81c0",
686 => x"f8335757",
687 => x"767626a2",
688 => x"3880c352",
689 => x"76518dab",
690 => x"3f800861",
691 => x"2e8aec38",
692 => x"81177081",
693 => x"ff0681c0",
694 => x"f8335858",
695 => x"58757727",
696 => x"e0387960",
697 => x"29627054",
698 => x"71535b59",
699 => x"99be3f80",
700 => x"0840787a",
701 => x"31708729",
702 => x"80083180",
703 => x"088a0581",
704 => x"c0f43381",
705 => x"c0f0085e",
706 => x"5b525a56",
707 => x"7780c12e",
708 => x"8ad8387b",
709 => x"f738811b",
710 => x"5b80e2b0",
711 => x"087b25fd",
712 => x"af3881c0",
713 => x"e451b98c",
714 => x"3f0b0b80",
715 => x"d5fc51f5",
716 => x"fd3f0b0b",
717 => x"80ded451",
718 => x"f5f43f0b",
719 => x"0b80d68c",
720 => x"51f5eb3f",
721 => x"0b0b80de",
722 => x"d451f5e2",
723 => x"3f81c0f0",
724 => x"08520b0b",
725 => x"80d6c451",
726 => x"f5d43f85",
727 => x"520b0b80",
728 => x"d6e051f5",
729 => x"c93f81c2",
730 => x"d008520b",
731 => x"0b80d6fc",
732 => x"51f5bb3f",
733 => x"81520b0b",
734 => x"80d6e051",
735 => x"f5b03f81",
736 => x"c0f43352",
737 => x"0b0b80d7",
738 => x"9851f5a2",
739 => x"3f80c152",
740 => x"0b0b80d7",
741 => x"b451f596",
742 => x"3f81c0f8",
743 => x"33520b0b",
744 => x"80d7d051",
745 => x"f5883f80",
746 => x"c2520b0b",
747 => x"80d7b451",
748 => x"f4fc3f81",
749 => x"c1a80852",
750 => x"0b0b80d7",
751 => x"ec51f4ee",
752 => x"3f87520b",
753 => x"0b80d6e0",
754 => x"51f4e33f",
755 => x"80ffb008",
756 => x"520b0b80",
757 => x"d88851f4",
758 => x"d53f0b0b",
759 => x"80d8a451",
760 => x"f4cc3f0b",
761 => x"0b80d8d0",
762 => x"51f4c33f",
763 => x"81c0fc08",
764 => x"7008535a",
765 => x"0b0b80d8",
766 => x"dc51f4b2",
767 => x"3f0b0b80",
768 => x"d8f851f4",
769 => x"a93f81c0",
770 => x"fc088411",
771 => x"0853560b",
772 => x"0b80d9ac",
773 => x"51f4973f",
774 => x"80520b0b",
775 => x"80d6e051",
776 => x"f48c3f81",
777 => x"c0fc0888",
778 => x"11085358",
779 => x"0b0b80d9",
780 => x"c851f3fa",
781 => x"3f82520b",
782 => x"0b80d6e0",
783 => x"51f3ef3f",
784 => x"81c0fc08",
785 => x"8c110853",
786 => x"570b0b80",
787 => x"d9e451f3",
788 => x"dd3f9152",
789 => x"0b0b80d6",
790 => x"e051f3d2",
791 => x"3f81c0fc",
792 => x"08900552",
793 => x"0b0b80da",
794 => x"8051f3c2",
795 => x"3f0b0b80",
796 => x"da9c51f3",
797 => x"b93f0b0b",
798 => x"80dad451",
799 => x"f3b03f81",
800 => x"c0ec0870",
801 => x"08535f0b",
802 => x"0b80d8dc",
803 => x"51f39f3f",
804 => x"0b0b80da",
805 => x"e851f396",
806 => x"3f81c0ec",
807 => x"08841108",
808 => x"535b0b0b",
809 => x"80d9ac51",
810 => x"f3843f80",
811 => x"520b0b80",
812 => x"d6e051f2",
813 => x"f93f81c0",
814 => x"ec088811",
815 => x"08535c0b",
816 => x"0b80d9c8",
817 => x"51f2e73f",
818 => x"81520b0b",
819 => x"80d6e051",
820 => x"f2dc3f81",
821 => x"c0ec088c",
822 => x"1108535a",
823 => x"0b0b80d9",
824 => x"e451f2ca",
825 => x"3f92520b",
826 => x"0b80d6e0",
827 => x"51f2bf3f",
828 => x"81c0ec08",
829 => x"9005520b",
830 => x"0b80da80",
831 => x"51f2af3f",
832 => x"0b0b80da",
833 => x"9c51f2a6",
834 => x"3f7f520b",
835 => x"0b80dba8",
836 => x"51f29b3f",
837 => x"85520b0b",
838 => x"80d6e051",
839 => x"f2903f78",
840 => x"520b0b80",
841 => x"dbc451f2",
842 => x"853f8d52",
843 => x"0b0b80d6",
844 => x"e051f1fa",
845 => x"3f61520b",
846 => x"0b80dbe0",
847 => x"51f1ef3f",
848 => x"87520b0b",
849 => x"80d6e051",
850 => x"f1e43f60",
851 => x"520b0b80",
852 => x"dbfc51f1",
853 => x"d93f8152",
854 => x"0b0b80d6",
855 => x"e051f1ce",
856 => x"3f7d520b",
857 => x"0b80dc98",
858 => x"51f1c33f",
859 => x"0b0b80dc",
860 => x"b451f1ba",
861 => x"3f7c520b",
862 => x"0b80dcec",
863 => x"51f1af3f",
864 => x"0b0b80dd",
865 => x"8851f1a6",
866 => x"3f0b0b80",
867 => x"ded451f1",
868 => x"9d3f81c0",
869 => x"e40881c0",
870 => x"e80880f2",
871 => x"cc0880f2",
872 => x"d0087271",
873 => x"31707426",
874 => x"75743170",
875 => x"723180f2",
876 => x"c40c4444",
877 => x"80f2c80c",
878 => x"80f2c808",
879 => x"560b0b80",
880 => x"ddc0555c",
881 => x"595758f0",
882 => x"e53f80f2",
883 => x"c4085680",
884 => x"762582b1",
885 => x"3880e2b0",
886 => x"0870719f",
887 => x"2c9a3d53",
888 => x"565680f2",
889 => x"c40880f2",
890 => x"c8084153",
891 => x"7f547052",
892 => x"5a8a8d3f",
893 => x"66685f80",
894 => x"f2b40c7d",
895 => x"80f2b80c",
896 => x"80e2b008",
897 => x"709f2c58",
898 => x"568058bd",
899 => x"84c07855",
900 => x"55765275",
901 => x"53795187",
902 => x"f33f953d",
903 => x"80f2c408",
904 => x"80f2c808",
905 => x"41557f56",
906 => x"67694053",
907 => x"7e547052",
908 => x"5c89cd3f",
909 => x"64665e80",
910 => x"f2bc0c7c",
911 => x"80f2c00c",
912 => x"80e2b008",
913 => x"709f2c40",
914 => x"58805783",
915 => x"dceb9480",
916 => x"7755557e",
917 => x"5277537b",
918 => x"5187b13f",
919 => x"64665d5b",
920 => x"805e8ddd",
921 => x"7e555580",
922 => x"f2c40880",
923 => x"f2c80859",
924 => x"52775379",
925 => x"5187953f",
926 => x"66684054",
927 => x"7e557a52",
928 => x"7b53a93d",
929 => x"ffa80551",
930 => x"88f63f62",
931 => x"645e81c1",
932 => x"800c7c81",
933 => x"c1840c0b",
934 => x"0b80ddd0",
935 => x"51ef8f3f",
936 => x"80f2b808",
937 => x"520b0b80",
938 => x"de8051ef",
939 => x"813f0b0b",
940 => x"80de8851",
941 => x"eef83f80",
942 => x"f2c00852",
943 => x"0b0b80de",
944 => x"8051eeea",
945 => x"3f81c184",
946 => x"08520b0b",
947 => x"80deb851",
948 => x"eedc3f0b",
949 => x"0b80ded4",
950 => x"51eed33f",
951 => x"800b800c",
952 => x"a93d0d04",
953 => x"0b0b80de",
954 => x"d851f5b0",
955 => x"39770857",
956 => x"b0537652",
957 => x"77519fe0",
958 => x"3f80c10b",
959 => x"81c0f833",
960 => x"5757f7b8",
961 => x"39758a38",
962 => x"80f2c808",
963 => x"8126fdc5",
964 => x"380b0b80",
965 => x"df8851ee",
966 => x"953f0b0b",
967 => x"80dfc051",
968 => x"ee8c3f0b",
969 => x"0b80ded4",
970 => x"51ee833f",
971 => x"80e2b008",
972 => x"70719f2c",
973 => x"9a3d5356",
974 => x"5680f2c4",
975 => x"0880f2c8",
976 => x"0841537f",
977 => x"5470525a",
978 => x"87b63f66",
979 => x"685f80f2",
980 => x"b40c7d80",
981 => x"f2b80c80",
982 => x"e2b00870",
983 => x"9f2c5856",
984 => x"8058bd84",
985 => x"c0785555",
986 => x"76527553",
987 => x"7951859c",
988 => x"3f953d80",
989 => x"f2c40880",
990 => x"f2c80841",
991 => x"557f5667",
992 => x"6940537e",
993 => x"5470525c",
994 => x"86f63f64",
995 => x"665e80f2",
996 => x"bc0c7c80",
997 => x"f2c00c80",
998 => x"e2b00870",
999 => x"9f2c4058",
1000 => x"805783dc",
1001 => x"eb948077",
1002 => x"55557e52",
1003 => x"77537b51",
1004 => x"84da3f64",
1005 => x"665d5b80",
1006 => x"5e8ddd7e",
1007 => x"555580f2",
1008 => x"c40880f2",
1009 => x"c8085952",
1010 => x"77537951",
1011 => x"84be3f66",
1012 => x"6840547e",
1013 => x"557a527b",
1014 => x"53a93dff",
1015 => x"a8055186",
1016 => x"9f3f6264",
1017 => x"5e81c180",
1018 => x"0c7c81c1",
1019 => x"840c0b0b",
1020 => x"80ddd051",
1021 => x"ecb83f80",
1022 => x"f2b80852",
1023 => x"0b0b80de",
1024 => x"8051ecaa",
1025 => x"3f0b0b80",
1026 => x"de8851ec",
1027 => x"a13f80f2",
1028 => x"c008520b",
1029 => x"0b80de80",
1030 => x"51ec933f",
1031 => x"81c18408",
1032 => x"520b0b80",
1033 => x"deb851ec",
1034 => x"853f0b0b",
1035 => x"80ded451",
1036 => x"ebfc3f80",
1037 => x"0b800ca9",
1038 => x"3d0d04a9",
1039 => x"3dffa005",
1040 => x"52805180",
1041 => x"d43f9f53",
1042 => x"0b0b80df",
1043 => x"e0527c51",
1044 => x"9d863f7a",
1045 => x"7b81c0f0",
1046 => x"0c811870",
1047 => x"81ff0681",
1048 => x"c0f83359",
1049 => x"59595af4",
1050 => x"f439ff16",
1051 => x"707b3160",
1052 => x"0c5c800b",
1053 => x"811c5c5c",
1054 => x"80e2b008",
1055 => x"7b25f2d0",
1056 => x"38f59f39",
1057 => x"ff3d0d73",
1058 => x"82327030",
1059 => x"70720780",
1060 => x"25800c52",
1061 => x"52833d0d",
1062 => x"04fe3d0d",
1063 => x"74767153",
1064 => x"54527182",
1065 => x"2e833883",
1066 => x"5171812e",
1067 => x"9a388172",
1068 => x"269f3871",
1069 => x"822eb838",
1070 => x"71842ea9",
1071 => x"3870730c",
1072 => x"70800c84",
1073 => x"3d0d0480",
1074 => x"e40b81c0",
1075 => x"f008258b",
1076 => x"3880730c",
1077 => x"70800c84",
1078 => x"3d0d0483",
1079 => x"730c7080",
1080 => x"0c843d0d",
1081 => x"0482730c",
1082 => x"70800c84",
1083 => x"3d0d0481",
1084 => x"730c7080",
1085 => x"0c843d0d",
1086 => x"04803d0d",
1087 => x"74741482",
1088 => x"05710c80",
1089 => x"0c823d0d",
1090 => x"04f73d0d",
1091 => x"7b7d7f61",
1092 => x"85127082",
1093 => x"2b751170",
1094 => x"74717084",
1095 => x"05530c5a",
1096 => x"5a5d5b76",
1097 => x"0c7980f8",
1098 => x"180c7986",
1099 => x"12525758",
1100 => x"5a5a7676",
1101 => x"24993876",
1102 => x"b329822b",
1103 => x"79115153",
1104 => x"76737084",
1105 => x"05550c81",
1106 => x"14547574",
1107 => x"25f23876",
1108 => x"81cc2919",
1109 => x"fc110881",
1110 => x"05fc120c",
1111 => x"7a197008",
1112 => x"9fa0130c",
1113 => x"5856850b",
1114 => x"81c0f00c",
1115 => x"75800c8b",
1116 => x"3d0d04fe",
1117 => x"3d0d0293",
1118 => x"05335180",
1119 => x"02840597",
1120 => x"05335452",
1121 => x"70732e88",
1122 => x"3871800c",
1123 => x"843d0d04",
1124 => x"7081c0f4",
1125 => x"34810b80",
1126 => x"0c843d0d",
1127 => x"04f83d0d",
1128 => x"7a7c5956",
1129 => x"820b8319",
1130 => x"55557416",
1131 => x"70337533",
1132 => x"5b515372",
1133 => x"792e80c6",
1134 => x"3880c10b",
1135 => x"81168116",
1136 => x"56565782",
1137 => x"7525e338",
1138 => x"ffa91770",
1139 => x"81ff0655",
1140 => x"59738226",
1141 => x"83388755",
1142 => x"81537680",
1143 => x"d22e9838",
1144 => x"77527551",
1145 => x"9bc43f80",
1146 => x"53728008",
1147 => x"25893887",
1148 => x"1581c0f0",
1149 => x"0c815372",
1150 => x"800c8a3d",
1151 => x"0d047281",
1152 => x"c0f43482",
1153 => x"7525ffa2",
1154 => x"38ffbd39",
1155 => x"ef3d0d63",
1156 => x"65675b42",
1157 => x"79436769",
1158 => x"59407741",
1159 => x"5a805d80",
1160 => x"5e617083",
1161 => x"ffff0671",
1162 => x"902a6270",
1163 => x"83ffff06",
1164 => x"71902a74",
1165 => x"72297473",
1166 => x"29757329",
1167 => x"77742973",
1168 => x"902a0572",
1169 => x"11515856",
1170 => x"535f5a57",
1171 => x"5a585558",
1172 => x"73732786",
1173 => x"38848080",
1174 => x"16567390",
1175 => x"2a165b78",
1176 => x"83ffff06",
1177 => x"74848080",
1178 => x"29055c7a",
1179 => x"7c5a5d78",
1180 => x"5e777f29",
1181 => x"61782905",
1182 => x"7d055d7c",
1183 => x"7e567a0c",
1184 => x"74841b0c",
1185 => x"79800c93",
1186 => x"3d0d04f9",
1187 => x"3d0d797b",
1188 => x"7d545872",
1189 => x"59773079",
1190 => x"70307072",
1191 => x"079f2a73",
1192 => x"71315a52",
1193 => x"59777956",
1194 => x"730c5373",
1195 => x"84130c54",
1196 => x"800c893d",
1197 => x"0d04f93d",
1198 => x"0d797b7d",
1199 => x"7f565452",
1200 => x"5472802e",
1201 => x"a0387057",
1202 => x"7158a073",
1203 => x"31528072",
1204 => x"25a13877",
1205 => x"70742b57",
1206 => x"70732a78",
1207 => x"752b0756",
1208 => x"51747653",
1209 => x"5170740c",
1210 => x"7184150c",
1211 => x"73800c89",
1212 => x"3d0d0480",
1213 => x"56777230",
1214 => x"2b557476",
1215 => x"5351e639",
1216 => x"e43d0d6e",
1217 => x"a13d08a3",
1218 => x"3d085957",
1219 => x"5f80764d",
1220 => x"774ea33d",
1221 => x"08a53d08",
1222 => x"574b754c",
1223 => x"5e7d6c24",
1224 => x"86fb3880",
1225 => x"6a24878f",
1226 => x"38696b58",
1227 => x"566b6d5d",
1228 => x"467b4775",
1229 => x"44764564",
1230 => x"6468685c",
1231 => x"5c565674",
1232 => x"81e73878",
1233 => x"762782c7",
1234 => x"387581ff",
1235 => x"26832b55",
1236 => x"83ffff76",
1237 => x"278c3890",
1238 => x"55fe800a",
1239 => x"76278338",
1240 => x"98557575",
1241 => x"2a80e080",
1242 => x"057033a0",
1243 => x"77317131",
1244 => x"57555774",
1245 => x"802e9538",
1246 => x"75752ba0",
1247 => x"76317a77",
1248 => x"2b7c722a",
1249 => x"077c782b",
1250 => x"5d5b5956",
1251 => x"75902a76",
1252 => x"83ffff06",
1253 => x"71547a53",
1254 => x"59578880",
1255 => x"3f80085b",
1256 => x"87ea3f80",
1257 => x"08800879",
1258 => x"297c902b",
1259 => x"7c902a07",
1260 => x"56565973",
1261 => x"75279438",
1262 => x"8008ff05",
1263 => x"76155559",
1264 => x"75742687",
1265 => x"38747426",
1266 => x"87b93876",
1267 => x"52737531",
1268 => x"5187c93f",
1269 => x"80085587",
1270 => x"b33f8008",
1271 => x"80087929",
1272 => x"7b83ffff",
1273 => x"0677902b",
1274 => x"07565957",
1275 => x"73782796",
1276 => x"388008ff",
1277 => x"05761555",
1278 => x"57757426",
1279 => x"89387774",
1280 => x"26777131",
1281 => x"58567890",
1282 => x"2b770758",
1283 => x"805b7a40",
1284 => x"77417f61",
1285 => x"56547d80",
1286 => x"d938737f",
1287 => x"0c747f84",
1288 => x"050c7e80",
1289 => x"0c9e3d0d",
1290 => x"0480705c",
1291 => x"58747926",
1292 => x"dd387481",
1293 => x"ff26832b",
1294 => x"577483ff",
1295 => x"ff2682a5",
1296 => x"3874772a",
1297 => x"80e08005",
1298 => x"7033a079",
1299 => x"31713159",
1300 => x"5c5d7682",
1301 => x"b3387654",
1302 => x"74792783",
1303 => x"38815479",
1304 => x"76277407",
1305 => x"59815878",
1306 => x"ffa23876",
1307 => x"58805bff",
1308 => x"9d397352",
1309 => x"74539e3d",
1310 => x"e80551fc",
1311 => x"8e3f6769",
1312 => x"567f0c74",
1313 => x"7f84050c",
1314 => x"7e800c9e",
1315 => x"3d0d0475",
1316 => x"802e81c4",
1317 => x"387581ff",
1318 => x"26832b55",
1319 => x"83ffff76",
1320 => x"278c3890",
1321 => x"55fe800a",
1322 => x"76278338",
1323 => x"98557575",
1324 => x"2a80e080",
1325 => x"057033a0",
1326 => x"77317131",
1327 => x"575e5474",
1328 => x"84913878",
1329 => x"76315481",
1330 => x"76902a77",
1331 => x"83ffff06",
1332 => x"5f5d5b7b",
1333 => x"52735185",
1334 => x"c33f8008",
1335 => x"5785ad3f",
1336 => x"80088008",
1337 => x"7e297890",
1338 => x"2b7c902a",
1339 => x"07565659",
1340 => x"73752794",
1341 => x"388008ff",
1342 => x"05761555",
1343 => x"59757426",
1344 => x"87387474",
1345 => x"2684f338",
1346 => x"7b527375",
1347 => x"3151858c",
1348 => x"3f800855",
1349 => x"84f63f80",
1350 => x"0880087e",
1351 => x"297b83ff",
1352 => x"ff067790",
1353 => x"2b075659",
1354 => x"57737827",
1355 => x"96388008",
1356 => x"ff057615",
1357 => x"55577574",
1358 => x"26893877",
1359 => x"74267771",
1360 => x"31585a78",
1361 => x"902b7707",
1362 => x"7b41417f",
1363 => x"6156547d",
1364 => x"802efdc6",
1365 => x"38fe9b39",
1366 => x"75528151",
1367 => x"84ae3f80",
1368 => x"0856feb1",
1369 => x"399057fe",
1370 => x"800a7527",
1371 => x"fdd33898",
1372 => x"75712a80",
1373 => x"e0800570",
1374 => x"33a07331",
1375 => x"7131535d",
1376 => x"5e577680",
1377 => x"2efdcf38",
1378 => x"a0773175",
1379 => x"782b7772",
1380 => x"2a077779",
1381 => x"2b7b7a2b",
1382 => x"7d742a07",
1383 => x"7d7b2b73",
1384 => x"902a7483",
1385 => x"ffff0671",
1386 => x"597f772a",
1387 => x"585e5c41",
1388 => x"5f585c54",
1389 => x"83e63f80",
1390 => x"085483d0",
1391 => x"3f800880",
1392 => x"08792975",
1393 => x"902b7e90",
1394 => x"2a075656",
1395 => x"59737527",
1396 => x"99388008",
1397 => x"ff057b15",
1398 => x"55597a74",
1399 => x"268c3873",
1400 => x"75278738",
1401 => x"ff197b15",
1402 => x"55597652",
1403 => x"73753151",
1404 => x"83aa3f80",
1405 => x"08558394",
1406 => x"3f800880",
1407 => x"0879297d",
1408 => x"83ffff06",
1409 => x"77902b07",
1410 => x"56595773",
1411 => x"78279938",
1412 => x"8008ff05",
1413 => x"7b155557",
1414 => x"7a74268c",
1415 => x"38737827",
1416 => x"8738ff17",
1417 => x"7b155557",
1418 => x"73783179",
1419 => x"902b7807",
1420 => x"7083ffff",
1421 => x"0671902a",
1422 => x"7983ffff",
1423 => x"067a902a",
1424 => x"73722973",
1425 => x"73297473",
1426 => x"29767429",
1427 => x"73902a05",
1428 => x"72055755",
1429 => x"435f5b58",
1430 => x"5a57595a",
1431 => x"747c2786",
1432 => x"38848080",
1433 => x"17577490",
1434 => x"2a177983",
1435 => x"ffff0676",
1436 => x"84808029",
1437 => x"05575776",
1438 => x"7a269a38",
1439 => x"767a3270",
1440 => x"30707207",
1441 => x"8025565a",
1442 => x"5b7c7627",
1443 => x"fafe3873",
1444 => x"802efaf8",
1445 => x"38ff1858",
1446 => x"805bfaf2",
1447 => x"39ff7653",
1448 => x"77549f3d",
1449 => x"e805525e",
1450 => x"f7e13f67",
1451 => x"69574c75",
1452 => x"4d698025",
1453 => x"f8f3387d",
1454 => x"096a6c5c",
1455 => x"537a549f",
1456 => x"3de80552",
1457 => x"5ef7c43f",
1458 => x"6769714c",
1459 => x"704d5856",
1460 => x"f8db39a0",
1461 => x"75317676",
1462 => x"2b7a772b",
1463 => x"7c732a07",
1464 => x"7c782b72",
1465 => x"902a7383",
1466 => x"ffff0671",
1467 => x"587e762a",
1468 => x"5742405d",
1469 => x"5d575881",
1470 => x"a33f8008",
1471 => x"57818d3f",
1472 => x"80088008",
1473 => x"7e297890",
1474 => x"2b7d902a",
1475 => x"07565659",
1476 => x"73752799",
1477 => x"388008ff",
1478 => x"05761555",
1479 => x"59757426",
1480 => x"8c387375",
1481 => x"278738ff",
1482 => x"19761555",
1483 => x"597b5273",
1484 => x"75315180",
1485 => x"e73f8008",
1486 => x"5580d13f",
1487 => x"80088008",
1488 => x"7e297c83",
1489 => x"ffff0670",
1490 => x"78902b07",
1491 => x"51565858",
1492 => x"73772799",
1493 => x"388008ff",
1494 => x"05761555",
1495 => x"58757426",
1496 => x"8c387377",
1497 => x"278738ff",
1498 => x"18761555",
1499 => x"5878902b",
1500 => x"78077478",
1501 => x"31555bfa",
1502 => x"da39ff19",
1503 => x"76155559",
1504 => x"fb8639ff",
1505 => x"19761555",
1506 => x"59f8c039",
1507 => x"fe3d0d80",
1508 => x"53755274",
1509 => x"5181913f",
1510 => x"843d0d04",
1511 => x"fe3d0d81",
1512 => x"53755274",
1513 => x"5181813f",
1514 => x"843d0d04",
1515 => x"fb3d0d77",
1516 => x"79555580",
1517 => x"56757524",
1518 => x"ab388074",
1519 => x"249d3880",
1520 => x"53735274",
1521 => x"5180e13f",
1522 => x"80085475",
1523 => x"802e8538",
1524 => x"80083054",
1525 => x"73800c87",
1526 => x"3d0d0473",
1527 => x"30768132",
1528 => x"5754dc39",
1529 => x"74305581",
1530 => x"56738025",
1531 => x"d238ec39",
1532 => x"fa3d0d78",
1533 => x"7a575580",
1534 => x"57767524",
1535 => x"a438759f",
1536 => x"2c548153",
1537 => x"75743274",
1538 => x"31527451",
1539 => x"9b3f8008",
1540 => x"5476802e",
1541 => x"85388008",
1542 => x"30547380",
1543 => x"0c883d0d",
1544 => x"04743055",
1545 => x"8157d739",
1546 => x"fc3d0d76",
1547 => x"78535481",
1548 => x"53807473",
1549 => x"26525572",
1550 => x"802e9838",
1551 => x"70802eab",
1552 => x"38807224",
1553 => x"a6387110",
1554 => x"73107572",
1555 => x"26535452",
1556 => x"72ea3873",
1557 => x"51788338",
1558 => x"74517080",
1559 => x"0c863d0d",
1560 => x"04720a10",
1561 => x"0a720a10",
1562 => x"0a535372",
1563 => x"802ee438",
1564 => x"717426ed",
1565 => x"38737231",
1566 => x"75740774",
1567 => x"0a100a74",
1568 => x"0a100a55",
1569 => x"555654e3",
1570 => x"39ff3d0d",
1571 => x"735280ea",
1572 => x"fc085196",
1573 => x"3f833d0d",
1574 => x"04ff3d0d",
1575 => x"735280ea",
1576 => x"fc085190",
1577 => x"cc3f833d",
1578 => x"0d04f43d",
1579 => x"0d7e608b",
1580 => x"1170f806",
1581 => x"5b55555d",
1582 => x"72962683",
1583 => x"38905880",
1584 => x"78247479",
1585 => x"26075580",
1586 => x"5474742e",
1587 => x"09810680",
1588 => x"ca387c51",
1589 => x"8d9e3f77",
1590 => x"83f72680",
1591 => x"c5387783",
1592 => x"2a701010",
1593 => x"1080e2f4",
1594 => x"058c1108",
1595 => x"58585475",
1596 => x"772e81f0",
1597 => x"38841608",
1598 => x"fc068c17",
1599 => x"08881808",
1600 => x"718c120c",
1601 => x"88120c5b",
1602 => x"76058411",
1603 => x"08810784",
1604 => x"120c537c",
1605 => x"518cde3f",
1606 => x"88165473",
1607 => x"800c8e3d",
1608 => x"0d047789",
1609 => x"2a78832a",
1610 => x"58547380",
1611 => x"2ebf3877",
1612 => x"862ab805",
1613 => x"57847427",
1614 => x"b43880db",
1615 => x"14579474",
1616 => x"27ab3877",
1617 => x"8c2a80ee",
1618 => x"055780d4",
1619 => x"74279e38",
1620 => x"778f2a80",
1621 => x"f7055782",
1622 => x"d4742791",
1623 => x"3877922a",
1624 => x"80fc0557",
1625 => x"8ad47427",
1626 => x"843880fe",
1627 => x"57761010",
1628 => x"1080e2f4",
1629 => x"058c1108",
1630 => x"56537473",
1631 => x"2ea33884",
1632 => x"1508fc06",
1633 => x"70793155",
1634 => x"56738f24",
1635 => x"88e43873",
1636 => x"802588e6",
1637 => x"388c1508",
1638 => x"5574732e",
1639 => x"098106df",
1640 => x"38811759",
1641 => x"80e38408",
1642 => x"567580e2",
1643 => x"fc2e82cc",
1644 => x"38841608",
1645 => x"fc067079",
1646 => x"31555573",
1647 => x"8f24bb38",
1648 => x"80e2fc0b",
1649 => x"80e3880c",
1650 => x"80e2fc0b",
1651 => x"80e3840c",
1652 => x"80742480",
1653 => x"db387416",
1654 => x"84110881",
1655 => x"0784120c",
1656 => x"53feb039",
1657 => x"88168c11",
1658 => x"08575975",
1659 => x"792e0981",
1660 => x"06fe8238",
1661 => x"821459ff",
1662 => x"ab397716",
1663 => x"78810784",
1664 => x"180c7080",
1665 => x"e3880c70",
1666 => x"80e3840c",
1667 => x"80e2fc0b",
1668 => x"8c120c8c",
1669 => x"11088812",
1670 => x"0c748107",
1671 => x"84120c74",
1672 => x"0574710c",
1673 => x"5b7c518a",
1674 => x"cc3f8816",
1675 => x"54fdec39",
1676 => x"83ff7527",
1677 => x"83913874",
1678 => x"892a7583",
1679 => x"2a545473",
1680 => x"802ebf38",
1681 => x"74862ab8",
1682 => x"05538474",
1683 => x"27b43880",
1684 => x"db145394",
1685 => x"7427ab38",
1686 => x"748c2a80",
1687 => x"ee055380",
1688 => x"d474279e",
1689 => x"38748f2a",
1690 => x"80f70553",
1691 => x"82d47427",
1692 => x"91387492",
1693 => x"2a80fc05",
1694 => x"538ad474",
1695 => x"27843880",
1696 => x"fe537210",
1697 => x"101080e2",
1698 => x"f4058811",
1699 => x"08555773",
1700 => x"772e868b",
1701 => x"38841408",
1702 => x"fc065b74",
1703 => x"7b278d38",
1704 => x"88140854",
1705 => x"73772e09",
1706 => x"8106ea38",
1707 => x"8c140880",
1708 => x"e2f40b84",
1709 => x"0508718c",
1710 => x"190c7588",
1711 => x"190c7788",
1712 => x"130c5c57",
1713 => x"758c150c",
1714 => x"78538079",
1715 => x"24839838",
1716 => x"72822c81",
1717 => x"712b5656",
1718 => x"747b2680",
1719 => x"ca387a75",
1720 => x"06577682",
1721 => x"a33878fc",
1722 => x"06840559",
1723 => x"7410707c",
1724 => x"06555573",
1725 => x"82923884",
1726 => x"1959f139",
1727 => x"80e2f40b",
1728 => x"84050879",
1729 => x"545b7880",
1730 => x"25c63882",
1731 => x"da397409",
1732 => x"7b067080",
1733 => x"e2f40b84",
1734 => x"050c5b74",
1735 => x"1055747b",
1736 => x"26853874",
1737 => x"85bc3880",
1738 => x"e2f40b88",
1739 => x"05087084",
1740 => x"1208fc06",
1741 => x"707b317b",
1742 => x"72268f72",
1743 => x"25075d57",
1744 => x"5c5c5578",
1745 => x"802e80d9",
1746 => x"38791580",
1747 => x"e2ec0819",
1748 => x"90115954",
1749 => x"5680e2e8",
1750 => x"08ff2e88",
1751 => x"38a08f13",
1752 => x"e0800657",
1753 => x"76527c51",
1754 => x"888c3f80",
1755 => x"08548008",
1756 => x"ff2e9038",
1757 => x"80087627",
1758 => x"82a73874",
1759 => x"80e2f42e",
1760 => x"829f3880",
1761 => x"e2f40b88",
1762 => x"05085584",
1763 => x"1508fc06",
1764 => x"70793179",
1765 => x"72268f72",
1766 => x"25075d55",
1767 => x"5a7a83f2",
1768 => x"38778107",
1769 => x"84160c77",
1770 => x"157080e2",
1771 => x"f40b8805",
1772 => x"0c748107",
1773 => x"84120c56",
1774 => x"7c5187b9",
1775 => x"3f881554",
1776 => x"73800c8e",
1777 => x"3d0d0474",
1778 => x"832a7054",
1779 => x"54807424",
1780 => x"819b3872",
1781 => x"822c8171",
1782 => x"2b80e2f8",
1783 => x"08077080",
1784 => x"e2f40b84",
1785 => x"050c7510",
1786 => x"101080e2",
1787 => x"f4058811",
1788 => x"08718c1b",
1789 => x"0c70881b",
1790 => x"0c798813",
1791 => x"0c57555c",
1792 => x"55758c15",
1793 => x"0cfdc139",
1794 => x"78791010",
1795 => x"1080e2f4",
1796 => x"0570565b",
1797 => x"5c8c1408",
1798 => x"5675742e",
1799 => x"a3388416",
1800 => x"08fc0670",
1801 => x"79315853",
1802 => x"768f2483",
1803 => x"f1387680",
1804 => x"2584af38",
1805 => x"8c160856",
1806 => x"75742e09",
1807 => x"8106df38",
1808 => x"8814811a",
1809 => x"70830655",
1810 => x"5a5472c9",
1811 => x"387b8306",
1812 => x"5675802e",
1813 => x"fdb838ff",
1814 => x"1cf81b5b",
1815 => x"5c881a08",
1816 => x"7a2eea38",
1817 => x"fdb53983",
1818 => x"1953fce4",
1819 => x"39831470",
1820 => x"822c8171",
1821 => x"2b80e2f8",
1822 => x"08077080",
1823 => x"e2f40b84",
1824 => x"050c7610",
1825 => x"101080e2",
1826 => x"f4058811",
1827 => x"08718c1c",
1828 => x"0c70881c",
1829 => x"0c7a8813",
1830 => x"0c58535d",
1831 => x"5653fee1",
1832 => x"3980e2b8",
1833 => x"08175980",
1834 => x"08762e81",
1835 => x"8b3880e2",
1836 => x"e808ff2e",
1837 => x"848e3873",
1838 => x"76311980",
1839 => x"e2b80c73",
1840 => x"87067056",
1841 => x"5372802e",
1842 => x"88388873",
1843 => x"31701555",
1844 => x"5576149f",
1845 => x"ff06a080",
1846 => x"71311670",
1847 => x"547e5351",
1848 => x"5385933f",
1849 => x"80085680",
1850 => x"08ff2e81",
1851 => x"9e3880e2",
1852 => x"b8081370",
1853 => x"80e2b80c",
1854 => x"747580e2",
1855 => x"f40b8805",
1856 => x"0c777631",
1857 => x"15810755",
1858 => x"56597a80",
1859 => x"e2f42e83",
1860 => x"c038798f",
1861 => x"2682ef38",
1862 => x"810b8415",
1863 => x"0c841508",
1864 => x"fc067079",
1865 => x"31797226",
1866 => x"8f722507",
1867 => x"5d555a7a",
1868 => x"802efced",
1869 => x"3880db39",
1870 => x"80089fff",
1871 => x"065574fe",
1872 => x"ed387880",
1873 => x"e2b80c80",
1874 => x"e2f40b88",
1875 => x"05087a18",
1876 => x"81078412",
1877 => x"0c5580e2",
1878 => x"e4087927",
1879 => x"86387880",
1880 => x"e2e40c80",
1881 => x"e2e00879",
1882 => x"27fca038",
1883 => x"7880e2e0",
1884 => x"0c841508",
1885 => x"fc067079",
1886 => x"31797226",
1887 => x"8f722507",
1888 => x"5d555a7a",
1889 => x"802efc99",
1890 => x"38883980",
1891 => x"745753fe",
1892 => x"dd397c51",
1893 => x"83df3f80",
1894 => x"0b800c8e",
1895 => x"3d0d0480",
1896 => x"7324a538",
1897 => x"72822c81",
1898 => x"712b80e2",
1899 => x"f8080770",
1900 => x"80e2f40b",
1901 => x"84050c5c",
1902 => x"5a768c17",
1903 => x"0c738817",
1904 => x"0c758818",
1905 => x"0cf9fd39",
1906 => x"83137082",
1907 => x"2c81712b",
1908 => x"80e2f808",
1909 => x"077080e2",
1910 => x"f40b8405",
1911 => x"0c5d5b53",
1912 => x"d8397a75",
1913 => x"065c7bfc",
1914 => x"9f388419",
1915 => x"75105659",
1916 => x"f139ff17",
1917 => x"810559f7",
1918 => x"ab398c15",
1919 => x"08881608",
1920 => x"718c120c",
1921 => x"88120c59",
1922 => x"75158411",
1923 => x"08810784",
1924 => x"120c587c",
1925 => x"5182de3f",
1926 => x"881554fb",
1927 => x"a3397716",
1928 => x"78810784",
1929 => x"180c8c17",
1930 => x"08881808",
1931 => x"718c120c",
1932 => x"88120c5c",
1933 => x"7080e388",
1934 => x"0c7080e3",
1935 => x"840c80e2",
1936 => x"fc0b8c12",
1937 => x"0c8c1108",
1938 => x"88120c77",
1939 => x"81078412",
1940 => x"0c770577",
1941 => x"710c557c",
1942 => x"51829a3f",
1943 => x"881654f5",
1944 => x"ba397216",
1945 => x"84110881",
1946 => x"0784120c",
1947 => x"588c1608",
1948 => x"88170871",
1949 => x"8c120c88",
1950 => x"120c577c",
1951 => x"5181f63f",
1952 => x"881654f5",
1953 => x"96397284",
1954 => x"150cf41a",
1955 => x"f8067084",
1956 => x"1d088106",
1957 => x"07841d0c",
1958 => x"701c5556",
1959 => x"850b8415",
1960 => x"0c850b88",
1961 => x"150c8f76",
1962 => x"27fdab38",
1963 => x"881b527c",
1964 => x"5184be3f",
1965 => x"80e2f40b",
1966 => x"88050880",
1967 => x"e2b8085a",
1968 => x"55fd9339",
1969 => x"7880e2b8",
1970 => x"0c7380e2",
1971 => x"e80cfbef",
1972 => x"39728415",
1973 => x"0cfcff39",
1974 => x"fb3d0d77",
1975 => x"707a7c58",
1976 => x"5553568f",
1977 => x"752780e6",
1978 => x"38727607",
1979 => x"83065170",
1980 => x"80dc3875",
1981 => x"73525470",
1982 => x"70840552",
1983 => x"08747084",
1984 => x"05560c73",
1985 => x"71708405",
1986 => x"53087170",
1987 => x"8405530c",
1988 => x"71708405",
1989 => x"53087170",
1990 => x"8405530c",
1991 => x"71708405",
1992 => x"53087170",
1993 => x"8405530c",
1994 => x"f0165654",
1995 => x"748f26c7",
1996 => x"38837527",
1997 => x"95387070",
1998 => x"84055208",
1999 => x"74708405",
2000 => x"560cfc15",
2001 => x"55748326",
2002 => x"ed387371",
2003 => x"5452ff15",
2004 => x"5170ff2e",
2005 => x"98387270",
2006 => x"81055433",
2007 => x"72708105",
2008 => x"5434ff11",
2009 => x"5170ff2e",
2010 => x"098106ea",
2011 => x"3875800c",
2012 => x"873d0d04",
2013 => x"0404fd3d",
2014 => x"0d800b81",
2015 => x"c2d40c76",
2016 => x"5187ca3f",
2017 => x"80085380",
2018 => x"08ff2e88",
2019 => x"3872800c",
2020 => x"853d0d04",
2021 => x"81c2d408",
2022 => x"5473802e",
2023 => x"f0387574",
2024 => x"710c5272",
2025 => x"800c853d",
2026 => x"0d04fb3d",
2027 => x"0d777970",
2028 => x"72078306",
2029 => x"53545270",
2030 => x"93387173",
2031 => x"73085456",
2032 => x"54717308",
2033 => x"2e80c438",
2034 => x"73755452",
2035 => x"71337081",
2036 => x"ff065254",
2037 => x"70802e9d",
2038 => x"38723355",
2039 => x"70752e09",
2040 => x"81069538",
2041 => x"81128114",
2042 => x"71337081",
2043 => x"ff065456",
2044 => x"545270e5",
2045 => x"38723355",
2046 => x"7381ff06",
2047 => x"7581ff06",
2048 => x"71713180",
2049 => x"0c555287",
2050 => x"3d0d0471",
2051 => x"09f7fbfd",
2052 => x"ff1306f8",
2053 => x"84828180",
2054 => x"06527197",
2055 => x"38841484",
2056 => x"16710854",
2057 => x"56547175",
2058 => x"082ee038",
2059 => x"73755452",
2060 => x"ff9a3980",
2061 => x"0b800c87",
2062 => x"3d0d04fb",
2063 => x"3d0d7770",
2064 => x"5256feb0",
2065 => x"3f80e2f4",
2066 => x"0b880508",
2067 => x"841108fc",
2068 => x"06707b31",
2069 => x"9fef05e0",
2070 => x"8006e080",
2071 => x"05525555",
2072 => x"a0807524",
2073 => x"94388052",
2074 => x"7551fe8a",
2075 => x"3f80e2fc",
2076 => x"08145372",
2077 => x"80082e8f",
2078 => x"387551fd",
2079 => x"f83f8053",
2080 => x"72800c87",
2081 => x"3d0d0474",
2082 => x"30527551",
2083 => x"fde83f80",
2084 => x"08ff2ea8",
2085 => x"3880e2f4",
2086 => x"0b880508",
2087 => x"74763181",
2088 => x"0784120c",
2089 => x"5380e2b8",
2090 => x"08753180",
2091 => x"e2b80c75",
2092 => x"51fdc23f",
2093 => x"810b800c",
2094 => x"873d0d04",
2095 => x"80527551",
2096 => x"fdb43f80",
2097 => x"e2f40b88",
2098 => x"05088008",
2099 => x"71315454",
2100 => x"8f7325ff",
2101 => x"a4388008",
2102 => x"80e2e808",
2103 => x"3180e2b8",
2104 => x"0c728107",
2105 => x"84150c75",
2106 => x"51fd8a3f",
2107 => x"8053ff90",
2108 => x"39f73d0d",
2109 => x"7b7d545a",
2110 => x"72802e82",
2111 => x"83387951",
2112 => x"fcf23ff8",
2113 => x"13841108",
2114 => x"70fe0670",
2115 => x"13841108",
2116 => x"fc065c57",
2117 => x"58545780",
2118 => x"e2fc0874",
2119 => x"2e82de38",
2120 => x"7784150c",
2121 => x"80738106",
2122 => x"56597479",
2123 => x"2e81d538",
2124 => x"77148411",
2125 => x"08810656",
2126 => x"5374a038",
2127 => x"77165678",
2128 => x"81e63888",
2129 => x"14085574",
2130 => x"80e2fc2e",
2131 => x"82f9388c",
2132 => x"1408708c",
2133 => x"170c7588",
2134 => x"120c5875",
2135 => x"81078418",
2136 => x"0c751776",
2137 => x"710c5478",
2138 => x"81913883",
2139 => x"ff762781",
2140 => x"c8387589",
2141 => x"2a76832a",
2142 => x"54547380",
2143 => x"2ebf3875",
2144 => x"862ab805",
2145 => x"53847427",
2146 => x"b43880db",
2147 => x"14539474",
2148 => x"27ab3875",
2149 => x"8c2a80ee",
2150 => x"055380d4",
2151 => x"74279e38",
2152 => x"758f2a80",
2153 => x"f7055382",
2154 => x"d4742791",
2155 => x"3875922a",
2156 => x"80fc0553",
2157 => x"8ad47427",
2158 => x"843880fe",
2159 => x"53721010",
2160 => x"1080e2f4",
2161 => x"05881108",
2162 => x"55557375",
2163 => x"2e82bf38",
2164 => x"841408fc",
2165 => x"06597579",
2166 => x"278d3888",
2167 => x"14085473",
2168 => x"752e0981",
2169 => x"06ea388c",
2170 => x"1408708c",
2171 => x"190c7488",
2172 => x"190c7788",
2173 => x"120c5576",
2174 => x"8c150c79",
2175 => x"51faf63f",
2176 => x"8b3d0d04",
2177 => x"76087771",
2178 => x"31587605",
2179 => x"88180856",
2180 => x"567480e2",
2181 => x"fc2e80e0",
2182 => x"388c1708",
2183 => x"708c170c",
2184 => x"7588120c",
2185 => x"53fe8939",
2186 => x"8814088c",
2187 => x"1508708c",
2188 => x"130c5988",
2189 => x"190cfea3",
2190 => x"3975832a",
2191 => x"70545480",
2192 => x"74248198",
2193 => x"3872822c",
2194 => x"81712b80",
2195 => x"e2f80807",
2196 => x"80e2f40b",
2197 => x"84050c74",
2198 => x"10101080",
2199 => x"e2f40588",
2200 => x"1108718c",
2201 => x"1b0c7088",
2202 => x"1b0c7988",
2203 => x"130c565a",
2204 => x"55768c15",
2205 => x"0cff8439",
2206 => x"8159fdb4",
2207 => x"39771673",
2208 => x"81065455",
2209 => x"72983876",
2210 => x"08777131",
2211 => x"5875058c",
2212 => x"18088819",
2213 => x"08718c12",
2214 => x"0c88120c",
2215 => x"55557481",
2216 => x"0784180c",
2217 => x"7680e2f4",
2218 => x"0b88050c",
2219 => x"80e2f008",
2220 => x"7526fec7",
2221 => x"3880e2ec",
2222 => x"08527951",
2223 => x"fafd3f79",
2224 => x"51f9b23f",
2225 => x"feba3981",
2226 => x"778c170c",
2227 => x"7788170c",
2228 => x"758c190c",
2229 => x"7588190c",
2230 => x"59fd8039",
2231 => x"83147082",
2232 => x"2c81712b",
2233 => x"80e2f808",
2234 => x"0780e2f4",
2235 => x"0b84050c",
2236 => x"75101010",
2237 => x"80e2f405",
2238 => x"88110871",
2239 => x"8c1c0c70",
2240 => x"881c0c7a",
2241 => x"88130c57",
2242 => x"5b5653fe",
2243 => x"e4398073",
2244 => x"24a33872",
2245 => x"822c8171",
2246 => x"2b80e2f8",
2247 => x"080780e2",
2248 => x"f40b8405",
2249 => x"0c58748c",
2250 => x"180c7388",
2251 => x"180c7688",
2252 => x"160cfdc3",
2253 => x"39831370",
2254 => x"822c8171",
2255 => x"2b80e2f8",
2256 => x"080780e2",
2257 => x"f40b8405",
2258 => x"0c5953da",
2259 => x"39fe3d0d",
2260 => x"81c2d808",
2261 => x"51708a38",
2262 => x"81c2e070",
2263 => x"81c2d80c",
2264 => x"51741152",
2265 => x"ff537187",
2266 => x"fb808026",
2267 => x"88387181",
2268 => x"c2d80c70",
2269 => x"5372800c",
2270 => x"843d0d04",
2271 => x"fd3d0d80",
2272 => x"0b80e2a4",
2273 => x"08545472",
2274 => x"812e9b38",
2275 => x"7381c2dc",
2276 => x"0cc28e3f",
2277 => x"c0ea3f80",
2278 => x"f1fc5281",
2279 => x"51caf83f",
2280 => x"80085189",
2281 => x"a73f7281",
2282 => x"c2dc0cc1",
2283 => x"f43fc0d0",
2284 => x"3f80f1fc",
2285 => x"528151ca",
2286 => x"de3f8008",
2287 => x"51898d3f",
2288 => x"00ff3900",
2289 => x"ff39f53d",
2290 => x"0d7e6081",
2291 => x"c2dc0870",
2292 => x"5b585b5b",
2293 => x"7580c238",
2294 => x"777a25a1",
2295 => x"38771b70",
2296 => x"337081ff",
2297 => x"06585859",
2298 => x"758a2e98",
2299 => x"387681ff",
2300 => x"0651c18c",
2301 => x"3f811858",
2302 => x"797824e1",
2303 => x"3879800c",
2304 => x"8d3d0d04",
2305 => x"8d51c0f8",
2306 => x"3f783370",
2307 => x"81ff0652",
2308 => x"57c0ed3f",
2309 => x"811858e0",
2310 => x"3979557a",
2311 => x"547d5385",
2312 => x"528d3dfc",
2313 => x"0551c09a",
2314 => x"3f800856",
2315 => x"88973f7b",
2316 => x"80080c75",
2317 => x"800c8d3d",
2318 => x"0d04f63d",
2319 => x"0d7d7f81",
2320 => x"c2dc0870",
2321 => x"5a585a5a",
2322 => x"7580c338",
2323 => x"767925b1",
2324 => x"38761a58",
2325 => x"c08a3f80",
2326 => x"08783480",
2327 => x"0b800881",
2328 => x"ff065758",
2329 => x"758a2ea2",
2330 => x"38758d32",
2331 => x"70307080",
2332 => x"257a0751",
2333 => x"515675b8",
2334 => x"38811757",
2335 => x"787724d1",
2336 => x"38765675",
2337 => x"800c8c3d",
2338 => x"0d048158",
2339 => x"dc397855",
2340 => x"79547c53",
2341 => x"84528c3d",
2342 => x"fc0551ff",
2343 => x"bfa43f80",
2344 => x"085687a1",
2345 => x"3f7a8008",
2346 => x"0c75800c",
2347 => x"8c3d0d04",
2348 => x"811756cf",
2349 => x"39f93d0d",
2350 => x"795781c2",
2351 => x"dc08802e",
2352 => x"ad387651",
2353 => x"89b43f7b",
2354 => x"567a5580",
2355 => x"08810554",
2356 => x"76538252",
2357 => x"893dfc05",
2358 => x"51ffbee6",
2359 => x"3f800857",
2360 => x"86e33f77",
2361 => x"80080c76",
2362 => x"800c893d",
2363 => x"0d0486d5",
2364 => x"3f850b80",
2365 => x"080cff0b",
2366 => x"800c893d",
2367 => x"0d04fb3d",
2368 => x"0d81c2dc",
2369 => x"08705654",
2370 => x"73883874",
2371 => x"800c873d",
2372 => x"0d047753",
2373 => x"8352873d",
2374 => x"fc0551ff",
2375 => x"bea43f80",
2376 => x"085486a1",
2377 => x"3f758008",
2378 => x"0c73800c",
2379 => x"873d0d04",
2380 => x"ff0b800c",
2381 => x"04fb3d0d",
2382 => x"775581c2",
2383 => x"dc08802e",
2384 => x"a9387451",
2385 => x"88b43f80",
2386 => x"08810554",
2387 => x"74538752",
2388 => x"873dfc05",
2389 => x"51ffbdea",
2390 => x"3f800855",
2391 => x"85e73f75",
2392 => x"80080c74",
2393 => x"800c873d",
2394 => x"0d0485d9",
2395 => x"3f850b80",
2396 => x"080cff0b",
2397 => x"800c873d",
2398 => x"0d04fa3d",
2399 => x"0d81c2dc",
2400 => x"08802ea3",
2401 => x"387a5579",
2402 => x"54785386",
2403 => x"52883dfc",
2404 => x"0551ffbd",
2405 => x"ad3f8008",
2406 => x"5685aa3f",
2407 => x"7680080c",
2408 => x"75800c88",
2409 => x"3d0d0485",
2410 => x"9c3f9d0b",
2411 => x"80080cff",
2412 => x"0b800c88",
2413 => x"3d0d04f7",
2414 => x"3d0d7b7d",
2415 => x"5b59bc53",
2416 => x"80527951",
2417 => x"86aa3f80",
2418 => x"70565798",
2419 => x"56741970",
2420 => x"3370782b",
2421 => x"79078118",
2422 => x"f81a5a58",
2423 => x"59555884",
2424 => x"7524ea38",
2425 => x"767a2384",
2426 => x"19588070",
2427 => x"56579856",
2428 => x"74187033",
2429 => x"70782b79",
2430 => x"078118f8",
2431 => x"1a5a5859",
2432 => x"51548475",
2433 => x"24ea3876",
2434 => x"821b2388",
2435 => x"19588070",
2436 => x"56579856",
2437 => x"74187033",
2438 => x"70782b79",
2439 => x"078118f8",
2440 => x"1a5a5859",
2441 => x"51548475",
2442 => x"24ea3876",
2443 => x"841b0c8c",
2444 => x"19588070",
2445 => x"56579856",
2446 => x"74187033",
2447 => x"70782b79",
2448 => x"078118f8",
2449 => x"1a5a5859",
2450 => x"51548475",
2451 => x"24ea3876",
2452 => x"881b2390",
2453 => x"19588070",
2454 => x"56579856",
2455 => x"74187033",
2456 => x"70782b79",
2457 => x"078118f8",
2458 => x"1a5a5859",
2459 => x"51548475",
2460 => x"24ea3876",
2461 => x"8a1b2394",
2462 => x"19588070",
2463 => x"56579856",
2464 => x"74187033",
2465 => x"70782b79",
2466 => x"078118f8",
2467 => x"1a5a5859",
2468 => x"51548475",
2469 => x"24ea3876",
2470 => x"8c1b2398",
2471 => x"19588070",
2472 => x"56579856",
2473 => x"74187033",
2474 => x"70782b79",
2475 => x"078118f8",
2476 => x"1a5a5859",
2477 => x"51548475",
2478 => x"24ea3876",
2479 => x"8e1b239c",
2480 => x"19588070",
2481 => x"5657b856",
2482 => x"74187033",
2483 => x"70782b79",
2484 => x"078118f8",
2485 => x"1a5a5859",
2486 => x"5a548875",
2487 => x"24ea3876",
2488 => x"901b0c8b",
2489 => x"3d0d04e9",
2490 => x"3d0d6a81",
2491 => x"c2dc0857",
2492 => x"57759338",
2493 => x"80c0800b",
2494 => x"84180c75",
2495 => x"ac180c75",
2496 => x"800c993d",
2497 => x"0d04893d",
2498 => x"70556a54",
2499 => x"558a5299",
2500 => x"3dffbc05",
2501 => x"51ffbaaa",
2502 => x"3f800877",
2503 => x"53755256",
2504 => x"fd953f82",
2505 => x"a03f7780",
2506 => x"080c7580",
2507 => x"0c993d0d",
2508 => x"04e93d0d",
2509 => x"695781c2",
2510 => x"dc08802e",
2511 => x"b6387651",
2512 => x"84b83f89",
2513 => x"3d705680",
2514 => x"08810555",
2515 => x"7754568f",
2516 => x"52993dff",
2517 => x"bc0551ff",
2518 => x"b9e83f80",
2519 => x"086b5376",
2520 => x"5257fcd3",
2521 => x"3f81de3f",
2522 => x"7780080c",
2523 => x"76800c99",
2524 => x"3d0d0481",
2525 => x"d03f850b",
2526 => x"80080cff",
2527 => x"0b800c99",
2528 => x"3d0d04fc",
2529 => x"3d0d8154",
2530 => x"81c2dc08",
2531 => x"88387380",
2532 => x"0c863d0d",
2533 => x"04765397",
2534 => x"b952863d",
2535 => x"fc0551ff",
2536 => x"b9a03f80",
2537 => x"0854819d",
2538 => x"3f748008",
2539 => x"0c73800c",
2540 => x"863d0d04",
2541 => x"f43d0d7e",
2542 => x"80f2a808",
2543 => x"700881ff",
2544 => x"06913df8",
2545 => x"05545159",
2546 => x"59ffbac5",
2547 => x"3f775780",
2548 => x"5476557b",
2549 => x"7d585276",
2550 => x"538e3df0",
2551 => x"0551d6a0",
2552 => x"3f797b58",
2553 => x"790c7684",
2554 => x"1a0c7880",
2555 => x"0c8e3d0d",
2556 => x"04f43d0d",
2557 => x"7e80f2a8",
2558 => x"08700870",
2559 => x"81ff0692",
2560 => x"3df80555",
2561 => x"515a5759",
2562 => x"ffba863f",
2563 => x"7757800b",
2564 => x"8b3d5954",
2565 => x"76557b7d",
2566 => x"58527653",
2567 => x"7751d5e0",
2568 => x"3f8056bd",
2569 => x"84c07655",
2570 => x"55797b58",
2571 => x"52765377",
2572 => x"51d5cd3f",
2573 => x"7a577880",
2574 => x"2e843876",
2575 => x"790c7680",
2576 => x"0c8e3d0d",
2577 => x"0480eafc",
2578 => x"08800c04",
2579 => x"f73d0d7b",
2580 => x"80eafc08",
2581 => x"82c81108",
2582 => x"5a545a77",
2583 => x"802e80da",
2584 => x"38818818",
2585 => x"841908ff",
2586 => x"0581712b",
2587 => x"59555980",
2588 => x"742480ea",
2589 => x"38807424",
2590 => x"b5387382",
2591 => x"2b781188",
2592 => x"05565681",
2593 => x"80190877",
2594 => x"06537280",
2595 => x"2eb63878",
2596 => x"16700853",
2597 => x"53795174",
2598 => x"0853722d",
2599 => x"ff14fc17",
2600 => x"fc177981",
2601 => x"2c5a5757",
2602 => x"54738025",
2603 => x"d6387708",
2604 => x"5877ffad",
2605 => x"3880eafc",
2606 => x"0853bc13",
2607 => x"08a53879",
2608 => x"51f5fd3f",
2609 => x"74085372",
2610 => x"2dff14fc",
2611 => x"17fc1779",
2612 => x"812c5a57",
2613 => x"57547380",
2614 => x"25ffa838",
2615 => x"d1398057",
2616 => x"ff933972",
2617 => x"51bc1308",
2618 => x"54732d79",
2619 => x"51f5d13f",
2620 => x"fb3d0d77",
2621 => x"7a71028c",
2622 => x"05a30533",
2623 => x"58545456",
2624 => x"83732780",
2625 => x"d4387583",
2626 => x"06517080",
2627 => x"cc387488",
2628 => x"2b750770",
2629 => x"71902b07",
2630 => x"55518f73",
2631 => x"27a73873",
2632 => x"72708405",
2633 => x"540c7174",
2634 => x"71708405",
2635 => x"530c7471",
2636 => x"70840553",
2637 => x"0c747170",
2638 => x"8405530c",
2639 => x"f0145452",
2640 => x"728f26db",
2641 => x"38837327",
2642 => x"90387372",
2643 => x"70840554",
2644 => x"0cfc1353",
2645 => x"728326f2",
2646 => x"38ff1351",
2647 => x"70ff2e93",
2648 => x"38747270",
2649 => x"81055434",
2650 => x"ff115170",
2651 => x"ff2e0981",
2652 => x"06ef3875",
2653 => x"800c873d",
2654 => x"0d04fd3d",
2655 => x"0d757071",
2656 => x"83065355",
2657 => x"5270b438",
2658 => x"71700870",
2659 => x"09f7fbfd",
2660 => x"ff1206f8",
2661 => x"84828180",
2662 => x"06545253",
2663 => x"719b3884",
2664 => x"13700870",
2665 => x"09f7fbfd",
2666 => x"ff1206f8",
2667 => x"84828180",
2668 => x"06545253",
2669 => x"71802ee7",
2670 => x"38725271",
2671 => x"33537280",
2672 => x"2e8a3881",
2673 => x"12703354",
2674 => x"5272f838",
2675 => x"71743180",
2676 => x"0c853d0d",
2677 => x"04ff3d0d",
2678 => x"80f2840b",
2679 => x"fc057008",
2680 => x"525270ff",
2681 => x"2e913870",
2682 => x"2dfc1270",
2683 => x"08525270",
2684 => x"ff2e0981",
2685 => x"06f13883",
2686 => x"3d0d0404",
2687 => x"ffb7a63f",
2688 => x"04000000",
2689 => x"30313233",
2690 => x"34353637",
2691 => x"38390000",
2692 => x"44485259",
2693 => x"53544f4e",
2694 => x"45205052",
2695 => x"4f475241",
2696 => x"4d2c2053",
2697 => x"4f4d4520",
2698 => x"53545249",
2699 => x"4e470000",
2700 => x"44485259",
2701 => x"53544f4e",
2702 => x"45205052",
2703 => x"4f475241",
2704 => x"4d2c2031",
2705 => x"27535420",
2706 => x"53545249",
2707 => x"4e470000",
2708 => x"44687279",
2709 => x"73746f6e",
2710 => x"65204265",
2711 => x"6e63686d",
2712 => x"61726b2c",
2713 => x"20566572",
2714 => x"73696f6e",
2715 => x"20322e31",
2716 => x"20284c61",
2717 => x"6e677561",
2718 => x"67653a20",
2719 => x"43290a00",
2720 => x"50726f67",
2721 => x"72616d20",
2722 => x"636f6d70",
2723 => x"696c6564",
2724 => x"20776974",
2725 => x"68202772",
2726 => x"65676973",
2727 => x"74657227",
2728 => x"20617474",
2729 => x"72696275",
2730 => x"74650a00",
2731 => x"45786563",
2732 => x"7574696f",
2733 => x"6e207374",
2734 => x"61727473",
2735 => x"2c202564",
2736 => x"2072756e",
2737 => x"73207468",
2738 => x"726f7567",
2739 => x"68204468",
2740 => x"72797374",
2741 => x"6f6e650a",
2742 => x"00000000",
2743 => x"44485259",
2744 => x"53544f4e",
2745 => x"45205052",
2746 => x"4f475241",
2747 => x"4d2c2032",
2748 => x"274e4420",
2749 => x"53545249",
2750 => x"4e470000",
2751 => x"45786563",
2752 => x"7574696f",
2753 => x"6e20656e",
2754 => x"64730a00",
2755 => x"46696e61",
2756 => x"6c207661",
2757 => x"6c756573",
2758 => x"206f6620",
2759 => x"74686520",
2760 => x"76617269",
2761 => x"61626c65",
2762 => x"73207573",
2763 => x"65642069",
2764 => x"6e207468",
2765 => x"65206265",
2766 => x"6e63686d",
2767 => x"61726b3a",
2768 => x"0a000000",
2769 => x"496e745f",
2770 => x"476c6f62",
2771 => x"3a202020",
2772 => x"20202020",
2773 => x"20202020",
2774 => x"2025640a",
2775 => x"00000000",
2776 => x"20202020",
2777 => x"20202020",
2778 => x"73686f75",
2779 => x"6c642062",
2780 => x"653a2020",
2781 => x"2025640a",
2782 => x"00000000",
2783 => x"426f6f6c",
2784 => x"5f476c6f",
2785 => x"623a2020",
2786 => x"20202020",
2787 => x"20202020",
2788 => x"2025640a",
2789 => x"00000000",
2790 => x"43685f31",
2791 => x"5f476c6f",
2792 => x"623a2020",
2793 => x"20202020",
2794 => x"20202020",
2795 => x"2025630a",
2796 => x"00000000",
2797 => x"20202020",
2798 => x"20202020",
2799 => x"73686f75",
2800 => x"6c642062",
2801 => x"653a2020",
2802 => x"2025630a",
2803 => x"00000000",
2804 => x"43685f32",
2805 => x"5f476c6f",
2806 => x"623a2020",
2807 => x"20202020",
2808 => x"20202020",
2809 => x"2025630a",
2810 => x"00000000",
2811 => x"4172725f",
2812 => x"315f476c",
2813 => x"6f625b38",
2814 => x"5d3a2020",
2815 => x"20202020",
2816 => x"2025640a",
2817 => x"00000000",
2818 => x"4172725f",
2819 => x"325f476c",
2820 => x"6f625b38",
2821 => x"5d5b375d",
2822 => x"3a202020",
2823 => x"2025640a",
2824 => x"00000000",
2825 => x"20202020",
2826 => x"20202020",
2827 => x"73686f75",
2828 => x"6c642062",
2829 => x"653a2020",
2830 => x"204e756d",
2831 => x"6265725f",
2832 => x"4f665f52",
2833 => x"756e7320",
2834 => x"2b203130",
2835 => x"0a000000",
2836 => x"5074725f",
2837 => x"476c6f62",
2838 => x"2d3e0a00",
2839 => x"20205074",
2840 => x"725f436f",
2841 => x"6d703a20",
2842 => x"20202020",
2843 => x"20202020",
2844 => x"2025640a",
2845 => x"00000000",
2846 => x"20202020",
2847 => x"20202020",
2848 => x"73686f75",
2849 => x"6c642062",
2850 => x"653a2020",
2851 => x"2028696d",
2852 => x"706c656d",
2853 => x"656e7461",
2854 => x"74696f6e",
2855 => x"2d646570",
2856 => x"656e6465",
2857 => x"6e74290a",
2858 => x"00000000",
2859 => x"20204469",
2860 => x"7363723a",
2861 => x"20202020",
2862 => x"20202020",
2863 => x"20202020",
2864 => x"2025640a",
2865 => x"00000000",
2866 => x"2020456e",
2867 => x"756d5f43",
2868 => x"6f6d703a",
2869 => x"20202020",
2870 => x"20202020",
2871 => x"2025640a",
2872 => x"00000000",
2873 => x"2020496e",
2874 => x"745f436f",
2875 => x"6d703a20",
2876 => x"20202020",
2877 => x"20202020",
2878 => x"2025640a",
2879 => x"00000000",
2880 => x"20205374",
2881 => x"725f436f",
2882 => x"6d703a20",
2883 => x"20202020",
2884 => x"20202020",
2885 => x"2025730a",
2886 => x"00000000",
2887 => x"20202020",
2888 => x"20202020",
2889 => x"73686f75",
2890 => x"6c642062",
2891 => x"653a2020",
2892 => x"20444852",
2893 => x"5953544f",
2894 => x"4e452050",
2895 => x"524f4752",
2896 => x"414d2c20",
2897 => x"534f4d45",
2898 => x"20535452",
2899 => x"494e470a",
2900 => x"00000000",
2901 => x"4e657874",
2902 => x"5f507472",
2903 => x"5f476c6f",
2904 => x"622d3e0a",
2905 => x"00000000",
2906 => x"20202020",
2907 => x"20202020",
2908 => x"73686f75",
2909 => x"6c642062",
2910 => x"653a2020",
2911 => x"2028696d",
2912 => x"706c656d",
2913 => x"656e7461",
2914 => x"74696f6e",
2915 => x"2d646570",
2916 => x"656e6465",
2917 => x"6e74292c",
2918 => x"2073616d",
2919 => x"65206173",
2920 => x"2061626f",
2921 => x"76650a00",
2922 => x"496e745f",
2923 => x"315f4c6f",
2924 => x"633a2020",
2925 => x"20202020",
2926 => x"20202020",
2927 => x"2025640a",
2928 => x"00000000",
2929 => x"496e745f",
2930 => x"325f4c6f",
2931 => x"633a2020",
2932 => x"20202020",
2933 => x"20202020",
2934 => x"2025640a",
2935 => x"00000000",
2936 => x"496e745f",
2937 => x"335f4c6f",
2938 => x"633a2020",
2939 => x"20202020",
2940 => x"20202020",
2941 => x"2025640a",
2942 => x"00000000",
2943 => x"456e756d",
2944 => x"5f4c6f63",
2945 => x"3a202020",
2946 => x"20202020",
2947 => x"20202020",
2948 => x"2025640a",
2949 => x"00000000",
2950 => x"5374725f",
2951 => x"315f4c6f",
2952 => x"633a2020",
2953 => x"20202020",
2954 => x"20202020",
2955 => x"2025730a",
2956 => x"00000000",
2957 => x"20202020",
2958 => x"20202020",
2959 => x"73686f75",
2960 => x"6c642062",
2961 => x"653a2020",
2962 => x"20444852",
2963 => x"5953544f",
2964 => x"4e452050",
2965 => x"524f4752",
2966 => x"414d2c20",
2967 => x"31275354",
2968 => x"20535452",
2969 => x"494e470a",
2970 => x"00000000",
2971 => x"5374725f",
2972 => x"325f4c6f",
2973 => x"633a2020",
2974 => x"20202020",
2975 => x"20202020",
2976 => x"2025730a",
2977 => x"00000000",
2978 => x"20202020",
2979 => x"20202020",
2980 => x"73686f75",
2981 => x"6c642062",
2982 => x"653a2020",
2983 => x"20444852",
2984 => x"5953544f",
2985 => x"4e452050",
2986 => x"524f4752",
2987 => x"414d2c20",
2988 => x"32274e44",
2989 => x"20535452",
2990 => x"494e470a",
2991 => x"00000000",
2992 => x"55736572",
2993 => x"2074696d",
2994 => x"653a2025",
2995 => x"640a0000",
2996 => x"4d696372",
2997 => x"6f736563",
2998 => x"6f6e6473",
2999 => x"20666f72",
3000 => x"206f6e65",
3001 => x"2072756e",
3002 => x"20746872",
3003 => x"6f756768",
3004 => x"20446872",
3005 => x"7973746f",
3006 => x"6e653a20",
3007 => x"00000000",
3008 => x"2564200a",
3009 => x"00000000",
3010 => x"44687279",
3011 => x"73746f6e",
3012 => x"65732070",
3013 => x"65722053",
3014 => x"65636f6e",
3015 => x"643a2020",
3016 => x"20202020",
3017 => x"20202020",
3018 => x"20202020",
3019 => x"20202020",
3020 => x"20202020",
3021 => x"00000000",
3022 => x"56415820",
3023 => x"4d495053",
3024 => x"20726174",
3025 => x"696e6720",
3026 => x"2a203130",
3027 => x"3030203d",
3028 => x"20256420",
3029 => x"0a000000",
3030 => x"50726f67",
3031 => x"72616d20",
3032 => x"636f6d70",
3033 => x"696c6564",
3034 => x"20776974",
3035 => x"686f7574",
3036 => x"20277265",
3037 => x"67697374",
3038 => x"65722720",
3039 => x"61747472",
3040 => x"69627574",
3041 => x"650a0000",
3042 => x"4d656173",
3043 => x"75726564",
3044 => x"2074696d",
3045 => x"6520746f",
3046 => x"6f20736d",
3047 => x"616c6c20",
3048 => x"746f206f",
3049 => x"62746169",
3050 => x"6e206d65",
3051 => x"616e696e",
3052 => x"6766756c",
3053 => x"20726573",
3054 => x"756c7473",
3055 => x"0a000000",
3056 => x"506c6561",
3057 => x"73652069",
3058 => x"6e637265",
3059 => x"61736520",
3060 => x"6e756d62",
3061 => x"6572206f",
3062 => x"66207275",
3063 => x"6e730a00",
3064 => x"44485259",
3065 => x"53544f4e",
3066 => x"45205052",
3067 => x"4f475241",
3068 => x"4d2c2033",
3069 => x"27524420",
3070 => x"53545249",
3071 => x"4e470000",
3072 => x"00010202",
3073 => x"03030303",
3074 => x"04040404",
3075 => x"04040404",
3076 => x"05050505",
3077 => x"05050505",
3078 => x"05050505",
3079 => x"05050505",
3080 => x"06060606",
3081 => x"06060606",
3082 => x"06060606",
3083 => x"06060606",
3084 => x"06060606",
3085 => x"06060606",
3086 => x"06060606",
3087 => x"06060606",
3088 => x"07070707",
3089 => x"07070707",
3090 => x"07070707",
3091 => x"07070707",
3092 => x"07070707",
3093 => x"07070707",
3094 => x"07070707",
3095 => x"07070707",
3096 => x"07070707",
3097 => x"07070707",
3098 => x"07070707",
3099 => x"07070707",
3100 => x"07070707",
3101 => x"07070707",
3102 => x"07070707",
3103 => x"07070707",
3104 => x"08080808",
3105 => x"08080808",
3106 => x"08080808",
3107 => x"08080808",
3108 => x"08080808",
3109 => x"08080808",
3110 => x"08080808",
3111 => x"08080808",
3112 => x"08080808",
3113 => x"08080808",
3114 => x"08080808",
3115 => x"08080808",
3116 => x"08080808",
3117 => x"08080808",
3118 => x"08080808",
3119 => x"08080808",
3120 => x"08080808",
3121 => x"08080808",
3122 => x"08080808",
3123 => x"08080808",
3124 => x"08080808",
3125 => x"08080808",
3126 => x"08080808",
3127 => x"08080808",
3128 => x"08080808",
3129 => x"08080808",
3130 => x"08080808",
3131 => x"08080808",
3132 => x"08080808",
3133 => x"08080808",
3134 => x"08080808",
3135 => x"08080808",
3136 => x"43000000",
3137 => x"64756d6d",
3138 => x"792e6578",
3139 => x"65000000",
3140 => x"00ffffff",
3141 => x"ff00ffff",
3142 => x"ffff00ff",
3143 => x"ffffff00",
3144 => x"00000000",
3145 => x"00000000",
3146 => x"00000000",
3147 => x"0000390c",
3148 => x"000004d2", -- iterations 0x4d2=1234 
3149 => x"00000000",
3150 => x"00000000",
3151 => x"00000000",
3152 => x"00000000",
3153 => x"00000000",
3154 => x"00000000",
3155 => x"00000000",
3156 => x"00000000",
3157 => x"00000000",
3158 => x"00000000",
3159 => x"00000000",
3160 => x"00000000",
3161 => x"00000000",
3162 => x"ffffffff",
3163 => x"00000000",
3164 => x"00020000",
3165 => x"00000000",
3166 => x"00000000",
3167 => x"00003174",
3168 => x"00003174",
3169 => x"0000317c",
3170 => x"0000317c",
3171 => x"00003184",
3172 => x"00003184",
3173 => x"0000318c",
3174 => x"0000318c",
3175 => x"00003194",
3176 => x"00003194",
3177 => x"0000319c",
3178 => x"0000319c",
3179 => x"000031a4",
3180 => x"000031a4",
3181 => x"000031ac",
3182 => x"000031ac",
3183 => x"000031b4",
3184 => x"000031b4",
3185 => x"000031bc",
3186 => x"000031bc",
3187 => x"000031c4",
3188 => x"000031c4",
3189 => x"000031cc",
3190 => x"000031cc",
3191 => x"000031d4",
3192 => x"000031d4",
3193 => x"000031dc",
3194 => x"000031dc",
3195 => x"000031e4",
3196 => x"000031e4",
3197 => x"000031ec",
3198 => x"000031ec",
3199 => x"000031f4",
3200 => x"000031f4",
3201 => x"000031fc",
3202 => x"000031fc",
3203 => x"00003204",
3204 => x"00003204",
3205 => x"0000320c",
3206 => x"0000320c",
3207 => x"00003214",
3208 => x"00003214",
3209 => x"0000321c",
3210 => x"0000321c",
3211 => x"00003224",
3212 => x"00003224",
3213 => x"0000322c",
3214 => x"0000322c",
3215 => x"00003234",
3216 => x"00003234",
3217 => x"0000323c",
3218 => x"0000323c",
3219 => x"00003244",
3220 => x"00003244",
3221 => x"0000324c",
3222 => x"0000324c",
3223 => x"00003254",
3224 => x"00003254",
3225 => x"0000325c",
3226 => x"0000325c",
3227 => x"00003264",
3228 => x"00003264",
3229 => x"0000326c",
3230 => x"0000326c",
3231 => x"00003274",
3232 => x"00003274",
3233 => x"0000327c",
3234 => x"0000327c",
3235 => x"00003284",
3236 => x"00003284",
3237 => x"0000328c",
3238 => x"0000328c",
3239 => x"00003294",
3240 => x"00003294",
3241 => x"0000329c",
3242 => x"0000329c",
3243 => x"000032a4",
3244 => x"000032a4",
3245 => x"000032ac",
3246 => x"000032ac",
3247 => x"000032b4",
3248 => x"000032b4",
3249 => x"000032bc",
3250 => x"000032bc",
3251 => x"000032c4",
3252 => x"000032c4",
3253 => x"000032cc",
3254 => x"000032cc",
3255 => x"000032d4",
3256 => x"000032d4",
3257 => x"000032dc",
3258 => x"000032dc",
3259 => x"000032e4",
3260 => x"000032e4",
3261 => x"000032ec",
3262 => x"000032ec",
3263 => x"000032f4",
3264 => x"000032f4",
3265 => x"000032fc",
3266 => x"000032fc",
3267 => x"00003304",
3268 => x"00003304",
3269 => x"0000330c",
3270 => x"0000330c",
3271 => x"00003314",
3272 => x"00003314",
3273 => x"0000331c",
3274 => x"0000331c",
3275 => x"00003324",
3276 => x"00003324",
3277 => x"0000332c",
3278 => x"0000332c",
3279 => x"00003334",
3280 => x"00003334",
3281 => x"0000333c",
3282 => x"0000333c",
3283 => x"00003344",
3284 => x"00003344",
3285 => x"0000334c",
3286 => x"0000334c",
3287 => x"00003354",
3288 => x"00003354",
3289 => x"0000335c",
3290 => x"0000335c",
3291 => x"00003364",
3292 => x"00003364",
3293 => x"0000336c",
3294 => x"0000336c",
3295 => x"00003374",
3296 => x"00003374",
3297 => x"0000337c",
3298 => x"0000337c",
3299 => x"00003384",
3300 => x"00003384",
3301 => x"0000338c",
3302 => x"0000338c",
3303 => x"00003394",
3304 => x"00003394",
3305 => x"0000339c",
3306 => x"0000339c",
3307 => x"000033a4",
3308 => x"000033a4",
3309 => x"000033ac",
3310 => x"000033ac",
3311 => x"000033b4",
3312 => x"000033b4",
3313 => x"000033bc",
3314 => x"000033bc",
3315 => x"000033c4",
3316 => x"000033c4",
3317 => x"000033cc",
3318 => x"000033cc",
3319 => x"000033d4",
3320 => x"000033d4",
3321 => x"000033dc",
3322 => x"000033dc",
3323 => x"000033e4",
3324 => x"000033e4",
3325 => x"000033ec",
3326 => x"000033ec",
3327 => x"000033f4",
3328 => x"000033f4",
3329 => x"000033fc",
3330 => x"000033fc",
3331 => x"00003404",
3332 => x"00003404",
3333 => x"0000340c",
3334 => x"0000340c",
3335 => x"00003414",
3336 => x"00003414",
3337 => x"0000341c",
3338 => x"0000341c",
3339 => x"00003424",
3340 => x"00003424",
3341 => x"0000342c",
3342 => x"0000342c",
3343 => x"00003434",
3344 => x"00003434",
3345 => x"0000343c",
3346 => x"0000343c",
3347 => x"00003444",
3348 => x"00003444",
3349 => x"0000344c",
3350 => x"0000344c",
3351 => x"00003454",
3352 => x"00003454",
3353 => x"0000345c",
3354 => x"0000345c",
3355 => x"00003464",
3356 => x"00003464",
3357 => x"0000346c",
3358 => x"0000346c",
3359 => x"00003474",
3360 => x"00003474",
3361 => x"0000347c",
3362 => x"0000347c",
3363 => x"00003484",
3364 => x"00003484",
3365 => x"0000348c",
3366 => x"0000348c",
3367 => x"00003494",
3368 => x"00003494",
3369 => x"0000349c",
3370 => x"0000349c",
3371 => x"000034a4",
3372 => x"000034a4",
3373 => x"000034ac",
3374 => x"000034ac",
3375 => x"000034b4",
3376 => x"000034b4",
3377 => x"000034bc",
3378 => x"000034bc",
3379 => x"000034c4",
3380 => x"000034c4",
3381 => x"000034cc",
3382 => x"000034cc",
3383 => x"000034d4",
3384 => x"000034d4",
3385 => x"000034dc",
3386 => x"000034dc",
3387 => x"000034e4",
3388 => x"000034e4",
3389 => x"000034ec",
3390 => x"000034ec",
3391 => x"000034f4",
3392 => x"000034f4",
3393 => x"000034fc",
3394 => x"000034fc",
3395 => x"00003504",
3396 => x"00003504",
3397 => x"0000350c",
3398 => x"0000350c",
3399 => x"00003514",
3400 => x"00003514",
3401 => x"0000351c",
3402 => x"0000351c",
3403 => x"00003524",
3404 => x"00003524",
3405 => x"0000352c",
3406 => x"0000352c",
3407 => x"00003534",
3408 => x"00003534",
3409 => x"0000353c",
3410 => x"0000353c",
3411 => x"00003544",
3412 => x"00003544",
3413 => x"0000354c",
3414 => x"0000354c",
3415 => x"00003554",
3416 => x"00003554",
3417 => x"0000355c",
3418 => x"0000355c",
3419 => x"00003564",
3420 => x"00003564",
3421 => x"0000356c",
3422 => x"0000356c",
3423 => x"00003580",
3424 => x"00000000",
3425 => x"000037e8",
3426 => x"00003844",
3427 => x"000038a0",
3428 => x"00000000",
3429 => x"00000000",
3430 => x"00000000",
3431 => x"00000000",
3432 => x"00000000",
3433 => x"00000000",
3434 => x"00000000",
3435 => x"00000000",
3436 => x"00000000",
3437 => x"00003100",
3438 => x"00000000",
3439 => x"00000000",
3440 => x"00000000",
3441 => x"00000000",
3442 => x"00000000",
3443 => x"00000000",
3444 => x"00000000",
3445 => x"00000000",
3446 => x"00000000",
3447 => x"00000000",
3448 => x"00000000",
3449 => x"00000000",
3450 => x"00000000",
3451 => x"00000000",
3452 => x"00000000",
3453 => x"00000000",
3454 => x"00000000",
3455 => x"00000000",
3456 => x"00000000",
3457 => x"00000000",
3458 => x"00000000",
3459 => x"00000000",
3460 => x"00000000",
3461 => x"00000000",
3462 => x"00000000",
3463 => x"00000000",
3464 => x"00000000",
3465 => x"00000000",
3466 => x"00000001",
3467 => x"330eabcd",
3468 => x"1234e66d",
3469 => x"deec0005",
3470 => x"000b0000",
3471 => x"00000000",
3472 => x"00000000",
3473 => x"00000000",
3474 => x"00000000",
3475 => x"00000000",
3476 => x"00000000",
3477 => x"00000000",
3478 => x"00000000",
3479 => x"00000000",
3480 => x"00000000",
3481 => x"00000000",
3482 => x"00000000",
3483 => x"00000000",
3484 => x"00000000",
3485 => x"00000000",
3486 => x"00000000",
3487 => x"00000000",
3488 => x"00000000",
3489 => x"00000000",
3490 => x"00000000",
3491 => x"00000000",
3492 => x"00000000",
3493 => x"00000000",
3494 => x"00000000",
3495 => x"00000000",
3496 => x"00000000",
3497 => x"00000000",
3498 => x"00000000",
3499 => x"00000000",
3500 => x"00000000",
3501 => x"00000000",
3502 => x"00000000",
3503 => x"00000000",
3504 => x"00000000",
3505 => x"00000000",
3506 => x"00000000",
3507 => x"00000000",
3508 => x"00000000",
3509 => x"00000000",
3510 => x"00000000",
3511 => x"00000000",
3512 => x"00000000",
3513 => x"00000000",
3514 => x"00000000",
3515 => x"00000000",
3516 => x"00000000",
3517 => x"00000000",
3518 => x"00000000",
3519 => x"00000000",
3520 => x"00000000",
3521 => x"00000000",
3522 => x"00000000",
3523 => x"00000000",
3524 => x"00000000",
3525 => x"00000000",
3526 => x"00000000",
3527 => x"00000000",
3528 => x"00000000",
3529 => x"00000000",
3530 => x"00000000",
3531 => x"00000000",
3532 => x"00000000",
3533 => x"00000000",
3534 => x"00000000",
3535 => x"00000000",
3536 => x"00000000",
3537 => x"00000000",
3538 => x"00000000",
3539 => x"00000000",
3540 => x"00000000",
3541 => x"00000000",
3542 => x"00000000",
3543 => x"00000000",
3544 => x"00000000",
3545 => x"00000000",
3546 => x"00000000",
3547 => x"00000000",
3548 => x"00000000",
3549 => x"00000000",
3550 => x"00000000",
3551 => x"00000000",
3552 => x"00000000",
3553 => x"00000000",
3554 => x"00000000",
3555 => x"00000000",
3556 => x"00000000",
3557 => x"00000000",
3558 => x"00000000",
3559 => x"00000000",
3560 => x"00000000",
3561 => x"00000000",
3562 => x"00000000",
3563 => x"00000000",
3564 => x"00000000",
3565 => x"00000000",
3566 => x"00000000",
3567 => x"00000000",
3568 => x"00000000",
3569 => x"00000000",
3570 => x"00000000",
3571 => x"00000000",
3572 => x"00000000",
3573 => x"00000000",
3574 => x"00000000",
3575 => x"00000000",
3576 => x"00000000",
3577 => x"00000000",
3578 => x"00000000",
3579 => x"00000000",
3580 => x"00000000",
3581 => x"00000000",
3582 => x"00000000",
3583 => x"00000000",
3584 => x"00000000",
3585 => x"00000000",
3586 => x"00000000",
3587 => x"00000000",
3588 => x"00000000",
3589 => x"00000000",
3590 => x"00000000",
3591 => x"00000000",
3592 => x"00000000",
3593 => x"00000000",
3594 => x"00000000",
3595 => x"00000000",
3596 => x"00000000",
3597 => x"00000000",
3598 => x"00000000",
3599 => x"00000000",
3600 => x"00000000",
3601 => x"00000000",
3602 => x"00000000",
3603 => x"00000000",
3604 => x"00000000",
3605 => x"00000000",
3606 => x"00000000",
3607 => x"00000000",
3608 => x"00000000",
3609 => x"00000000",
3610 => x"00000000",
3611 => x"00000000",
3612 => x"00000000",
3613 => x"00000000",
3614 => x"00000000",
3615 => x"00000000",
3616 => x"00000000",
3617 => x"00000000",
3618 => x"00000000",
3619 => x"00000000",
3620 => x"00000000",
3621 => x"00000000",
3622 => x"00000000",
3623 => x"00000000",
3624 => x"00000000",
3625 => x"00000000",
3626 => x"00000000",
3627 => x"00000000",
3628 => x"00000000",
3629 => x"00000000",
3630 => x"00000000",
3631 => x"00000000",
3632 => x"00000000",
3633 => x"00000000",
3634 => x"00000000",
3635 => x"00000000",
3636 => x"00000000",
3637 => x"00000000",
3638 => x"00000000",
3639 => x"00000000",
3640 => x"00000000",
3641 => x"00000000",
3642 => x"00000000",
3643 => x"00000000",
3644 => x"00000000",
3645 => x"00000000",
3646 => x"00000000",
3647 => x"00003104",
3648 => x"ffffffff",
3649 => x"00000000",
3650 => x"ffffffff",
3651 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
