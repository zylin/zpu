-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80c3ac0c",
     3 => x"3a0b0b0b",
     4 => x"bce80400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0bbdad2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80c3",
   162 => x"98738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0bb7",
   171 => x"d32d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bb9",
   179 => x"852d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80c3a80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82803fb6",
   257 => x"cf3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"53510480",
   280 => x"c3a80880",
   281 => x"2ea43880",
   282 => x"c3ac0882",
   283 => x"2ebd3883",
   284 => x"80800b0b",
   285 => x"0b80cae0",
   286 => x"0c82a080",
   287 => x"0b80cae4",
   288 => x"0c829080",
   289 => x"0b80cae8",
   290 => x"0c04f880",
   291 => x"8080a40b",
   292 => x"0b0b80ca",
   293 => x"e00cf880",
   294 => x"8082800b",
   295 => x"80cae40c",
   296 => x"f8808084",
   297 => x"800b80ca",
   298 => x"e80c0480",
   299 => x"c0a8808c",
   300 => x"0b0b0b80",
   301 => x"cae00c80",
   302 => x"c0a88094",
   303 => x"0b80cae4",
   304 => x"0c0b0b0b",
   305 => x"bf800b80",
   306 => x"cae80c04",
   307 => x"ff3d0d80",
   308 => x"caec3351",
   309 => x"70a73880",
   310 => x"c3b40870",
   311 => x"08525270",
   312 => x"802e9438",
   313 => x"841280c3",
   314 => x"b40c702d",
   315 => x"80c3b408",
   316 => x"70085252",
   317 => x"70ee3881",
   318 => x"0b80caec",
   319 => x"34833d0d",
   320 => x"0404803d",
   321 => x"0d0b0b80",
   322 => x"cadc0880",
   323 => x"2e8e380b",
   324 => x"0b0b0b80",
   325 => x"0b802e09",
   326 => x"81068538",
   327 => x"823d0d04",
   328 => x"0b0b80ca",
   329 => x"dc510b0b",
   330 => x"0bf5d53f",
   331 => x"823d0d04",
   332 => x"04fd3d0d",
   333 => x"80c3c008",
   334 => x"76b0ea29",
   335 => x"94120c54",
   336 => x"850b9815",
   337 => x"0c981408",
   338 => x"70810651",
   339 => x"5372f638",
   340 => x"853d0d04",
   341 => x"ff3d0d80",
   342 => x"c3c00874",
   343 => x"10107510",
   344 => x"0594120c",
   345 => x"52850b98",
   346 => x"130c9812",
   347 => x"08708106",
   348 => x"515170f6",
   349 => x"38833d0d",
   350 => x"04803d0d",
   351 => x"72518071",
   352 => x"278738ff",
   353 => x"115170fb",
   354 => x"38823d0d",
   355 => x"04803d0d",
   356 => x"80c3c008",
   357 => x"51870b84",
   358 => x"120c823d",
   359 => x"0d04803d",
   360 => x"0d80c3c4",
   361 => x"0851b60b",
   362 => x"8c120c83",
   363 => x"0b88120c",
   364 => x"823d0d04",
   365 => x"ff3d0d80",
   366 => x"c3c40852",
   367 => x"84120870",
   368 => x"81065151",
   369 => x"70802ef4",
   370 => x"38710870",
   371 => x"81ff0680",
   372 => x"0c51833d",
   373 => x"0d04fe3d",
   374 => x"0d029305",
   375 => x"3380c3c4",
   376 => x"08535384",
   377 => x"12087089",
   378 => x"2a708106",
   379 => x"51515170",
   380 => x"f2387272",
   381 => x"0c843d0d",
   382 => x"04fe3d0d",
   383 => x"02930533",
   384 => x"53728a2e",
   385 => x"9c3880c3",
   386 => x"c4085284",
   387 => x"12087089",
   388 => x"2a708106",
   389 => x"51515170",
   390 => x"f2387272",
   391 => x"0c843d0d",
   392 => x"0480c3c4",
   393 => x"08528412",
   394 => x"0870892a",
   395 => x"70810651",
   396 => x"515170f2",
   397 => x"388d720c",
   398 => x"84120870",
   399 => x"892a7081",
   400 => x"06515151",
   401 => x"70c538d2",
   402 => x"39fd3d0d",
   403 => x"75703352",
   404 => x"5470802e",
   405 => x"a8387080",
   406 => x"c3c40853",
   407 => x"53811454",
   408 => x"728a2e9d",
   409 => x"38841208",
   410 => x"70892a70",
   411 => x"81065151",
   412 => x"5170f238",
   413 => x"72720c73",
   414 => x"335372e1",
   415 => x"38853d0d",
   416 => x"04841208",
   417 => x"70892a70",
   418 => x"81065151",
   419 => x"5170f238",
   420 => x"8d720c84",
   421 => x"12087089",
   422 => x"2a708106",
   423 => x"51515170",
   424 => x"c438d139",
   425 => x"f53d0d7e",
   426 => x"028405b7",
   427 => x"05338c3d",
   428 => x"5b55578b",
   429 => x"53bf8452",
   430 => x"7851ae93",
   431 => x"3f825673",
   432 => x"882e9638",
   433 => x"84567390",
   434 => x"2e8f3888",
   435 => x"5673a02e",
   436 => x"88387456",
   437 => x"74802ea7",
   438 => x"3802a505",
   439 => x"58768f06",
   440 => x"54738926",
   441 => x"80cc3875",
   442 => x"18b01555",
   443 => x"55737534",
   444 => x"76842aff",
   445 => x"177081ff",
   446 => x"06585557",
   447 => x"75df3878",
   448 => x"79335557",
   449 => x"73802ea6",
   450 => x"387380c3",
   451 => x"c4085656",
   452 => x"81175775",
   453 => x"8a2eb738",
   454 => x"84150870",
   455 => x"892a8106",
   456 => x"595477f4",
   457 => x"3875750c",
   458 => x"76335675",
   459 => x"e3388d3d",
   460 => x"0d047518",
   461 => x"b7155555",
   462 => x"73753476",
   463 => x"842aff17",
   464 => x"7081ff06",
   465 => x"58555775",
   466 => x"ff9338ff",
   467 => x"b2398415",
   468 => x"0870892a",
   469 => x"81065954",
   470 => x"77f4388d",
   471 => x"750c8415",
   472 => x"0870892a",
   473 => x"81065954",
   474 => x"77ffad38",
   475 => x"ffb739f8",
   476 => x"3d0d7a7c",
   477 => x"59538073",
   478 => x"56577673",
   479 => x"2480dc38",
   480 => x"7717548a",
   481 => x"527451a8",
   482 => x"a53f8008",
   483 => x"b0055372",
   484 => x"74348117",
   485 => x"578a5274",
   486 => x"51a7ee3f",
   487 => x"80085580",
   488 => x"08de3880",
   489 => x"08779f2a",
   490 => x"1870812c",
   491 => x"5b565680",
   492 => x"79259e38",
   493 => x"7717ff05",
   494 => x"55751870",
   495 => x"33555374",
   496 => x"33733473",
   497 => x"75348116",
   498 => x"ff165656",
   499 => x"787624e9",
   500 => x"38761856",
   501 => x"8076348a",
   502 => x"3d0d04ad",
   503 => x"78708105",
   504 => x"5a347230",
   505 => x"78185555",
   506 => x"8a527451",
   507 => x"a7c03f80",
   508 => x"08b00553",
   509 => x"72743481",
   510 => x"17578a52",
   511 => x"7451a789",
   512 => x"3f800855",
   513 => x"8008fef8",
   514 => x"38ff9839",
   515 => x"803d0d80",
   516 => x"c3bc0851",
   517 => x"81ff0b88",
   518 => x"120c823d",
   519 => x"0d04fa3d",
   520 => x"0d785788",
   521 => x"80e0870b",
   522 => x"80c3bc08",
   523 => x"80c3c008",
   524 => x"56575574",
   525 => x"84170c76",
   526 => x"802e9838",
   527 => x"afd7c20b",
   528 => x"94150c85",
   529 => x"0b98150c",
   530 => x"98140870",
   531 => x"81065153",
   532 => x"72f63874",
   533 => x"9f2a7510",
   534 => x"0755d839",
   535 => x"fd3d0d80",
   536 => x"c3bc0854",
   537 => x"80d50b84",
   538 => x"150c80c3",
   539 => x"c4085284",
   540 => x"12088106",
   541 => x"5170802e",
   542 => x"f6387108",
   543 => x"7081ff06",
   544 => x"f6115254",
   545 => x"5170ae26",
   546 => x"8c387010",
   547 => x"1080c1cc",
   548 => x"05517008",
   549 => x"04841208",
   550 => x"70892a70",
   551 => x"81065151",
   552 => x"5170f238",
   553 => x"ab720c72",
   554 => x"8a2ea638",
   555 => x"84120870",
   556 => x"892a7081",
   557 => x"06515151",
   558 => x"70f23872",
   559 => x"720c8412",
   560 => x"0870892a",
   561 => x"81065153",
   562 => x"72f438ad",
   563 => x"720cff9f",
   564 => x"39841208",
   565 => x"70892a70",
   566 => x"81065151",
   567 => x"5170f238",
   568 => x"8d720c84",
   569 => x"12087089",
   570 => x"2a708106",
   571 => x"51515170",
   572 => x"ffba38c7",
   573 => x"3981ff0b",
   574 => x"84150cfe",
   575 => x"f23980ff",
   576 => x"0b84150c",
   577 => x"fee939bf",
   578 => x"0b84150c",
   579 => x"fee1399f",
   580 => x"0b84150c",
   581 => x"fed9398f",
   582 => x"0b84150c",
   583 => x"fed13987",
   584 => x"0b84150c",
   585 => x"fec93983",
   586 => x"0b84150c",
   587 => x"fec13981",
   588 => x"0b84150c",
   589 => x"feb93980",
   590 => x"0b84150c",
   591 => x"feb139ff",
   592 => x"3d0d80c3",
   593 => x"bc085271",
   594 => x"08708f06",
   595 => x"7071842b",
   596 => x"0784150c",
   597 => x"51517108",
   598 => x"708f0670",
   599 => x"71842b07",
   600 => x"84150c51",
   601 => x"51e139d5",
   602 => x"3d0d80c3",
   603 => x"b80858ff",
   604 => x"0b84190c",
   605 => x"fdaad50b",
   606 => x"88190c85",
   607 => x"adaad5aa",
   608 => x"0b8c190c",
   609 => x"a4b40b94",
   610 => x"190c8186",
   611 => x"a10b9819",
   612 => x"0cbf900b",
   613 => x"bf903355",
   614 => x"5773802e",
   615 => x"a7387380",
   616 => x"c3c40856",
   617 => x"56811757",
   618 => x"758a2e8d",
   619 => x"a3388415",
   620 => x"0870892a",
   621 => x"81065159",
   622 => x"78f43875",
   623 => x"750c7633",
   624 => x"5675e238",
   625 => x"bfa40bbf",
   626 => x"a4335557",
   627 => x"73802ea7",
   628 => x"3880c3c4",
   629 => x"08745755",
   630 => x"81175775",
   631 => x"8a2e8d91",
   632 => x"38841508",
   633 => x"70892a81",
   634 => x"06515978",
   635 => x"f4387575",
   636 => x"0c763356",
   637 => x"75e23877",
   638 => x"08a63d5a",
   639 => x"568b53bf",
   640 => x"84527851",
   641 => x"a7c93f88",
   642 => x"02840581",
   643 => x"91055957",
   644 => x"758f0654",
   645 => x"7389268c",
   646 => x"f9387618",
   647 => x"b0155555",
   648 => x"73753475",
   649 => x"842aff18",
   650 => x"7081ff06",
   651 => x"59565676",
   652 => x"df387879",
   653 => x"33555773",
   654 => x"802ea738",
   655 => x"80c3c408",
   656 => x"74575581",
   657 => x"1757758a",
   658 => x"2e8ce338",
   659 => x"84150870",
   660 => x"892a8106",
   661 => x"595977f4",
   662 => x"3875750c",
   663 => x"76335675",
   664 => x"e238bfb4",
   665 => x"0bbfb433",
   666 => x"55577380",
   667 => x"2ea73880",
   668 => x"c3c40874",
   669 => x"57558117",
   670 => x"57758a2e",
   671 => x"8cd13884",
   672 => x"15087089",
   673 => x"2a810659",
   674 => x"5977f438",
   675 => x"75750c76",
   676 => x"335675e2",
   677 => x"3880c3b8",
   678 => x"08841108",
   679 => x"a43d5b57",
   680 => x"578b53bf",
   681 => x"84527851",
   682 => x"a6a53f88",
   683 => x"02840581",
   684 => x"85055957",
   685 => x"758f0654",
   686 => x"73892691",
   687 => x"ac387618",
   688 => x"b0155555",
   689 => x"73753475",
   690 => x"842aff18",
   691 => x"7081ff06",
   692 => x"59565676",
   693 => x"df387879",
   694 => x"33555773",
   695 => x"802ea738",
   696 => x"80c3c408",
   697 => x"74575581",
   698 => x"1757758a",
   699 => x"2e8c8138",
   700 => x"84150870",
   701 => x"892a8106",
   702 => x"595977f4",
   703 => x"3875750c",
   704 => x"76335675",
   705 => x"e238bfc4",
   706 => x"0bbfc433",
   707 => x"55577380",
   708 => x"2ea73880",
   709 => x"c3c40874",
   710 => x"57558117",
   711 => x"57758a2e",
   712 => x"8bef3884",
   713 => x"15087089",
   714 => x"2a810659",
   715 => x"5977f438",
   716 => x"75750c76",
   717 => x"335675e2",
   718 => x"3880c3b8",
   719 => x"08881108",
   720 => x"a13d5b57",
   721 => x"578b53bf",
   722 => x"84527851",
   723 => x"a5813f88",
   724 => x"02840580",
   725 => x"f9055957",
   726 => x"758f0654",
   727 => x"7389268f",
   728 => x"ff387618",
   729 => x"b0155555",
   730 => x"73753475",
   731 => x"842aff18",
   732 => x"7081ff06",
   733 => x"59565676",
   734 => x"df387879",
   735 => x"33555773",
   736 => x"802ea738",
   737 => x"80c3c408",
   738 => x"74575581",
   739 => x"1757758a",
   740 => x"2e8b9f38",
   741 => x"84150870",
   742 => x"892a8106",
   743 => x"595977f4",
   744 => x"3875750c",
   745 => x"76335675",
   746 => x"e238bfd4",
   747 => x"0bbfd433",
   748 => x"55577380",
   749 => x"2ea73880",
   750 => x"c3c40874",
   751 => x"57558117",
   752 => x"57758a2e",
   753 => x"8b8d3884",
   754 => x"15087089",
   755 => x"2a810659",
   756 => x"5977f438",
   757 => x"75750c76",
   758 => x"335675e2",
   759 => x"3880c3b8",
   760 => x"088c1108",
   761 => x"9e3d5b57",
   762 => x"578b53bf",
   763 => x"84527851",
   764 => x"a3dd3f88",
   765 => x"02840580",
   766 => x"ed055957",
   767 => x"758f0654",
   768 => x"7389268e",
   769 => x"d2387618",
   770 => x"b0155555",
   771 => x"73753475",
   772 => x"842aff18",
   773 => x"7081ff06",
   774 => x"59565676",
   775 => x"df387879",
   776 => x"33555773",
   777 => x"802ea738",
   778 => x"80c3c408",
   779 => x"74575581",
   780 => x"1757758a",
   781 => x"2e8abd38",
   782 => x"84150870",
   783 => x"892a8106",
   784 => x"595977f4",
   785 => x"3875750c",
   786 => x"76335675",
   787 => x"e238bfe4",
   788 => x"0bbfe433",
   789 => x"55577380",
   790 => x"2ea73880",
   791 => x"c3c40874",
   792 => x"57558117",
   793 => x"57758a2e",
   794 => x"8aab3884",
   795 => x"15087089",
   796 => x"2a810659",
   797 => x"5977f438",
   798 => x"75750c76",
   799 => x"335675e2",
   800 => x"3880c3b8",
   801 => x"08901108",
   802 => x"9b3d5b57",
   803 => x"578b53bf",
   804 => x"84527851",
   805 => x"a2b93f88",
   806 => x"02840580",
   807 => x"e1055957",
   808 => x"758f0654",
   809 => x"7389268d",
   810 => x"a5387618",
   811 => x"b0155555",
   812 => x"73753475",
   813 => x"842aff18",
   814 => x"7081ff06",
   815 => x"59565676",
   816 => x"df387879",
   817 => x"33555773",
   818 => x"802ea738",
   819 => x"80c3c408",
   820 => x"74575581",
   821 => x"1757758a",
   822 => x"2e89db38",
   823 => x"84150870",
   824 => x"892a8106",
   825 => x"595977f4",
   826 => x"3875750c",
   827 => x"76335675",
   828 => x"e238bff4",
   829 => x"0bbff433",
   830 => x"55577380",
   831 => x"2ea73880",
   832 => x"c3c40874",
   833 => x"57558117",
   834 => x"57758a2e",
   835 => x"89c93884",
   836 => x"15087089",
   837 => x"2a810659",
   838 => x"5977f438",
   839 => x"75750c76",
   840 => x"335675e2",
   841 => x"3880c3b8",
   842 => x"08941108",
   843 => x"983d5b57",
   844 => x"578b53bf",
   845 => x"84527851",
   846 => x"a1953f88",
   847 => x"02840580",
   848 => x"d5055957",
   849 => x"758f0654",
   850 => x"7389268b",
   851 => x"f8387618",
   852 => x"b0155555",
   853 => x"73753475",
   854 => x"842aff18",
   855 => x"7081ff06",
   856 => x"59565676",
   857 => x"df387879",
   858 => x"33555773",
   859 => x"802ea738",
   860 => x"80c3c408",
   861 => x"74575581",
   862 => x"1757758a",
   863 => x"2e88f938",
   864 => x"84150870",
   865 => x"892a8106",
   866 => x"595977f4",
   867 => x"3875750c",
   868 => x"76335675",
   869 => x"e23880c0",
   870 => x"840b80c0",
   871 => x"84335557",
   872 => x"73802ea7",
   873 => x"3880c3c4",
   874 => x"08745755",
   875 => x"81175775",
   876 => x"8a2e88e5",
   877 => x"38841508",
   878 => x"70892a81",
   879 => x"06595977",
   880 => x"f4387575",
   881 => x"0c763356",
   882 => x"75e23880",
   883 => x"c3b80898",
   884 => x"1108953d",
   885 => x"5b57578b",
   886 => x"53bf8452",
   887 => x"78519fef",
   888 => x"3f880284",
   889 => x"0580c905",
   890 => x"5957758f",
   891 => x"06547389",
   892 => x"268ac938",
   893 => x"7618b015",
   894 => x"55557375",
   895 => x"3475842a",
   896 => x"ff187081",
   897 => x"ff065956",
   898 => x"5676df38",
   899 => x"78793355",
   900 => x"5773802e",
   901 => x"a73880c3",
   902 => x"c4087457",
   903 => x"55811757",
   904 => x"758a2e88",
   905 => x"95388415",
   906 => x"0870892a",
   907 => x"81065959",
   908 => x"77f43875",
   909 => x"750c7633",
   910 => x"5675e238",
   911 => x"80c0940b",
   912 => x"80c09433",
   913 => x"55577380",
   914 => x"2ea73880",
   915 => x"c3c40874",
   916 => x"57558117",
   917 => x"57758a2e",
   918 => x"88813884",
   919 => x"15087089",
   920 => x"2a810659",
   921 => x"5977f438",
   922 => x"75750c76",
   923 => x"335675e2",
   924 => x"3880c3b8",
   925 => x"089c1108",
   926 => x"923d5b57",
   927 => x"578b53bf",
   928 => x"84527851",
   929 => x"9ec93f88",
   930 => x"028405bd",
   931 => x"05595775",
   932 => x"8f065473",
   933 => x"8926899b",
   934 => x"387618b0",
   935 => x"15555573",
   936 => x"75347584",
   937 => x"2aff1870",
   938 => x"81ff0659",
   939 => x"565676df",
   940 => x"38787933",
   941 => x"55577380",
   942 => x"2ea73880",
   943 => x"c3c40874",
   944 => x"57558117",
   945 => x"57758a2e",
   946 => x"87b23884",
   947 => x"15087089",
   948 => x"2a810659",
   949 => x"5977f438",
   950 => x"75750c76",
   951 => x"335675e2",
   952 => x"3880c0a4",
   953 => x"0b80c0a4",
   954 => x"33555773",
   955 => x"802ea738",
   956 => x"80c3c408",
   957 => x"74575581",
   958 => x"1757758a",
   959 => x"2e879e38",
   960 => x"84150870",
   961 => x"892a8106",
   962 => x"595977f4",
   963 => x"3875750c",
   964 => x"76335675",
   965 => x"e23880c3",
   966 => x"b808a011",
   967 => x"088f3d5b",
   968 => x"57578b53",
   969 => x"bf845278",
   970 => x"519da43f",
   971 => x"88028405",
   972 => x"b1055957",
   973 => x"758f0654",
   974 => x"73892687",
   975 => x"ed387618",
   976 => x"b0155555",
   977 => x"73753475",
   978 => x"842aff18",
   979 => x"7081ff06",
   980 => x"59565676",
   981 => x"df387879",
   982 => x"33555773",
   983 => x"802ea738",
   984 => x"80c3c408",
   985 => x"74575581",
   986 => x"1757758a",
   987 => x"2e86cf38",
   988 => x"84150870",
   989 => x"892a8106",
   990 => x"595977f4",
   991 => x"3875750c",
   992 => x"76335675",
   993 => x"e23880c0",
   994 => x"b40b80c0",
   995 => x"b4335557",
   996 => x"73802ea7",
   997 => x"3880c3c4",
   998 => x"08745755",
   999 => x"81175775",
  1000 => x"8a2e86bb",
  1001 => x"38841508",
  1002 => x"70892a81",
  1003 => x"06595977",
  1004 => x"f4387575",
  1005 => x"0c763356",
  1006 => x"75e23880",
  1007 => x"c3b808a4",
  1008 => x"11088c3d",
  1009 => x"5b57578b",
  1010 => x"53bf8452",
  1011 => x"78519bff",
  1012 => x"3f880284",
  1013 => x"05a50559",
  1014 => x"57758f06",
  1015 => x"54738926",
  1016 => x"86bf3876",
  1017 => x"18b01555",
  1018 => x"55737534",
  1019 => x"75842aff",
  1020 => x"187081ff",
  1021 => x"06595656",
  1022 => x"76df3878",
  1023 => x"79335557",
  1024 => x"73802e86",
  1025 => x"ed3880c3",
  1026 => x"c4087457",
  1027 => x"55811757",
  1028 => x"758a2e85",
  1029 => x"eb388415",
  1030 => x"0870892a",
  1031 => x"81065959",
  1032 => x"77f43875",
  1033 => x"750c7633",
  1034 => x"5675e238",
  1035 => x"84150870",
  1036 => x"892a8106",
  1037 => x"575875f4",
  1038 => x"388d750c",
  1039 => x"84150870",
  1040 => x"892a8106",
  1041 => x"555673f4",
  1042 => x"388a750c",
  1043 => x"ad3d0d04",
  1044 => x"84150870",
  1045 => x"892a8106",
  1046 => x"515473f4",
  1047 => x"388d750c",
  1048 => x"84150870",
  1049 => x"892a8106",
  1050 => x"515978f2",
  1051 => x"c138f2cb",
  1052 => x"39841508",
  1053 => x"70892a81",
  1054 => x"06515473",
  1055 => x"f4388d75",
  1056 => x"0c841508",
  1057 => x"70892a81",
  1058 => x"06515978",
  1059 => x"f2d338f2",
  1060 => x"dd397618",
  1061 => x"b7155555",
  1062 => x"73753475",
  1063 => x"842aff18",
  1064 => x"7081ff06",
  1065 => x"59565676",
  1066 => x"f2e638f3",
  1067 => x"85398415",
  1068 => x"0870892a",
  1069 => x"81065959",
  1070 => x"77f4388d",
  1071 => x"750c8415",
  1072 => x"0870892a",
  1073 => x"81065959",
  1074 => x"77f38138",
  1075 => x"f38b3984",
  1076 => x"15087089",
  1077 => x"2a810659",
  1078 => x"5977f438",
  1079 => x"8d750c84",
  1080 => x"15087089",
  1081 => x"2a810659",
  1082 => x"5977f393",
  1083 => x"38f39d39",
  1084 => x"84150870",
  1085 => x"892a8106",
  1086 => x"595977f4",
  1087 => x"388d750c",
  1088 => x"84150870",
  1089 => x"892a8106",
  1090 => x"595977f3",
  1091 => x"e338f3ed",
  1092 => x"39841508",
  1093 => x"70892a81",
  1094 => x"06595977",
  1095 => x"f4388d75",
  1096 => x"0c841508",
  1097 => x"70892a81",
  1098 => x"06595977",
  1099 => x"f3f538f3",
  1100 => x"ff398415",
  1101 => x"0870892a",
  1102 => x"81065959",
  1103 => x"77f4388d",
  1104 => x"750c8415",
  1105 => x"0870892a",
  1106 => x"81065959",
  1107 => x"77f4c538",
  1108 => x"f4cf3984",
  1109 => x"15087089",
  1110 => x"2a810659",
  1111 => x"5977f438",
  1112 => x"8d750c84",
  1113 => x"15087089",
  1114 => x"2a810659",
  1115 => x"5977f4d7",
  1116 => x"38f4e139",
  1117 => x"84150870",
  1118 => x"892a8106",
  1119 => x"595977f4",
  1120 => x"388d750c",
  1121 => x"84150870",
  1122 => x"892a8106",
  1123 => x"595977f5",
  1124 => x"a738f5b1",
  1125 => x"39841508",
  1126 => x"70892a81",
  1127 => x"06595977",
  1128 => x"f4388d75",
  1129 => x"0c841508",
  1130 => x"70892a81",
  1131 => x"06595977",
  1132 => x"f5b938f5",
  1133 => x"c3398415",
  1134 => x"0870892a",
  1135 => x"81065959",
  1136 => x"77f4388d",
  1137 => x"750c8415",
  1138 => x"0870892a",
  1139 => x"81065959",
  1140 => x"77f68938",
  1141 => x"f6933984",
  1142 => x"15087089",
  1143 => x"2a810659",
  1144 => x"5977f438",
  1145 => x"8d750c84",
  1146 => x"15087089",
  1147 => x"2a810659",
  1148 => x"5977f69b",
  1149 => x"38f6a539",
  1150 => x"84150870",
  1151 => x"892a8106",
  1152 => x"595977f4",
  1153 => x"388d750c",
  1154 => x"84150870",
  1155 => x"892a8106",
  1156 => x"595977f6",
  1157 => x"eb38f6f5",
  1158 => x"39841508",
  1159 => x"70892a81",
  1160 => x"06595977",
  1161 => x"f4388d75",
  1162 => x"0c841508",
  1163 => x"70892a81",
  1164 => x"06595977",
  1165 => x"f6ff38f7",
  1166 => x"89398415",
  1167 => x"0870892a",
  1168 => x"81065959",
  1169 => x"77f4388d",
  1170 => x"750c8415",
  1171 => x"0870892a",
  1172 => x"81065959",
  1173 => x"77f7cf38",
  1174 => x"f7d93984",
  1175 => x"15087089",
  1176 => x"2a810659",
  1177 => x"5977f438",
  1178 => x"8d750c84",
  1179 => x"15087089",
  1180 => x"2a810659",
  1181 => x"5977f7e3",
  1182 => x"38f7ed39",
  1183 => x"84150870",
  1184 => x"892a8106",
  1185 => x"595977f4",
  1186 => x"388d750c",
  1187 => x"84150870",
  1188 => x"892a8106",
  1189 => x"595977f8",
  1190 => x"b238f8bc",
  1191 => x"39841508",
  1192 => x"70892a81",
  1193 => x"06595977",
  1194 => x"f4388d75",
  1195 => x"0c841508",
  1196 => x"70892a81",
  1197 => x"06595977",
  1198 => x"f8c638f8",
  1199 => x"d0398415",
  1200 => x"0870892a",
  1201 => x"81065959",
  1202 => x"77f4388d",
  1203 => x"750c8415",
  1204 => x"0870892a",
  1205 => x"81065959",
  1206 => x"77f99538",
  1207 => x"f99f3984",
  1208 => x"15087089",
  1209 => x"2a810659",
  1210 => x"5977f438",
  1211 => x"8d750c84",
  1212 => x"15087089",
  1213 => x"2a810659",
  1214 => x"5977f9a9",
  1215 => x"38f9b339",
  1216 => x"84150870",
  1217 => x"892a8106",
  1218 => x"595977f4",
  1219 => x"388d750c",
  1220 => x"84150870",
  1221 => x"892a8106",
  1222 => x"595977f9",
  1223 => x"f938fa83",
  1224 => x"397618b7",
  1225 => x"155555f9",
  1226 => x"c0397618",
  1227 => x"b7155555",
  1228 => x"f8923976",
  1229 => x"18b71555",
  1230 => x"55f6e439",
  1231 => x"7618b715",
  1232 => x"5555f5b6",
  1233 => x"397618b7",
  1234 => x"155555f4",
  1235 => x"87397618",
  1236 => x"b7155555",
  1237 => x"f2da3976",
  1238 => x"18b71555",
  1239 => x"55f1ad39",
  1240 => x"7618b715",
  1241 => x"5555f080",
  1242 => x"397618b7",
  1243 => x"155555ee",
  1244 => x"d33980c3",
  1245 => x"c4088411",
  1246 => x"0870892a",
  1247 => x"81065859",
  1248 => x"5575f9a8",
  1249 => x"38f9b239",
  1250 => x"fc3d0d02",
  1251 => x"9a052202",
  1252 => x"84059e05",
  1253 => x"22028805",
  1254 => x"a2052280",
  1255 => x"c3b80855",
  1256 => x"56545590",
  1257 => x"12087083",
  1258 => x"2a708106",
  1259 => x"51515170",
  1260 => x"f2387490",
  1261 => x"2b738b2b",
  1262 => x"0774862b",
  1263 => x"07810790",
  1264 => x"130c863d",
  1265 => x"0d04fd3d",
  1266 => x"0d029605",
  1267 => x"22028405",
  1268 => x"9a052280",
  1269 => x"c3b80854",
  1270 => x"54549012",
  1271 => x"0870832a",
  1272 => x"70810651",
  1273 => x"515170f2",
  1274 => x"38738b2b",
  1275 => x"73862b07",
  1276 => x"82079013",
  1277 => x"0c901208",
  1278 => x"70832a81",
  1279 => x"06555173",
  1280 => x"f4389012",
  1281 => x"0870902a",
  1282 => x"800c5485",
  1283 => x"3d0d04e3",
  1284 => x"3d0d80c0",
  1285 => x"c40b80c0",
  1286 => x"c4335557",
  1287 => x"73802ea7",
  1288 => x"387380c3",
  1289 => x"c4085656",
  1290 => x"81175775",
  1291 => x"8a2e86a9",
  1292 => x"38841508",
  1293 => x"70892a81",
  1294 => x"065b5c79",
  1295 => x"f4387575",
  1296 => x"0c763356",
  1297 => x"75e2389f",
  1298 => x"0b9d3d02",
  1299 => x"880580ed",
  1300 => x"059c3d02",
  1301 => x"900580e1",
  1302 => x"059b3d99",
  1303 => x"3d029c05",
  1304 => x"80c90502",
  1305 => x"a00580d5",
  1306 => x"05434044",
  1307 => x"455e445f",
  1308 => x"435c80c0",
  1309 => x"d80b80c0",
  1310 => x"d8335557",
  1311 => x"73802ea7",
  1312 => x"3880c3c4",
  1313 => x"08745755",
  1314 => x"81175775",
  1315 => x"8a2e85ea",
  1316 => x"38841508",
  1317 => x"70892a81",
  1318 => x"0640587e",
  1319 => x"f4387575",
  1320 => x"0c763356",
  1321 => x"75e2387b",
  1322 => x"568b53bf",
  1323 => x"84526151",
  1324 => x"929d3f82",
  1325 => x"57758f06",
  1326 => x"54738926",
  1327 => x"85dd3876",
  1328 => x"1db01555",
  1329 => x"55737534",
  1330 => x"75842aff",
  1331 => x"187081ff",
  1332 => x"06595656",
  1333 => x"76df3861",
  1334 => x"62335557",
  1335 => x"73802ea7",
  1336 => x"3880c3c4",
  1337 => x"08745755",
  1338 => x"81175775",
  1339 => x"8a2e85c7",
  1340 => x"38841508",
  1341 => x"70892a81",
  1342 => x"0640587e",
  1343 => x"f4387575",
  1344 => x"0c763356",
  1345 => x"75e23880",
  1346 => x"7c83ffff",
  1347 => x"06405880",
  1348 => x"c0e80b80",
  1349 => x"c0e83355",
  1350 => x"5773802e",
  1351 => x"a93880c3",
  1352 => x"c4087457",
  1353 => x"55811757",
  1354 => x"758a2e85",
  1355 => x"ab388415",
  1356 => x"0870892a",
  1357 => x"70810651",
  1358 => x"515473f2",
  1359 => x"3875750c",
  1360 => x"76335675",
  1361 => x"e0387756",
  1362 => x"8b53bf84",
  1363 => x"52605190",
  1364 => x"fe3f8257",
  1365 => x"758f0654",
  1366 => x"73892686",
  1367 => x"eb38761a",
  1368 => x"b0155555",
  1369 => x"73753475",
  1370 => x"842aff18",
  1371 => x"7081ff06",
  1372 => x"59565676",
  1373 => x"df386061",
  1374 => x"33555773",
  1375 => x"802ea938",
  1376 => x"80c3c408",
  1377 => x"74575581",
  1378 => x"1757758a",
  1379 => x"2e84ee38",
  1380 => x"84150870",
  1381 => x"892a7081",
  1382 => x"06515154",
  1383 => x"73f23875",
  1384 => x"750c7633",
  1385 => x"5675e038",
  1386 => x"80c0f40b",
  1387 => x"80c0f433",
  1388 => x"55577380",
  1389 => x"2ea93880",
  1390 => x"c3c40874",
  1391 => x"57558117",
  1392 => x"57758a2e",
  1393 => x"84dc3884",
  1394 => x"15087089",
  1395 => x"2a708106",
  1396 => x"51515473",
  1397 => x"f2387575",
  1398 => x"0c763356",
  1399 => x"75e03877",
  1400 => x"83ffff06",
  1401 => x"80c3b808",
  1402 => x"56569015",
  1403 => x"0870832a",
  1404 => x"81065157",
  1405 => x"76f4387e",
  1406 => x"8b2b7686",
  1407 => x"2b078207",
  1408 => x"90160c90",
  1409 => x"15087083",
  1410 => x"2a810658",
  1411 => x"5476f438",
  1412 => x"90150870",
  1413 => x"902a5757",
  1414 => x"8b53bf84",
  1415 => x"527f518f",
  1416 => x"ae3f8457",
  1417 => x"758f0654",
  1418 => x"73892685",
  1419 => x"9238761b",
  1420 => x"b0155555",
  1421 => x"73753475",
  1422 => x"842aff18",
  1423 => x"7081ff06",
  1424 => x"59565676",
  1425 => x"df387f60",
  1426 => x"33555773",
  1427 => x"802ea938",
  1428 => x"80c3c408",
  1429 => x"74575581",
  1430 => x"1757758a",
  1431 => x"2e83e838",
  1432 => x"84150870",
  1433 => x"892a7081",
  1434 => x"06515154",
  1435 => x"73f23875",
  1436 => x"750c7633",
  1437 => x"5675e038",
  1438 => x"80c0f40b",
  1439 => x"80c0f433",
  1440 => x"55577380",
  1441 => x"2ea93880",
  1442 => x"c3c40874",
  1443 => x"57558117",
  1444 => x"57758a2e",
  1445 => x"83d63884",
  1446 => x"15087089",
  1447 => x"2a708106",
  1448 => x"51515473",
  1449 => x"f2387575",
  1450 => x"0c763356",
  1451 => x"75e03880",
  1452 => x"c3b80890",
  1453 => x"11085757",
  1454 => x"8b53bf84",
  1455 => x"527d518e",
  1456 => x"8e3f8857",
  1457 => x"758f0654",
  1458 => x"73892683",
  1459 => x"e9387619",
  1460 => x"b0155555",
  1461 => x"73753475",
  1462 => x"842aff18",
  1463 => x"7081ff06",
  1464 => x"59565676",
  1465 => x"df387d7e",
  1466 => x"33555773",
  1467 => x"802ea938",
  1468 => x"80c3c408",
  1469 => x"74575581",
  1470 => x"1757758a",
  1471 => x"2e839238",
  1472 => x"84150870",
  1473 => x"892a7081",
  1474 => x"06515154",
  1475 => x"73f23875",
  1476 => x"750c7633",
  1477 => x"5675e038",
  1478 => x"77862e83",
  1479 => x"b4388118",
  1480 => x"589f7827",
  1481 => x"fbe93881",
  1482 => x"1c5c9f7c",
  1483 => x"27fac338",
  1484 => x"80c3c408",
  1485 => x"55841508",
  1486 => x"70892a81",
  1487 => x"065e407c",
  1488 => x"f4388d75",
  1489 => x"0c841508",
  1490 => x"70892a81",
  1491 => x"06425960",
  1492 => x"f4388a75",
  1493 => x"0c9f3d0d",
  1494 => x"04841508",
  1495 => x"70892a81",
  1496 => x"06555973",
  1497 => x"f4388d75",
  1498 => x"0c841508",
  1499 => x"70892a81",
  1500 => x"065b5c79",
  1501 => x"f9bb38f9",
  1502 => x"c5398415",
  1503 => x"0870892a",
  1504 => x"81064058",
  1505 => x"7ef4388d",
  1506 => x"750c8415",
  1507 => x"0870892a",
  1508 => x"81064058",
  1509 => x"7ef9fa38",
  1510 => x"fa843976",
  1511 => x"1db71555",
  1512 => x"55737534",
  1513 => x"75842aff",
  1514 => x"187081ff",
  1515 => x"06595656",
  1516 => x"76fa8238",
  1517 => x"faa13984",
  1518 => x"15087089",
  1519 => x"2a810640",
  1520 => x"587ef438",
  1521 => x"8d750c84",
  1522 => x"15087089",
  1523 => x"2a810640",
  1524 => x"587efa9d",
  1525 => x"38faa739",
  1526 => x"84150870",
  1527 => x"892a7081",
  1528 => x"06515154",
  1529 => x"73f2388d",
  1530 => x"750c8415",
  1531 => x"0870892a",
  1532 => x"70810651",
  1533 => x"515473fa",
  1534 => x"b538fac1",
  1535 => x"39841508",
  1536 => x"70892a70",
  1537 => x"81065151",
  1538 => x"5473f238",
  1539 => x"8d750c84",
  1540 => x"15087089",
  1541 => x"2a708106",
  1542 => x"51515473",
  1543 => x"faf238fa",
  1544 => x"fe398415",
  1545 => x"0870892a",
  1546 => x"70810651",
  1547 => x"515473f2",
  1548 => x"388d750c",
  1549 => x"84150870",
  1550 => x"892a7081",
  1551 => x"06515154",
  1552 => x"73fb8438",
  1553 => x"fb903984",
  1554 => x"15087089",
  1555 => x"2a708106",
  1556 => x"51515473",
  1557 => x"f2388d75",
  1558 => x"0c841508",
  1559 => x"70892a70",
  1560 => x"81065151",
  1561 => x"5473fbf8",
  1562 => x"38fc8439",
  1563 => x"84150870",
  1564 => x"892a7081",
  1565 => x"06515154",
  1566 => x"73f2388d",
  1567 => x"750c8415",
  1568 => x"0870892a",
  1569 => x"70810651",
  1570 => x"515473fc",
  1571 => x"8a38fc96",
  1572 => x"39841508",
  1573 => x"70892a70",
  1574 => x"81065151",
  1575 => x"5473f238",
  1576 => x"8d750c84",
  1577 => x"15087089",
  1578 => x"2a708106",
  1579 => x"51515473",
  1580 => x"fcce38fc",
  1581 => x"da397619",
  1582 => x"b7155555",
  1583 => x"fc963976",
  1584 => x"1bb71555",
  1585 => x"55faed39",
  1586 => x"761ab715",
  1587 => x"5555f994",
  1588 => x"399058f8",
  1589 => x"ba39fd3d",
  1590 => x"0d80c3bc",
  1591 => x"0854810b",
  1592 => x"84150c80",
  1593 => x"52fa8080",
  1594 => x"82805380",
  1595 => x"e4723173",
  1596 => x"70840555",
  1597 => x"0c811252",
  1598 => x"80c07226",
  1599 => x"ee38830b",
  1600 => x"84150cfa",
  1601 => x"80808280",
  1602 => x"0bfa8080",
  1603 => x"80840cb0",
  1604 => x"c00b850a",
  1605 => x"0c80c3b8",
  1606 => x"0852850a",
  1607 => x"0b94130c",
  1608 => x"91720c80",
  1609 => x"f59751ff",
  1610 => x"b5115170",
  1611 => x"8025f838",
  1612 => x"870b8415",
  1613 => x"0c850a08",
  1614 => x"708b2a84",
  1615 => x"160c5185",
  1616 => x"0a08708b",
  1617 => x"2a810653",
  1618 => x"5171f438",
  1619 => x"850a0870",
  1620 => x"8b2a8416",
  1621 => x"0c53853d",
  1622 => x"0d04fa3d",
  1623 => x"0d80c3bc",
  1624 => x"08700881",
  1625 => x"0a0680c3",
  1626 => x"c0085658",
  1627 => x"53870b84",
  1628 => x"150c80c3",
  1629 => x"c40854b6",
  1630 => x"0b8c150c",
  1631 => x"830b8815",
  1632 => x"0c81ff0b",
  1633 => x"88140c80",
  1634 => x"c0f80b80",
  1635 => x"c0f83354",
  1636 => x"5672802e",
  1637 => x"a4387255",
  1638 => x"81165674",
  1639 => x"8a2e81f1",
  1640 => x"38841408",
  1641 => x"70892a70",
  1642 => x"81065151",
  1643 => x"5372f238",
  1644 => x"74740c75",
  1645 => x"335574e0",
  1646 => x"3880c0fc",
  1647 => x"0b80c0fc",
  1648 => x"33545672",
  1649 => x"802ea438",
  1650 => x"72558116",
  1651 => x"56748a2e",
  1652 => x"81e43884",
  1653 => x"14087089",
  1654 => x"2a708106",
  1655 => x"51515372",
  1656 => x"f2387474",
  1657 => x"0c753355",
  1658 => x"74e03876",
  1659 => x"802e82b5",
  1660 => x"3880c188",
  1661 => x"0b80c188",
  1662 => x"33545672",
  1663 => x"802ea438",
  1664 => x"72558116",
  1665 => x"56748a2e",
  1666 => x"81d13884",
  1667 => x"14087089",
  1668 => x"2a708106",
  1669 => x"51515372",
  1670 => x"f2387474",
  1671 => x"0c753355",
  1672 => x"74e03880",
  1673 => x"c1980b80",
  1674 => x"c1983354",
  1675 => x"5672802e",
  1676 => x"a4387255",
  1677 => x"81165674",
  1678 => x"8a2e81c4",
  1679 => x"38841408",
  1680 => x"70892a70",
  1681 => x"81065151",
  1682 => x"5372f238",
  1683 => x"74740c75",
  1684 => x"335574e0",
  1685 => x"38fcff3f",
  1686 => x"8880e087",
  1687 => x"0b80c3bc",
  1688 => x"0880c3c0",
  1689 => x"08565755",
  1690 => x"7484170c",
  1691 => x"76802e98",
  1692 => x"38afd7c2",
  1693 => x"0b94150c",
  1694 => x"850b9815",
  1695 => x"0c981408",
  1696 => x"70810651",
  1697 => x"5372f638",
  1698 => x"749f2a75",
  1699 => x"100755d8",
  1700 => x"39841408",
  1701 => x"70892a70",
  1702 => x"81065151",
  1703 => x"5372f238",
  1704 => x"8d740c84",
  1705 => x"14087089",
  1706 => x"2a708106",
  1707 => x"51515372",
  1708 => x"fdef38fd",
  1709 => x"fb398414",
  1710 => x"0870892a",
  1711 => x"70810651",
  1712 => x"515372f2",
  1713 => x"388d740c",
  1714 => x"84140870",
  1715 => x"892a7081",
  1716 => x"06515153",
  1717 => x"72fdfc38",
  1718 => x"fe883984",
  1719 => x"14087089",
  1720 => x"2a708106",
  1721 => x"51515372",
  1722 => x"f2388d74",
  1723 => x"0c841408",
  1724 => x"70892a70",
  1725 => x"81065151",
  1726 => x"5372fe8f",
  1727 => x"38fe9b39",
  1728 => x"84140870",
  1729 => x"892a7081",
  1730 => x"06515153",
  1731 => x"72f2388d",
  1732 => x"740c8414",
  1733 => x"0870892a",
  1734 => x"70810651",
  1735 => x"515372fe",
  1736 => x"9c38fea8",
  1737 => x"3980c1bc",
  1738 => x"0b80c1bc",
  1739 => x"33545672",
  1740 => x"802efdef",
  1741 => x"38728117",
  1742 => x"5755748a",
  1743 => x"2ea73884",
  1744 => x"14087089",
  1745 => x"2a708106",
  1746 => x"51515372",
  1747 => x"f2387474",
  1748 => x"0c753355",
  1749 => x"74802efd",
  1750 => x"ca388116",
  1751 => x"56748a2e",
  1752 => x"098106db",
  1753 => x"38841408",
  1754 => x"70892a70",
  1755 => x"81065151",
  1756 => x"5372f238",
  1757 => x"8d740c84",
  1758 => x"14087089",
  1759 => x"2a708106",
  1760 => x"51515372",
  1761 => x"ffb938c6",
  1762 => x"398c0802",
  1763 => x"8c0cfd3d",
  1764 => x"0d80538c",
  1765 => x"088c0508",
  1766 => x"528c0888",
  1767 => x"05085182",
  1768 => x"de3f8008",
  1769 => x"70800c54",
  1770 => x"853d0d8c",
  1771 => x"0c048c08",
  1772 => x"028c0cfd",
  1773 => x"3d0d8153",
  1774 => x"8c088c05",
  1775 => x"08528c08",
  1776 => x"88050851",
  1777 => x"82b93f80",
  1778 => x"0870800c",
  1779 => x"54853d0d",
  1780 => x"8c0c048c",
  1781 => x"08028c0c",
  1782 => x"f93d0d80",
  1783 => x"0b8c08fc",
  1784 => x"050c8c08",
  1785 => x"88050880",
  1786 => x"25ab388c",
  1787 => x"08880508",
  1788 => x"308c0888",
  1789 => x"050c800b",
  1790 => x"8c08f405",
  1791 => x"0c8c08fc",
  1792 => x"05088838",
  1793 => x"810b8c08",
  1794 => x"f4050c8c",
  1795 => x"08f40508",
  1796 => x"8c08fc05",
  1797 => x"0c8c088c",
  1798 => x"05088025",
  1799 => x"ab388c08",
  1800 => x"8c050830",
  1801 => x"8c088c05",
  1802 => x"0c800b8c",
  1803 => x"08f0050c",
  1804 => x"8c08fc05",
  1805 => x"08883881",
  1806 => x"0b8c08f0",
  1807 => x"050c8c08",
  1808 => x"f005088c",
  1809 => x"08fc050c",
  1810 => x"80538c08",
  1811 => x"8c050852",
  1812 => x"8c088805",
  1813 => x"085181a7",
  1814 => x"3f800870",
  1815 => x"8c08f805",
  1816 => x"0c548c08",
  1817 => x"fc050880",
  1818 => x"2e8c388c",
  1819 => x"08f80508",
  1820 => x"308c08f8",
  1821 => x"050c8c08",
  1822 => x"f8050870",
  1823 => x"800c5489",
  1824 => x"3d0d8c0c",
  1825 => x"048c0802",
  1826 => x"8c0cfb3d",
  1827 => x"0d800b8c",
  1828 => x"08fc050c",
  1829 => x"8c088805",
  1830 => x"08802593",
  1831 => x"388c0888",
  1832 => x"0508308c",
  1833 => x"0888050c",
  1834 => x"810b8c08",
  1835 => x"fc050c8c",
  1836 => x"088c0508",
  1837 => x"80258c38",
  1838 => x"8c088c05",
  1839 => x"08308c08",
  1840 => x"8c050c81",
  1841 => x"538c088c",
  1842 => x"0508528c",
  1843 => x"08880508",
  1844 => x"51ad3f80",
  1845 => x"08708c08",
  1846 => x"f8050c54",
  1847 => x"8c08fc05",
  1848 => x"08802e8c",
  1849 => x"388c08f8",
  1850 => x"0508308c",
  1851 => x"08f8050c",
  1852 => x"8c08f805",
  1853 => x"0870800c",
  1854 => x"54873d0d",
  1855 => x"8c0c048c",
  1856 => x"08028c0c",
  1857 => x"fd3d0d81",
  1858 => x"0b8c08fc",
  1859 => x"050c800b",
  1860 => x"8c08f805",
  1861 => x"0c8c088c",
  1862 => x"05088c08",
  1863 => x"88050827",
  1864 => x"ac388c08",
  1865 => x"fc050880",
  1866 => x"2ea33880",
  1867 => x"0b8c088c",
  1868 => x"05082499",
  1869 => x"388c088c",
  1870 => x"0508108c",
  1871 => x"088c050c",
  1872 => x"8c08fc05",
  1873 => x"08108c08",
  1874 => x"fc050cc9",
  1875 => x"398c08fc",
  1876 => x"0508802e",
  1877 => x"80c9388c",
  1878 => x"088c0508",
  1879 => x"8c088805",
  1880 => x"0826a138",
  1881 => x"8c088805",
  1882 => x"088c088c",
  1883 => x"0508318c",
  1884 => x"0888050c",
  1885 => x"8c08f805",
  1886 => x"088c08fc",
  1887 => x"0508078c",
  1888 => x"08f8050c",
  1889 => x"8c08fc05",
  1890 => x"08812a8c",
  1891 => x"08fc050c",
  1892 => x"8c088c05",
  1893 => x"08812a8c",
  1894 => x"088c050c",
  1895 => x"ffaf398c",
  1896 => x"08900508",
  1897 => x"802e8f38",
  1898 => x"8c088805",
  1899 => x"08708c08",
  1900 => x"f4050c51",
  1901 => x"8d398c08",
  1902 => x"f8050870",
  1903 => x"8c08f405",
  1904 => x"0c518c08",
  1905 => x"f4050880",
  1906 => x"0c853d0d",
  1907 => x"8c0c04fc",
  1908 => x"3d0d7670",
  1909 => x"797b5555",
  1910 => x"55558f72",
  1911 => x"278c3872",
  1912 => x"75078306",
  1913 => x"5170802e",
  1914 => x"a738ff12",
  1915 => x"5271ff2e",
  1916 => x"98387270",
  1917 => x"81055433",
  1918 => x"74708105",
  1919 => x"5634ff12",
  1920 => x"5271ff2e",
  1921 => x"098106ea",
  1922 => x"3874800c",
  1923 => x"863d0d04",
  1924 => x"74517270",
  1925 => x"84055408",
  1926 => x"71708405",
  1927 => x"530c7270",
  1928 => x"84055408",
  1929 => x"71708405",
  1930 => x"530c7270",
  1931 => x"84055408",
  1932 => x"71708405",
  1933 => x"530c7270",
  1934 => x"84055408",
  1935 => x"71708405",
  1936 => x"530cf012",
  1937 => x"52718f26",
  1938 => x"c9388372",
  1939 => x"27953872",
  1940 => x"70840554",
  1941 => x"08717084",
  1942 => x"05530cfc",
  1943 => x"12527183",
  1944 => x"26ed3870",
  1945 => x"54ff8339",
  1946 => x"fd3d0d80",
  1947 => x"0b80c3ac",
  1948 => x"08545472",
  1949 => x"812e9a38",
  1950 => x"7380caf0",
  1951 => x"0ccbe03f",
  1952 => x"cafe3f80",
  1953 => x"c3c85281",
  1954 => x"51f5cf3f",
  1955 => x"800851a0",
  1956 => x"3f7280ca",
  1957 => x"f00ccbc7",
  1958 => x"3fcae53f",
  1959 => x"80c3c852",
  1960 => x"8151f5b6",
  1961 => x"3f800851",
  1962 => x"873f00ff",
  1963 => x"3900ff39",
  1964 => x"f73d0d7b",
  1965 => x"80c3cc08",
  1966 => x"82c81108",
  1967 => x"5a545a77",
  1968 => x"802e80da",
  1969 => x"38818818",
  1970 => x"841908ff",
  1971 => x"0581712b",
  1972 => x"59555980",
  1973 => x"742480ea",
  1974 => x"38807424",
  1975 => x"b5387382",
  1976 => x"2b781188",
  1977 => x"05565681",
  1978 => x"80190877",
  1979 => x"06537280",
  1980 => x"2eb63878",
  1981 => x"16700853",
  1982 => x"53795174",
  1983 => x"0853722d",
  1984 => x"ff14fc17",
  1985 => x"fc177981",
  1986 => x"2c5a5757",
  1987 => x"54738025",
  1988 => x"d6387708",
  1989 => x"5877ffad",
  1990 => x"3880c3cc",
  1991 => x"0853bc13",
  1992 => x"08a53879",
  1993 => x"51ff833f",
  1994 => x"74085372",
  1995 => x"2dff14fc",
  1996 => x"17fc1779",
  1997 => x"812c5a57",
  1998 => x"57547380",
  1999 => x"25ffa838",
  2000 => x"d1398057",
  2001 => x"ff933972",
  2002 => x"51bc1308",
  2003 => x"53722d79",
  2004 => x"51fed73f",
  2005 => x"ff3d0d80",
  2006 => x"cad00bfc",
  2007 => x"05700852",
  2008 => x"5270ff2e",
  2009 => x"9138702d",
  2010 => x"fc127008",
  2011 => x"525270ff",
  2012 => x"2e098106",
  2013 => x"f138833d",
  2014 => x"0d0404ca",
  2015 => x"cf3f0400",
  2016 => x"00000040",
  2017 => x"30782020",
  2018 => x"20202020",
  2019 => x"20200000",
  2020 => x"0a677265",
  2021 => x"74682072",
  2022 => x"65676973",
  2023 => x"74657273",
  2024 => x"3a000000",
  2025 => x"0a636f6e",
  2026 => x"74726f6c",
  2027 => x"3a202020",
  2028 => x"20202000",
  2029 => x"0a737461",
  2030 => x"7475733a",
  2031 => x"20202020",
  2032 => x"20202000",
  2033 => x"0a6d6163",
  2034 => x"5f6d7362",
  2035 => x"3a202020",
  2036 => x"20202000",
  2037 => x"0a6d6163",
  2038 => x"5f6c7362",
  2039 => x"3a202020",
  2040 => x"20202000",
  2041 => x"0a6d6469",
  2042 => x"6f5f636f",
  2043 => x"6e74726f",
  2044 => x"6c3a2000",
  2045 => x"0a74785f",
  2046 => x"706f696e",
  2047 => x"7465723a",
  2048 => x"20202000",
  2049 => x"0a72785f",
  2050 => x"706f696e",
  2051 => x"7465723a",
  2052 => x"20202000",
  2053 => x"0a656463",
  2054 => x"6c5f6970",
  2055 => x"3a202020",
  2056 => x"20202000",
  2057 => x"0a686173",
  2058 => x"685f6d73",
  2059 => x"623a2020",
  2060 => x"20202000",
  2061 => x"0a686173",
  2062 => x"685f6c73",
  2063 => x"623a2020",
  2064 => x"20202000",
  2065 => x"0a6d6469",
  2066 => x"6f207068",
  2067 => x"79207265",
  2068 => x"67697374",
  2069 => x"65727300",
  2070 => x"0a206d64",
  2071 => x"696f2070",
  2072 => x"68793a20",
  2073 => x"00000000",
  2074 => x"0a202072",
  2075 => x"65673a20",
  2076 => x"00000000",
  2077 => x"2d3e2000",
  2078 => x"0a0a0000",
  2079 => x"5a505520",
  2080 => x"74657374",
  2081 => x"20000000",
  2082 => x"286f6e20",
  2083 => x"73696d75",
  2084 => x"6c61746f",
  2085 => x"72290a00",
  2086 => x"636f6d70",
  2087 => x"696c6564",
  2088 => x"3a204175",
  2089 => x"67202039",
  2090 => x"20323031",
  2091 => x"30202031",
  2092 => x"383a3034",
  2093 => x"3a30390a",
  2094 => x"00000000",
  2095 => x"286f6e20",
  2096 => x"68617264",
  2097 => x"77617265",
  2098 => x"290a0000",
  2099 => x"0000086f",
  2100 => x"00000895",
  2101 => x"00000895",
  2102 => x"0000086f",
  2103 => x"00000895",
  2104 => x"00000895",
  2105 => x"00000895",
  2106 => x"00000895",
  2107 => x"00000895",
  2108 => x"00000895",
  2109 => x"00000895",
  2110 => x"00000895",
  2111 => x"00000895",
  2112 => x"00000895",
  2113 => x"00000895",
  2114 => x"00000895",
  2115 => x"00000895",
  2116 => x"00000895",
  2117 => x"00000895",
  2118 => x"00000895",
  2119 => x"00000895",
  2120 => x"00000895",
  2121 => x"00000895",
  2122 => x"00000895",
  2123 => x"00000895",
  2124 => x"00000895",
  2125 => x"00000895",
  2126 => x"00000895",
  2127 => x"00000895",
  2128 => x"00000895",
  2129 => x"00000895",
  2130 => x"00000895",
  2131 => x"00000895",
  2132 => x"00000895",
  2133 => x"00000895",
  2134 => x"00000895",
  2135 => x"00000895",
  2136 => x"00000895",
  2137 => x"00000937",
  2138 => x"0000092f",
  2139 => x"00000927",
  2140 => x"0000091f",
  2141 => x"00000917",
  2142 => x"0000090f",
  2143 => x"00000907",
  2144 => x"000008fe",
  2145 => x"000008f5",
  2146 => x"64756d6d",
  2147 => x"792e6578",
  2148 => x"65000000",
  2149 => x"43000000",
  2150 => x"00ffffff",
  2151 => x"ff00ffff",
  2152 => x"ffff00ff",
  2153 => x"ffffff00",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00002558",
  2158 => x"80000c00",
  2159 => x"80000800",
  2160 => x"80000200",
  2161 => x"80000100",
  2162 => x"00002188",
  2163 => x"000021d0",
  2164 => x"00000000",
  2165 => x"00002438",
  2166 => x"00002494",
  2167 => x"000024f0",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00002194",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000001",
  2207 => x"330eabcd",
  2208 => x"1234e66d",
  2209 => x"deec0005",
  2210 => x"000b0000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"00000000",
  2265 => x"00000000",
  2266 => x"00000000",
  2267 => x"00000000",
  2268 => x"00000000",
  2269 => x"00000000",
  2270 => x"00000000",
  2271 => x"00000000",
  2272 => x"00000000",
  2273 => x"00000000",
  2274 => x"00000000",
  2275 => x"00000000",
  2276 => x"00000000",
  2277 => x"00000000",
  2278 => x"00000000",
  2279 => x"00000000",
  2280 => x"00000000",
  2281 => x"00000000",
  2282 => x"00000000",
  2283 => x"00000000",
  2284 => x"00000000",
  2285 => x"00000000",
  2286 => x"00000000",
  2287 => x"00000000",
  2288 => x"00000000",
  2289 => x"00000000",
  2290 => x"00000000",
  2291 => x"00000000",
  2292 => x"00000000",
  2293 => x"00000000",
  2294 => x"00000000",
  2295 => x"00000000",
  2296 => x"00000000",
  2297 => x"00000000",
  2298 => x"00000000",
  2299 => x"00000000",
  2300 => x"00000000",
  2301 => x"00000000",
  2302 => x"00000000",
  2303 => x"00000000",
  2304 => x"00000000",
  2305 => x"00000000",
  2306 => x"00000000",
  2307 => x"00000000",
  2308 => x"00000000",
  2309 => x"00000000",
  2310 => x"00000000",
  2311 => x"00000000",
  2312 => x"00000000",
  2313 => x"00000000",
  2314 => x"00000000",
  2315 => x"00000000",
  2316 => x"00000000",
  2317 => x"00000000",
  2318 => x"00000000",
  2319 => x"00000000",
  2320 => x"00000000",
  2321 => x"00000000",
  2322 => x"00000000",
  2323 => x"00000000",
  2324 => x"00000000",
  2325 => x"00000000",
  2326 => x"00000000",
  2327 => x"00000000",
  2328 => x"00000000",
  2329 => x"00000000",
  2330 => x"00000000",
  2331 => x"00000000",
  2332 => x"00000000",
  2333 => x"00000000",
  2334 => x"00000000",
  2335 => x"00000000",
  2336 => x"00000000",
  2337 => x"00000000",
  2338 => x"00000000",
  2339 => x"00000000",
  2340 => x"00000000",
  2341 => x"00000000",
  2342 => x"00000000",
  2343 => x"00000000",
  2344 => x"00000000",
  2345 => x"00000000",
  2346 => x"00000000",
  2347 => x"00000000",
  2348 => x"00000000",
  2349 => x"00000000",
  2350 => x"00000000",
  2351 => x"00000000",
  2352 => x"00000000",
  2353 => x"00000000",
  2354 => x"00000000",
  2355 => x"00000000",
  2356 => x"00000000",
  2357 => x"00000000",
  2358 => x"00000000",
  2359 => x"00000000",
  2360 => x"00000000",
  2361 => x"00000000",
  2362 => x"00000000",
  2363 => x"00000000",
  2364 => x"00000000",
  2365 => x"00000000",
  2366 => x"00000000",
  2367 => x"00000000",
  2368 => x"00000000",
  2369 => x"00000000",
  2370 => x"00000000",
  2371 => x"00000000",
  2372 => x"00000000",
  2373 => x"00000000",
  2374 => x"00000000",
  2375 => x"00000000",
  2376 => x"00000000",
  2377 => x"00000000",
  2378 => x"00000000",
  2379 => x"00000000",
  2380 => x"00000000",
  2381 => x"00000000",
  2382 => x"00000000",
  2383 => x"00000000",
  2384 => x"00000000",
  2385 => x"00000000",
  2386 => x"00000000",
  2387 => x"ffffffff",
  2388 => x"00000000",
  2389 => x"ffffffff",
  2390 => x"00000000",
  2391 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
