-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80e2980c",
     3 => x"3a0b0b80",
     4 => x"d2890400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80d2d22d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80e2",
   162 => x"84738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80cc",
   171 => x"f42d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80ce",
   179 => x"a62d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80e2940c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"cbf33f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80e29408",
   281 => x"802ea438",
   282 => x"80e29808",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80e9",
   286 => x"d40c82a0",
   287 => x"800b80e9",
   288 => x"d80c8290",
   289 => x"800b80e9",
   290 => x"dc0c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"e9d40cf8",
   294 => x"80808280",
   295 => x"0b80e9d8",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"e9dc0c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80e9d40c",
   302 => x"80c0a880",
   303 => x"940b80e9",
   304 => x"d80c0b0b",
   305 => x"80d4a80b",
   306 => x"80e9dc0c",
   307 => x"04ff3d0d",
   308 => x"80e9e033",
   309 => x"5170a738",
   310 => x"80e2a008",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"e2a00c70",
   315 => x"2d80e2a0",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80e9",
   319 => x"e034833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80e9d008",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"e9d0510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404fb3d",
   333 => x"0d775680",
   334 => x"55747627",
   335 => x"81993880",
   336 => x"e2b40854",
   337 => x"bfa9bc0b",
   338 => x"94150c85",
   339 => x"0b98150c",
   340 => x"98140870",
   341 => x"81065153",
   342 => x"72f638bf",
   343 => x"a9bc0b94",
   344 => x"150c850b",
   345 => x"98150c98",
   346 => x"14087081",
   347 => x"06515372",
   348 => x"f638bfa9",
   349 => x"bc0b9415",
   350 => x"0c850b98",
   351 => x"150c9814",
   352 => x"08708106",
   353 => x"515372f6",
   354 => x"38bfa9bc",
   355 => x"0b94150c",
   356 => x"850b9815",
   357 => x"0c981408",
   358 => x"70810651",
   359 => x"5372f638",
   360 => x"bfa9bc0b",
   361 => x"94150c85",
   362 => x"0b98150c",
   363 => x"98140870",
   364 => x"81065153",
   365 => x"72f638bf",
   366 => x"a9bc0b94",
   367 => x"150c850b",
   368 => x"98150c98",
   369 => x"14087081",
   370 => x"06515372",
   371 => x"f6388115",
   372 => x"55757526",
   373 => x"feee3887",
   374 => x"3d0d0480",
   375 => x"3d0d80e2",
   376 => x"b4085187",
   377 => x"0b84120c",
   378 => x"823d0d04",
   379 => x"f83d0d7a",
   380 => x"7c595380",
   381 => x"73565776",
   382 => x"732480de",
   383 => x"38771754",
   384 => x"8a527451",
   385 => x"80c0c83f",
   386 => x"8008b005",
   387 => x"53727434",
   388 => x"8117578a",
   389 => x"52745180",
   390 => x"c0903f80",
   391 => x"08558008",
   392 => x"dc388008",
   393 => x"779f2a18",
   394 => x"70812c5b",
   395 => x"56568079",
   396 => x"259e3877",
   397 => x"17ff0555",
   398 => x"75187033",
   399 => x"55537433",
   400 => x"73347375",
   401 => x"348116ff",
   402 => x"16565678",
   403 => x"7624e938",
   404 => x"76185680",
   405 => x"76348a3d",
   406 => x"0d04ad78",
   407 => x"7081055a",
   408 => x"34723078",
   409 => x"1855558a",
   410 => x"527451bf",
   411 => x"e23f8008",
   412 => x"b0055372",
   413 => x"74348117",
   414 => x"578a5274",
   415 => x"51bfab3f",
   416 => x"80085580",
   417 => x"08fef638",
   418 => x"ff9839f9",
   419 => x"3d0d7970",
   420 => x"71337081",
   421 => x"ff065455",
   422 => x"55557080",
   423 => x"2eb13880",
   424 => x"e2b80852",
   425 => x"7281ff06",
   426 => x"81155553",
   427 => x"728a2e80",
   428 => x"f5388412",
   429 => x"0870822a",
   430 => x"81065257",
   431 => x"70802ef2",
   432 => x"3872720c",
   433 => x"73337081",
   434 => x"ff065953",
   435 => x"77d63874",
   436 => x"75335256",
   437 => x"70802e80",
   438 => x"c9387080",
   439 => x"e2b00859",
   440 => x"53811680",
   441 => x"e9e83370",
   442 => x"81ff0670",
   443 => x"10101180",
   444 => x"e9ec3370",
   445 => x"81ff0672",
   446 => x"90291170",
   447 => x"882b7a07",
   448 => x"7f0c5359",
   449 => x"59545458",
   450 => x"56728a2e",
   451 => x"be387380",
   452 => x"cf2eb838",
   453 => x"81155372",
   454 => x"80e9ec34",
   455 => x"75335372",
   456 => x"c038893d",
   457 => x"0d048412",
   458 => x"0870822a",
   459 => x"81065758",
   460 => x"75802ef2",
   461 => x"388d720c",
   462 => x"84120870",
   463 => x"822a8106",
   464 => x"52577080",
   465 => x"2efeeb38",
   466 => x"fef73971",
   467 => x"a3269938",
   468 => x"81175271",
   469 => x"80e9e834",
   470 => x"800b80e9",
   471 => x"ec347533",
   472 => x"5372fefd",
   473 => x"38ffbb39",
   474 => x"800b80e9",
   475 => x"e834800b",
   476 => x"80e9ec34",
   477 => x"e939fd3d",
   478 => x"0d80e2ac",
   479 => x"085480d5",
   480 => x"0b84150c",
   481 => x"80e2b808",
   482 => x"52841208",
   483 => x"81065170",
   484 => x"802ef638",
   485 => x"71087081",
   486 => x"ff06f611",
   487 => x"52545170",
   488 => x"ae268c38",
   489 => x"70101080",
   490 => x"e0840551",
   491 => x"70080484",
   492 => x"12087082",
   493 => x"2a708106",
   494 => x"51515170",
   495 => x"802ef038",
   496 => x"ab720c72",
   497 => x"8a2eaa38",
   498 => x"84120870",
   499 => x"822a7081",
   500 => x"06515151",
   501 => x"70802ef0",
   502 => x"3872720c",
   503 => x"84120870",
   504 => x"822a8106",
   505 => x"51537280",
   506 => x"2ef238ad",
   507 => x"720cff99",
   508 => x"39841208",
   509 => x"70822a70",
   510 => x"81065151",
   511 => x"5170802e",
   512 => x"f0388d72",
   513 => x"0c841208",
   514 => x"70822a70",
   515 => x"81065151",
   516 => x"5170802e",
   517 => x"ffb238c1",
   518 => x"3981ff0b",
   519 => x"84150cfe",
   520 => x"e83980ff",
   521 => x"0b84150c",
   522 => x"fedf39bf",
   523 => x"0b84150c",
   524 => x"fed7399f",
   525 => x"0b84150c",
   526 => x"fecf398f",
   527 => x"0b84150c",
   528 => x"fec73987",
   529 => x"0b84150c",
   530 => x"febf3983",
   531 => x"0b84150c",
   532 => x"feb73981",
   533 => x"0b84150c",
   534 => x"feaf3980",
   535 => x"0b84150c",
   536 => x"fea739d7",
   537 => x"3d0d80e2",
   538 => x"b0085580",
   539 => x"0b84160c",
   540 => x"fe800a0b",
   541 => x"88160c80",
   542 => x"0b80e9e8",
   543 => x"34800b80",
   544 => x"e9ec34a6",
   545 => x"3d705380",
   546 => x"e2a8088c",
   547 => x"11085355",
   548 => x"5bfad93f",
   549 => x"80d7d40b",
   550 => x"80d7d433",
   551 => x"555a7380",
   552 => x"2e80cc38",
   553 => x"80e2b008",
   554 => x"74575c81",
   555 => x"1a80e9e8",
   556 => x"337081ff",
   557 => x"06701010",
   558 => x"1180e9ec",
   559 => x"337081ff",
   560 => x"06729029",
   561 => x"1170882b",
   562 => x"7d07630c",
   563 => x"445c5c42",
   564 => x"575a5a75",
   565 => x"8a2e87bc",
   566 => x"387680cf",
   567 => x"2e87b538",
   568 => x"81185776",
   569 => x"80e9ec34",
   570 => x"79335675",
   571 => x"ffbd387a",
   572 => x"7b33555a",
   573 => x"73802e80",
   574 => x"cc3880e2",
   575 => x"b0087457",
   576 => x"5b811a80",
   577 => x"e9e83370",
   578 => x"81ff0670",
   579 => x"10101180",
   580 => x"e9ec3370",
   581 => x"81ff0672",
   582 => x"90291170",
   583 => x"882b7d07",
   584 => x"620c465c",
   585 => x"5c44575a",
   586 => x"5a758a2e",
   587 => x"87843876",
   588 => x"80cf2e86",
   589 => x"fd388118",
   590 => x"597880e9",
   591 => x"ec347933",
   592 => x"5675ffbd",
   593 => x"3880d7ec",
   594 => x"0b80d7ec",
   595 => x"33555a73",
   596 => x"802e80cc",
   597 => x"3880e2b0",
   598 => x"0874575b",
   599 => x"811a80e9",
   600 => x"e8337081",
   601 => x"ff067010",
   602 => x"101180e9",
   603 => x"ec337081",
   604 => x"ff067290",
   605 => x"29117088",
   606 => x"2b7d0762",
   607 => x"0c495c5c",
   608 => x"57575a5a",
   609 => x"758a2e85",
   610 => x"ed387680",
   611 => x"cf2e85e6",
   612 => x"3881185d",
   613 => x"7c80e9ec",
   614 => x"34793356",
   615 => x"75ffbd38",
   616 => x"80e2a808",
   617 => x"7008a53d",
   618 => x"5b575a8b",
   619 => x"5380d4ac",
   620 => x"527851bd",
   621 => x"bb3f8202",
   622 => x"84058189",
   623 => x"05595775",
   624 => x"8f065473",
   625 => x"89268592",
   626 => x"387618b0",
   627 => x"15555573",
   628 => x"75347584",
   629 => x"2aff1870",
   630 => x"81ff0659",
   631 => x"5c5676df",
   632 => x"38787933",
   633 => x"555a7380",
   634 => x"2e80cc38",
   635 => x"80e2b008",
   636 => x"74575b81",
   637 => x"1a80e9e8",
   638 => x"337081ff",
   639 => x"06701010",
   640 => x"1180e9ec",
   641 => x"337081ff",
   642 => x"06729029",
   643 => x"1170882b",
   644 => x"7d07620c",
   645 => x"455c5c5f",
   646 => x"575a5a75",
   647 => x"8a2e87f3",
   648 => x"387680cf",
   649 => x"2e87ec38",
   650 => x"81185776",
   651 => x"80e9ec34",
   652 => x"79335675",
   653 => x"ffbd3880",
   654 => x"d7f80b80",
   655 => x"d7f83355",
   656 => x"5a73802e",
   657 => x"80cc3880",
   658 => x"e2b00874",
   659 => x"575b811a",
   660 => x"80e9e833",
   661 => x"7081ff06",
   662 => x"70101011",
   663 => x"80e9ec33",
   664 => x"7081ff06",
   665 => x"72902911",
   666 => x"70882b7d",
   667 => x"07620c47",
   668 => x"5c5c4557",
   669 => x"5a5a758a",
   670 => x"2e87b638",
   671 => x"7680cf2e",
   672 => x"87af3881",
   673 => x"18597880",
   674 => x"e9ec3479",
   675 => x"335675ff",
   676 => x"bd38805f",
   677 => x"890a5cac",
   678 => x"3d087f2e",
   679 => x"09810687",
   680 => x"ca387ea1",
   681 => x"3d028805",
   682 => x"80fd0540",
   683 => x"415d7cbf",
   684 => x"06436285",
   685 => x"d43880d7",
   686 => x"cc0b80d7",
   687 => x"cc33555a",
   688 => x"73802e80",
   689 => x"cc3880e2",
   690 => x"b0087457",
   691 => x"5b811a80",
   692 => x"e9e83370",
   693 => x"81ff0670",
   694 => x"10101180",
   695 => x"e9ec3370",
   696 => x"81ff0672",
   697 => x"90291170",
   698 => x"882b7d07",
   699 => x"620c475c",
   700 => x"5c45575a",
   701 => x"5a758a2e",
   702 => x"848a3876",
   703 => x"80cf2e84",
   704 => x"83388118",
   705 => x"567580e9",
   706 => x"ec347933",
   707 => x"5675ffbd",
   708 => x"387b568b",
   709 => x"5380d4ac",
   710 => x"527f51ba",
   711 => x"d33f8857",
   712 => x"758f0654",
   713 => x"73892683",
   714 => x"d238761e",
   715 => x"b0155555",
   716 => x"73753475",
   717 => x"842aff18",
   718 => x"7081ff06",
   719 => x"595b5676",
   720 => x"df387f60",
   721 => x"33555a73",
   722 => x"802e85bf",
   723 => x"3880e2b0",
   724 => x"0874575b",
   725 => x"811a80e9",
   726 => x"e8337081",
   727 => x"ff067010",
   728 => x"101180e9",
   729 => x"ec337081",
   730 => x"ff067290",
   731 => x"29117088",
   732 => x"2b7d0762",
   733 => x"0c5a5c5c",
   734 => x"44575a5a",
   735 => x"758a2e83",
   736 => x"bf387680",
   737 => x"cf2e83b8",
   738 => x"38811859",
   739 => x"7880e9ec",
   740 => x"34793356",
   741 => x"75ffbd38",
   742 => x"80d7fc0b",
   743 => x"80d7fc33",
   744 => x"555a7380",
   745 => x"2e80c738",
   746 => x"7356811a",
   747 => x"80e9e833",
   748 => x"7081ff06",
   749 => x"70101011",
   750 => x"80e9ec33",
   751 => x"7081ff06",
   752 => x"72902911",
   753 => x"70882b7d",
   754 => x"07620c49",
   755 => x"5c5c5757",
   756 => x"5a5a758a",
   757 => x"2e82cb38",
   758 => x"7680cf2e",
   759 => x"82c43881",
   760 => x"18557480",
   761 => x"e9ec3479",
   762 => x"335675ff",
   763 => x"bd387b08",
   764 => x"7c327030",
   765 => x"7107709f",
   766 => x"2a7081ff",
   767 => x"06b01170",
   768 => x"81ff0680",
   769 => x"e9e83370",
   770 => x"81ff0670",
   771 => x"10101180",
   772 => x"e9ec3370",
   773 => x"81ff0672",
   774 => x"90291170",
   775 => x"882b7707",
   776 => x"670c4e58",
   777 => x"595c535f",
   778 => x"465a5259",
   779 => x"5b58608a",
   780 => x"2e83a438",
   781 => x"7680cf2e",
   782 => x"839d3881",
   783 => x"18416080",
   784 => x"e9ec3479",
   785 => x"1f841d81",
   786 => x"1f5f5d5f",
   787 => x"8fff7d27",
   788 => x"fcdc387e",
   789 => x"800cab3d",
   790 => x"0d047618",
   791 => x"b7155555",
   792 => x"73753475",
   793 => x"842aff18",
   794 => x"7081ff06",
   795 => x"595c5676",
   796 => x"facd38fa",
   797 => x"ec3974a3",
   798 => x"2680f138",
   799 => x"81195574",
   800 => x"80e9e834",
   801 => x"800b80e9",
   802 => x"ec347933",
   803 => x"5675f9cc",
   804 => x"38fa8d39",
   805 => x"74a32680",
   806 => x"c4388119",
   807 => x"567580e9",
   808 => x"e834800b",
   809 => x"80e9ec34",
   810 => x"79335675",
   811 => x"f7fd38f8",
   812 => x"be3974a3",
   813 => x"26993881",
   814 => x"19587780",
   815 => x"e9e83480",
   816 => x"0b80e9ec",
   817 => x"34793356",
   818 => x"75f8b638",
   819 => x"f8f73980",
   820 => x"0b80e9e8",
   821 => x"34800b80",
   822 => x"e9ec34e9",
   823 => x"39800b80",
   824 => x"e9e83480",
   825 => x"0b80e9ec",
   826 => x"34ffbd39",
   827 => x"800b80e9",
   828 => x"e834800b",
   829 => x"80e9ec34",
   830 => x"ff903976",
   831 => x"1eb71555",
   832 => x"55fcad39",
   833 => x"74a32680",
   834 => x"f1388119",
   835 => x"557480e9",
   836 => x"e834800b",
   837 => x"80e9ec34",
   838 => x"79335675",
   839 => x"fbaf38fb",
   840 => x"f03974a3",
   841 => x"2680c438",
   842 => x"81195877",
   843 => x"80e9e834",
   844 => x"800b80e9",
   845 => x"ec347933",
   846 => x"5675fcee",
   847 => x"38fdaf39",
   848 => x"74a32699",
   849 => x"38811957",
   850 => x"7680e9e8",
   851 => x"34800b80",
   852 => x"e9ec3479",
   853 => x"335675fb",
   854 => x"fb38fcbc",
   855 => x"39800b80",
   856 => x"e9e83480",
   857 => x"0b80e9ec",
   858 => x"34e93980",
   859 => x"0b80e9e8",
   860 => x"34800b80",
   861 => x"e9ec34ff",
   862 => x"bd39800b",
   863 => x"80e9e834",
   864 => x"800b80e9",
   865 => x"ec34ff90",
   866 => x"3980e2b0",
   867 => x"087c087d",
   868 => x"32703071",
   869 => x"07709f2a",
   870 => x"7081ff06",
   871 => x"b0117081",
   872 => x"ff0680e9",
   873 => x"e8337081",
   874 => x"ff067010",
   875 => x"101180e9",
   876 => x"ec337081",
   877 => x"ff067290",
   878 => x"29117088",
   879 => x"2b77077d",
   880 => x"0c4f5859",
   881 => x"5d534047",
   882 => x"5b525a5c",
   883 => x"595b608a",
   884 => x"2e098106",
   885 => x"fcde3875",
   886 => x"a326a238",
   887 => x"81195b7a",
   888 => x"80e9e834",
   889 => x"800b80e9",
   890 => x"ec34791f",
   891 => x"841d811f",
   892 => x"5f5d5f8f",
   893 => x"ff7d27f9",
   894 => x"b538fcd7",
   895 => x"39800b80",
   896 => x"e9e83480",
   897 => x"0b80e9ec",
   898 => x"34e03980",
   899 => x"e2b0085b",
   900 => x"fb863974",
   901 => x"a32680c4",
   902 => x"38811956",
   903 => x"7580e9e8",
   904 => x"34800b80",
   905 => x"e9ec3479",
   906 => x"335675f7",
   907 => x"c638f887",
   908 => x"3974a326",
   909 => x"99388119",
   910 => x"587780e9",
   911 => x"e834800b",
   912 => x"80e9ec34",
   913 => x"79335675",
   914 => x"f88438f8",
   915 => x"c539800b",
   916 => x"80e9e834",
   917 => x"800b80e9",
   918 => x"ec34e939",
   919 => x"800b80e9",
   920 => x"e834800b",
   921 => x"80e9ec34",
   922 => x"ffbd397b",
   923 => x"7f9f3d02",
   924 => x"8c0580f1",
   925 => x"05983d02",
   926 => x"940580cd",
   927 => x"05454245",
   928 => x"43445d80",
   929 => x"d7cc0b80",
   930 => x"d7cc3355",
   931 => x"5a73802e",
   932 => x"80cc3880",
   933 => x"e2b00874",
   934 => x"575b811a",
   935 => x"80e9e833",
   936 => x"7081ff06",
   937 => x"70101011",
   938 => x"80e9ec33",
   939 => x"7081ff06",
   940 => x"72902911",
   941 => x"70882b7d",
   942 => x"07620c5a",
   943 => x"5c5c5f57",
   944 => x"5a5a758a",
   945 => x"2e848338",
   946 => x"7680cf2e",
   947 => x"83fc3881",
   948 => x"18577680",
   949 => x"e9ec3479",
   950 => x"335675ff",
   951 => x"bd387c56",
   952 => x"8b5380d4",
   953 => x"ac526051",
   954 => x"b3863f88",
   955 => x"57758f06",
   956 => x"54738926",
   957 => x"83cb3861",
   958 => x"17b01555",
   959 => x"55737534",
   960 => x"75842aff",
   961 => x"187081ff",
   962 => x"06595b56",
   963 => x"76df3860",
   964 => x"6133555a",
   965 => x"73802e84",
   966 => x"e33880e2",
   967 => x"b0087457",
   968 => x"5b811a80",
   969 => x"e9e83370",
   970 => x"81ff0670",
   971 => x"10101180",
   972 => x"e9ec3370",
   973 => x"81ff0672",
   974 => x"90291170",
   975 => x"882b7d07",
   976 => x"620c425c",
   977 => x"5c57575a",
   978 => x"5a758a2e",
   979 => x"839a3876",
   980 => x"80cf2e83",
   981 => x"93388118",
   982 => x"597880e9",
   983 => x"ec347933",
   984 => x"5675ffbd",
   985 => x"3880e9e8",
   986 => x"337081ff",
   987 => x"06701010",
   988 => x"1180e9ec",
   989 => x"337081ff",
   990 => x"06729029",
   991 => x"1170882b",
   992 => x"a007610c",
   993 => x"41595a56",
   994 => x"57587480",
   995 => x"cf2e84a0",
   996 => x"38811756",
   997 => x"7580e9ec",
   998 => x"347c0870",
   999 => x"585ca353",
  1000 => x"80d4b852",
  1001 => x"7d51b1c8",
  1002 => x"3fa0567f",
  1003 => x"1677b106",
  1004 => x"b0075659",
  1005 => x"74793476",
  1006 => x"0a100aff",
  1007 => x"177081ff",
  1008 => x"06585957",
  1009 => x"75e5387d",
  1010 => x"7e33555a",
  1011 => x"73802e84",
  1012 => x"883880e2",
  1013 => x"b0087457",
  1014 => x"5b811a80",
  1015 => x"e9e83370",
  1016 => x"81ff0670",
  1017 => x"10101180",
  1018 => x"e9ec3370",
  1019 => x"81ff0672",
  1020 => x"90291170",
  1021 => x"882b7d07",
  1022 => x"620c535c",
  1023 => x"5c57575a",
  1024 => x"5a758a2e",
  1025 => x"82803876",
  1026 => x"80cf2e81",
  1027 => x"f9388118",
  1028 => x"567580e9",
  1029 => x"ec347933",
  1030 => x"5675ffbd",
  1031 => x"3880e9e8",
  1032 => x"337081ff",
  1033 => x"06701010",
  1034 => x"1180e9ec",
  1035 => x"337081ff",
  1036 => x"06729029",
  1037 => x"1170882b",
  1038 => x"a007610c",
  1039 => x"5a5e5a56",
  1040 => x"57587980",
  1041 => x"cf2e83c5",
  1042 => x"38811758",
  1043 => x"7780e9ec",
  1044 => x"347c7c2e",
  1045 => x"83d43880",
  1046 => x"d8800b80",
  1047 => x"d8803355",
  1048 => x"5a73802e",
  1049 => x"80c73873",
  1050 => x"56811a80",
  1051 => x"e9e83370",
  1052 => x"81ff0670",
  1053 => x"10101180",
  1054 => x"e9ec3370",
  1055 => x"81ff0672",
  1056 => x"90291170",
  1057 => x"882b7d07",
  1058 => x"620c425c",
  1059 => x"5c57575a",
  1060 => x"5a758a2e",
  1061 => x"818d3876",
  1062 => x"80cf2e81",
  1063 => x"86388118",
  1064 => x"577680e9",
  1065 => x"ec347933",
  1066 => x"5675ffbd",
  1067 => x"38841d63",
  1068 => x"8105445d",
  1069 => x"9f6327fb",
  1070 => x"ca387e80",
  1071 => x"0cab3d0d",
  1072 => x"046117b7",
  1073 => x"155555fc",
  1074 => x"b43974a3",
  1075 => x"26818038",
  1076 => x"81195675",
  1077 => x"80e9e834",
  1078 => x"800b80e9",
  1079 => x"ec347933",
  1080 => x"5675fbb6",
  1081 => x"38fbf739",
  1082 => x"74a32680",
  1083 => x"f1388119",
  1084 => x"587780e9",
  1085 => x"e834800b",
  1086 => x"80e9ec34",
  1087 => x"79335675",
  1088 => x"fc9f38fc",
  1089 => x"e03974a3",
  1090 => x"26b73881",
  1091 => x"19577680",
  1092 => x"e9e83480",
  1093 => x"0b80e9ec",
  1094 => x"34793356",
  1095 => x"75fdba38",
  1096 => x"fdfb3974",
  1097 => x"a32680c5",
  1098 => x"38811955",
  1099 => x"7480e9e8",
  1100 => x"34800b80",
  1101 => x"e9ec3479",
  1102 => x"335675fe",
  1103 => x"ac38feed",
  1104 => x"39800b80",
  1105 => x"e9e83480",
  1106 => x"0b80e9ec",
  1107 => x"34cb3980",
  1108 => x"0b80e9e8",
  1109 => x"34800b80",
  1110 => x"e9ec34ff",
  1111 => x"8139800b",
  1112 => x"80e9e834",
  1113 => x"800b80e9",
  1114 => x"ec34ff90",
  1115 => x"39800b80",
  1116 => x"e9e83480",
  1117 => x"0b80e9ec",
  1118 => x"34ffbc39",
  1119 => x"80e2b008",
  1120 => x"80e9e833",
  1121 => x"7081ff06",
  1122 => x"70101011",
  1123 => x"80e9ec33",
  1124 => x"7081ff06",
  1125 => x"72902911",
  1126 => x"70882ba0",
  1127 => x"07770c42",
  1128 => x"5a5b5758",
  1129 => x"595b7480",
  1130 => x"cf2e0981",
  1131 => x"06fbe238",
  1132 => x"75a32682",
  1133 => x"b8388118",
  1134 => x"5b7a80e9",
  1135 => x"e834800b",
  1136 => x"80e9ec34",
  1137 => x"7c087058",
  1138 => x"5ca35380",
  1139 => x"d4b8527d",
  1140 => x"51ad9d3f",
  1141 => x"a056fbd3",
  1142 => x"3980e2b0",
  1143 => x"0880e9e8",
  1144 => x"337081ff",
  1145 => x"06701010",
  1146 => x"1180e9ec",
  1147 => x"337081ff",
  1148 => x"06729029",
  1149 => x"1170882b",
  1150 => x"a007770c",
  1151 => x"5b5f5b57",
  1152 => x"58595b79",
  1153 => x"80cf2e09",
  1154 => x"8106fcbd",
  1155 => x"3875a326",
  1156 => x"81cc3881",
  1157 => x"18577680",
  1158 => x"e9e83480",
  1159 => x"0b80e9ec",
  1160 => x"347c7c2e",
  1161 => x"098106fc",
  1162 => x"ae3880d8",
  1163 => x"880b80d8",
  1164 => x"8833555a",
  1165 => x"73802efc",
  1166 => x"f4387381",
  1167 => x"1b80e9e8",
  1168 => x"337081ff",
  1169 => x"06701010",
  1170 => x"1180e9ec",
  1171 => x"337081ff",
  1172 => x"06729029",
  1173 => x"1170882b",
  1174 => x"7807630c",
  1175 => x"5b5d5d40",
  1176 => x"585b5b56",
  1177 => x"758a2e80",
  1178 => x"ca387680",
  1179 => x"cf2e80c3",
  1180 => x"38811859",
  1181 => x"7880e9ec",
  1182 => x"34793356",
  1183 => x"75802efc",
  1184 => x"ac38811a",
  1185 => x"80e9e833",
  1186 => x"7081ff06",
  1187 => x"70101011",
  1188 => x"80e9ec33",
  1189 => x"7081ff06",
  1190 => x"72902911",
  1191 => x"70882b7d",
  1192 => x"07620c5a",
  1193 => x"5c5c5f57",
  1194 => x"5a5a758a",
  1195 => x"2e098106",
  1196 => x"ffb83874",
  1197 => x"a3269938",
  1198 => x"81195675",
  1199 => x"80e9e834",
  1200 => x"800b80e9",
  1201 => x"ec347933",
  1202 => x"5675ffb6",
  1203 => x"38fbde39",
  1204 => x"800b80e9",
  1205 => x"e834800b",
  1206 => x"80e9ec34",
  1207 => x"e939800b",
  1208 => x"80e9e834",
  1209 => x"800b80e9",
  1210 => x"ec34feb5",
  1211 => x"39800b80",
  1212 => x"e9e83480",
  1213 => x"0b80e9ec",
  1214 => x"34fdc939",
  1215 => x"d93d0d80",
  1216 => x"d89051e7",
  1217 => x"863f80e2",
  1218 => x"a4087008",
  1219 => x"80d8a053",
  1220 => x"5d55e6f7",
  1221 => x"3fa63d70",
  1222 => x"537c81ff",
  1223 => x"ff06525d",
  1224 => x"e5ca3f7c",
  1225 => x"51e6e43f",
  1226 => x"80d8b451",
  1227 => x"e6dd3f7b",
  1228 => x"8f2a8106",
  1229 => x"a43d5a56",
  1230 => x"8b5380d4",
  1231 => x"ac527851",
  1232 => x"aaae3f82",
  1233 => x"02840581",
  1234 => x"89055957",
  1235 => x"758f0654",
  1236 => x"73892687",
  1237 => x"fc387618",
  1238 => x"b0155555",
  1239 => x"73753475",
  1240 => x"842aff18",
  1241 => x"7081ff06",
  1242 => x"595b5676",
  1243 => x"df387879",
  1244 => x"33555773",
  1245 => x"802ea938",
  1246 => x"7380e2b8",
  1247 => x"08565681",
  1248 => x"1757758a",
  1249 => x"2e87e638",
  1250 => x"84150870",
  1251 => x"822a8106",
  1252 => x"5b5b7980",
  1253 => x"2ef23875",
  1254 => x"750c7633",
  1255 => x"5675e038",
  1256 => x"78793355",
  1257 => x"5a73802e",
  1258 => x"80cc3873",
  1259 => x"80e2b008",
  1260 => x"5c56811a",
  1261 => x"80e9e833",
  1262 => x"7081ff06",
  1263 => x"70101011",
  1264 => x"80e9ec33",
  1265 => x"7081ff06",
  1266 => x"72902911",
  1267 => x"70882b7d",
  1268 => x"07620c53",
  1269 => x"5c5c5757",
  1270 => x"5a5a758a",
  1271 => x"2e87cf38",
  1272 => x"7680cf2e",
  1273 => x"87c83881",
  1274 => x"18577680",
  1275 => x"e9ec3479",
  1276 => x"335675ff",
  1277 => x"bd3880d8",
  1278 => x"c851e58f",
  1279 => x"3f7b902a",
  1280 => x"8106a13d",
  1281 => x"5a568b53",
  1282 => x"80d4ac52",
  1283 => x"7851a8e0",
  1284 => x"3f820284",
  1285 => x"0580fd05",
  1286 => x"5957758f",
  1287 => x"06547389",
  1288 => x"2686ef38",
  1289 => x"7618b015",
  1290 => x"55557375",
  1291 => x"3475842a",
  1292 => x"ff187081",
  1293 => x"ff065956",
  1294 => x"5676df38",
  1295 => x"78793355",
  1296 => x"5773802e",
  1297 => x"a93880e2",
  1298 => x"b8087457",
  1299 => x"55811757",
  1300 => x"758a2e87",
  1301 => x"84388415",
  1302 => x"0870822a",
  1303 => x"81065558",
  1304 => x"73802ef2",
  1305 => x"3875750c",
  1306 => x"76335675",
  1307 => x"e0387879",
  1308 => x"33555a73",
  1309 => x"802e80cc",
  1310 => x"3880e2b0",
  1311 => x"0874575b",
  1312 => x"811a80e9",
  1313 => x"e8337081",
  1314 => x"ff067010",
  1315 => x"101180e9",
  1316 => x"ec337081",
  1317 => x"ff067290",
  1318 => x"29117088",
  1319 => x"2b7d0762",
  1320 => x"0c535c5c",
  1321 => x"57575a5a",
  1322 => x"758a2e93",
  1323 => x"bb387680",
  1324 => x"cf2e93b4",
  1325 => x"38811857",
  1326 => x"7680e9ec",
  1327 => x"34793356",
  1328 => x"75ffbd38",
  1329 => x"80d8dc51",
  1330 => x"e3c13f7b",
  1331 => x"952a8306",
  1332 => x"5473812e",
  1333 => x"95993881",
  1334 => x"742694ff",
  1335 => x"3873822e",
  1336 => x"95ab3873",
  1337 => x"832e90d7",
  1338 => x"3880d8f0",
  1339 => x"51e39c3f",
  1340 => x"7c527b97",
  1341 => x"2a870683",
  1342 => x"0581712b",
  1343 => x"525ae1ec",
  1344 => x"3f7c51e3",
  1345 => x"863f80d9",
  1346 => x"8451e2ff",
  1347 => x"3f80d98c",
  1348 => x"51e2f83f",
  1349 => x"7c527b9a",
  1350 => x"2a810681",
  1351 => x"0551e1cc",
  1352 => x"3f7c51e2",
  1353 => x"e63f80d9",
  1354 => x"a051e2df",
  1355 => x"3f7c527b",
  1356 => x"9b2a8706",
  1357 => x"830551e1",
  1358 => x"b33f7c51",
  1359 => x"e2cd3f80",
  1360 => x"d9b451e2",
  1361 => x"c63f7c52",
  1362 => x"7b9e2a82",
  1363 => x"0751e19c",
  1364 => x"3f7c51e2",
  1365 => x"b63f80d9",
  1366 => x"c851e2af",
  1367 => x"3f7b9f2a",
  1368 => x"9e3d5a56",
  1369 => x"8b5380d4",
  1370 => x"ac527851",
  1371 => x"a6823f82",
  1372 => x"02840580",
  1373 => x"f1055957",
  1374 => x"758f0654",
  1375 => x"73892690",
  1376 => x"d7387618",
  1377 => x"b0155555",
  1378 => x"73753475",
  1379 => x"842aff18",
  1380 => x"7081ff06",
  1381 => x"595d5676",
  1382 => x"df387879",
  1383 => x"33555773",
  1384 => x"802ea938",
  1385 => x"80e2b808",
  1386 => x"74575581",
  1387 => x"1757758a",
  1388 => x"2e84cb38",
  1389 => x"84150870",
  1390 => x"822a8106",
  1391 => x"59547780",
  1392 => x"2ef23875",
  1393 => x"750c7633",
  1394 => x"5675e038",
  1395 => x"78793355",
  1396 => x"5a73802e",
  1397 => x"80cc3880",
  1398 => x"e2b00874",
  1399 => x"575b811a",
  1400 => x"80e9e833",
  1401 => x"7081ff06",
  1402 => x"70101011",
  1403 => x"80e9ec33",
  1404 => x"7081ff06",
  1405 => x"72902911",
  1406 => x"70882b7d",
  1407 => x"07620c5a",
  1408 => x"5c5c5f57",
  1409 => x"5a5a758a",
  1410 => x"2e91b738",
  1411 => x"7680cf2e",
  1412 => x"91b03881",
  1413 => x"18577680",
  1414 => x"e9ec3479",
  1415 => x"335675ff",
  1416 => x"bd3880e2",
  1417 => x"a4088411",
  1418 => x"0880d9dc",
  1419 => x"535658e0",
  1420 => x"da3f7c52",
  1421 => x"749fff06",
  1422 => x"51dfb13f",
  1423 => x"7c51e0cb",
  1424 => x"3f80d9f0",
  1425 => x"51e0c43f",
  1426 => x"7c52748c",
  1427 => x"2a870683",
  1428 => x"0581712b",
  1429 => x"525bdf94",
  1430 => x"3f7c51e0",
  1431 => x"ae3f80da",
  1432 => x"8451e0a7",
  1433 => x"3f748f2a",
  1434 => x"81069b3d",
  1435 => x"5a568b53",
  1436 => x"80d4ac52",
  1437 => x"7851a3f8",
  1438 => x"3f820284",
  1439 => x"0580e505",
  1440 => x"5957758f",
  1441 => x"06547389",
  1442 => x"268efa38",
  1443 => x"7618b015",
  1444 => x"55557375",
  1445 => x"3475842a",
  1446 => x"ff187081",
  1447 => x"ff065955",
  1448 => x"5676df38",
  1449 => x"78793355",
  1450 => x"5773802e",
  1451 => x"a93880e2",
  1452 => x"b8087457",
  1453 => x"55811757",
  1454 => x"758a2e82",
  1455 => x"e6388415",
  1456 => x"0870822a",
  1457 => x"8106595c",
  1458 => x"77802ef2",
  1459 => x"3875750c",
  1460 => x"76335675",
  1461 => x"e0387879",
  1462 => x"33555a73",
  1463 => x"802e80cc",
  1464 => x"3880e2b0",
  1465 => x"0874575b",
  1466 => x"811a80e9",
  1467 => x"e8337081",
  1468 => x"ff067010",
  1469 => x"101180e9",
  1470 => x"ec337081",
  1471 => x"ff067290",
  1472 => x"29117088",
  1473 => x"2b7d0762",
  1474 => x"0c425c5c",
  1475 => x"57575a5a",
  1476 => x"758a2e8d",
  1477 => x"f9387680",
  1478 => x"cf2e8df2",
  1479 => x"38811857",
  1480 => x"7680e9ec",
  1481 => x"34793356",
  1482 => x"75ffbd38",
  1483 => x"80e2a408",
  1484 => x"88110880",
  1485 => x"da985356",
  1486 => x"59ded03f",
  1487 => x"74870654",
  1488 => x"73862682",
  1489 => x"83387310",
  1490 => x"1080e1c0",
  1491 => x"055b7a08",
  1492 => x"047618b7",
  1493 => x"15555573",
  1494 => x"75347584",
  1495 => x"2aff1870",
  1496 => x"81ff0659",
  1497 => x"5b5676f7",
  1498 => x"e338f882",
  1499 => x"39841508",
  1500 => x"70822a81",
  1501 => x"06595477",
  1502 => x"802ef238",
  1503 => x"8d750c84",
  1504 => x"15087082",
  1505 => x"2a81065b",
  1506 => x"5b79802e",
  1507 => x"f7fa38f8",
  1508 => x"86397618",
  1509 => x"b7155555",
  1510 => x"73753475",
  1511 => x"842aff18",
  1512 => x"7081ff06",
  1513 => x"59565676",
  1514 => x"f8f038f9",
  1515 => x"8f3974a3",
  1516 => x"26993881",
  1517 => x"19567580",
  1518 => x"e9e83480",
  1519 => x"0b80e9ec",
  1520 => x"34793356",
  1521 => x"75f7eb38",
  1522 => x"f8ac3980",
  1523 => x"0b80e9e8",
  1524 => x"34800b80",
  1525 => x"e9ec34e9",
  1526 => x"39841508",
  1527 => x"70822a81",
  1528 => x"065b5b79",
  1529 => x"802ef238",
  1530 => x"8d750c84",
  1531 => x"15087082",
  1532 => x"2a810655",
  1533 => x"5873802e",
  1534 => x"f8dc38f8",
  1535 => x"e8398415",
  1536 => x"0870822a",
  1537 => x"8106555a",
  1538 => x"73802ef2",
  1539 => x"388d750c",
  1540 => x"84150870",
  1541 => x"822a8106",
  1542 => x"59547780",
  1543 => x"2efb9538",
  1544 => x"fba13984",
  1545 => x"15087082",
  1546 => x"2a81065d",
  1547 => x"5a7b802e",
  1548 => x"f2388d75",
  1549 => x"0c841508",
  1550 => x"70822a81",
  1551 => x"06595c77",
  1552 => x"802efcfa",
  1553 => x"38fd8639",
  1554 => x"80daac51",
  1555 => x"dcbd3f80",
  1556 => x"dab451dc",
  1557 => x"b63f80da",
  1558 => x"bc51dcaf",
  1559 => x"3f74832a",
  1560 => x"83065473",
  1561 => x"812e8dfd",
  1562 => x"38817426",
  1563 => x"8de33873",
  1564 => x"822e8e85",
  1565 => x"3873832e",
  1566 => x"89973880",
  1567 => x"dad051dc",
  1568 => x"8a3f80da",
  1569 => x"d451dc83",
  1570 => x"3f74852a",
  1571 => x"87065473",
  1572 => x"812e89a1",
  1573 => x"38817426",
  1574 => x"8dad3873",
  1575 => x"822e8de3",
  1576 => x"3873832e",
  1577 => x"88e13880",
  1578 => x"dae851db",
  1579 => x"de3f7490",
  1580 => x"2a870654",
  1581 => x"7385268c",
  1582 => x"38731010",
  1583 => x"80e1dc05",
  1584 => x"54730804",
  1585 => x"80daac51",
  1586 => x"dbc13f80",
  1587 => x"dafc51db",
  1588 => x"ba3f7c52",
  1589 => x"74932a83",
  1590 => x"06820751",
  1591 => x"da8e3f7c",
  1592 => x"51dba83f",
  1593 => x"80db9051",
  1594 => x"dba13f7c",
  1595 => x"5274942a",
  1596 => x"8f0651d9",
  1597 => x"f73f7c51",
  1598 => x"db913f80",
  1599 => x"dba451db",
  1600 => x"8a3f7c52",
  1601 => x"74982a81",
  1602 => x"06810551",
  1603 => x"d9de3f7c",
  1604 => x"51daf83f",
  1605 => x"80dbb851",
  1606 => x"daf13f7c",
  1607 => x"52749e2a",
  1608 => x"820751d9",
  1609 => x"c73f7c51",
  1610 => x"dae13f80",
  1611 => x"dbcc51da",
  1612 => x"da3f749f",
  1613 => x"2a983d5a",
  1614 => x"568b5380",
  1615 => x"d4ac5278",
  1616 => x"519ead3f",
  1617 => x"82028405",
  1618 => x"80d90559",
  1619 => x"57758f06",
  1620 => x"54738926",
  1621 => x"89a63876",
  1622 => x"18b01555",
  1623 => x"55737534",
  1624 => x"75842aff",
  1625 => x"187081ff",
  1626 => x"06595e56",
  1627 => x"76df3878",
  1628 => x"79335557",
  1629 => x"73802ea9",
  1630 => x"3880e2b8",
  1631 => x"08745755",
  1632 => x"81175775",
  1633 => x"8a2e85eb",
  1634 => x"38841508",
  1635 => x"70822a81",
  1636 => x"065d5d7b",
  1637 => x"802ef238",
  1638 => x"75750c76",
  1639 => x"335675e0",
  1640 => x"38787933",
  1641 => x"555a7380",
  1642 => x"2e80cc38",
  1643 => x"80e2b008",
  1644 => x"74575b81",
  1645 => x"1a80e9e8",
  1646 => x"337081ff",
  1647 => x"06701010",
  1648 => x"1180e9ec",
  1649 => x"337081ff",
  1650 => x"06729029",
  1651 => x"1170882b",
  1652 => x"7d07620c",
  1653 => x"5a5c5c40",
  1654 => x"575a5a75",
  1655 => x"8a2e88ea",
  1656 => x"387680cf",
  1657 => x"2e88e338",
  1658 => x"81185675",
  1659 => x"80e9ec34",
  1660 => x"79335675",
  1661 => x"ffbd3880",
  1662 => x"e2a40890",
  1663 => x"110880db",
  1664 => x"e0535859",
  1665 => x"d9853f76",
  1666 => x"953d5a56",
  1667 => x"8b5380d4",
  1668 => x"ac527851",
  1669 => x"9cda3f88",
  1670 => x"02840580",
  1671 => x"cd055957",
  1672 => x"758f0654",
  1673 => x"73892687",
  1674 => x"ca387618",
  1675 => x"b0155555",
  1676 => x"73753475",
  1677 => x"842aff18",
  1678 => x"7081ff06",
  1679 => x"595c5676",
  1680 => x"df387879",
  1681 => x"33555773",
  1682 => x"802ea938",
  1683 => x"80e2b808",
  1684 => x"74575581",
  1685 => x"1757758a",
  1686 => x"2e84bd38",
  1687 => x"84150870",
  1688 => x"822a8106",
  1689 => x"555b7380",
  1690 => x"2ef23875",
  1691 => x"750c7633",
  1692 => x"5675e038",
  1693 => x"78793355",
  1694 => x"5a73802e",
  1695 => x"80cc3880",
  1696 => x"e2b00874",
  1697 => x"575b811a",
  1698 => x"80e9e833",
  1699 => x"7081ff06",
  1700 => x"70101011",
  1701 => x"80e9ec33",
  1702 => x"7081ff06",
  1703 => x"72902911",
  1704 => x"70882b7d",
  1705 => x"07620c5a",
  1706 => x"5c5c4057",
  1707 => x"5a5a758a",
  1708 => x"2e86f938",
  1709 => x"7680cf2e",
  1710 => x"86f23881",
  1711 => x"18567580",
  1712 => x"e9ec3479",
  1713 => x"335675ff",
  1714 => x"bd3880e2",
  1715 => x"a4089411",
  1716 => x"0880dbf4",
  1717 => x"535859d7",
  1718 => x"b23f7692",
  1719 => x"3d5a568b",
  1720 => x"5380d4ac",
  1721 => x"5278519b",
  1722 => x"873f8802",
  1723 => x"840580c1",
  1724 => x"05595775",
  1725 => x"8f065473",
  1726 => x"892685ee",
  1727 => x"387618b0",
  1728 => x"15555573",
  1729 => x"75347584",
  1730 => x"2aff1870",
  1731 => x"81ff0659",
  1732 => x"5b5676df",
  1733 => x"38787933",
  1734 => x"55577380",
  1735 => x"2ea93880",
  1736 => x"e2b80874",
  1737 => x"57558117",
  1738 => x"57758a2e",
  1739 => x"838f3884",
  1740 => x"15087082",
  1741 => x"2a810655",
  1742 => x"5a73802e",
  1743 => x"f2387575",
  1744 => x"0c763356",
  1745 => x"75e03878",
  1746 => x"7933555a",
  1747 => x"73802e80",
  1748 => x"cc3880e2",
  1749 => x"b0087457",
  1750 => x"5b811a80",
  1751 => x"e9e83370",
  1752 => x"81ff0670",
  1753 => x"10101180",
  1754 => x"e9ec3370",
  1755 => x"81ff0672",
  1756 => x"90291170",
  1757 => x"882b7d07",
  1758 => x"620c5a5c",
  1759 => x"5c40575a",
  1760 => x"5a758a2e",
  1761 => x"869e3876",
  1762 => x"80cf2e86",
  1763 => x"97388118",
  1764 => x"567580e9",
  1765 => x"ec347933",
  1766 => x"5675ffbd",
  1767 => x"3880e2a4",
  1768 => x"08981108",
  1769 => x"80dc8853",
  1770 => x"5859d5df",
  1771 => x"3f768f3d",
  1772 => x"5a568b53",
  1773 => x"80d4ac52",
  1774 => x"785199b4",
  1775 => x"3f880284",
  1776 => x"05b50559",
  1777 => x"57758f06",
  1778 => x"54738926",
  1779 => x"84933876",
  1780 => x"18b01555",
  1781 => x"55737534",
  1782 => x"75842aff",
  1783 => x"187081ff",
  1784 => x"06595c56",
  1785 => x"76df3878",
  1786 => x"79335557",
  1787 => x"73802ea9",
  1788 => x"3880e2b8",
  1789 => x"08745755",
  1790 => x"81175775",
  1791 => x"8a2e81e2",
  1792 => x"38841508",
  1793 => x"70822a81",
  1794 => x"06555b73",
  1795 => x"802ef238",
  1796 => x"75750c76",
  1797 => x"335675e0",
  1798 => x"38787933",
  1799 => x"555a7380",
  1800 => x"2e80cc38",
  1801 => x"80e2b008",
  1802 => x"74575b81",
  1803 => x"1a80e9e8",
  1804 => x"337081ff",
  1805 => x"06701010",
  1806 => x"1180e9ec",
  1807 => x"337081ff",
  1808 => x"06729029",
  1809 => x"1170882b",
  1810 => x"7d07620c",
  1811 => x"5a5c5c40",
  1812 => x"575a5a75",
  1813 => x"8a2e84ae",
  1814 => x"387680cf",
  1815 => x"2e84a738",
  1816 => x"81185675",
  1817 => x"80e9ec34",
  1818 => x"79335675",
  1819 => x"ffbd38a9",
  1820 => x"3d0d0484",
  1821 => x"15087082",
  1822 => x"2a81065c",
  1823 => x"587a802e",
  1824 => x"f2388d75",
  1825 => x"0c841508",
  1826 => x"70822a81",
  1827 => x"065d5d7b",
  1828 => x"802ef9f5",
  1829 => x"38fa8139",
  1830 => x"84150870",
  1831 => x"822a8106",
  1832 => x"5b5c7980",
  1833 => x"2ef2388d",
  1834 => x"750c8415",
  1835 => x"0870822a",
  1836 => x"8106555b",
  1837 => x"73802efb",
  1838 => x"a338fbaf",
  1839 => x"39841508",
  1840 => x"70822a81",
  1841 => x"06595c77",
  1842 => x"802ef238",
  1843 => x"8d750c84",
  1844 => x"15087082",
  1845 => x"2a810655",
  1846 => x"5a73802e",
  1847 => x"fcd138fc",
  1848 => x"dd398415",
  1849 => x"0870822a",
  1850 => x"8106595c",
  1851 => x"77802ef2",
  1852 => x"388d750c",
  1853 => x"84150870",
  1854 => x"822a8106",
  1855 => x"555b7380",
  1856 => x"2efdfe38",
  1857 => x"fe8a3980",
  1858 => x"dc9c51d2",
  1859 => x"fe3ff797",
  1860 => x"3980dca0",
  1861 => x"51d2f43f",
  1862 => x"80dad051",
  1863 => x"d2ed3f80",
  1864 => x"dad451d2",
  1865 => x"e63f7485",
  1866 => x"2a870654",
  1867 => x"73812e09",
  1868 => x"8106f6e1",
  1869 => x"3880dca4",
  1870 => x"51d2d03f",
  1871 => x"f6e93980",
  1872 => x"dcac51d2",
  1873 => x"c63f80d8",
  1874 => x"f051d2bf",
  1875 => x"3f7c527b",
  1876 => x"972a8706",
  1877 => x"83058171",
  1878 => x"2b525ad1",
  1879 => x"8f3f7c51",
  1880 => x"d2a93f80",
  1881 => x"d98451d2",
  1882 => x"a23f80d9",
  1883 => x"8c51d29b",
  1884 => x"3f7c527b",
  1885 => x"9a2a8106",
  1886 => x"810551d0",
  1887 => x"ef3f7c51",
  1888 => x"d2893f80",
  1889 => x"d9a051d2",
  1890 => x"823f7c52",
  1891 => x"7b9b2a87",
  1892 => x"06830551",
  1893 => x"d0d63f7c",
  1894 => x"51d1f03f",
  1895 => x"80d9b451",
  1896 => x"d1e93f7c",
  1897 => x"527b9e2a",
  1898 => x"820751d0",
  1899 => x"bf3f7c51",
  1900 => x"d1d93f80",
  1901 => x"d9c851d1",
  1902 => x"d23f7b9f",
  1903 => x"2a9e3d5a",
  1904 => x"568b5380",
  1905 => x"d4ac5278",
  1906 => x"5195a53f",
  1907 => x"82028405",
  1908 => x"80f10559",
  1909 => x"57efa139",
  1910 => x"7618b715",
  1911 => x"5555efa8",
  1912 => x"397618b7",
  1913 => x"155555fb",
  1914 => x"ec397618",
  1915 => x"b7155555",
  1916 => x"fa913976",
  1917 => x"18b71555",
  1918 => x"55f8b539",
  1919 => x"7618b715",
  1920 => x"5555f6d9",
  1921 => x"397618b7",
  1922 => x"155555f1",
  1923 => x"853974a3",
  1924 => x"2682a538",
  1925 => x"81195675",
  1926 => x"80e9e834",
  1927 => x"800b80e9",
  1928 => x"ec347933",
  1929 => x"5675f1c0",
  1930 => x"38f28139",
  1931 => x"74a32681",
  1932 => x"f8388119",
  1933 => x"557480e9",
  1934 => x"e834800b",
  1935 => x"80e9ec34",
  1936 => x"79335675",
  1937 => x"f8c038f9",
  1938 => x"813974a3",
  1939 => x"2681cb38",
  1940 => x"81195574",
  1941 => x"80e9e834",
  1942 => x"800b80e9",
  1943 => x"ec347933",
  1944 => x"5675f6cf",
  1945 => x"38f79039",
  1946 => x"74a32681",
  1947 => x"9e388119",
  1948 => x"567580e9",
  1949 => x"e834800b",
  1950 => x"80e9ec34",
  1951 => x"79335675",
  1952 => x"ebfe38ec",
  1953 => x"bf3974a3",
  1954 => x"2680f138",
  1955 => x"81195574",
  1956 => x"80e9e834",
  1957 => x"800b80e9",
  1958 => x"ec347933",
  1959 => x"5675fb8b",
  1960 => x"38fbcc39",
  1961 => x"74a32680",
  1962 => x"c4388119",
  1963 => x"557480e9",
  1964 => x"e834800b",
  1965 => x"80e9ec34",
  1966 => x"79335675",
  1967 => x"f99b38f9",
  1968 => x"dc3974a3",
  1969 => x"26993881",
  1970 => x"19567580",
  1971 => x"e9e83480",
  1972 => x"0b80e9ec",
  1973 => x"34793356",
  1974 => x"75ee8338",
  1975 => x"eec43980",
  1976 => x"0b80e9e8",
  1977 => x"34800b80",
  1978 => x"e9ec34e9",
  1979 => x"39800b80",
  1980 => x"e9e83480",
  1981 => x"0b80e9ec",
  1982 => x"34ffbd39",
  1983 => x"800b80e9",
  1984 => x"e834800b",
  1985 => x"80e9ec34",
  1986 => x"ff903980",
  1987 => x"0b80e9e8",
  1988 => x"34800b80",
  1989 => x"e9ec34fe",
  1990 => x"e339800b",
  1991 => x"80e9e834",
  1992 => x"800b80e9",
  1993 => x"ec34feb6",
  1994 => x"39800b80",
  1995 => x"e9e83480",
  1996 => x"0b80e9ec",
  1997 => x"34fe8939",
  1998 => x"800b80e9",
  1999 => x"e834800b",
  2000 => x"80e9ec34",
  2001 => x"fddc3980",
  2002 => x"dcb451ce",
  2003 => x"be3ff2d7",
  2004 => x"3980dcbc",
  2005 => x"51ceb43f",
  2006 => x"fbbe3980",
  2007 => x"dcc051ce",
  2008 => x"aa3ffbe2",
  2009 => x"3980dcc8",
  2010 => x"51cea03f",
  2011 => x"fbaa3980",
  2012 => x"dccc51ce",
  2013 => x"963ffbce",
  2014 => x"3980dcd4",
  2015 => x"51ce8c3f",
  2016 => x"fb963980",
  2017 => x"dcd851ce",
  2018 => x"823ff29b",
  2019 => x"3980dcdc",
  2020 => x"51cdf83f",
  2021 => x"fbb03980",
  2022 => x"dce451f1",
  2023 => x"af3980dc",
  2024 => x"d851f1a8",
  2025 => x"3980dce8",
  2026 => x"51f1a139",
  2027 => x"80dcec51",
  2028 => x"f19a3980",
  2029 => x"dcf051cd",
  2030 => x"d23f80da",
  2031 => x"fc51cdcb",
  2032 => x"3f7c5274",
  2033 => x"932a8306",
  2034 => x"820751cc",
  2035 => x"9f3f7c51",
  2036 => x"cdb93f80",
  2037 => x"db9051cd",
  2038 => x"b23f7c52",
  2039 => x"74942a8f",
  2040 => x"0651cc88",
  2041 => x"3f7c51cd",
  2042 => x"a23f80db",
  2043 => x"a451cd9b",
  2044 => x"3f7c5274",
  2045 => x"982a8106",
  2046 => x"810551cb",
  2047 => x"ef3f7c51",
  2048 => x"cd893f80",
  2049 => x"dbb851cd",
  2050 => x"823f7c52",
  2051 => x"749e2a82",
  2052 => x"0751cbd8",
  2053 => x"3f7c51cc",
  2054 => x"f23f80db",
  2055 => x"cc51cceb",
  2056 => x"3f749f2a",
  2057 => x"983d5a56",
  2058 => x"8b5380d4",
  2059 => x"ac527851",
  2060 => x"90be3f82",
  2061 => x"02840580",
  2062 => x"d9055957",
  2063 => x"f28f3980",
  2064 => x"dd8051cc",
  2065 => x"c63f80da",
  2066 => x"fc51ccbf",
  2067 => x"3f7c5274",
  2068 => x"932a8306",
  2069 => x"820751cb",
  2070 => x"933f7c51",
  2071 => x"ccad3f80",
  2072 => x"db9051cc",
  2073 => x"a63f7c52",
  2074 => x"74942a8f",
  2075 => x"0651cafc",
  2076 => x"3f7c51cc",
  2077 => x"963f80db",
  2078 => x"a451cc8f",
  2079 => x"3f7c5274",
  2080 => x"982a8106",
  2081 => x"810551ca",
  2082 => x"e33f7c51",
  2083 => x"cbfd3f80",
  2084 => x"dbb851cb",
  2085 => x"f63f7c52",
  2086 => x"749e2a82",
  2087 => x"0751cacc",
  2088 => x"3f7c51cb",
  2089 => x"e63f80db",
  2090 => x"cc51cbdf",
  2091 => x"3f749f2a",
  2092 => x"983d5a56",
  2093 => x"8b5380d4",
  2094 => x"ac527851",
  2095 => x"8fb23f82",
  2096 => x"02840580",
  2097 => x"d9055957",
  2098 => x"f1833980",
  2099 => x"dd8c51cb",
  2100 => x"ba3f80da",
  2101 => x"fc51cbb3",
  2102 => x"3f7c5274",
  2103 => x"932a8306",
  2104 => x"820751ca",
  2105 => x"873f7c51",
  2106 => x"cba13f80",
  2107 => x"db9051cb",
  2108 => x"9a3f7c52",
  2109 => x"74942a8f",
  2110 => x"0651c9f0",
  2111 => x"3f7c51cb",
  2112 => x"8a3f80db",
  2113 => x"a451cb83",
  2114 => x"3f7c5274",
  2115 => x"982a8106",
  2116 => x"810551c9",
  2117 => x"d73f7c51",
  2118 => x"caf13f80",
  2119 => x"dbb851ca",
  2120 => x"ea3f7c52",
  2121 => x"749e2a82",
  2122 => x"0751c9c0",
  2123 => x"3f7c51ca",
  2124 => x"da3f80db",
  2125 => x"cc51cad3",
  2126 => x"3f749f2a",
  2127 => x"983d5a56",
  2128 => x"8b5380d4",
  2129 => x"ac527851",
  2130 => x"8ea63f82",
  2131 => x"02840580",
  2132 => x"d9055957",
  2133 => x"eff73980",
  2134 => x"dd9c51ca",
  2135 => x"ae3f80da",
  2136 => x"fc51caa7",
  2137 => x"3f7c5274",
  2138 => x"932a8306",
  2139 => x"820751c8",
  2140 => x"fb3f7c51",
  2141 => x"ca953f80",
  2142 => x"db9051ca",
  2143 => x"8e3f7c52",
  2144 => x"74942a8f",
  2145 => x"0651c8e4",
  2146 => x"3f7c51c9",
  2147 => x"fe3f80db",
  2148 => x"a451c9f7",
  2149 => x"3f7c5274",
  2150 => x"982a8106",
  2151 => x"810551c8",
  2152 => x"cb3f7c51",
  2153 => x"c9e53f80",
  2154 => x"dbb851c9",
  2155 => x"de3f7c52",
  2156 => x"749e2a82",
  2157 => x"0751c8b4",
  2158 => x"3f7c51c9",
  2159 => x"ce3f80db",
  2160 => x"cc51c9c7",
  2161 => x"3f749f2a",
  2162 => x"983d5a56",
  2163 => x"8b5380d4",
  2164 => x"ac527851",
  2165 => x"8d9a3f82",
  2166 => x"02840580",
  2167 => x"d9055957",
  2168 => x"eeeb3980",
  2169 => x"dda851c9",
  2170 => x"a23f80da",
  2171 => x"fc51c99b",
  2172 => x"3f7c5274",
  2173 => x"932a8306",
  2174 => x"820751c7",
  2175 => x"ef3f7c51",
  2176 => x"c9893f80",
  2177 => x"db9051c9",
  2178 => x"823f7c52",
  2179 => x"74942a8f",
  2180 => x"0651c7d8",
  2181 => x"3f7c51c8",
  2182 => x"f23f80db",
  2183 => x"a451c8eb",
  2184 => x"3f7c5274",
  2185 => x"982a8106",
  2186 => x"810551c7",
  2187 => x"bf3f7c51",
  2188 => x"c8d93f80",
  2189 => x"dbb851c8",
  2190 => x"d23f7c52",
  2191 => x"749e2a82",
  2192 => x"0751c7a8",
  2193 => x"3f7c51c8",
  2194 => x"c23f80db",
  2195 => x"cc51c8bb",
  2196 => x"3f749f2a",
  2197 => x"983d5a56",
  2198 => x"8b5380d4",
  2199 => x"ac527851",
  2200 => x"8c8e3f82",
  2201 => x"02840580",
  2202 => x"d9055957",
  2203 => x"eddf39ea",
  2204 => x"3d0d80e2",
  2205 => x"a4088411",
  2206 => x"08709fff",
  2207 => x"06515454",
  2208 => x"8a54bb73",
  2209 => x"2783388f",
  2210 => x"54725287",
  2211 => x"e851879a",
  2212 => x"3f8008fd",
  2213 => x"05742970",
  2214 => x"83ffff06",
  2215 => x"5a558070",
  2216 => x"80e2a808",
  2217 => x"7b30575a",
  2218 => x"5d5d8c18",
  2219 => x"08567376",
  2220 => x"24963880",
  2221 => x"0b84190c",
  2222 => x"77085776",
  2223 => x"ed387708",
  2224 => x"5776802e",
  2225 => x"f338e339",
  2226 => x"7b307c07",
  2227 => x"7080257e",
  2228 => x"81320754",
  2229 => x"5472802e",
  2230 => x"80fb388c",
  2231 => x"18085574",
  2232 => x"792480f1",
  2233 => x"38805789",
  2234 => x"0a558fff",
  2235 => x"56740875",
  2236 => x"32703070",
  2237 => x"7207709f",
  2238 => x"2a7a0584",
  2239 => x"19ff1b5b",
  2240 => x"595a5154",
  2241 => x"54758025",
  2242 => x"e4387683",
  2243 => x"ffff067c",
  2244 => x"81325454",
  2245 => x"73923881",
  2246 => x"70740657",
  2247 => x"5575802e",
  2248 => x"8738748c",
  2249 => x"19085b5c",
  2250 => x"73802e92",
  2251 => x"3881707d",
  2252 => x"06565474",
  2253 => x"802e8738",
  2254 => x"738c1908",
  2255 => x"5c5d800b",
  2256 => x"88190c77",
  2257 => x"085776fe",
  2258 => x"ff387708",
  2259 => x"5776802e",
  2260 => x"f238fef4",
  2261 => x"39739f2a",
  2262 => x"537c802e",
  2263 => x"82893872",
  2264 => x"802e8283",
  2265 => x"387a7a31",
  2266 => x"709f2a11",
  2267 => x"70812c7d",
  2268 => x"71318c1c",
  2269 => x"08707231",
  2270 => x"525b525b",
  2271 => x"55568074",
  2272 => x"259938ff",
  2273 => x"1454800b",
  2274 => x"84190c77",
  2275 => x"085372ee",
  2276 => x"38770853",
  2277 => x"72802ef3",
  2278 => x"38e43980",
  2279 => x"0b80e2b0",
  2280 => x"08565473",
  2281 => x"882b750c",
  2282 => x"81145497",
  2283 => x"907426f3",
  2284 => x"38800b80",
  2285 => x"e9e83480",
  2286 => x"0b80e9ec",
  2287 => x"3480d7cc",
  2288 => x"51c5c83f",
  2289 => x"7b802e81",
  2290 => x"af3880dd",
  2291 => x"f851c5bb",
  2292 => x"3f80d7cc",
  2293 => x"51c5b43f",
  2294 => x"7c802e81",
  2295 => x"a23880de",
  2296 => x"8451c5a7",
  2297 => x"3f80de90",
  2298 => x"51c5a03f",
  2299 => x"933d7053",
  2300 => x"7a525cc3",
  2301 => x"f73f7b51",
  2302 => x"c5913f80",
  2303 => x"dea051c5",
  2304 => x"8a3f7b52",
  2305 => x"7a51c3e4",
  2306 => x"3f7b51c4",
  2307 => x"fe3f80d7",
  2308 => x"cc51c4f7",
  2309 => x"3f80deb0",
  2310 => x"51c4f03f",
  2311 => x"7b527551",
  2312 => x"c3ca3f7b",
  2313 => x"51c4e43f",
  2314 => x"80dec051",
  2315 => x"c4dd3f7b",
  2316 => x"52759f2a",
  2317 => x"1670812c",
  2318 => x"525bc3b0",
  2319 => x"3f7b51c4",
  2320 => x"ca3f80d7",
  2321 => x"cc51c4c3",
  2322 => x"3f80df80",
  2323 => x"51c4bc3f",
  2324 => x"7b5280e2",
  2325 => x"a8088c11",
  2326 => x"08525ac3",
  2327 => x"8f3f7b51",
  2328 => x"c4a93f98",
  2329 => x"3d0d048b",
  2330 => x"7b7b318c",
  2331 => x"1a087073",
  2332 => x"31535957",
  2333 => x"54fe8739",
  2334 => x"80dfa851",
  2335 => x"fed03980",
  2336 => x"df9851fe",
  2337 => x"dd39f73d",
  2338 => x"0d800b80",
  2339 => x"e2ac0870",
  2340 => x"08810a06",
  2341 => x"80e9e40c",
  2342 => x"5555c2bf",
  2343 => x"3f80e2b8",
  2344 => x"0852b60b",
  2345 => x"8c130c83",
  2346 => x"0b88130c",
  2347 => x"80e2a408",
  2348 => x"54fac98e",
  2349 => x"868b740c",
  2350 => x"73087084",
  2351 => x"2a810651",
  2352 => x"5372f538",
  2353 => x"80e2b008",
  2354 => x"7384120c",
  2355 => x"54fe800a",
  2356 => x"0b88150c",
  2357 => x"7280e9e8",
  2358 => x"347280e9",
  2359 => x"ec3480df",
  2360 => x"b851c3a7",
  2361 => x"3f80e9e4",
  2362 => x"08802e82",
  2363 => x"b63880df",
  2364 => x"c051c397",
  2365 => x"3f80dfd0",
  2366 => x"51c3903f",
  2367 => x"890a5283",
  2368 => x"ffff5371",
  2369 => x"720c8412",
  2370 => x"ff145452",
  2371 => x"728025f3",
  2372 => x"3880d79c",
  2373 => x"51c2f43f",
  2374 => x"800b80e2",
  2375 => x"b0085553",
  2376 => x"72882b74",
  2377 => x"0c811353",
  2378 => x"97907326",
  2379 => x"f338800b",
  2380 => x"80e9e834",
  2381 => x"800b80e9",
  2382 => x"ec34dbc0",
  2383 => x"3f8551ff",
  2384 => x"bff03ffa",
  2385 => x"aa3f8a51",
  2386 => x"ffbfe73f",
  2387 => x"800b80e2",
  2388 => x"b0085553",
  2389 => x"72882b74",
  2390 => x"0c811353",
  2391 => x"97907326",
  2392 => x"f338800b",
  2393 => x"80e9e834",
  2394 => x"800b80e9",
  2395 => x"ec347451",
  2396 => x"c5f13f80",
  2397 => x"e2ac0870",
  2398 => x"0870872a",
  2399 => x"81065155",
  2400 => x"5373802e",
  2401 => x"8b3880e2",
  2402 => x"a8085280",
  2403 => x"0b84130c",
  2404 => x"72087084",
  2405 => x"2a810651",
  2406 => x"5473802e",
  2407 => x"8b3880e2",
  2408 => x"a8085280",
  2409 => x"0b88130c",
  2410 => x"72087085",
  2411 => x"2a810651",
  2412 => x"5473802e",
  2413 => x"b63880e2",
  2414 => x"a40853fa",
  2415 => x"c98e868b",
  2416 => x"730c7208",
  2417 => x"70842a81",
  2418 => x"06515271",
  2419 => x"f538f99f",
  2420 => x"3f890a52",
  2421 => x"83ffff53",
  2422 => x"71720c84",
  2423 => x"12ff1454",
  2424 => x"52728025",
  2425 => x"f33880e2",
  2426 => x"ac085372",
  2427 => x"0870862a",
  2428 => x"81065452",
  2429 => x"72802efe",
  2430 => x"f538800b",
  2431 => x"80e2b008",
  2432 => x"55537288",
  2433 => x"2b740c81",
  2434 => x"13539790",
  2435 => x"7326f338",
  2436 => x"800b80e9",
  2437 => x"e834800b",
  2438 => x"80e9ec34",
  2439 => x"74813255",
  2440 => x"fecc3980",
  2441 => x"dff451fd",
  2442 => x"c9398c08",
  2443 => x"028c0cfd",
  2444 => x"3d0d8053",
  2445 => x"8c088c05",
  2446 => x"08528c08",
  2447 => x"88050851",
  2448 => x"82de3f80",
  2449 => x"0870800c",
  2450 => x"54853d0d",
  2451 => x"8c0c048c",
  2452 => x"08028c0c",
  2453 => x"fd3d0d81",
  2454 => x"538c088c",
  2455 => x"0508528c",
  2456 => x"08880508",
  2457 => x"5182b93f",
  2458 => x"80087080",
  2459 => x"0c54853d",
  2460 => x"0d8c0c04",
  2461 => x"8c08028c",
  2462 => x"0cf93d0d",
  2463 => x"800b8c08",
  2464 => x"fc050c8c",
  2465 => x"08880508",
  2466 => x"8025ab38",
  2467 => x"8c088805",
  2468 => x"08308c08",
  2469 => x"88050c80",
  2470 => x"0b8c08f4",
  2471 => x"050c8c08",
  2472 => x"fc050888",
  2473 => x"38810b8c",
  2474 => x"08f4050c",
  2475 => x"8c08f405",
  2476 => x"088c08fc",
  2477 => x"050c8c08",
  2478 => x"8c050880",
  2479 => x"25ab388c",
  2480 => x"088c0508",
  2481 => x"308c088c",
  2482 => x"050c800b",
  2483 => x"8c08f005",
  2484 => x"0c8c08fc",
  2485 => x"05088838",
  2486 => x"810b8c08",
  2487 => x"f0050c8c",
  2488 => x"08f00508",
  2489 => x"8c08fc05",
  2490 => x"0c80538c",
  2491 => x"088c0508",
  2492 => x"528c0888",
  2493 => x"05085181",
  2494 => x"a73f8008",
  2495 => x"708c08f8",
  2496 => x"050c548c",
  2497 => x"08fc0508",
  2498 => x"802e8c38",
  2499 => x"8c08f805",
  2500 => x"08308c08",
  2501 => x"f8050c8c",
  2502 => x"08f80508",
  2503 => x"70800c54",
  2504 => x"893d0d8c",
  2505 => x"0c048c08",
  2506 => x"028c0cfb",
  2507 => x"3d0d800b",
  2508 => x"8c08fc05",
  2509 => x"0c8c0888",
  2510 => x"05088025",
  2511 => x"93388c08",
  2512 => x"88050830",
  2513 => x"8c088805",
  2514 => x"0c810b8c",
  2515 => x"08fc050c",
  2516 => x"8c088c05",
  2517 => x"0880258c",
  2518 => x"388c088c",
  2519 => x"0508308c",
  2520 => x"088c050c",
  2521 => x"81538c08",
  2522 => x"8c050852",
  2523 => x"8c088805",
  2524 => x"0851ad3f",
  2525 => x"8008708c",
  2526 => x"08f8050c",
  2527 => x"548c08fc",
  2528 => x"0508802e",
  2529 => x"8c388c08",
  2530 => x"f8050830",
  2531 => x"8c08f805",
  2532 => x"0c8c08f8",
  2533 => x"05087080",
  2534 => x"0c54873d",
  2535 => x"0d8c0c04",
  2536 => x"8c08028c",
  2537 => x"0cfd3d0d",
  2538 => x"810b8c08",
  2539 => x"fc050c80",
  2540 => x"0b8c08f8",
  2541 => x"050c8c08",
  2542 => x"8c05088c",
  2543 => x"08880508",
  2544 => x"27ac388c",
  2545 => x"08fc0508",
  2546 => x"802ea338",
  2547 => x"800b8c08",
  2548 => x"8c050824",
  2549 => x"99388c08",
  2550 => x"8c050810",
  2551 => x"8c088c05",
  2552 => x"0c8c08fc",
  2553 => x"0508108c",
  2554 => x"08fc050c",
  2555 => x"c9398c08",
  2556 => x"fc050880",
  2557 => x"2e80c938",
  2558 => x"8c088c05",
  2559 => x"088c0888",
  2560 => x"050826a1",
  2561 => x"388c0888",
  2562 => x"05088c08",
  2563 => x"8c050831",
  2564 => x"8c088805",
  2565 => x"0c8c08f8",
  2566 => x"05088c08",
  2567 => x"fc050807",
  2568 => x"8c08f805",
  2569 => x"0c8c08fc",
  2570 => x"0508812a",
  2571 => x"8c08fc05",
  2572 => x"0c8c088c",
  2573 => x"0508812a",
  2574 => x"8c088c05",
  2575 => x"0cffaf39",
  2576 => x"8c089005",
  2577 => x"08802e8f",
  2578 => x"388c0888",
  2579 => x"0508708c",
  2580 => x"08f4050c",
  2581 => x"518d398c",
  2582 => x"08f80508",
  2583 => x"708c08f4",
  2584 => x"050c518c",
  2585 => x"08f40508",
  2586 => x"800c853d",
  2587 => x"0d8c0c04",
  2588 => x"fc3d0d76",
  2589 => x"70797b55",
  2590 => x"5555558f",
  2591 => x"72278c38",
  2592 => x"72750783",
  2593 => x"06517080",
  2594 => x"2ea738ff",
  2595 => x"125271ff",
  2596 => x"2e983872",
  2597 => x"70810554",
  2598 => x"33747081",
  2599 => x"055634ff",
  2600 => x"125271ff",
  2601 => x"2e098106",
  2602 => x"ea387480",
  2603 => x"0c863d0d",
  2604 => x"04745172",
  2605 => x"70840554",
  2606 => x"08717084",
  2607 => x"05530c72",
  2608 => x"70840554",
  2609 => x"08717084",
  2610 => x"05530c72",
  2611 => x"70840554",
  2612 => x"08717084",
  2613 => x"05530c72",
  2614 => x"70840554",
  2615 => x"08717084",
  2616 => x"05530cf0",
  2617 => x"1252718f",
  2618 => x"26c93883",
  2619 => x"72279538",
  2620 => x"72708405",
  2621 => x"54087170",
  2622 => x"8405530c",
  2623 => x"fc125271",
  2624 => x"8326ed38",
  2625 => x"7054ff83",
  2626 => x"39fd3d0d",
  2627 => x"800b80e2",
  2628 => x"98085454",
  2629 => x"72812e9c",
  2630 => x"387380e9",
  2631 => x"f00cffb6",
  2632 => x"bf3fffb5",
  2633 => x"db3f80e2",
  2634 => x"bc528151",
  2635 => x"f6d83f80",
  2636 => x"0851a23f",
  2637 => x"7280e9f0",
  2638 => x"0cffb6a4",
  2639 => x"3fffb5c0",
  2640 => x"3f80e2bc",
  2641 => x"528151f6",
  2642 => x"bd3f8008",
  2643 => x"51873f00",
  2644 => x"ff3900ff",
  2645 => x"39f73d0d",
  2646 => x"7b80e2c0",
  2647 => x"0882c811",
  2648 => x"085a545a",
  2649 => x"77802e80",
  2650 => x"da388188",
  2651 => x"18841908",
  2652 => x"ff058171",
  2653 => x"2b595559",
  2654 => x"80742480",
  2655 => x"ea388074",
  2656 => x"24b53873",
  2657 => x"822b7811",
  2658 => x"88055656",
  2659 => x"81801908",
  2660 => x"77065372",
  2661 => x"802eb638",
  2662 => x"78167008",
  2663 => x"53537951",
  2664 => x"74085372",
  2665 => x"2dff14fc",
  2666 => x"17fc1779",
  2667 => x"812c5a57",
  2668 => x"57547380",
  2669 => x"25d63877",
  2670 => x"085877ff",
  2671 => x"ad3880e2",
  2672 => x"c00853bc",
  2673 => x"1308a538",
  2674 => x"7951ff83",
  2675 => x"3f740853",
  2676 => x"722dff14",
  2677 => x"fc17fc17",
  2678 => x"79812c5a",
  2679 => x"57575473",
  2680 => x"8025ffa8",
  2681 => x"38d13980",
  2682 => x"57ff9339",
  2683 => x"7251bc13",
  2684 => x"0853722d",
  2685 => x"7951fed7",
  2686 => x"3fff3d0d",
  2687 => x"80e9c40b",
  2688 => x"fc057008",
  2689 => x"525270ff",
  2690 => x"2e913870",
  2691 => x"2dfc1270",
  2692 => x"08525270",
  2693 => x"ff2e0981",
  2694 => x"06f13883",
  2695 => x"3d0d0404",
  2696 => x"ffb5aa3f",
  2697 => x"04000000",
  2698 => x"00000040",
  2699 => x"30782020",
  2700 => x"20202020",
  2701 => x"20200000",
  2702 => x"30622020",
  2703 => x"20202020",
  2704 => x"20202020",
  2705 => x"20202020",
  2706 => x"20202020",
  2707 => x"20202020",
  2708 => x"20202020",
  2709 => x"20202020",
  2710 => x"20200000",
  2711 => x"0a677265",
  2712 => x"74682072",
  2713 => x"65676973",
  2714 => x"74657273",
  2715 => x"3a000000",
  2716 => x"0a636f6e",
  2717 => x"74726f6c",
  2718 => x"3a202020",
  2719 => x"20202000",
  2720 => x"0a737461",
  2721 => x"7475733a",
  2722 => x"20202020",
  2723 => x"20202000",
  2724 => x"0a6d6163",
  2725 => x"5f6d7362",
  2726 => x"3a202020",
  2727 => x"20202000",
  2728 => x"0a6d6163",
  2729 => x"5f6c7362",
  2730 => x"3a202020",
  2731 => x"20202000",
  2732 => x"0a6d6469",
  2733 => x"6f5f636f",
  2734 => x"6e74726f",
  2735 => x"6c3a2000",
  2736 => x"0a74785f",
  2737 => x"706f696e",
  2738 => x"7465723a",
  2739 => x"20202000",
  2740 => x"0a72785f",
  2741 => x"706f696e",
  2742 => x"7465723a",
  2743 => x"20202000",
  2744 => x"0a656463",
  2745 => x"6c5f6970",
  2746 => x"3a202020",
  2747 => x"20202000",
  2748 => x"0a686173",
  2749 => x"685f6d73",
  2750 => x"623a2020",
  2751 => x"20202000",
  2752 => x"0a686173",
  2753 => x"685f6c73",
  2754 => x"623a2020",
  2755 => x"20202000",
  2756 => x"0a6d6469",
  2757 => x"6f207068",
  2758 => x"79207265",
  2759 => x"67697374",
  2760 => x"65727300",
  2761 => x"0a206d64",
  2762 => x"696f2070",
  2763 => x"68793a20",
  2764 => x"00000000",
  2765 => x"0a202072",
  2766 => x"65673a20",
  2767 => x"00000000",
  2768 => x"2d3e2000",
  2769 => x"0a677265",
  2770 => x"74682d3e",
  2771 => x"636f6e74",
  2772 => x"726f6c20",
  2773 => x"3a000000",
  2774 => x"0a677265",
  2775 => x"74682d3e",
  2776 => x"73746174",
  2777 => x"75732020",
  2778 => x"3a000000",
  2779 => x"0a646573",
  2780 => x"63722d3e",
  2781 => x"636f6e74",
  2782 => x"726f6c20",
  2783 => x"3a000000",
  2784 => x"77726974",
  2785 => x"65206164",
  2786 => x"64726573",
  2787 => x"733a2000",
  2788 => x"20206c65",
  2789 => x"6e677468",
  2790 => x"3a200000",
  2791 => x"0a0a0000",
  2792 => x"72656164",
  2793 => x"20206164",
  2794 => x"64726573",
  2795 => x"733a2000",
  2796 => x"20206578",
  2797 => x"70656374",
  2798 => x"3a200000",
  2799 => x"2020676f",
  2800 => x"743a2000",
  2801 => x"20657272",
  2802 => x"6f720000",
  2803 => x"0a000000",
  2804 => x"206f6b00",
  2805 => x"70686173",
  2806 => x"65207368",
  2807 => x"69667420",
  2808 => x"202d2020",
  2809 => x"76616c75",
  2810 => x"653a2000",
  2811 => x"20207374",
  2812 => x"61747573",
  2813 => x"3a200000",
  2814 => x"20202020",
  2815 => x"20000000",
  2816 => x"4641494c",
  2817 => x"00000000",
  2818 => x"6f6b2020",
  2819 => x"00000000",
  2820 => x"44445220",
  2821 => x"6d656d6f",
  2822 => x"72792069",
  2823 => x"6e666f00",
  2824 => x"0a0a6175",
  2825 => x"746f2074",
  2826 => x"5f524552",
  2827 => x"45534820",
  2828 => x"3a000000",
  2829 => x"0a636c6f",
  2830 => x"636b2065",
  2831 => x"6e61626c",
  2832 => x"6520203a",
  2833 => x"00000000",
  2834 => x"0a696e69",
  2835 => x"74616c69",
  2836 => x"7a652020",
  2837 => x"2020203a",
  2838 => x"00000000",
  2839 => x"0a636f6c",
  2840 => x"756d6e20",
  2841 => x"73697a65",
  2842 => x"2020203a",
  2843 => x"00000000",
  2844 => x"0a62616e",
  2845 => x"6b73697a",
  2846 => x"65202020",
  2847 => x"2020203a",
  2848 => x"00000000",
  2849 => x"4d627974",
  2850 => x"65000000",
  2851 => x"0a745f52",
  2852 => x"43442020",
  2853 => x"20202020",
  2854 => x"2020203a",
  2855 => x"00000000",
  2856 => x"0a745f52",
  2857 => x"46432020",
  2858 => x"20202020",
  2859 => x"2020203a",
  2860 => x"00000000",
  2861 => x"0a745f52",
  2862 => x"50202020",
  2863 => x"20202020",
  2864 => x"2020203a",
  2865 => x"00000000",
  2866 => x"0a726566",
  2867 => x"72657368",
  2868 => x"20656e2e",
  2869 => x"2020203a",
  2870 => x"00000000",
  2871 => x"0a0a4444",
  2872 => x"52206672",
  2873 => x"65717565",
  2874 => x"6e637920",
  2875 => x"3a000000",
  2876 => x"0a444452",
  2877 => x"20646174",
  2878 => x"61207769",
  2879 => x"6474683a",
  2880 => x"00000000",
  2881 => x"0a6d6f62",
  2882 => x"696c6520",
  2883 => x"73757070",
  2884 => x"6f72743a",
  2885 => x"00000000",
  2886 => x"0a0a7365",
  2887 => x"6c662072",
  2888 => x"65667265",
  2889 => x"73682020",
  2890 => x"3a000000",
  2891 => x"756e6b6e",
  2892 => x"6f776e00",
  2893 => x"20617272",
  2894 => x"61790000",
  2895 => x"0a74656d",
  2896 => x"702d636f",
  2897 => x"6d702072",
  2898 => x"6566723a",
  2899 => x"00000000",
  2900 => x"c2b04300",
  2901 => x"0a647269",
  2902 => x"76652073",
  2903 => x"7472656e",
  2904 => x"6774683a",
  2905 => x"00000000",
  2906 => x"0a706f77",
  2907 => x"65722073",
  2908 => x"6176696e",
  2909 => x"6720203a",
  2910 => x"00000000",
  2911 => x"0a745f58",
  2912 => x"50202020",
  2913 => x"20202020",
  2914 => x"2020203a",
  2915 => x"00000000",
  2916 => x"0a745f58",
  2917 => x"53522020",
  2918 => x"20202020",
  2919 => x"2020203a",
  2920 => x"00000000",
  2921 => x"0a745f43",
  2922 => x"4b452020",
  2923 => x"20202020",
  2924 => x"2020203a",
  2925 => x"00000000",
  2926 => x"0a434153",
  2927 => x"206c6174",
  2928 => x"656e6379",
  2929 => x"2020203a",
  2930 => x"00000000",
  2931 => x"0a6d6f62",
  2932 => x"696c6520",
  2933 => x"656e6162",
  2934 => x"6c65643a",
  2935 => x"00000000",
  2936 => x"0a0a7374",
  2937 => x"61747573",
  2938 => x"20726561",
  2939 => x"64202020",
  2940 => x"3a000000",
  2941 => x"0a0a7068",
  2942 => x"7920636f",
  2943 => x"6e666967",
  2944 => x"20302020",
  2945 => x"3a000000",
  2946 => x"0a0a7068",
  2947 => x"7920636f",
  2948 => x"6e666967",
  2949 => x"20312020",
  2950 => x"3a000000",
  2951 => x"332f3400",
  2952 => x"38350000",
  2953 => x"68616c66",
  2954 => x"00000000",
  2955 => x"34303639",
  2956 => x"00000000",
  2957 => x"66756c6c",
  2958 => x"00000000",
  2959 => x"37300000",
  2960 => x"20353132",
  2961 => x"00000000",
  2962 => x"34350000",
  2963 => x"31303234",
  2964 => x"00000000",
  2965 => x"31350000",
  2966 => x"312f3400",
  2967 => x"32303438",
  2968 => x"00000000",
  2969 => x"312f3800",
  2970 => x"312f3200",
  2971 => x"312f3100",
  2972 => x"64656570",
  2973 => x"20706f77",
  2974 => x"65722064",
  2975 => x"6f776e00",
  2976 => x"636c6f63",
  2977 => x"6b207374",
  2978 => x"6f700000",
  2979 => x"73656c66",
  2980 => x"20726566",
  2981 => x"72657368",
  2982 => x"00000000",
  2983 => x"706f7765",
  2984 => x"7220646f",
  2985 => x"776e0000",
  2986 => x"6e6f6e65",
  2987 => x"00000000",
  2988 => x"61646472",
  2989 => x"6573733a",
  2990 => x"20000000",
  2991 => x"20646174",
  2992 => x"613a2000",
  2993 => x"0a0a4443",
  2994 => x"4d207068",
  2995 => x"61736520",
  2996 => x"73686966",
  2997 => x"74207465",
  2998 => x"7374696e",
  2999 => x"67000000",
  3000 => x"0a696e69",
  3001 => x"7469616c",
  3002 => x"3a200000",
  3003 => x"09000000",
  3004 => x"20202020",
  3005 => x"00000000",
  3006 => x"6c6f7720",
  3007 => x"666f756e",
  3008 => x"64000000",
  3009 => x"68696768",
  3010 => x"20666f75",
  3011 => x"6e640000",
  3012 => x"0a6c6f77",
  3013 => x"3a202020",
  3014 => x"20202020",
  3015 => x"20200000",
  3016 => x"0a686967",
  3017 => x"683a2020",
  3018 => x"20202020",
  3019 => x"20200000",
  3020 => x"0a646966",
  3021 => x"663a2020",
  3022 => x"20202020",
  3023 => x"20200000",
  3024 => x"0a646966",
  3025 => x"662f323a",
  3026 => x"20202020",
  3027 => x"20200000",
  3028 => x"0a6d696e",
  3029 => x"5f657272",
  3030 => x"3a202020",
  3031 => x"20200000",
  3032 => x"0a6d696e",
  3033 => x"5f657272",
  3034 => x"5f706f73",
  3035 => x"3a200000",
  3036 => x"676f206d",
  3037 => x"696e5f65",
  3038 => x"72726f72",
  3039 => x"00000000",
  3040 => x"0a66696e",
  3041 => x"616c3a20",
  3042 => x"20202020",
  3043 => x"20200000",
  3044 => x"676f207a",
  3045 => x"65726f00",
  3046 => x"68696768",
  3047 => x"204e4f54",
  3048 => x"20666f75",
  3049 => x"6e640000",
  3050 => x"6c6f7720",
  3051 => x"4e4f5420",
  3052 => x"666f756e",
  3053 => x"64000000",
  3054 => x"74657374",
  3055 => x"2e632000",
  3056 => x"286f6e20",
  3057 => x"73696d75",
  3058 => x"6c61746f",
  3059 => x"72290a00",
  3060 => x"636f6d70",
  3061 => x"696c6564",
  3062 => x"3a204f63",
  3063 => x"74203231",
  3064 => x"20323031",
  3065 => x"30202031",
  3066 => x"363a3032",
  3067 => x"3a31340a",
  3068 => x"00000000",
  3069 => x"286f6e20",
  3070 => x"68617264",
  3071 => x"77617265",
  3072 => x"290a0000",
  3073 => x"00000789",
  3074 => x"000007af",
  3075 => x"000007af",
  3076 => x"00000789",
  3077 => x"000007af",
  3078 => x"000007af",
  3079 => x"000007af",
  3080 => x"000007af",
  3081 => x"000007af",
  3082 => x"000007af",
  3083 => x"000007af",
  3084 => x"000007af",
  3085 => x"000007af",
  3086 => x"000007af",
  3087 => x"000007af",
  3088 => x"000007af",
  3089 => x"000007af",
  3090 => x"000007af",
  3091 => x"000007af",
  3092 => x"000007af",
  3093 => x"000007af",
  3094 => x"000007af",
  3095 => x"000007af",
  3096 => x"000007af",
  3097 => x"000007af",
  3098 => x"000007af",
  3099 => x"000007af",
  3100 => x"000007af",
  3101 => x"000007af",
  3102 => x"000007af",
  3103 => x"000007af",
  3104 => x"000007af",
  3105 => x"000007af",
  3106 => x"000007af",
  3107 => x"000007af",
  3108 => x"000007af",
  3109 => x"000007af",
  3110 => x"000007af",
  3111 => x"0000085b",
  3112 => x"00000853",
  3113 => x"0000084b",
  3114 => x"00000843",
  3115 => x"0000083b",
  3116 => x"00000833",
  3117 => x"0000082b",
  3118 => x"00000822",
  3119 => x"00000819",
  3120 => x"00001fac",
  3121 => x"00001fa5",
  3122 => x"00001f9e",
  3123 => x"00001848",
  3124 => x"00001848",
  3125 => x"00001f97",
  3126 => x"00001f97",
  3127 => x"000021e3",
  3128 => x"00002157",
  3129 => x"000020cb",
  3130 => x"000018c4",
  3131 => x"0000203f",
  3132 => x"00001fb3",
  3133 => x"64756d6d",
  3134 => x"792e6578",
  3135 => x"65000000",
  3136 => x"43000000",
  3137 => x"00ffffff",
  3138 => x"ff00ffff",
  3139 => x"ffff00ff",
  3140 => x"ffffff00",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"000034cc",
  3145 => x"fff00000",
  3146 => x"80000e00",
  3147 => x"80000800",
  3148 => x"80000600",
  3149 => x"80000200",
  3150 => x"80000100",
  3151 => x"000030f4",
  3152 => x"00003144",
  3153 => x"00000000",
  3154 => x"000033ac",
  3155 => x"00003408",
  3156 => x"00003464",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"00000000",
  3161 => x"00000000",
  3162 => x"00000000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"00000000",
  3166 => x"00003100",
  3167 => x"00000000",
  3168 => x"00000000",
  3169 => x"00000000",
  3170 => x"00000000",
  3171 => x"00000000",
  3172 => x"00000000",
  3173 => x"00000000",
  3174 => x"00000000",
  3175 => x"00000000",
  3176 => x"00000000",
  3177 => x"00000000",
  3178 => x"00000000",
  3179 => x"00000000",
  3180 => x"00000000",
  3181 => x"00000000",
  3182 => x"00000000",
  3183 => x"00000000",
  3184 => x"00000000",
  3185 => x"00000000",
  3186 => x"00000000",
  3187 => x"00000000",
  3188 => x"00000000",
  3189 => x"00000000",
  3190 => x"00000000",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00000000",
  3195 => x"00000001",
  3196 => x"330eabcd",
  3197 => x"1234e66d",
  3198 => x"deec0005",
  3199 => x"000b0000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"00000000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000000",
  3246 => x"00000000",
  3247 => x"00000000",
  3248 => x"00000000",
  3249 => x"00000000",
  3250 => x"00000000",
  3251 => x"00000000",
  3252 => x"00000000",
  3253 => x"00000000",
  3254 => x"00000000",
  3255 => x"00000000",
  3256 => x"00000000",
  3257 => x"00000000",
  3258 => x"00000000",
  3259 => x"00000000",
  3260 => x"00000000",
  3261 => x"00000000",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00000000",
  3265 => x"00000000",
  3266 => x"00000000",
  3267 => x"00000000",
  3268 => x"00000000",
  3269 => x"00000000",
  3270 => x"00000000",
  3271 => x"00000000",
  3272 => x"00000000",
  3273 => x"00000000",
  3274 => x"00000000",
  3275 => x"00000000",
  3276 => x"00000000",
  3277 => x"00000000",
  3278 => x"00000000",
  3279 => x"00000000",
  3280 => x"00000000",
  3281 => x"00000000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"00000000",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00000000",
  3288 => x"00000000",
  3289 => x"00000000",
  3290 => x"00000000",
  3291 => x"00000000",
  3292 => x"00000000",
  3293 => x"00000000",
  3294 => x"00000000",
  3295 => x"00000000",
  3296 => x"00000000",
  3297 => x"00000000",
  3298 => x"00000000",
  3299 => x"00000000",
  3300 => x"00000000",
  3301 => x"00000000",
  3302 => x"00000000",
  3303 => x"00000000",
  3304 => x"00000000",
  3305 => x"00000000",
  3306 => x"00000000",
  3307 => x"00000000",
  3308 => x"00000000",
  3309 => x"00000000",
  3310 => x"00000000",
  3311 => x"00000000",
  3312 => x"00000000",
  3313 => x"00000000",
  3314 => x"00000000",
  3315 => x"00000000",
  3316 => x"00000000",
  3317 => x"00000000",
  3318 => x"00000000",
  3319 => x"00000000",
  3320 => x"00000000",
  3321 => x"00000000",
  3322 => x"00000000",
  3323 => x"00000000",
  3324 => x"00000000",
  3325 => x"00000000",
  3326 => x"00000000",
  3327 => x"00000000",
  3328 => x"00000000",
  3329 => x"00000000",
  3330 => x"00000000",
  3331 => x"00000000",
  3332 => x"00000000",
  3333 => x"00000000",
  3334 => x"00000000",
  3335 => x"00000000",
  3336 => x"00000000",
  3337 => x"00000000",
  3338 => x"00000000",
  3339 => x"00000000",
  3340 => x"00000000",
  3341 => x"00000000",
  3342 => x"00000000",
  3343 => x"00000000",
  3344 => x"00000000",
  3345 => x"00000000",
  3346 => x"00000000",
  3347 => x"00000000",
  3348 => x"00000000",
  3349 => x"00000000",
  3350 => x"00000000",
  3351 => x"00000000",
  3352 => x"00000000",
  3353 => x"00000000",
  3354 => x"00000000",
  3355 => x"00000000",
  3356 => x"00000000",
  3357 => x"00000000",
  3358 => x"00000000",
  3359 => x"00000000",
  3360 => x"00000000",
  3361 => x"00000000",
  3362 => x"00000000",
  3363 => x"00000000",
  3364 => x"00000000",
  3365 => x"00000000",
  3366 => x"00000000",
  3367 => x"00000000",
  3368 => x"00000000",
  3369 => x"00000000",
  3370 => x"00000000",
  3371 => x"00000000",
  3372 => x"00000000",
  3373 => x"00000000",
  3374 => x"00000000",
  3375 => x"00000000",
  3376 => x"ffffffff",
  3377 => x"00000000",
  3378 => x"ffffffff",
  3379 => x"00000000",
  3380 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
