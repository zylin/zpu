library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"82f4e00c",
3 => x"3a0b0b81",
4 => x"e48c0400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"81e4fd2d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c9040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88ac",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b82f4",
162 => x"cc738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88af0400",
166 => x"00000000",
167 => x"00000000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0b8e",
171 => x"c42d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0b90",
179 => x"8d2d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"82f4dc0c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"0b0b0b83",
257 => x"e93f0b0b",
258 => x"82e4cc3f",
259 => x"04101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101010",
266 => x"10101010",
267 => x"53510473",
268 => x"81ff0673",
269 => x"83060981",
270 => x"05830510",
271 => x"10102b07",
272 => x"72fc060c",
273 => x"5151043c",
274 => x"04727280",
275 => x"728106ff",
276 => x"05097206",
277 => x"05711052",
278 => x"720a100a",
279 => x"5372ed38",
280 => x"51515351",
281 => x"04fe3d0d",
282 => x"0b0b8384",
283 => x"e8085384",
284 => x"13087088",
285 => x"2a708106",
286 => x"51525270",
287 => x"802e0b0b",
288 => x"0b0bec38",
289 => x"7181ff06",
290 => x"800c843d",
291 => x"0d04ff3d",
292 => x"0d0b0b83",
293 => x"84e80852",
294 => x"71087088",
295 => x"2a813270",
296 => x"81065151",
297 => x"51700b0b",
298 => x"0b0bed38",
299 => x"73720c83",
300 => x"3d0d040b",
301 => x"0b82f4dc",
302 => x"08802e0b",
303 => x"0b0b0bae",
304 => x"380b0b82",
305 => x"f4e00882",
306 => x"2e0b0b0b",
307 => x"80c53883",
308 => x"80800b0b",
309 => x"0b8384e8",
310 => x"0c82a080",
311 => x"0b0b0b83",
312 => x"84ec0c82",
313 => x"90800b0b",
314 => x"0b8384f0",
315 => x"0c04f880",
316 => x"8080a40b",
317 => x"0b0b8384",
318 => x"e80cf880",
319 => x"8082800b",
320 => x"0b0b8384",
321 => x"ec0cf880",
322 => x"8084800b",
323 => x"0b0b8384",
324 => x"f00c0480",
325 => x"c0a8808c",
326 => x"0b0b0b83",
327 => x"84e80c80",
328 => x"c0a88094",
329 => x"0b0b0b83",
330 => x"84ec0c0b",
331 => x"0b82ed90",
332 => x"0b0b0b83",
333 => x"84f00c04",
334 => x"f23d0d60",
335 => x"0b0b8384",
336 => x"ec08565d",
337 => x"82750c80",
338 => x"59805a80",
339 => x"0b8f3d5d",
340 => x"5b7a1010",
341 => x"15700871",
342 => x"08719f2c",
343 => x"7e852b58",
344 => x"55557d53",
345 => x"59570b0b",
346 => x"0b81d13f",
347 => x"7d7f7a72",
348 => x"077c7207",
349 => x"71716081",
350 => x"05415f5d",
351 => x"5b595755",
352 => x"817b270b",
353 => x"0b0b0b8f",
354 => x"38767d0c",
355 => x"77841e0c",
356 => x"7c800c90",
357 => x"3d0d040b",
358 => x"0b8384ec",
359 => x"08550b0b",
360 => x"0bffae39",
361 => x"70700b0b",
362 => x"8384f433",
363 => x"51700b0b",
364 => x"0b0bb738",
365 => x"0b0b82f4",
366 => x"e8087008",
367 => x"52527080",
368 => x"2e0b0b0b",
369 => x"0b9c3884",
370 => x"120b0b82",
371 => x"f4e80c70",
372 => x"2d0b0b82",
373 => x"f4e80870",
374 => x"08525270",
375 => x"0b0b0b0b",
376 => x"e638810b",
377 => x"0b0b8384",
378 => x"f4345050",
379 => x"0404700b",
380 => x"0b8384e4",
381 => x"08802e0b",
382 => x"0b0b0b92",
383 => x"380b0b0b",
384 => x"0b800b80",
385 => x"2e098106",
386 => x"0b0b0b0b",
387 => x"83385004",
388 => x"0b0b8384",
389 => x"e4510b0b",
390 => x"0bf3e53f",
391 => x"5004048c",
392 => x"08028c0c",
393 => x"ff3d0d0b",
394 => x"0b82ed94",
395 => x"510b0b0b",
396 => x"88ab3f71",
397 => x"800c833d",
398 => x"0d8c0c04",
399 => x"8c08028c",
400 => x"0cf53d0d",
401 => x"8c089405",
402 => x"080b0b0b",
403 => x"0ba0388c",
404 => x"088c0508",
405 => x"8c089005",
406 => x"088c0888",
407 => x"05085856",
408 => x"5473760c",
409 => x"7484170c",
410 => x"0b0b0b81",
411 => x"ca39800b",
412 => x"8c08f005",
413 => x"0c800b8c",
414 => x"08f4050c",
415 => x"8c088c05",
416 => x"088c0890",
417 => x"05085654",
418 => x"738c08f0",
419 => x"050c748c",
420 => x"08f4050c",
421 => x"8c08f805",
422 => x"8c08f005",
423 => x"56568870",
424 => x"54755376",
425 => x"52540b0b",
426 => x"0b85e03f",
427 => x"a00b8c08",
428 => x"94050831",
429 => x"8c08ec05",
430 => x"0c8c08ec",
431 => x"05088024",
432 => x"0b0b0b0b",
433 => x"a138800b",
434 => x"8c08f405",
435 => x"0c8c08ec",
436 => x"0508308c",
437 => x"08fc0508",
438 => x"712b8c08",
439 => x"f0050c54",
440 => x"0b0b0b0b",
441 => x"b9398c08",
442 => x"fc05088c",
443 => x"08ec0508",
444 => x"2a8c08e8",
445 => x"050c8c08",
446 => x"fc05088c",
447 => x"08940508",
448 => x"2b8c08f4",
449 => x"050c8c08",
450 => x"f805088c",
451 => x"08940508",
452 => x"2b708c08",
453 => x"e8050807",
454 => x"8c08f005",
455 => x"0c548c08",
456 => x"f005088c",
457 => x"08f40508",
458 => x"8c088805",
459 => x"08585654",
460 => x"73760c74",
461 => x"84170c8c",
462 => x"08880508",
463 => x"800c8d3d",
464 => x"0d8c0c04",
465 => x"8c08028c",
466 => x"0cf93d0d",
467 => x"800b8c08",
468 => x"fc050c8c",
469 => x"08880508",
470 => x"80250b0b",
471 => x"0b0baf38",
472 => x"8c088805",
473 => x"08308c08",
474 => x"88050c80",
475 => x"0b8c08f4",
476 => x"050c8c08",
477 => x"fc05080b",
478 => x"0b0b0b88",
479 => x"38810b8c",
480 => x"08f4050c",
481 => x"8c08f405",
482 => x"088c08fc",
483 => x"050c8c08",
484 => x"8c050880",
485 => x"250b0b0b",
486 => x"0baf388c",
487 => x"088c0508",
488 => x"308c088c",
489 => x"050c800b",
490 => x"8c08f005",
491 => x"0c8c08fc",
492 => x"05080b0b",
493 => x"0b0b8838",
494 => x"810b8c08",
495 => x"f0050c8c",
496 => x"08f00508",
497 => x"8c08fc05",
498 => x"0c80538c",
499 => x"088c0508",
500 => x"528c0888",
501 => x"0508510b",
502 => x"0b0b81bb",
503 => x"3f800870",
504 => x"8c08f805",
505 => x"0c548c08",
506 => x"fc050880",
507 => x"2e0b0b0b",
508 => x"0b8c388c",
509 => x"08f80508",
510 => x"308c08f8",
511 => x"050c8c08",
512 => x"f8050870",
513 => x"800c5489",
514 => x"3d0d8c0c",
515 => x"048c0802",
516 => x"8c0cfb3d",
517 => x"0d800b8c",
518 => x"08fc050c",
519 => x"8c088805",
520 => x"0880250b",
521 => x"0b0b0b93",
522 => x"388c0888",
523 => x"0508308c",
524 => x"0888050c",
525 => x"810b8c08",
526 => x"fc050c8c",
527 => x"088c0508",
528 => x"80250b0b",
529 => x"0b0b8c38",
530 => x"8c088c05",
531 => x"08308c08",
532 => x"8c050c81",
533 => x"538c088c",
534 => x"0508528c",
535 => x"08880508",
536 => x"510b0b0b",
537 => x"0bb13f80",
538 => x"08708c08",
539 => x"f8050c54",
540 => x"8c08fc05",
541 => x"08802e0b",
542 => x"0b0b0b8c",
543 => x"388c08f8",
544 => x"0508308c",
545 => x"08f8050c",
546 => x"8c08f805",
547 => x"0870800c",
548 => x"54873d0d",
549 => x"8c0c048c",
550 => x"08028c0c",
551 => x"70707070",
552 => x"810b8c08",
553 => x"fc050c80",
554 => x"0b8c08f8",
555 => x"050c8c08",
556 => x"8c05088c",
557 => x"08880508",
558 => x"270b0b0b",
559 => x"0bb8388c",
560 => x"08fc0508",
561 => x"802e0b0b",
562 => x"0b0bab38",
563 => x"800b8c08",
564 => x"8c050824",
565 => x"0b0b0b0b",
566 => x"9d388c08",
567 => x"8c050810",
568 => x"8c088c05",
569 => x"0c8c08fc",
570 => x"0508108c",
571 => x"08fc050c",
572 => x"0b0b0bff",
573 => x"b9398c08",
574 => x"fc050880",
575 => x"2e0b0b0b",
576 => x"80d0388c",
577 => x"088c0508",
578 => x"8c088805",
579 => x"08260b0b",
580 => x"0b0ba138",
581 => x"8c088805",
582 => x"088c088c",
583 => x"0508318c",
584 => x"0888050c",
585 => x"8c08f805",
586 => x"088c08fc",
587 => x"0508078c",
588 => x"08f8050c",
589 => x"8c08fc05",
590 => x"08812a8c",
591 => x"08fc050c",
592 => x"8c088c05",
593 => x"08812a8c",
594 => x"088c050c",
595 => x"0b0b0bff",
596 => x"a5398c08",
597 => x"90050880",
598 => x"2e0b0b0b",
599 => x"0b93388c",
600 => x"08880508",
601 => x"708c08f4",
602 => x"050c510b",
603 => x"0b0b0b8d",
604 => x"398c08f8",
605 => x"0508708c",
606 => x"08f4050c",
607 => x"518c08f4",
608 => x"0508800c",
609 => x"50505050",
610 => x"8c0c04fc",
611 => x"3d0d7670",
612 => x"797b5555",
613 => x"55558f72",
614 => x"270b0b0b",
615 => x"0b903872",
616 => x"75078306",
617 => x"5170802e",
618 => x"0b0b0b0b",
619 => x"af38ff12",
620 => x"5271ff2e",
621 => x"0b0b0b0b",
622 => x"9c387270",
623 => x"81055433",
624 => x"74708105",
625 => x"5634ff12",
626 => x"5271ff2e",
627 => x"0981060b",
628 => x"0b0b0be6",
629 => x"3874800c",
630 => x"863d0d04",
631 => x"74517270",
632 => x"84055408",
633 => x"71708405",
634 => x"530c7270",
635 => x"84055408",
636 => x"71708405",
637 => x"530c7270",
638 => x"84055408",
639 => x"71708405",
640 => x"530c7270",
641 => x"84055408",
642 => x"71708405",
643 => x"530cf012",
644 => x"52718f26",
645 => x"0b0b0b0b",
646 => x"c5388372",
647 => x"270b0b0b",
648 => x"0b993872",
649 => x"70840554",
650 => x"08717084",
651 => x"05530cfc",
652 => x"12527183",
653 => x"260b0b0b",
654 => x"0be93870",
655 => x"540b0b0b",
656 => x"feec39fb",
657 => x"3d0d7789",
658 => x"3d880555",
659 => x"79548811",
660 => x"0853510b",
661 => x"0b0b80e3",
662 => x"3f873d0d",
663 => x"04fc3d0d",
664 => x"873d7070",
665 => x"84055208",
666 => x"56537452",
667 => x"0b0b82f4",
668 => x"ec088811",
669 => x"0852540b",
670 => x"0b0bb4a2",
671 => x"3f863d0d",
672 => x"04707070",
673 => x"70768811",
674 => x"08545472",
675 => x"0b0b0b0b",
676 => x"8d387284",
677 => x"150c7280",
678 => x"0c505050",
679 => x"50047352",
680 => x"75510b0b",
681 => x"80fcfe3f",
682 => x"800b8815",
683 => x"0c800b84",
684 => x"150c8008",
685 => x"800c5050",
686 => x"505004fc",
687 => x"c43d0d83",
688 => x"bf3d0883",
689 => x"c13d0883",
690 => x"c33d0883",
691 => x"c53d0848",
692 => x"5e484b0b",
693 => x"0b8186f6",
694 => x"3f800808",
695 => x"4c800b83",
696 => x"bb3d0c80",
697 => x"0b83bc3d",
698 => x"0c807071",
699 => x"698c0522",
700 => x"70832a81",
701 => x"32708106",
702 => x"515d5d4c",
703 => x"4f4d786d",
704 => x"2e098106",
705 => x"0b0b0b0b",
706 => x"90386690",
707 => x"05086d2e",
708 => x"0981060b",
709 => x"0b0b0b98",
710 => x"3866510b",
711 => x"0b0bbfc8",
712 => x"3fff5980",
713 => x"080b0b0b",
714 => x"82893866",
715 => x"8c05225a",
716 => x"799a0659",
717 => x"788a2e0b",
718 => x"0b0b80ce",
719 => x"387b83a6",
720 => x"3d707183",
721 => x"b93d0c5e",
722 => x"475d800b",
723 => x"83b83d0c",
724 => x"800b83b7",
725 => x"3d0c8049",
726 => x"7c5e807d",
727 => x"337081ff",
728 => x"065b5b5b",
729 => x"787b2e0b",
730 => x"0b0b0b83",
731 => x"38815b78",
732 => x"a52e0b0b",
733 => x"0b81c438",
734 => x"7a802e0b",
735 => x"0b0b81bb",
736 => x"38811d5d",
737 => x"0b0b0b0b",
738 => x"d139668e",
739 => x"05227090",
740 => x"2b5a5b80",
741 => x"79240b0b",
742 => x"0bffa238",
743 => x"79fd0659",
744 => x"7882ba3d",
745 => x"237a0284",
746 => x"0589e205",
747 => x"23669c05",
748 => x"0882be3d",
749 => x"0c66a405",
750 => x"0882c03d",
751 => x"0cb63d70",
752 => x"82b83d0c",
753 => x"82bb3d0c",
754 => x"88800b82",
755 => x"b93d0c88",
756 => x"800b82bc",
757 => x"3d0c800b",
758 => x"82bd3d0c",
759 => x"64537b52",
760 => x"82b63d70",
761 => x"52590b0b",
762 => x"0bb1b33f",
763 => x"80085a80",
764 => x"0b800824",
765 => x"0b0b0b0b",
766 => x"95387851",
767 => x"0b0b80ec",
768 => x"bf3f8008",
769 => x"802e0b0b",
770 => x"0b0b8338",
771 => x"ff5a82b9",
772 => x"3d227086",
773 => x"2a708106",
774 => x"515a5b78",
775 => x"802e0b0b",
776 => x"0b0b8e38",
777 => x"668c0522",
778 => x"80c00759",
779 => x"78678c05",
780 => x"23795978",
781 => x"800c83be",
782 => x"3d0d047c",
783 => x"7e315b7a",
784 => x"802e0b0b",
785 => x"0b0bb138",
786 => x"7d7c0c7a",
787 => x"841d0c83",
788 => x"b73d081b",
789 => x"83b83d0c",
790 => x"881c83b7",
791 => x"3d088111",
792 => x"83b93d0c",
793 => x"8111515a",
794 => x"5c788724",
795 => x"0b0b0b80",
796 => x"cb38681b",
797 => x"7d335b49",
798 => x"7981ff06",
799 => x"5978802e",
800 => x"0b0b0bae",
801 => x"df38811d",
802 => x"5d807071",
803 => x"4a4543ff",
804 => x"416283be",
805 => x"3d347c33",
806 => x"5a7981ff",
807 => x"06811e5e",
808 => x"407fe005",
809 => x"597880d8",
810 => x"260b0b0b",
811 => x"88a83878",
812 => x"10100b0b",
813 => x"82edc405",
814 => x"59780804",
815 => x"83be3ddc",
816 => x"05526651",
817 => x"0b0b0bfb",
818 => x"b83f8008",
819 => x"0b0b0b8b",
820 => x"b3386569",
821 => x"1c7e335c",
822 => x"4a5c0b0b",
823 => x"0bff9939",
824 => x"62900743",
825 => x"62842a70",
826 => x"81065159",
827 => x"780b0b0b",
828 => x"9e873862",
829 => x"862a7081",
830 => x"06515978",
831 => x"802e0b0b",
832 => x"0b9df638",
833 => x"64658405",
834 => x"8212225d",
835 => x"4659815f",
836 => x"800b83be",
837 => x"3d346044",
838 => x"8061240b",
839 => x"0b0b0b86",
840 => x"3862feff",
841 => x"0643657b",
842 => x"30707d07",
843 => x"9f2a6630",
844 => x"7068079f",
845 => x"2a720752",
846 => x"5c515b5e",
847 => x"79802e0b",
848 => x"0b0b98fd",
849 => x"387e812e",
850 => x"0b0b0b8c",
851 => x"8438817f",
852 => x"250b0b0b",
853 => x"a0eb387e",
854 => x"822e0b0b",
855 => x"0b8cc038",
856 => x"0b0b82f0",
857 => x"a85e7d51",
858 => x"0b0b81c0",
859 => x"ae3f8008",
860 => x"5f7e427e",
861 => x"64250b0b",
862 => x"0b0b8338",
863 => x"634283bd",
864 => x"3d337081",
865 => x"ff065a5b",
866 => x"78802e0b",
867 => x"0b0b9488",
868 => x"38618105",
869 => x"42628184",
870 => x"0641600b",
871 => x"0b0b8186",
872 => x"38676231",
873 => x"5a807a25",
874 => x"0b0b0b80",
875 => x"f938907a",
876 => x"250b0b0b",
877 => x"0bbd380b",
878 => x"0b82eda4",
879 => x"7c0c900b",
880 => x"841d0c83",
881 => x"b73d0890",
882 => x"0583b83d",
883 => x"0c881c83",
884 => x"b73d0881",
885 => x"1183b93d",
886 => x"0c811151",
887 => x"5a5c7887",
888 => x"240b0b0b",
889 => x"868e38f0",
890 => x"1a5a7990",
891 => x"240b0b0b",
892 => x"0bc5380b",
893 => x"0b82eda4",
894 => x"7c0c7984",
895 => x"1d0c83b7",
896 => x"3d081a83",
897 => x"b83d0c88",
898 => x"1c83b73d",
899 => x"08811183",
900 => x"b93d0c81",
901 => x"11515a5c",
902 => x"7887240b",
903 => x"0b0b96fe",
904 => x"3883bd3d",
905 => x"335b7a81",
906 => x"ff065978",
907 => x"802e0b0b",
908 => x"0b938138",
909 => x"83be3dfc",
910 => x"057c0c81",
911 => x"0b841d0c",
912 => x"83b73d08",
913 => x"810583b8",
914 => x"3d0c881c",
915 => x"83b73d08",
916 => x"811183b9",
917 => x"3d0c8111",
918 => x"515a5c78",
919 => x"87240b0b",
920 => x"0b879f38",
921 => x"6081802e",
922 => x"0b0b0b85",
923 => x"c938637f",
924 => x"315a807a",
925 => x"250b0b0b",
926 => x"818c3890",
927 => x"7a250b0b",
928 => x"0b0bbd38",
929 => x"0b0b82ed",
930 => x"b47c0c90",
931 => x"0b841d0c",
932 => x"83b73d08",
933 => x"900583b8",
934 => x"3d0c881c",
935 => x"83b73d08",
936 => x"811183b9",
937 => x"3d0c8111",
938 => x"515a5c78",
939 => x"87240b0b",
940 => x"0b84e238",
941 => x"f01a5a79",
942 => x"90240b0b",
943 => x"0b0bc538",
944 => x"0b0b82ed",
945 => x"b47c0c79",
946 => x"841d0c83",
947 => x"b73d081a",
948 => x"83b83d0c",
949 => x"881c83b7",
950 => x"3d088111",
951 => x"83b93d0c",
952 => x"8111515a",
953 => x"5c877925",
954 => x"0b0b0b0b",
955 => x"993883be",
956 => x"3ddc0552",
957 => x"66510b0b",
958 => x"0bf7863f",
959 => x"80080b0b",
960 => x"0b878138",
961 => x"655c6288",
962 => x"2a813270",
963 => x"81065159",
964 => x"78802e0b",
965 => x"0b0b91f3",
966 => x"387d7c0c",
967 => x"7e841d0c",
968 => x"83b73d08",
969 => x"1f83b83d",
970 => x"0c881c83",
971 => x"b73d0881",
972 => x"1183b93d",
973 => x"0c811151",
974 => x"5a5c7887",
975 => x"240b0b0b",
976 => x"868c3862",
977 => x"822a7081",
978 => x"06515978",
979 => x"802e0b0b",
980 => x"0b819438",
981 => x"6762315a",
982 => x"807a250b",
983 => x"0b0b8187",
984 => x"38907a25",
985 => x"0b0b0b0b",
986 => x"bd380b0b",
987 => x"82eda47c",
988 => x"0c900b84",
989 => x"1d0c83b7",
990 => x"3d089005",
991 => x"83b83d0c",
992 => x"881c83b7",
993 => x"3d088111",
994 => x"83b93d0c",
995 => x"8111515a",
996 => x"5c788724",
997 => x"0b0b0b85",
998 => x"9438f01a",
999 => x"5a799024",
1000 => x"0b0b0b0b",
1001 => x"c5380b0b",
1002 => x"82eda47c",
1003 => x"0c79841d",
1004 => x"0c83b73d",
1005 => x"081a83b8",
1006 => x"3d0c83b6",
1007 => x"3d088111",
1008 => x"83b83d0c",
1009 => x"81115159",
1010 => x"8779250b",
1011 => x"0b0b0b97",
1012 => x"3883be3d",
1013 => x"dc055266",
1014 => x"510b0b0b",
1015 => x"f5a33f80",
1016 => x"080b0b0b",
1017 => x"859e3861",
1018 => x"59616825",
1019 => x"0b0b0b0b",
1020 => x"83386759",
1021 => x"68194983",
1022 => x"b73d080b",
1023 => x"0b0b84ec",
1024 => x"38800b83",
1025 => x"b73d0c65",
1026 => x"5c69802e",
1027 => x"0b0b0bf6",
1028 => x"c7386951",
1029 => x"0b0b80ff",
1030 => x"953f807d",
1031 => x"5f4a0b0b",
1032 => x"0bf6b739",
1033 => x"62900743",
1034 => x"62842a70",
1035 => x"81065159",
1036 => x"780b0b0b",
1037 => x"97d43862",
1038 => x"862a7081",
1039 => x"06515978",
1040 => x"802e0b0b",
1041 => x"0b97c338",
1042 => x"64658405",
1043 => x"8212225d",
1044 => x"4659805f",
1045 => x"800b83be",
1046 => x"3d340b0b",
1047 => x"0bf9b739",
1048 => x"62900743",
1049 => x"62842a70",
1050 => x"81065159",
1051 => x"780b0b0b",
1052 => x"97a93862",
1053 => x"862a7081",
1054 => x"06515978",
1055 => x"802e0b0b",
1056 => x"0b979838",
1057 => x"64658405",
1058 => x"7108902b",
1059 => x"70902c51",
1060 => x"5d465980",
1061 => x"7b240b0b",
1062 => x"0b8bdf38",
1063 => x"815f0b0b",
1064 => x"0bf8f339",
1065 => x"64658405",
1066 => x"71084a46",
1067 => x"59678025",
1068 => x"0b0b0bf7",
1069 => x"e1386730",
1070 => x"48628407",
1071 => x"7d335b43",
1072 => x"0b0b0bf7",
1073 => x"d439811d",
1074 => x"5d629007",
1075 => x"7d335b43",
1076 => x"0b0b0bf7",
1077 => x"c4397f80",
1078 => x"2e0b0b0b",
1079 => x"a6863882",
1080 => x"ce3d5e7f",
1081 => x"7e34815f",
1082 => x"800b83be",
1083 => x"3d340b0b",
1084 => x"0bf8fe39",
1085 => x"83be3ddc",
1086 => x"05526651",
1087 => x"0b0b0bf3",
1088 => x"803f8008",
1089 => x"0b0b0b82",
1090 => x"fb3865f0",
1091 => x"1b5b5c0b",
1092 => x"0b0bf9d6",
1093 => x"3983be3d",
1094 => x"dc055266",
1095 => x"510b0b0b",
1096 => x"f2df3f80",
1097 => x"080b0b0b",
1098 => x"82da3865",
1099 => x"f01b5b5c",
1100 => x"0b0b0bfb",
1101 => x"82396762",
1102 => x"315a807a",
1103 => x"250b0b0b",
1104 => x"faac3890",
1105 => x"7a250b0b",
1106 => x"0b0bbd38",
1107 => x"0b0b82ed",
1108 => x"b47c0c90",
1109 => x"0b841d0c",
1110 => x"83b73d08",
1111 => x"900583b8",
1112 => x"3d0c881c",
1113 => x"83b73d08",
1114 => x"811183b9",
1115 => x"3d0c8111",
1116 => x"515a5c78",
1117 => x"87240b0b",
1118 => x"0b80e638",
1119 => x"f01a5a79",
1120 => x"90240b0b",
1121 => x"0b0bc538",
1122 => x"0b0b82ed",
1123 => x"b47c0c79",
1124 => x"841d0c83",
1125 => x"b73d081a",
1126 => x"83b83d0c",
1127 => x"881c83b7",
1128 => x"3d088111",
1129 => x"83b93d0c",
1130 => x"8111515a",
1131 => x"5c877925",
1132 => x"0b0b0bf9",
1133 => x"b93883be",
1134 => x"3ddc0552",
1135 => x"66510b0b",
1136 => x"0bf1be3f",
1137 => x"80080b0b",
1138 => x"0b81b938",
1139 => x"65646031",
1140 => x"5b5c7980",
1141 => x"240b0b0b",
1142 => x"f9a1380b",
1143 => x"0b0bfaa6",
1144 => x"3983be3d",
1145 => x"dc055266",
1146 => x"510b0b0b",
1147 => x"f1933f80",
1148 => x"080b0b0b",
1149 => x"818e3865",
1150 => x"f01b5b5c",
1151 => x"0b0b0bfe",
1152 => x"fe3983be",
1153 => x"3ddc0552",
1154 => x"66510b0b",
1155 => x"0bf0f23f",
1156 => x"80080b0b",
1157 => x"0b80ed38",
1158 => x"655c6081",
1159 => x"802e0981",
1160 => x"060b0b0b",
1161 => x"f8c8380b",
1162 => x"0b0bfe8a",
1163 => x"3983be3d",
1164 => x"dc055266",
1165 => x"510b0b0b",
1166 => x"f0c73f80",
1167 => x"080b0b0b",
1168 => x"80c23865",
1169 => x"f01b5b5c",
1170 => x"0b0b0bfa",
1171 => x"d03983be",
1172 => x"3ddc0552",
1173 => x"66510b0b",
1174 => x"0bf0a63f",
1175 => x"80080b0b",
1176 => x"0b0ba138",
1177 => x"655c0b0b",
1178 => x"0bf9d839",
1179 => x"83be3ddc",
1180 => x"05526651",
1181 => x"0b0b0bf0",
1182 => x"883f8008",
1183 => x"802e0b0b",
1184 => x"0bfafe38",
1185 => x"69802e0b",
1186 => x"0b0b0b89",
1187 => x"3869510b",
1188 => x"0b80fa9a",
1189 => x"3f668c05",
1190 => x"2270862a",
1191 => x"7081066b",
1192 => x"5d515a47",
1193 => x"78802e0b",
1194 => x"0b0bf385",
1195 => x"38ff590b",
1196 => x"0b0bf2ff",
1197 => x"397c3370",
1198 => x"81ff065a",
1199 => x"5a7880ec",
1200 => x"2e0b0b0b",
1201 => x"fc803862",
1202 => x"90077a81",
1203 => x"ff06811f",
1204 => x"5f41430b",
1205 => x"0b0bf3c9",
1206 => x"397c7081",
1207 => x"055e3340",
1208 => x"7faa2e0b",
1209 => x"0b0ba2f9",
1210 => x"388060d0",
1211 => x"0571435a",
1212 => x"5a788926",
1213 => x"0b0b0bf3",
1214 => x"a8387910",
1215 => x"10107a10",
1216 => x"056005d0",
1217 => x"057d7081",
1218 => x"055f33d0",
1219 => x"115b415a",
1220 => x"8979270b",
1221 => x"0b0b0be2",
1222 => x"38794179",
1223 => x"ff250b0b",
1224 => x"0bf2fe38",
1225 => x"ff410b0b",
1226 => x"0bf2f639",
1227 => x"64658405",
1228 => x"71085d46",
1229 => x"59820b0b",
1230 => x"0b82f0c4",
1231 => x"64720745",
1232 => x"4f5f80f8",
1233 => x"40800b83",
1234 => x"be3d340b",
1235 => x"0b0bf3c6",
1236 => x"39897b27",
1237 => x"0b0b0b0b",
1238 => x"ac38ff1e",
1239 => x"5e8a527a",
1240 => x"510b0b82",
1241 => x"9e803f80",
1242 => x"08b00559",
1243 => x"787e348a",
1244 => x"527a510b",
1245 => x"0b829dc4",
1246 => x"3f80085b",
1247 => x"7a89260b",
1248 => x"0b0b0bd6",
1249 => x"38ff1eb0",
1250 => x"1c5a5e78",
1251 => x"7e3483be",
1252 => x"3d707f31",
1253 => x"ff9c0540",
1254 => x"5b0b0b0b",
1255 => x"f3d339ff",
1256 => x"1e7b8f06",
1257 => x"6f055a5e",
1258 => x"78337e34",
1259 => x"7a842a5b",
1260 => x"7a802e0b",
1261 => x"0b0b0bd6",
1262 => x"38ff1e7b",
1263 => x"8f066f05",
1264 => x"5a5e7833",
1265 => x"7e347a84",
1266 => x"2a5b7a0b",
1267 => x"0b0b0bcf",
1268 => x"380b0b0b",
1269 => x"ffb83962",
1270 => x"80c0077d",
1271 => x"335b430b",
1272 => x"0b0bf1b5",
1273 => x"3960ff2e",
1274 => x"0b0b0b9f",
1275 => x"a0387f80",
1276 => x"e7327030",
1277 => x"70720780",
1278 => x"256280c7",
1279 => x"32703070",
1280 => x"72078025",
1281 => x"73075354",
1282 => x"5e515b59",
1283 => x"79802e0b",
1284 => x"0b0b0b8a",
1285 => x"38600b0b",
1286 => x"0b0b8338",
1287 => x"81416465",
1288 => x"88058412",
1289 => x"08720870",
1290 => x"83bf3d0c",
1291 => x"7183c03d",
1292 => x"0c545446",
1293 => x"590b0b81",
1294 => x"adad3f80",
1295 => x"08802e0b",
1296 => x"0b0b95db",
1297 => x"38805980",
1298 => x"79545483",
1299 => x"ba3d0883",
1300 => x"bc3d085b",
1301 => x"5179520b",
1302 => x"0b8290c9",
1303 => x"3f800b80",
1304 => x"08240b0b",
1305 => x"0b85f138",
1306 => x"0b0b82f0",
1307 => x"d85e835f",
1308 => x"0b0b0bf1",
1309 => x"fc3982ce",
1310 => x"3d5e7f80",
1311 => x"c32e0b0b",
1312 => x"0b0b9238",
1313 => x"62842a70",
1314 => x"81065159",
1315 => x"78802e0b",
1316 => x"0b0b83d3",
1317 => x"38885380",
1318 => x"52b43d70",
1319 => x"52590b0b",
1320 => x"8188f23f",
1321 => x"78546465",
1322 => x"84057108",
1323 => x"557f546c",
1324 => x"5346590b",
1325 => x"0b0ba0b1",
1326 => x"3f80085f",
1327 => x"8008ff2e",
1328 => x"0b0b0bfb",
1329 => x"bf38800b",
1330 => x"83be3d34",
1331 => x"0b0b0bf1",
1332 => x"a0390b0b",
1333 => x"82f0dc63",
1334 => x"842a7081",
1335 => x"06515a4e",
1336 => x"780b0b0b",
1337 => x"82ca3862",
1338 => x"862a7081",
1339 => x"06515978",
1340 => x"802e0b0b",
1341 => x"0b82b938",
1342 => x"64658405",
1343 => x"8212225d",
1344 => x"46598263",
1345 => x"81065a5f",
1346 => x"7a802e0b",
1347 => x"0b0bf080",
1348 => x"3878802e",
1349 => x"0b0b0bef",
1350 => x"f738627f",
1351 => x"0743800b",
1352 => x"83be3d34",
1353 => x"0b0b0bef",
1354 => x"ed39800b",
1355 => x"83be3d34",
1356 => x"64658405",
1357 => x"71084046",
1358 => x"597d802e",
1359 => x"0b0b0b9c",
1360 => x"d4387f80",
1361 => x"d32e0b0b",
1362 => x"0b82c038",
1363 => x"62842a70",
1364 => x"81065159",
1365 => x"780b0b0b",
1366 => x"82b13880",
1367 => x"61240b0b",
1368 => x"0bf08338",
1369 => x"60537852",
1370 => x"7d510b0b",
1371 => x"8183e73f",
1372 => x"605f8008",
1373 => x"802e0b0b",
1374 => x"0beff638",
1375 => x"80087e31",
1376 => x"5f607f25",
1377 => x"0b0b0bef",
1378 => x"e838605f",
1379 => x"0b0b0bef",
1380 => x"e0396284",
1381 => x"2a708106",
1382 => x"5159780b",
1383 => x"0b0b908d",
1384 => x"3862862a",
1385 => x"70810651",
1386 => x"5978802e",
1387 => x"0b0b0b8f",
1388 => x"fc386465",
1389 => x"84057108",
1390 => x"52465968",
1391 => x"79237c5e",
1392 => x"0b0b0beb",
1393 => x"9539ab0b",
1394 => x"83be3d34",
1395 => x"7c335a0b",
1396 => x"0b0bedc5",
1397 => x"39805a79",
1398 => x"1010107a",
1399 => x"10056005",
1400 => x"d0057d70",
1401 => x"81055f33",
1402 => x"d0115b41",
1403 => x"5a897927",
1404 => x"0b0b0b0b",
1405 => x"e2387948",
1406 => x"0b0b0bed",
1407 => x"a4396281",
1408 => x"80077d33",
1409 => x"5b430b0b",
1410 => x"0bed8e39",
1411 => x"6288077d",
1412 => x"335b430b",
1413 => x"0b0bed81",
1414 => x"390b0b82",
1415 => x"f0c46384",
1416 => x"2a708106",
1417 => x"515a4e78",
1418 => x"802e0b0b",
1419 => x"0bfdb838",
1420 => x"64658405",
1421 => x"71085d46",
1422 => x"590b0b0b",
1423 => x"fdc43962",
1424 => x"81077d33",
1425 => x"5b430b0b",
1426 => x"0becce39",
1427 => x"83bd3d33",
1428 => x"59780b0b",
1429 => x"0becbf38",
1430 => x"a00b83be",
1431 => x"3d347c33",
1432 => x"5a0b0b0b",
1433 => x"ecb33964",
1434 => x"65840546",
1435 => x"59831933",
1436 => x"7e34815f",
1437 => x"0b0b0bf4",
1438 => x"ef397a30",
1439 => x"5bad0b83",
1440 => x"be3d3481",
1441 => x"5f0b0b0b",
1442 => x"ed8c397d",
1443 => x"a23d0c80",
1444 => x"705c5f88",
1445 => x"537e52a6",
1446 => x"3d70525a",
1447 => x"0b0b8184",
1448 => x"f43f7e61",
1449 => x"240b0b0b",
1450 => x"81c2387a",
1451 => x"1010a23d",
1452 => x"08055978",
1453 => x"08802e0b",
1454 => x"0b0b0bbd",
1455 => x"38795478",
1456 => x"085383be",
1457 => x"3dfcc005",
1458 => x"526a510b",
1459 => x"0b0b9c99",
1460 => x"3f8008ff",
1461 => x"2e0b0b0b",
1462 => x"f7aa3880",
1463 => x"081f5978",
1464 => x"61240b0b",
1465 => x"0b0b9238",
1466 => x"811b7940",
1467 => x"5b78612e",
1468 => x"0981060b",
1469 => x"0b0bffb3",
1470 => x"387e802e",
1471 => x"0b0b0bec",
1472 => x"f038811f",
1473 => x"526a510b",
1474 => x"0b80f1b6",
1475 => x"3f80084a",
1476 => x"8008802e",
1477 => x"0b0b0bf6",
1478 => x"fc388853",
1479 => x"80527951",
1480 => x"0b0b8183",
1481 => x"f03f7955",
1482 => x"7e5483be",
1483 => x"3df38c05",
1484 => x"5369526a",
1485 => x"510b0b0b",
1486 => x"9cb03f80",
1487 => x"087f2e09",
1488 => x"81060b0b",
1489 => x"0bf6bd38",
1490 => x"696a8008",
1491 => x"055a5e80",
1492 => x"79340b0b",
1493 => x"0bec9a39",
1494 => x"ad0b83be",
1495 => x"3d340b0b",
1496 => x"82f0d85e",
1497 => x"835f0b0b",
1498 => x"0bec8639",
1499 => x"79557e54",
1500 => x"83be3df3",
1501 => x"8c05537e",
1502 => x"526a510b",
1503 => x"0b0b9bea",
1504 => x"3f80085f",
1505 => x"8008ff2e",
1506 => x"0b0b0bf5",
1507 => x"f7387da2",
1508 => x"3d0c0b0b",
1509 => x"0bfee239",
1510 => x"620a100a",
1511 => x"70810651",
1512 => x"5978802e",
1513 => x"0b0b0beb",
1514 => x"ec386182",
1515 => x"05420b0b",
1516 => x"0bebe239",
1517 => x"620a100a",
1518 => x"70810651",
1519 => x"5978802e",
1520 => x"0b0b0bed",
1521 => x"9f38b00b",
1522 => x"82ce3d34",
1523 => x"7f028405",
1524 => x"8ab10534",
1525 => x"83be3dfc",
1526 => x"bc057c0c",
1527 => x"820b841d",
1528 => x"0c83b73d",
1529 => x"08820583",
1530 => x"b83d0c88",
1531 => x"1c83b73d",
1532 => x"08811183",
1533 => x"b93d0c81",
1534 => x"11515a5c",
1535 => x"8779250b",
1536 => x"0b0bece0",
1537 => x"380b0b0b",
1538 => x"f3f83980",
1539 => x"e560250b",
1540 => x"0b0b83da",
1541 => x"38805980",
1542 => x"79545483",
1543 => x"ba3d0883",
1544 => x"bc3d085b",
1545 => x"5179520b",
1546 => x"0b8282bd",
1547 => x"3f80080b",
1548 => x"0b0b87ff",
1549 => x"380b0b82",
1550 => x"f0f07c0c",
1551 => x"810b841d",
1552 => x"0c83b73d",
1553 => x"08810583",
1554 => x"b83d0c88",
1555 => x"1c83b73d",
1556 => x"08811183",
1557 => x"b93d0c81",
1558 => x"11515a5c",
1559 => x"7887240b",
1560 => x"0b0b81ce",
1561 => x"38a43d08",
1562 => x"5b7aa63d",
1563 => x"08240b0b",
1564 => x"0b0b8e38",
1565 => x"62810659",
1566 => x"78802e0b",
1567 => x"0b0bedc3",
1568 => x"386b7c0c",
1569 => x"810b841d",
1570 => x"0c83b73d",
1571 => x"08810583",
1572 => x"b83d0c88",
1573 => x"1c83b73d",
1574 => x"08811183",
1575 => x"b93d0c81",
1576 => x"11515a5c",
1577 => x"7887240b",
1578 => x"0b0b81c5",
1579 => x"38ff1b5a",
1580 => x"807a250b",
1581 => x"0b0bed8b",
1582 => x"38907a25",
1583 => x"0b0b0b0b",
1584 => x"bd380b0b",
1585 => x"82edb47c",
1586 => x"0c900b84",
1587 => x"1d0c83b7",
1588 => x"3d089005",
1589 => x"83b83d0c",
1590 => x"881c83b7",
1591 => x"3d088111",
1592 => x"83b93d0c",
1593 => x"8111515a",
1594 => x"5c788724",
1595 => x"0b0b0b80",
1596 => x"df38f01a",
1597 => x"5a799024",
1598 => x"0b0b0b0b",
1599 => x"c5380b0b",
1600 => x"82edb47c",
1601 => x"0c79841d",
1602 => x"0c83b73d",
1603 => x"081a83b8",
1604 => x"3d0c881c",
1605 => x"83b73d08",
1606 => x"811183b9",
1607 => x"3d0c8111",
1608 => x"515a5c87",
1609 => x"79250b0b",
1610 => x"0bec9838",
1611 => x"0b0b0bf2",
1612 => x"9d3983be",
1613 => x"3ddc0552",
1614 => x"66510b0b",
1615 => x"0be2c23f",
1616 => x"80080b0b",
1617 => x"0bf2bd38",
1618 => x"655c0b0b",
1619 => x"0bfe9639",
1620 => x"83be3ddc",
1621 => x"05526651",
1622 => x"0b0b0be2",
1623 => x"a43f8008",
1624 => x"0b0b0bf2",
1625 => x"9f3865f0",
1626 => x"1b5b5c0b",
1627 => x"0b0bff85",
1628 => x"3983be3d",
1629 => x"dc055266",
1630 => x"510b0b0b",
1631 => x"e2833f80",
1632 => x"080b0b0b",
1633 => x"f1fe3865",
1634 => x"a53d08ff",
1635 => x"055b5c79",
1636 => x"80240b0b",
1637 => x"0bfea238",
1638 => x"0b0b0beb",
1639 => x"a63983be",
1640 => x"3ddc0552",
1641 => x"66510b0b",
1642 => x"0be1d63f",
1643 => x"80080b0b",
1644 => x"0bf1d138",
1645 => x"6583be3d",
1646 => x"335c5c0b",
1647 => x"0b0be8e6",
1648 => x"397e0b0b",
1649 => x"0bf3c738",
1650 => x"62810659",
1651 => x"78802e0b",
1652 => x"0b0bf3ba",
1653 => x"38028d8f",
1654 => x"055eb07e",
1655 => x"3483be3d",
1656 => x"707f31ff",
1657 => x"9c05405b",
1658 => x"0b0b0be7",
1659 => x"8439a43d",
1660 => x"085b817b",
1661 => x"250b0b0b",
1662 => x"83bc387d",
1663 => x"7081055f",
1664 => x"3382ce3d",
1665 => x"34ae0284",
1666 => x"058ab105",
1667 => x"3483be3d",
1668 => x"fcbc057c",
1669 => x"0c820b84",
1670 => x"1d0c83b7",
1671 => x"3d088205",
1672 => x"83b83d0c",
1673 => x"881c83b7",
1674 => x"3d088111",
1675 => x"83b93d0c",
1676 => x"8111515a",
1677 => x"5c788724",
1678 => x"0b0b0b81",
1679 => x"8b388059",
1680 => x"80795454",
1681 => x"83ba3d08",
1682 => x"83bc3d08",
1683 => x"5b517952",
1684 => x"0b0b8280",
1685 => x"a83f8008",
1686 => x"802e0b0b",
1687 => x"0b81a538",
1688 => x"7d7c0cff",
1689 => x"1b841d0c",
1690 => x"83b73d08",
1691 => x"1bff0583",
1692 => x"b83d0c88",
1693 => x"1c83b73d",
1694 => x"08811183",
1695 => x"b93d0c81",
1696 => x"11515a5c",
1697 => x"7887240b",
1698 => x"0b0b81f7",
1699 => x"3883be3d",
1700 => x"e8057c0c",
1701 => x"6c841d0c",
1702 => x"83b73d08",
1703 => x"6d0583b8",
1704 => x"3d0c881c",
1705 => x"83b73d08",
1706 => x"811183b9",
1707 => x"3d0c8111",
1708 => x"515a5c87",
1709 => x"79250b0b",
1710 => x"0be98838",
1711 => x"83be3ddc",
1712 => x"05520b0b",
1713 => x"0bef8d39",
1714 => x"83be3ddc",
1715 => x"05526651",
1716 => x"0b0b0bdf",
1717 => x"ac3f8008",
1718 => x"0b0b0bef",
1719 => x"a73865a5",
1720 => x"3d085c5c",
1721 => x"80598079",
1722 => x"545483ba",
1723 => x"3d0883bc",
1724 => x"3d085b51",
1725 => x"79520b0b",
1726 => x"81ff823f",
1727 => x"80080b0b",
1728 => x"0bfedd38",
1729 => x"ff1b5a80",
1730 => x"7a250b0b",
1731 => x"0bfefe38",
1732 => x"907a250b",
1733 => x"0b0b0bbd",
1734 => x"380b0b82",
1735 => x"edb47c0c",
1736 => x"900b841d",
1737 => x"0c83b73d",
1738 => x"08900583",
1739 => x"b83d0c88",
1740 => x"1c83b73d",
1741 => x"08811183",
1742 => x"b93d0c81",
1743 => x"11515a5c",
1744 => x"7887240b",
1745 => x"0b0b84c4",
1746 => x"38f01a5a",
1747 => x"7990240b",
1748 => x"0b0b0bc5",
1749 => x"380b0b82",
1750 => x"edb47c0c",
1751 => x"79841d0c",
1752 => x"83b73d08",
1753 => x"1a83b83d",
1754 => x"0c881c83",
1755 => x"b73d0881",
1756 => x"1183b93d",
1757 => x"0c811151",
1758 => x"5a5c8779",
1759 => x"250b0b0b",
1760 => x"fe8b3883",
1761 => x"be3ddc05",
1762 => x"5266510b",
1763 => x"0b0bddf1",
1764 => x"3f80080b",
1765 => x"0b0bedec",
1766 => x"386583bf",
1767 => x"3de80571",
1768 => x"0c6d8412",
1769 => x"0c83b83d",
1770 => x"086e0583",
1771 => x"b93d0c5c",
1772 => x"0b0b0bfd",
1773 => x"ed396281",
1774 => x"0659780b",
1775 => x"0b0bfcbb",
1776 => x"387d7c0c",
1777 => x"810b841d",
1778 => x"0c83b73d",
1779 => x"08810583",
1780 => x"b83d0c88",
1781 => x"1c83b73d",
1782 => x"08811183",
1783 => x"b93d0c81",
1784 => x"11515a5c",
1785 => x"8779250b",
1786 => x"0b0bfda1",
1787 => x"3883be3d",
1788 => x"dc05520b",
1789 => x"0b0bff91",
1790 => x"39646584",
1791 => x"0571085d",
1792 => x"4659815f",
1793 => x"0b0b0be2",
1794 => x"87396465",
1795 => x"84057108",
1796 => x"5d465980",
1797 => x"5f0b0b0b",
1798 => x"e8ba3964",
1799 => x"65840571",
1800 => x"085d4659",
1801 => x"7a80250b",
1802 => x"0b0be8f0",
1803 => x"380b0b0b",
1804 => x"f4c839a5",
1805 => x"3d085a80",
1806 => x"7a250b0b",
1807 => x"0b8bbd38",
1808 => x"a43d085b",
1809 => x"7a7a240b",
1810 => x"0b0b83b5",
1811 => x"387d7c0c",
1812 => x"7a841d0c",
1813 => x"83b73d08",
1814 => x"1b83b83d",
1815 => x"0c881c83",
1816 => x"b73d0881",
1817 => x"1183b93d",
1818 => x"0c811151",
1819 => x"5a5c7887",
1820 => x"240b0b0b",
1821 => x"81e33879",
1822 => x"7b315a80",
1823 => x"7a250b0b",
1824 => x"0b818c38",
1825 => x"907a250b",
1826 => x"0b0b0bbd",
1827 => x"380b0b82",
1828 => x"edb47c0c",
1829 => x"900b841d",
1830 => x"0c83b73d",
1831 => x"08900583",
1832 => x"b83d0c88",
1833 => x"1c83b73d",
1834 => x"08811183",
1835 => x"b93d0c81",
1836 => x"11515a5c",
1837 => x"7887240b",
1838 => x"0b0b80fc",
1839 => x"38f01a5a",
1840 => x"7990240b",
1841 => x"0b0b0bc5",
1842 => x"380b0b82",
1843 => x"edb47c0c",
1844 => x"79841d0c",
1845 => x"83b73d08",
1846 => x"1a83b83d",
1847 => x"0c881c83",
1848 => x"b73d0881",
1849 => x"1183b93d",
1850 => x"0c811151",
1851 => x"5a5c8779",
1852 => x"250b0b0b",
1853 => x"0b993883",
1854 => x"be3ddc05",
1855 => x"5266510b",
1856 => x"0b0bdafd",
1857 => x"3f80080b",
1858 => x"0b0beaf8",
1859 => x"38655c62",
1860 => x"81065978",
1861 => x"802e0b0b",
1862 => x"0be4a838",
1863 => x"0b0b82f0",
1864 => x"f47c0c81",
1865 => x"0b841d0c",
1866 => x"83b73d08",
1867 => x"810583b8",
1868 => x"3d0c0b0b",
1869 => x"0bfaeb39",
1870 => x"83be3ddc",
1871 => x"05526651",
1872 => x"0b0b0bda",
1873 => x"bc3f8008",
1874 => x"0b0b0bea",
1875 => x"b73865f0",
1876 => x"1b5b5c0b",
1877 => x"0b0bfee8",
1878 => x"3983be3d",
1879 => x"dc055266",
1880 => x"510b0b0b",
1881 => x"da9b3f80",
1882 => x"080b0b0b",
1883 => x"ea963865",
1884 => x"a63d08a6",
1885 => x"3d087171",
1886 => x"31525d5b",
1887 => x"5c798024",
1888 => x"0b0b0bfd",
1889 => x"ff380b0b",
1890 => x"0bff8439",
1891 => x"83be3ddc",
1892 => x"05526651",
1893 => x"0b0b0bd9",
1894 => x"e83f8008",
1895 => x"0b0b0be9",
1896 => x"e33865f0",
1897 => x"1b5b5c0b",
1898 => x"0b0bfba0",
1899 => x"39646584",
1900 => x"0571086b",
1901 => x"710c527e",
1902 => x"4046590b",
1903 => x"0b0bdb9a",
1904 => x"397e0b0b",
1905 => x"0bdf9938",
1906 => x"ff1e7bb7",
1907 => x"06b0075b",
1908 => x"5e797e34",
1909 => x"7a832a5b",
1910 => x"7a0b0b0b",
1911 => x"0bea3862",
1912 => x"81065978",
1913 => x"802e0b0b",
1914 => x"0beba338",
1915 => x"79b02e0b",
1916 => x"0b0beb9a",
1917 => x"38ff1e5e",
1918 => x"b07e340b",
1919 => x"0b0bf7dd",
1920 => x"397d7c0c",
1921 => x"79841d0c",
1922 => x"83b73d08",
1923 => x"1a83b83d",
1924 => x"0c881c83",
1925 => x"b73d0881",
1926 => x"1183b93d",
1927 => x"0c811151",
1928 => x"5a5c7887",
1929 => x"240b0b0b",
1930 => x"81a03879",
1931 => x"1e0b0b82",
1932 => x"f0f47d0c",
1933 => x"5e810b84",
1934 => x"1d0c83b7",
1935 => x"3d088105",
1936 => x"83b83d0c",
1937 => x"881c83b7",
1938 => x"3d088111",
1939 => x"83b93d0c",
1940 => x"8111515a",
1941 => x"5c788724",
1942 => x"0b0b0b0b",
1943 => x"b6387d7c",
1944 => x"0ca43d08",
1945 => x"7a317084",
1946 => x"1e0c83b8",
1947 => x"3d080583",
1948 => x"b83d0c88",
1949 => x"1c83b73d",
1950 => x"08811183",
1951 => x"b93d0c81",
1952 => x"11515a5c",
1953 => x"8779250b",
1954 => x"0b0be1b7",
1955 => x"380b0b0b",
1956 => x"e7bc3983",
1957 => x"be3ddc05",
1958 => x"5266510b",
1959 => x"0b0bd7e1",
1960 => x"3f80080b",
1961 => x"0b0be7dc",
1962 => x"3865a63d",
1963 => x"087f720c",
1964 => x"a63d0871",
1965 => x"31708414",
1966 => x"0c83ba3d",
1967 => x"080583ba",
1968 => x"3d0c5b5c",
1969 => x"0b0b0bff",
1970 => x"aa3983be",
1971 => x"3ddc0552",
1972 => x"66510b0b",
1973 => x"0bd7aa3f",
1974 => x"80080b0b",
1975 => x"0be7a538",
1976 => x"65a63d08",
1977 => x"7f110b0b",
1978 => x"82f0f473",
1979 => x"0c405b5c",
1980 => x"810b841d",
1981 => x"0c83b73d",
1982 => x"08810583",
1983 => x"b83d0c88",
1984 => x"1c83b73d",
1985 => x"08811183",
1986 => x"b93d0c81",
1987 => x"11515a5c",
1988 => x"8779250b",
1989 => x"0b0bfec6",
1990 => x"380b0b0b",
1991 => x"fef53983",
1992 => x"ba3d0883",
1993 => x"bc3d085b",
1994 => x"5179520b",
1995 => x"0b8197ea",
1996 => x"3f0b0b82",
1997 => x"f0f85e83",
1998 => x"5f80080b",
1999 => x"0b0bdcb1",
2000 => x"38628280",
2001 => x"0783bb3d",
2002 => x"0883bd3d",
2003 => x"086383c0",
2004 => x"3daa3da5",
2005 => x"3d0c5f45",
2006 => x"415f4383",
2007 => x"0ba13d0c",
2008 => x"7f80e62e",
2009 => x"0b0b0b0b",
2010 => x"b1388008",
2011 => x"5a7f80e5",
2012 => x"2e0b0b0b",
2013 => x"83ea3880",
2014 => x"08597f80",
2015 => x"c52e0b0b",
2016 => x"0b83f038",
2017 => x"79790759",
2018 => x"78802e0b",
2019 => x"0b0b0b85",
2020 => x"38608105",
2021 => x"42820ba1",
2022 => x"3d0c7db3",
2023 => x"3d0c7eb4",
2024 => x"3d0c800b",
2025 => x"b33d0824",
2026 => x"0b0b0b88",
2027 => x"ef38807b",
2028 => x"3483be3d",
2029 => x"f3941159",
2030 => x"f3900557",
2031 => x"6e566155",
2032 => x"6f547d52",
2033 => x"7e536a51",
2034 => x"0b0b0b9b",
2035 => x"b03f8008",
2036 => x"6080e732",
2037 => x"70307072",
2038 => x"079f2a51",
2039 => x"5b5ba13d",
2040 => x"0c7f80c7",
2041 => x"2e0b0b0b",
2042 => x"0b883878",
2043 => x"0b0b0b81",
2044 => x"e4386281",
2045 => x"0659780b",
2046 => x"0b0b81d9",
2047 => x"38a33d08",
2048 => x"5978a13d",
2049 => x"0831a53d",
2050 => x"0c6f6080",
2051 => x"e7327030",
2052 => x"70720780",
2053 => x"256380c7",
2054 => x"32703070",
2055 => x"72078025",
2056 => x"73075354",
2057 => x"5f515c5a",
2058 => x"5e79802e",
2059 => x"0b0b0b86",
2060 => x"f238a53d",
2061 => x"085afc7a",
2062 => x"250b0b0b",
2063 => x"0b8a3860",
2064 => x"7a250b0b",
2065 => x"0b82cc38",
2066 => x"80e5597f",
2067 => x"80e72e0b",
2068 => x"0b0b0b84",
2069 => x"3880c559",
2070 => x"78407f80",
2071 => x"e5240b0b",
2072 => x"0b86ca38",
2073 => x"ff1a70a7",
2074 => x"3d0c83b9",
2075 => x"3d715d43",
2076 => x"5a7f6234",
2077 => x"028ddd05",
2078 => x"5f807a24",
2079 => x"0b0b0b87",
2080 => x"c138ab7f",
2081 => x"34028dde",
2082 => x"05b33d70",
2083 => x"5c425f89",
2084 => x"7b250b0b",
2085 => x"0b818738",
2086 => x"ff1a8a7c",
2087 => x"36b0055a",
2088 => x"5a787a34",
2089 => x"8a7b355b",
2090 => x"7a89240b",
2091 => x"0b0b0be8",
2092 => x"38ff1ab0",
2093 => x"1c5a5a78",
2094 => x"7a347961",
2095 => x"270b0b0b",
2096 => x"80ed3879",
2097 => x"7081055b",
2098 => x"337f7081",
2099 => x"0541340b",
2100 => x"0b0b0be6",
2101 => x"39800862",
2102 => x"055b7f80",
2103 => x"e62e0b0b",
2104 => x"0b819838",
2105 => x"80598079",
2106 => x"54547d51",
2107 => x"7e520b0b",
2108 => x"81f0f63f",
2109 => x"80080b0b",
2110 => x"0b0b8538",
2111 => x"7aa43d0c",
2112 => x"a33d0859",
2113 => x"787b270b",
2114 => x"0b0bfdf5",
2115 => x"38b07934",
2116 => x"a33d0881",
2117 => x"05a43d0c",
2118 => x"0b0b0b0b",
2119 => x"e339b07f",
2120 => x"70810541",
2121 => x"34b01b59",
2122 => x"787f7081",
2123 => x"0541347e",
2124 => x"6231a53d",
2125 => x"08701241",
2126 => x"5a4d8179",
2127 => x"250b0b0b",
2128 => x"81a43881",
2129 => x"1f5f83bc",
2130 => x"3d335978",
2131 => x"802e0b0b",
2132 => x"0bd89e38",
2133 => x"ad0b83be",
2134 => x"3d340b0b",
2135 => x"0bd89239",
2136 => x"810b8008",
2137 => x"5a5a7f80",
2138 => x"c52e0981",
2139 => x"060b0b0b",
2140 => x"fc923881",
2141 => x"590b0b0b",
2142 => x"fc8a3980",
2143 => x"08335978",
2144 => x"b02e0b0b",
2145 => x"0b0bb438",
2146 => x"6e087b05",
2147 => x"5b0b0b0b",
2148 => x"fed23980",
2149 => x"e740a43d",
2150 => x"0859787a",
2151 => x"240b0b0b",
2152 => x"85883879",
2153 => x"6381065a",
2154 => x"5f78802e",
2155 => x"0b0b0bff",
2156 => x"9538811a",
2157 => x"5f0b0b0b",
2158 => x"ff8c3980",
2159 => x"59807954",
2160 => x"547d517e",
2161 => x"520b0b81",
2162 => x"f1b33f80",
2163 => x"08802e0b",
2164 => x"0b0bffb4",
2165 => x"38816231",
2166 => x"70a13d08",
2167 => x"0c7b055b",
2168 => x"0b0b0bfd",
2169 => x"ff396281",
2170 => x"06597880",
2171 => x"2e0b0b0b",
2172 => x"fed43881",
2173 => x"1f5f0b0b",
2174 => x"0bfecb39",
2175 => x"0b0b82f0",
2176 => x"f07c0c81",
2177 => x"0b841d0c",
2178 => x"83b73d08",
2179 => x"810583b8",
2180 => x"3d0c881c",
2181 => x"83b73d08",
2182 => x"811183b9",
2183 => x"3d0c8111",
2184 => x"515a5c78",
2185 => x"87240b0b",
2186 => x"0b829238",
2187 => x"790b0b0b",
2188 => x"0b8c38a4",
2189 => x"3d08802e",
2190 => x"0b0b0bda",
2191 => x"86386b7c",
2192 => x"0c810b84",
2193 => x"1d0c83b7",
2194 => x"3d088105",
2195 => x"83b83d0c",
2196 => x"881c83b7",
2197 => x"3d088111",
2198 => x"83b93d0c",
2199 => x"8111515a",
2200 => x"5c788724",
2201 => x"0b0b0b81",
2202 => x"f6387930",
2203 => x"5a807a25",
2204 => x"0b0b0b81",
2205 => x"8c38907a",
2206 => x"250b0b0b",
2207 => x"0bbd380b",
2208 => x"0b82edb4",
2209 => x"7c0c900b",
2210 => x"841d0c83",
2211 => x"b73d0890",
2212 => x"0583b83d",
2213 => x"0c881c83",
2214 => x"b73d0881",
2215 => x"1183b93d",
2216 => x"0c811151",
2217 => x"5a5c7887",
2218 => x"240b0b0b",
2219 => x"80ee38f0",
2220 => x"1a5a7990",
2221 => x"240b0b0b",
2222 => x"0bc5380b",
2223 => x"0b82edb4",
2224 => x"7c0c7984",
2225 => x"1d0c83b7",
2226 => x"3d081a83",
2227 => x"b83d0c88",
2228 => x"1c83b73d",
2229 => x"08811183",
2230 => x"b93d0c81",
2231 => x"11515a5c",
2232 => x"8779250b",
2233 => x"0b0b0b99",
2234 => x"3883be3d",
2235 => x"dc055266",
2236 => x"510b0b0b",
2237 => x"cf8b3f80",
2238 => x"080b0b0b",
2239 => x"df863865",
2240 => x"5c7d7c0c",
2241 => x"a43d0884",
2242 => x"1d0c83b7",
2243 => x"3d08a53d",
2244 => x"080583b8",
2245 => x"3d0c0b0b",
2246 => x"0bef8739",
2247 => x"83be3ddc",
2248 => x"05526651",
2249 => x"0b0b0bce",
2250 => x"d83f8008",
2251 => x"0b0b0bde",
2252 => x"d33865f0",
2253 => x"1b5b5c0b",
2254 => x"0b0bfef6",
2255 => x"3983be3d",
2256 => x"dc055266",
2257 => x"510b0b0b",
2258 => x"ceb73f80",
2259 => x"080b0b0b",
2260 => x"deb23865",
2261 => x"a63d085b",
2262 => x"5c0b0b0b",
2263 => x"fdce3983",
2264 => x"be3ddc05",
2265 => x"5266510b",
2266 => x"0b0bce95",
2267 => x"3f80080b",
2268 => x"0b0bde90",
2269 => x"3865a63d",
2270 => x"08703051",
2271 => x"5b5c7980",
2272 => x"240b0b0b",
2273 => x"fdf0380b",
2274 => x"0b0bfef5",
2275 => x"3986410b",
2276 => x"0b0be18a",
2277 => x"390b0b82",
2278 => x"f0fc5e86",
2279 => x"5f0b0b0b",
2280 => x"d3cf39a5",
2281 => x"3d085a0b",
2282 => x"0b0bf9ae",
2283 => x"397f80e6",
2284 => x"2e098106",
2285 => x"0b0b0bfb",
2286 => x"dd38807a",
2287 => x"250b0b0b",
2288 => x"81bc3879",
2289 => x"5f600b0b",
2290 => x"0b0b8e38",
2291 => x"62810659",
2292 => x"78802e0b",
2293 => x"0b0bfaee",
2294 => x"38601a81",
2295 => x"055f0b0b",
2296 => x"0bfae339",
2297 => x"83b73d08",
2298 => x"0b0b0b0b",
2299 => x"8d38800b",
2300 => x"83b73d0c",
2301 => x"0b0b0bdd",
2302 => x"8b3983be",
2303 => x"3ddc0552",
2304 => x"66510b0b",
2305 => x"0bccfa3f",
2306 => x"80080b0b",
2307 => x"0bdcf538",
2308 => x"800b83b7",
2309 => x"3d0c0b0b",
2310 => x"0bdce939",
2311 => x"7d810a32",
2312 => x"5ead7b34",
2313 => x"0b0b0bf7",
2314 => x"8839787a",
2315 => x"3182055f",
2316 => x"807a250b",
2317 => x"0b0bfa8e",
2318 => x"3881195f",
2319 => x"0b0b0bfa",
2320 => x"85397930",
2321 => x"5bad7f34",
2322 => x"028dde05",
2323 => x"b33d705c",
2324 => x"425f897b",
2325 => x"250b0b0b",
2326 => x"f9c4380b",
2327 => x"0b0bf8b8",
2328 => x"39646584",
2329 => x"05710843",
2330 => x"46596080",
2331 => x"250b0b0b",
2332 => x"d0a438ff",
2333 => x"7d335b41",
2334 => x"0b0b0bd0",
2335 => x"9c39600b",
2336 => x"0b0b0b90",
2337 => x"38628106",
2338 => x"59815f78",
2339 => x"802e0b0b",
2340 => x"0bf9b338",
2341 => x"6082055f",
2342 => x"0b0b0bf9",
2343 => x"a939fc3d",
2344 => x"0d0b0b82",
2345 => x"f4ec0855",
2346 => x"b8150880",
2347 => x"2e0b0b0b",
2348 => x"0b983878",
2349 => x"54775376",
2350 => x"520b0b82",
2351 => x"f4ec0851",
2352 => x"0b0b0bcb",
2353 => x"f63f863d",
2354 => x"0d047451",
2355 => x"0b0b0bbe",
2356 => x"8e3f7854",
2357 => x"77537652",
2358 => x"0b0b82f4",
2359 => x"ec08510b",
2360 => x"0b0bcbd7",
2361 => x"3f863d0d",
2362 => x"04f63d0d",
2363 => x"7c7e6159",
2364 => x"56588056",
2365 => x"74762e0b",
2366 => x"0b0b0ba3",
2367 => x"3876547e",
2368 => x"53745277",
2369 => x"510b0b0b",
2370 => x"83823f80",
2371 => x"08558008",
2372 => x"ff2e0b0b",
2373 => x"0b0ba938",
2374 => x"74800c8c",
2375 => x"3d0d0476",
2376 => x"5475538c",
2377 => x"3df40552",
2378 => x"77510b0b",
2379 => x"0b82dd3f",
2380 => x"80085580",
2381 => x"08ff2e09",
2382 => x"81060b0b",
2383 => x"0b0bd938",
2384 => x"80770c81",
2385 => x"8a780c74",
2386 => x"800c8c3d",
2387 => x"0d047070",
2388 => x"70707754",
2389 => x"76537552",
2390 => x"0b0b82f4",
2391 => x"ec08510b",
2392 => x"0b0bff85",
2393 => x"3f505050",
2394 => x"5004ec3d",
2395 => x"0d66686a",
2396 => x"6c6e735c",
2397 => x"405d4242",
2398 => x"4260802e",
2399 => x"0b0b0b81",
2400 => x"b2388060",
2401 => x"085a5d7c",
2402 => x"7a270b0b",
2403 => x"0b819b38",
2404 => x"933d5b7b",
2405 => x"08841d08",
2406 => x"7d567a08",
2407 => x"557c5463",
2408 => x"53405e0b",
2409 => x"0b0bfec1",
2410 => x"3f800858",
2411 => x"8008ff2e",
2412 => x"0b0b0b81",
2413 => x"9538807a",
2414 => x"80083156",
2415 => x"567c7526",
2416 => x"0b0b0b0b",
2417 => x"83388156",
2418 => x"80087a27",
2419 => x"0b0b0b80",
2420 => x"ea387580",
2421 => x"2e0b0b0b",
2422 => x"80e13880",
2423 => x"081d5d60",
2424 => x"802e0b0b",
2425 => x"0b0baa38",
2426 => x"80567580",
2427 => x"08250b0b",
2428 => x"0b0b9838",
2429 => x"751b5574",
2430 => x"33777081",
2431 => x"05593481",
2432 => x"16567776",
2433 => x"240b0b0b",
2434 => x"0bea387f",
2435 => x"08840560",
2436 => x"0c787084",
2437 => x"055a0855",
2438 => x"74802e0b",
2439 => x"0b0b0bb9",
2440 => x"38797d26",
2441 => x"0b0b0bfe",
2442 => x"ea387c55",
2443 => x"74800c96",
2444 => x"3d0d04ff",
2445 => x"5a0b0b0b",
2446 => x"fec8397d",
2447 => x"7c0c7e84",
2448 => x"1d0c7c55",
2449 => x"0b0b0b0b",
2450 => x"e339818a",
2451 => x"620c807c",
2452 => x"0c800880",
2453 => x"0c963d0d",
2454 => x"0460802e",
2455 => x"0b0b0b0b",
2456 => x"84387460",
2457 => x"0c747c0c",
2458 => x"ff1d800c",
2459 => x"963d0d04",
2460 => x"fc3d0d79",
2461 => x"55785477",
2462 => x"5376520b",
2463 => x"0b82f4ec",
2464 => x"08510b0b",
2465 => x"0bfde33f",
2466 => x"863d0d04",
2467 => x"f83d0d7b",
2468 => x"7d7f0b0b",
2469 => x"82fbec54",
2470 => x"5957550b",
2471 => x"0b818dfb",
2472 => x"3f800881",
2473 => x"260b0b0b",
2474 => x"0b983874",
2475 => x"5474802e",
2476 => x"0b0b0b0b",
2477 => x"86387575",
2478 => x"34815473",
2479 => x"800c8a3d",
2480 => x"0d040b0b",
2481 => x"82f18452",
2482 => x"0b0b82fb",
2483 => x"ec510b0b",
2484 => x"818c953f",
2485 => x"80080b0b",
2486 => x"0b81d838",
2487 => x"80085474",
2488 => x"802e0b0b",
2489 => x"0b0bd438",
2490 => x"80ff7625",
2491 => x"0b0b0b0b",
2492 => x"c538ff80",
2493 => x"16538eff",
2494 => x"73270b0b",
2495 => x"0b85e338",
2496 => x"f0801653",
2497 => x"83efff73",
2498 => x"270b0b0b",
2499 => x"82d838fc",
2500 => x"80801653",
2501 => x"80fbffff",
2502 => x"73270b0b",
2503 => x"0b85e838",
2504 => x"8fff0a16",
2505 => x"53f7c00a",
2506 => x"73270b0b",
2507 => x"0b86a638",
2508 => x"ff54c00a",
2509 => x"76250b0b",
2510 => x"0bff8038",
2511 => x"75820a06",
2512 => x"709e2c70",
2513 => x"fc075151",
2514 => x"53727570",
2515 => x"81055734",
2516 => x"7581fc0a",
2517 => x"0670982a",
2518 => x"ff800751",
2519 => x"53727570",
2520 => x"81055734",
2521 => x"7587f080",
2522 => x"80067092",
2523 => x"2aff8007",
2524 => x"51537275",
2525 => x"70810557",
2526 => x"34758fe0",
2527 => x"8006708c",
2528 => x"2aff8007",
2529 => x"51537275",
2530 => x"70810557",
2531 => x"34759fc0",
2532 => x"0670862a",
2533 => x"ff800751",
2534 => x"53727570",
2535 => x"81055734",
2536 => x"75ffbf06",
2537 => x"ff800753",
2538 => x"72753486",
2539 => x"0b800c8a",
2540 => x"3d0d040b",
2541 => x"0b82f18c",
2542 => x"520b0b82",
2543 => x"fbec510b",
2544 => x"0b818aa4",
2545 => x"3f80080b",
2546 => x"0b0b81f7",
2547 => x"387581ff",
2548 => x"0676882c",
2549 => x"7081ff06",
2550 => x"80085759",
2551 => x"54587480",
2552 => x"2e0b0b0b",
2553 => x"fdd53876",
2554 => x"802e0b0b",
2555 => x"0bfdbc38",
2556 => x"800880ff",
2557 => x"187081ff",
2558 => x"06515456",
2559 => x"729e260b",
2560 => x"0b0b0b83",
2561 => x"38815680",
2562 => x"08a01870",
2563 => x"81ff0651",
2564 => x"5454728f",
2565 => x"260b0b0b",
2566 => x"0b833881",
2567 => x"54757407",
2568 => x"5372802e",
2569 => x"0b0b0b0b",
2570 => x"b5388008",
2571 => x"c0195456",
2572 => x"72be260b",
2573 => x"0b0b0b83",
2574 => x"38815680",
2575 => x"08ff8019",
2576 => x"7081ff06",
2577 => x"51545472",
2578 => x"80fc260b",
2579 => x"0b0b0b83",
2580 => x"38815475",
2581 => x"74075372",
2582 => x"0b0b0b80",
2583 => x"d338ff0b",
2584 => x"800c8a3d",
2585 => x"0d04fcd0",
2586 => x"801653ff",
2587 => x"548fff73",
2588 => x"270b0b0b",
2589 => x"fcc53875",
2590 => x"83e08006",
2591 => x"708c2ae0",
2592 => x"07515372",
2593 => x"75708105",
2594 => x"5734759f",
2595 => x"c0067086",
2596 => x"2aff8007",
2597 => x"51537275",
2598 => x"70810557",
2599 => x"3475ffbf",
2600 => x"06ff8007",
2601 => x"53727534",
2602 => x"830b800c",
2603 => x"8a3d0d04",
2604 => x"76757081",
2605 => x"05573477",
2606 => x"75348254",
2607 => x"73800c8a",
2608 => x"3d0d040b",
2609 => x"0b82f194",
2610 => x"520b0b82",
2611 => x"fbec510b",
2612 => x"0b818894",
2613 => x"3f80080b",
2614 => x"0b0b80f8",
2615 => x"387581ff",
2616 => x"0676882c",
2617 => x"7081ff06",
2618 => x"80085759",
2619 => x"54587480",
2620 => x"2e0b0b0b",
2621 => x"fbc53876",
2622 => x"802e0b0b",
2623 => x"0bfbac38",
2624 => x"80085381",
2625 => x"a077270b",
2626 => x"0b0b0b83",
2627 => x"38815376",
2628 => x"81ff2e0b",
2629 => x"0b0bfec6",
2630 => x"38817074",
2631 => x"06545472",
2632 => x"802e0b0b",
2633 => x"0bfeb738",
2634 => x"80085381",
2635 => x"a078270b",
2636 => x"0b0b0b83",
2637 => x"38735377",
2638 => x"81ff2e0b",
2639 => x"0b0bfe9e",
2640 => x"38727406",
2641 => x"5372802e",
2642 => x"0b0b0bfe",
2643 => x"91380b0b",
2644 => x"0bfedd39",
2645 => x"0b0b82f1",
2646 => x"9c520b0b",
2647 => x"82fbec51",
2648 => x"0b0b8187",
2649 => x"833f8008",
2650 => x"0b0b0bfa",
2651 => x"be388008",
2652 => x"7681ff06",
2653 => x"77882c70",
2654 => x"81ff0659",
2655 => x"55595981",
2656 => x"5474802e",
2657 => x"0b0b0bfa",
2658 => x"b2387580",
2659 => x"2e0b0b0b",
2660 => x"82a538df",
2661 => x"16537280",
2662 => x"dd260b0b",
2663 => x"0bfdbf38",
2664 => x"df185372",
2665 => x"80dd260b",
2666 => x"0b0bfdb2",
2667 => x"3876080b",
2668 => x"0b0b0b9c",
2669 => x"3873770c",
2670 => x"9b757081",
2671 => x"055734a4",
2672 => x"75708105",
2673 => x"573480c2",
2674 => x"75708105",
2675 => x"57348359",
2676 => x"75757081",
2677 => x"05573477",
2678 => x"75348219",
2679 => x"800c8a3d",
2680 => x"0d04758f",
2681 => x"c0067086",
2682 => x"2ac00751",
2683 => x"53727570",
2684 => x"81055734",
2685 => x"75ffbf06",
2686 => x"ff800753",
2687 => x"72753482",
2688 => x"540b0b0b",
2689 => x"fdb63975",
2690 => x"80f08080",
2691 => x"0670922a",
2692 => x"f0075153",
2693 => x"72757081",
2694 => x"05573475",
2695 => x"8fe08006",
2696 => x"708c2aff",
2697 => x"80075153",
2698 => x"72757081",
2699 => x"05573475",
2700 => x"9fc00670",
2701 => x"862aff80",
2702 => x"07515372",
2703 => x"75708105",
2704 => x"573475ff",
2705 => x"bf06ff80",
2706 => x"07537275",
2707 => x"34840b80",
2708 => x"0c8a3d0d",
2709 => x"047581c0",
2710 => x"0a067098",
2711 => x"2af80751",
2712 => x"53727570",
2713 => x"81055734",
2714 => x"7587f080",
2715 => x"80067092",
2716 => x"2aff8007",
2717 => x"51537275",
2718 => x"70810557",
2719 => x"34758fe0",
2720 => x"8006708c",
2721 => x"2aff8007",
2722 => x"51537275",
2723 => x"70810557",
2724 => x"34759fc0",
2725 => x"0670862a",
2726 => x"ff800751",
2727 => x"53727570",
2728 => x"81055734",
2729 => x"75ffbf06",
2730 => x"ff800753",
2731 => x"72753485",
2732 => x"0b800c8a",
2733 => x"3d0d0476",
2734 => x"08802e0b",
2735 => x"0b0b0b9d",
2736 => x"38800877",
2737 => x"0c9b7570",
2738 => x"81055734",
2739 => x"a8757081",
2740 => x"05573480",
2741 => x"c2757081",
2742 => x"05573483",
2743 => x"59777534",
2744 => x"8119800c",
2745 => x"8a3d0d04",
2746 => x"fa3d0d78",
2747 => x"0b0b82f4",
2748 => x"ec085455",
2749 => x"b8130880",
2750 => x"2e0b0b0b",
2751 => x"81dc388c",
2752 => x"15227083",
2753 => x"ffff0670",
2754 => x"832a8132",
2755 => x"70810651",
2756 => x"55555672",
2757 => x"802e0b0b",
2758 => x"0b80f038",
2759 => x"73842a81",
2760 => x"32810657",
2761 => x"ff53760b",
2762 => x"0b0b8193",
2763 => x"3873822a",
2764 => x"70810651",
2765 => x"5372802e",
2766 => x"0b0b0b80",
2767 => x"c638b015",
2768 => x"08547380",
2769 => x"2e0b0b0b",
2770 => x"0ba53880",
2771 => x"c0155373",
2772 => x"732e0b0b",
2773 => x"0b0b9438",
2774 => x"73520b0b",
2775 => x"82f4ec08",
2776 => x"510b0b0b",
2777 => x"b5d23f8c",
2778 => x"15225676",
2779 => x"b0160c75",
2780 => x"db065372",
2781 => x"8c162380",
2782 => x"0b84160c",
2783 => x"90150875",
2784 => x"0c725675",
2785 => x"88075372",
2786 => x"8c162390",
2787 => x"1508802e",
2788 => x"0b0b0b80",
2789 => x"d3388c15",
2790 => x"22708106",
2791 => x"5553730b",
2792 => x"0b0b0ba2",
2793 => x"38720a10",
2794 => x"0a708106",
2795 => x"5153720b",
2796 => x"0b0b0b85",
2797 => x"38941508",
2798 => x"54738816",
2799 => x"0c805372",
2800 => x"800c883d",
2801 => x"0d04800b",
2802 => x"88160c94",
2803 => x"15083098",
2804 => x"160c8053",
2805 => x"0b0b0b0b",
2806 => x"e6397251",
2807 => x"0b0b0baf",
2808 => x"fe3f0b0b",
2809 => x"0bfe9839",
2810 => x"74510b0b",
2811 => x"80c4ef3f",
2812 => x"8c152270",
2813 => x"81065553",
2814 => x"73802e0b",
2815 => x"0b0bffa5",
2816 => x"380b0b0b",
2817 => x"0bc039ef",
2818 => x"3d0d6365",
2819 => x"9011085e",
2820 => x"40408053",
2821 => x"7b609005",
2822 => x"08240b0b",
2823 => x"0b81d038",
2824 => x"941f70ff",
2825 => x"1e70822b",
2826 => x"73116494",
2827 => x"05705c43",
2828 => x"5f610570",
2829 => x"087f0881",
2830 => x"0557555c",
2831 => x"5e42570b",
2832 => x"0b81ebf8",
2833 => x"3f80085d",
2834 => x"80080b0b",
2835 => x"0b81a738",
2836 => x"7e527f51",
2837 => x"0b0b80e9",
2838 => x"803f800b",
2839 => x"8008240b",
2840 => x"0b0b8189",
2841 => x"38811d5d",
2842 => x"80707f63",
2843 => x"5a585b58",
2844 => x"76708405",
2845 => x"58087083",
2846 => x"ffff067b",
2847 => x"0571902a",
2848 => x"71902a05",
2849 => x"70902a5d",
2850 => x"5283ffff",
2851 => x"06821822",
2852 => x"7072311b",
2853 => x"585b5483",
2854 => x"ffff0676",
2855 => x"22707231",
2856 => x"77902c05",
2857 => x"70902c5b",
2858 => x"52435372",
2859 => x"76237482",
2860 => x"17238416",
2861 => x"567a7727",
2862 => x"0b0b0bff",
2863 => x"b3387b10",
2864 => x"101e5978",
2865 => x"080b0b0b",
2866 => x"0ba338fc",
2867 => x"19597d79",
2868 => x"270b0b0b",
2869 => x"0b923878",
2870 => x"080b0b0b",
2871 => x"0b8a38ff",
2872 => x"1c5c0b0b",
2873 => x"0b0be439",
2874 => x"7b609005",
2875 => x"0c7c5372",
2876 => x"800c933d",
2877 => x"0d048070",
2878 => x"5b587670",
2879 => x"84055808",
2880 => x"7083ffff",
2881 => x"06707f29",
2882 => x"1c72902a",
2883 => x"60297190",
2884 => x"2a057090",
2885 => x"2a5e5283",
2886 => x"ffff0682",
2887 => x"19227072",
2888 => x"311c5945",
2889 => x"5283ffff",
2890 => x"06772270",
2891 => x"72317890",
2892 => x"2c057090",
2893 => x"2c5c5256",
2894 => x"51537276",
2895 => x"23748217",
2896 => x"23841656",
2897 => x"7a77270b",
2898 => x"0b0bffae",
2899 => x"3878080b",
2900 => x"0b0bfdfc",
2901 => x"38fc1959",
2902 => x"7d79270b",
2903 => x"0b0b0b92",
2904 => x"3878080b",
2905 => x"0b0b0b8a",
2906 => x"38ff1c5c",
2907 => x"0b0b0b0b",
2908 => x"e4397b60",
2909 => x"90050c0b",
2910 => x"0b0bfdd4",
2911 => x"398c08c8",
2912 => x"3d0dbc3d",
2913 => x"0880c03d",
2914 => x"0880c23d",
2915 => x"0880c53d",
2916 => x"0880c73d",
2917 => x"088c0c5d",
2918 => x"4b434080",
2919 => x"0bbe3d08",
2920 => x"80c03d08",
2921 => x"5bba3d0c",
2922 => x"79bb3d0c",
2923 => x"6080c005",
2924 => x"08574875",
2925 => x"682e0981",
2926 => x"060b0b0b",
2927 => x"80ea38b8",
2928 => x"3d085780",
2929 => x"77240b0b",
2930 => x"0b818c38",
2931 => x"677a0c76",
2932 => x"9ffe0a06",
2933 => x"56759ffe",
2934 => x"0a2e0b0b",
2935 => x"0b819838",
2936 => x"b83d08ba",
2937 => x"3d085a58",
2938 => x"80568076",
2939 => x"54547751",
2940 => x"78520b0b",
2941 => x"81d6f23f",
2942 => x"80080b0b",
2943 => x"0b81c638",
2944 => x"80c13d08",
2945 => x"5881780c",
2946 => x"0b0b82f0",
2947 => x"f05f8c08",
2948 => x"802e0b0b",
2949 => x"0b0b8638",
2950 => x"811f8c08",
2951 => x"0c7e5675",
2952 => x"800cba3d",
2953 => x"0d8c0c04",
2954 => x"7f80c405",
2955 => x"0884170c",
2956 => x"816080c4",
2957 => x"05082b88",
2958 => x"170c7552",
2959 => x"7f510b0b",
2960 => x"80d8ad3f",
2961 => x"676080c0",
2962 => x"050cb83d",
2963 => x"08577680",
2964 => x"250b0b0b",
2965 => x"fef63881",
2966 => x"7a0c76fe",
2967 => x"0a0670ba",
2968 => x"3d0c709f",
2969 => x"fe0a0657",
2970 => x"57759ffe",
2971 => x"0a2e0981",
2972 => x"060b0b0b",
2973 => x"feea3880",
2974 => x"c13d0856",
2975 => x"80ce8f76",
2976 => x"0cb93d08",
2977 => x"0b0b0b84",
2978 => x"c93876bf",
2979 => x"ffff060b",
2980 => x"0b82f1a4",
2981 => x"4056750b",
2982 => x"0b0b84b6",
2983 => x"388c0880",
2984 => x"2e0b0b0b",
2985 => x"fef73883",
2986 => x"1f337f88",
2987 => x"05585675",
2988 => x"0b0b0b0b",
2989 => x"8438831f",
2990 => x"57768c08",
2991 => x"0c7e560b",
2992 => x"0b0bfedb",
2993 => x"39ba3dff",
2994 => x"b41156ff",
2995 => x"b0055477",
2996 => x"5278537f",
2997 => x"510b0b80",
2998 => x"eaa43f80",
2999 => x"08b93d08",
3000 => x"70942a8f",
3001 => x"ff065e59",
3002 => x"417b0b0b",
3003 => x"0b83ef38",
3004 => x"a73d08a7",
3005 => x"3d080588",
3006 => x"b2115d56",
3007 => x"a07c250b",
3008 => x"0b0b8ff4",
3009 => x"3880c07c",
3010 => x"31889217",
3011 => x"79722bbc",
3012 => x"3d08722a",
3013 => x"07b53d71",
3014 => x"5670555d",
3015 => x"5157570b",
3016 => x"0b81dfa9",
3017 => x"3fb23d08",
3018 => x"b43d08b2",
3019 => x"3d5d5a58",
3020 => x"8076240b",
3021 => x"0b0b93f5",
3022 => x"3877b73d",
3023 => x"0c78b83d",
3024 => x"0cb63d08",
3025 => x"90ff0a05",
3026 => x"b73d0cf7",
3027 => x"cd1c5c81",
3028 => x"4ebffc0a",
3029 => x"56807655",
3030 => x"55b63d08",
3031 => x"b83d0858",
3032 => x"5276537a",
3033 => x"510b0b81",
3034 => x"a2803f83",
3035 => x"feca8fa7",
3036 => x"56869bbd",
3037 => x"86e17655",
3038 => x"55b03d08",
3039 => x"b23d0858",
3040 => x"52765379",
3041 => x"510b0b81",
3042 => x"a3933f83",
3043 => x"fe9a94a8",
3044 => x"56f8db83",
3045 => x"91b37655",
3046 => x"55b23d08",
3047 => x"b43d0858",
3048 => x"527653ba",
3049 => x"3dd00551",
3050 => x"0b0b81a0",
3051 => x"963fae3d",
3052 => x"08b03d08",
3053 => x"7d54ae3d",
3054 => x"535a580b",
3055 => x"0b81de8d",
3056 => x"3faa3d4c",
3057 => x"83fecd88",
3058 => x"93568584",
3059 => x"fdf3fb76",
3060 => x"5555ac3d",
3061 => x"08ae3d08",
3062 => x"58527653",
3063 => x"6b510b0b",
3064 => x"81a2ba3f",
3065 => x"a83dab3d",
3066 => x"08ad3d08",
3067 => x"59557756",
3068 => x"78537954",
3069 => x"7052450b",
3070 => x"0b819fc7",
3071 => x"3fa83d08",
3072 => x"aa3d0871",
3073 => x"5370545f",
3074 => x"5d0b0b81",
3075 => x"dfdf3f80",
3076 => x"08438056",
3077 => x"80765454",
3078 => x"7c517d52",
3079 => x"0b0b81d9",
3080 => x"843f800b",
3081 => x"8008240b",
3082 => x"0b0b8eae",
3083 => x"38810ba2",
3084 => x"3d0c6296",
3085 => x"260b0b0b",
3086 => x"0bb23862",
3087 => x"1010100b",
3088 => x"0b82f2d8",
3089 => x"05841108",
3090 => x"71085555",
3091 => x"b93d08bb",
3092 => x"3d085952",
3093 => x"5676520b",
3094 => x"0b81d8c9",
3095 => x"3f800b80",
3096 => x"08246371",
3097 => x"31445680",
3098 => x"0ba23d0c",
3099 => x"a73d087c",
3100 => x"31ff055a",
3101 => x"807a454b",
3102 => x"6a7a240b",
3103 => x"0b0b8da9",
3104 => x"38806324",
3105 => x"0b0b0ba0",
3106 => x"8b38800b",
3107 => x"a63d0c62",
3108 => x"4f636305",
3109 => x"44896227",
3110 => x"0b0b0b0b",
3111 => x"83388042",
3112 => x"81588562",
3113 => x"250b0b0b",
3114 => x"0b873861",
3115 => x"fc054280",
3116 => x"58810ba1",
3117 => x"3d0cff70",
3118 => x"a53d0c46",
3119 => x"6185260b",
3120 => x"0b0b82bd",
3121 => x"38611010",
3122 => x"0b0b82f1",
3123 => x"b0055675",
3124 => x"08040b0b",
3125 => x"82f0f85f",
3126 => x"0b0b0bfb",
3127 => x"c039b83d",
3128 => x"08ba3d08",
3129 => x"58b73d0c",
3130 => x"76b83d0c",
3131 => x"b63d08fc",
3132 => x"0a069ffc",
3133 => x"0a07b73d",
3134 => x"0cf8811c",
3135 => x"5c804eb2",
3136 => x"3db13d5c",
3137 => x"5abffc0a",
3138 => x"56807655",
3139 => x"55b63d08",
3140 => x"b83d0858",
3141 => x"5276537a",
3142 => x"510b0b81",
3143 => x"9ecc3f83",
3144 => x"feca8fa7",
3145 => x"56869bbd",
3146 => x"86e17655",
3147 => x"55b03d08",
3148 => x"b23d0858",
3149 => x"52765379",
3150 => x"510b0b81",
3151 => x"9fdf3f83",
3152 => x"fe9a94a8",
3153 => x"56f8db83",
3154 => x"91b37655",
3155 => x"55b23d08",
3156 => x"b43d0858",
3157 => x"527653ba",
3158 => x"3dd00551",
3159 => x"0b0b819c",
3160 => x"e23fae3d",
3161 => x"08b03d08",
3162 => x"7d54ae3d",
3163 => x"535a580b",
3164 => x"0b81dad9",
3165 => x"3faa3d4c",
3166 => x"83fecd88",
3167 => x"93568584",
3168 => x"fdf3fb76",
3169 => x"5555ac3d",
3170 => x"08ae3d08",
3171 => x"58527653",
3172 => x"6b510b0b",
3173 => x"819f863f",
3174 => x"a83dab3d",
3175 => x"08ad3d08",
3176 => x"59557756",
3177 => x"78537954",
3178 => x"7052450b",
3179 => x"0b819c93",
3180 => x"3fa83d08",
3181 => x"aa3d0871",
3182 => x"5370545f",
3183 => x"5d0b0b81",
3184 => x"dcab3f80",
3185 => x"08438056",
3186 => x"80765454",
3187 => x"7c517d52",
3188 => x"0b0b81d5",
3189 => x"d03f8008",
3190 => x"80250b0b",
3191 => x"0bfcce38",
3192 => x"0b0b0b8a",
3193 => x"f539800b",
3194 => x"a13d0c68",
3195 => x"63058111",
3196 => x"70485da4",
3197 => x"3d0c7b80",
3198 => x"240b0b0b",
3199 => x"0b833881",
3200 => x"5c845a80",
3201 => x"6080c405",
3202 => x"0c987c26",
3203 => x"0b0b0b0b",
3204 => x"9b388057",
3205 => x"81177a10",
3206 => x"9411585b",
3207 => x"577b7627",
3208 => x"0b0b0b0b",
3209 => x"ef387660",
3210 => x"80c4050c",
3211 => x"7f80c405",
3212 => x"08527f51",
3213 => x"0b0b80cf",
3214 => x"903f8008",
3215 => x"6080c005",
3216 => x"0c800880",
3217 => x"088e6827",
3218 => x"58404d77",
3219 => x"802e0b0b",
3220 => x"0b86fd38",
3221 => x"75802e0b",
3222 => x"0b0b86f4",
3223 => x"38b83d08",
3224 => x"ba3d0871",
3225 => x"b93d0c70",
3226 => x"ba3d0c64",
3227 => x"a53d0c67",
3228 => x"a73d0c5a",
3229 => x"58825c80",
3230 => x"63250b0b",
3231 => x"0b8cae38",
3232 => x"62832b80",
3233 => x"f8060b0b",
3234 => x"82f2d811",
3235 => x"080b0b82",
3236 => x"f2dc1208",
3237 => x"65842c70",
3238 => x"842a7081",
3239 => x"0651545d",
3240 => x"405e5675",
3241 => x"0b0b0b8a",
3242 => x"8a387980",
3243 => x"2e0b0b0b",
3244 => x"0ba8380b",
3245 => x"0b82f2b0",
3246 => x"58798106",
3247 => x"56750b0b",
3248 => x"0b88f138",
3249 => x"79812c88",
3250 => x"19595a79",
3251 => x"0b0b0b0b",
3252 => x"e838b83d",
3253 => x"08ba3d08",
3254 => x"5a587c54",
3255 => x"7d557752",
3256 => x"78536451",
3257 => x"0b0b81bb",
3258 => x"b43fa83d",
3259 => x"08aa3d08",
3260 => x"71bb3d0c",
3261 => x"70bc3d0c",
3262 => x"5a58a13d",
3263 => x"08802e0b",
3264 => x"0b0b80eb",
3265 => x"38805a9f",
3266 => x"fc0a5680",
3267 => x"76545477",
3268 => x"5178520b",
3269 => x"0b81d38d",
3270 => x"3f798008",
3271 => x"240b0b0b",
3272 => x"8def3880",
3273 => x"66250b0b",
3274 => x"0b80c438",
3275 => x"79802e0b",
3276 => x"0b0b0bbb",
3277 => x"38800ba4",
3278 => x"3d08250b",
3279 => x"0b0b84f8",
3280 => x"38a33d08",
3281 => x"63ff0544",
3282 => x"4680c882",
3283 => x"0a568076",
3284 => x"55557752",
3285 => x"78536451",
3286 => x"0b0b819b",
3287 => x"c03fa83d",
3288 => x"08aa3d08",
3289 => x"5ab93d0c",
3290 => x"78ba3d0c",
3291 => x"811c5c7b",
3292 => x"5264510b",
3293 => x"0b81d6d5",
3294 => x"3fb83d08",
3295 => x"ba3d0858",
3296 => x"547655a8",
3297 => x"3d08aa3d",
3298 => x"08585276",
3299 => x"536b510b",
3300 => x"0b819b89",
3301 => x"3f80f082",
3302 => x"0a568076",
3303 => x"5555aa3d",
3304 => x"08ac3d08",
3305 => x"58527653",
3306 => x"ac3d510b",
3307 => x"0b819893",
3308 => x"3fac3d08",
3309 => x"ae3d0858",
3310 => x"b53d0c76",
3311 => x"b63d0cb4",
3312 => x"3d0886bf",
3313 => x"0a05b53d",
3314 => x"0c65802e",
3315 => x"0b0b0b9b",
3316 => x"c9386f80",
3317 => x"2e0b0b0b",
3318 => x"99e23865",
3319 => x"1010100b",
3320 => x"0b82f2d0",
3321 => x"05841108",
3322 => x"71085656",
3323 => x"568ffc0a",
3324 => x"56807653",
3325 => x"5364510b",
3326 => x"0b81b9a1",
3327 => x"3fb43d08",
3328 => x"b63d0858",
3329 => x"547655a8",
3330 => x"3d08aa3d",
3331 => x"08585276",
3332 => x"536b510b",
3333 => x"0b8198d2",
3334 => x"3faa3d08",
3335 => x"ac3d0858",
3336 => x"b53d0c76",
3337 => x"b63d0c80",
3338 => x"0bb93d08",
3339 => x"bb3d085b",
3340 => x"595c80c8",
3341 => x"820a5d80",
3342 => x"5e775178",
3343 => x"520b0b81",
3344 => x"d7ab3f80",
3345 => x"08800853",
3346 => x"65525a0b",
3347 => x"0b81d4fd",
3348 => x"3fa83d08",
3349 => x"aa3d0858",
3350 => x"547655b8",
3351 => x"3d08ba3d",
3352 => x"08585276",
3353 => x"536b510b",
3354 => x"0b8197fe",
3355 => x"3faa3d08",
3356 => x"ac3d085a",
3357 => x"b93d0c78",
3358 => x"ba3d0cb0",
3359 => x"1a56757f",
3360 => x"70810541",
3361 => x"34b83d08",
3362 => x"ba3d08b6",
3363 => x"3d08b83d",
3364 => x"085a5578",
3365 => x"56715370",
3366 => x"545a580b",
3367 => x"0b81d085",
3368 => x"3f800b80",
3369 => x"08240b0b",
3370 => x"0b87d438",
3371 => x"77547855",
3372 => x"9ffc0a56",
3373 => x"80765353",
3374 => x"64510b0b",
3375 => x"8197ab3f",
3376 => x"b43d08b6",
3377 => x"3d087155",
3378 => x"7056aa3d",
3379 => x"08ac3d08",
3380 => x"5a537854",
3381 => x"5a580b0b",
3382 => x"81cfca3f",
3383 => x"800b8008",
3384 => x"240b0b0b",
3385 => x"86e63881",
3386 => x"1c5c7b66",
3387 => x"250b0b0b",
3388 => x"81c6387c",
3389 => x"547d5577",
3390 => x"5278536b",
3391 => x"510b0b81",
3392 => x"989b3faa",
3393 => x"3d08ac3d",
3394 => x"0858b53d",
3395 => x"0c76b63d",
3396 => x"0c7c547d",
3397 => x"55b83d08",
3398 => x"ba3d0858",
3399 => x"52765364",
3400 => x"510b0b81",
3401 => x"97f73fa8",
3402 => x"3d08aa3d",
3403 => x"0871bb3d",
3404 => x"0c70bc3d",
3405 => x"0c5a580b",
3406 => x"0b0bfdfd",
3407 => x"398ffc0a",
3408 => x"58807855",
3409 => x"7056b53d",
3410 => x"08b73d08",
3411 => x"59537754",
3412 => x"6552590b",
3413 => x"0b8194eb",
3414 => x"3fa83d08",
3415 => x"aa3d0858",
3416 => x"537654b8",
3417 => x"3d08ba3d",
3418 => x"08585176",
3419 => x"520b0b81",
3420 => x"cc9f3f80",
3421 => x"0880240b",
3422 => x"0b0b85d0",
3423 => x"38b43d08",
3424 => x"b63d0858",
3425 => x"54765577",
3426 => x"5278536b",
3427 => x"510b0b81",
3428 => x"95d83faa",
3429 => x"3d08ac3d",
3430 => x"08585376",
3431 => x"54b83d08",
3432 => x"ba3d0858",
3433 => x"5176520b",
3434 => x"0b81cdf9",
3435 => x"3f800b80",
3436 => x"08240b0b",
3437 => x"0b97cb38",
3438 => x"6cb73d08",
3439 => x"b93d085b",
3440 => x"ba3d0c79",
3441 => x"bb3d0ca3",
3442 => x"3d08a63d",
3443 => x"0848445f",
3444 => x"800ba73d",
3445 => x"08575877",
3446 => x"76240b0b",
3447 => x"0b0b8338",
3448 => x"81588078",
3449 => x"0657628e",
3450 => x"240b0b0b",
3451 => x"89ad3881",
3452 => x"70790658",
3453 => x"5976802e",
3454 => x"0b0b0b89",
3455 => x"9e386210",
3456 => x"10100b0b",
3457 => x"82f2d805",
3458 => x"70088412",
3459 => x"08806c24",
3460 => x"53405e56",
3461 => x"8066250b",
3462 => x"0b0b86c9",
3463 => x"38810bb9",
3464 => x"3d08bb3d",
3465 => x"085b595c",
3466 => x"7c547d55",
3467 => x"77527853",
3468 => x"64510b0b",
3469 => x"81b4e63f",
3470 => x"a83d08aa",
3471 => x"3d085851",
3472 => x"76520b0b",
3473 => x"81d3a63f",
3474 => x"80088008",
3475 => x"5365525a",
3476 => x"0b0b81d0",
3477 => x"f83f7c54",
3478 => x"7d55a83d",
3479 => x"08aa3d08",
3480 => x"58527653",
3481 => x"6b510b0b",
3482 => x"8195b23f",
3483 => x"aa3d08ac",
3484 => x"3d085854",
3485 => x"7655b83d",
3486 => x"08ba3d08",
3487 => x"58527653",
3488 => x"ac3d510b",
3489 => x"0b8193e2",
3490 => x"3fac3d08",
3491 => x"ae3d085a",
3492 => x"b93d0c78",
3493 => x"ba3d0cb0",
3494 => x"1a56757f",
3495 => x"70810541",
3496 => x"347b662e",
3497 => x"0b0b0b82",
3498 => x"c23880c8",
3499 => x"820a5680",
3500 => x"765555b8",
3501 => x"3d08ba3d",
3502 => x"08585276",
3503 => x"5364510b",
3504 => x"0b8194d9",
3505 => x"3fa83d08",
3506 => x"aa3d0871",
3507 => x"bb3d0c70",
3508 => x"bc3d0c5a",
3509 => x"58805680",
3510 => x"76545477",
3511 => x"5178520b",
3512 => x"0b81c585",
3513 => x"3f800880",
3514 => x"2e0b0b0b",
3515 => x"83913881",
3516 => x"1c5c0b0b",
3517 => x"0bfeb139",
3518 => x"a07c31ba",
3519 => x"3d08712b",
3520 => x"b43d7155",
3521 => x"70545c51",
3522 => x"560b0b81",
3523 => x"cfbf3fb2",
3524 => x"3d08b43d",
3525 => x"08b23d5d",
3526 => x"5a587580",
3527 => x"250b0b0b",
3528 => x"f097380b",
3529 => x"0b0b8485",
3530 => x"3979304b",
3531 => x"80440b0b",
3532 => x"0bf2ce39",
3533 => x"811c7808",
3534 => x"841a0859",
3535 => x"5577567d",
3536 => x"537e5465",
3537 => x"525c0b0b",
3538 => x"8193d23f",
3539 => x"a83d08aa",
3540 => x"3d085f5d",
3541 => x"0b0b0bf6",
3542 => x"eb396252",
3543 => x"64510b0b",
3544 => x"81ceea3f",
3545 => x"7c537d54",
3546 => x"a83d08aa",
3547 => x"3d085851",
3548 => x"76520b0b",
3549 => x"81c6863f",
3550 => x"80083070",
3551 => x"8008079f",
3552 => x"2a647131",
3553 => x"4551560b",
3554 => x"0b0bf1a1",
3555 => x"39800ba1",
3556 => x"3d0c8069",
3557 => x"250b0b0b",
3558 => x"84e73868",
3559 => x"69a53d0c",
3560 => x"69475c0b",
3561 => x"0b0bf4d9",
3562 => x"39925c80",
3563 => x"490b0b0b",
3564 => x"f4cf3979",
3565 => x"8f060b0b",
3566 => x"82f2d008",
3567 => x"0b0b82f2",
3568 => x"d4085955",
3569 => x"77567853",
3570 => x"79546552",
3571 => x"5a0b0b81",
3572 => x"b1cb3fa8",
3573 => x"3d08aa3d",
3574 => x"0871bb3d",
3575 => x"0c70bc3d",
3576 => x"0c5a5883",
3577 => x"5c0b0b0b",
3578 => x"f5c039b8",
3579 => x"3d08ba3d",
3580 => x"08715670",
3581 => x"57585276",
3582 => x"5364510b",
3583 => x"0b818fc3",
3584 => x"3fa83d08",
3585 => x"aa3d0871",
3586 => x"bb3d0c70",
3587 => x"bc3d0c7e",
3588 => x"557f5671",
3589 => x"5370545a",
3590 => x"580b0b81",
3591 => x"c6f33f80",
3592 => x"0880240b",
3593 => x"0b0b0ba4",
3594 => x"387c537d",
3595 => x"54775178",
3596 => x"520b0b81",
3597 => x"c2b33f80",
3598 => x"080b0b0b",
3599 => x"80c13879",
3600 => x"81065675",
3601 => x"802e0b0b",
3602 => x"0b0bb438",
3603 => x"ff1f7033",
3604 => x"575f75b9",
3605 => x"2e098106",
3606 => x"0b0b0b0b",
3607 => x"94387e6d",
3608 => x"2e098106",
3609 => x"0b0b0b0b",
3610 => x"e3386281",
3611 => x"0543b06d",
3612 => x"347e7f81",
3613 => x"05713381",
3614 => x"05584057",
3615 => x"75773460",
3616 => x"527f510b",
3617 => x"0b80c3e8",
3618 => x"3f807f34",
3619 => x"80c13d08",
3620 => x"63810571",
3621 => x"0c568c08",
3622 => x"802e0b0b",
3623 => x"0b0b8538",
3624 => x"7e8c080c",
3625 => x"6c800cba",
3626 => x"3d0d8c0c",
3627 => x"0462305b",
3628 => x"7a802e0b",
3629 => x"0b0bf4c2",
3630 => x"387a832b",
3631 => x"80f8060b",
3632 => x"0b82f2dc",
3633 => x"11080b0b",
3634 => x"82f2d812",
3635 => x"08565678",
3636 => x"53795465",
3637 => x"52560b0b",
3638 => x"8190c23f",
3639 => x"a83d08aa",
3640 => x"3d0871bb",
3641 => x"3d0c70bc",
3642 => x"3d0c7c84",
3643 => x"2c5c5a58",
3644 => x"79802e0b",
3645 => x"0b0bf482",
3646 => x"380b0b82",
3647 => x"f2b07a81",
3648 => x"06575b75",
3649 => x"0b0b0b82",
3650 => x"90387981",
3651 => x"2c881c5c",
3652 => x"5a79802e",
3653 => x"0b0b0bf3",
3654 => x"e1387981",
3655 => x"06567580",
3656 => x"2e0b0b0b",
3657 => x"0be4380b",
3658 => x"0b0b81ed",
3659 => x"399f820a",
3660 => x"56807655",
3661 => x"55775278",
3662 => x"537a510b",
3663 => x"0b818d83",
3664 => x"3fb03d08",
3665 => x"b23d085a",
3666 => x"b73d0c78",
3667 => x"b83d0cb6",
3668 => x"3d0890ff",
3669 => x"0a05b73d",
3670 => x"0cf7cd1c",
3671 => x"5c814e0b",
3672 => x"0b0bebed",
3673 => x"39757906",
3674 => x"5675802e",
3675 => x"0b0b0bf9",
3676 => x"ac388070",
3677 => x"484a6966",
3678 => x"240b0b0b",
3679 => x"82943880",
3680 => x"d0820a56",
3681 => x"80765555",
3682 => x"7c527d53",
3683 => x"64510b0b",
3684 => x"818f8a3f",
3685 => x"a83d08aa",
3686 => x"3d085853",
3687 => x"7654b83d",
3688 => x"08ba3d08",
3689 => x"58517652",
3690 => x"0b0b81c8",
3691 => x"8c3f6980",
3692 => x"08250b0b",
3693 => x"0b81db38",
3694 => x"6c5fb17f",
3695 => x"70810541",
3696 => x"34628105",
3697 => x"4366527f",
3698 => x"510b0b80",
3699 => x"c1a23f69",
3700 => x"802e0b0b",
3701 => x"0bfda838",
3702 => x"67307069",
3703 => x"079f2a51",
3704 => x"56676a2e",
3705 => x"0b0b0b0b",
3706 => x"8838750b",
3707 => x"0b0b80e5",
3708 => x"3869527f",
3709 => x"510b0b80",
3710 => x"c0f63f0b",
3711 => x"0b0bfcff",
3712 => x"39817071",
3713 => x"a63d0c71",
3714 => x"485d490b",
3715 => x"0b0beff1",
3716 => x"39815a0b",
3717 => x"0b0bf28b",
3718 => x"39811c7b",
3719 => x"08841d08",
3720 => x"59557756",
3721 => x"78537954",
3722 => x"65525c0b",
3723 => x"0b818ded",
3724 => x"3fa83d08",
3725 => x"aa3d0871",
3726 => x"bb3d0c70",
3727 => x"bc3d0c7b",
3728 => x"812c881e",
3729 => x"5e5c5a58",
3730 => x"790b0b0b",
3731 => x"fdcc380b",
3732 => x"0b0bf1a6",
3733 => x"3967527f",
3734 => x"510b0b80",
3735 => x"c0923f69",
3736 => x"527f510b",
3737 => x"0b80c088",
3738 => x"3f0b0b0b",
3739 => x"fc913977",
3740 => x"810a3253",
3741 => x"78547951",
3742 => x"7a520b0b",
3743 => x"81c4a63f",
3744 => x"80088025",
3745 => x"0b0b0bf6",
3746 => x"af3879b9",
3747 => x"3d0c7aba",
3748 => x"3d0c6809",
3749 => x"430b0b0b",
3750 => x"feab396a",
3751 => x"a63d0878",
3752 => x"794b4c59",
3753 => x"596f802e",
3754 => x"0b0b0b80",
3755 => x"d0388162",
3756 => x"250b0b0b",
3757 => x"8ec73865",
3758 => x"ff05a63d",
3759 => x"08713159",
3760 => x"5aa53d08",
3761 => x"7a250b0b",
3762 => x"0b0b9438",
3763 => x"79a63d08",
3764 => x"316f11a1",
3765 => x"3d0ca63d",
3766 => x"0805a63d",
3767 => x"0c765865",
3768 => x"5c806624",
3769 => x"0b0b0b84",
3770 => x"cb386a1c",
3771 => x"641d454b",
3772 => x"81527f51",
3773 => x"0b0b80c4",
3774 => x"de3f8008",
3775 => x"4a788024",
3776 => x"56806425",
3777 => x"0b0b0b0b",
3778 => x"a3387580",
3779 => x"2e0b0b0b",
3780 => x"0b9a3863",
3781 => x"5c786425",
3782 => x"0b0b0b0b",
3783 => x"8338785c",
3784 => x"6a7c3179",
3785 => x"7d31657e",
3786 => x"31465a4b",
3787 => x"800ba63d",
3788 => x"08250b0b",
3789 => x"0b80cb38",
3790 => x"6f802e0b",
3791 => x"0b0b8ae5",
3792 => x"38807825",
3793 => x"0b0b0b0b",
3794 => x"ac387753",
3795 => x"69527f51",
3796 => x"0b0b80c7",
3797 => x"943f8008",
3798 => x"61548008",
3799 => x"5360524a",
3800 => x"0b0b80c4",
3801 => x"8e3f8008",
3802 => x"61536052",
3803 => x"560b0b0b",
3804 => x"bdfe3f75",
3805 => x"41a53d08",
3806 => x"78315a79",
3807 => x"0b0b0b83",
3808 => x"9e388152",
3809 => x"7f510b0b",
3810 => x"80c3cc3f",
3811 => x"80084780",
3812 => x"6f250b0b",
3813 => x"0b0b9138",
3814 => x"6e538008",
3815 => x"527f510b",
3816 => x"0b80c6c5",
3817 => x"3f800847",
3818 => x"80588162",
3819 => x"250b0b0b",
3820 => x"829b3863",
3821 => x"81059f06",
3822 => x"5c6e0b0b",
3823 => x"0b81ee38",
3824 => x"7b802e0b",
3825 => x"0b0b0b85",
3826 => x"38a07c31",
3827 => x"5c847c25",
3828 => x"0b0b0b88",
3829 => x"c238fc1c",
3830 => x"6b11711b",
3831 => x"5b4c6405",
3832 => x"44806b25",
3833 => x"0b0b0b0b",
3834 => x"90386a53",
3835 => x"60527f51",
3836 => x"0b0b80c7",
3837 => x"f23f8008",
3838 => x"41806425",
3839 => x"0b0b0b0b",
3840 => x"90386353",
3841 => x"66527f51",
3842 => x"0b0b80c7",
3843 => x"da3f8008",
3844 => x"47a13d08",
3845 => x"0b0b0b80",
3846 => x"da388066",
3847 => x"25568262",
3848 => x"250b0b0b",
3849 => x"82c73875",
3850 => x"802e0b0b",
3851 => x"0b82be38",
3852 => x"8066240b",
3853 => x"0b0bfcda",
3854 => x"38805485",
3855 => x"5366527f",
3856 => x"510b0b0b",
3857 => x"bcce3f80",
3858 => x"08800853",
3859 => x"6152470b",
3860 => x"0b80c985",
3861 => x"3f800b80",
3862 => x"08250b0b",
3863 => x"0bfcb338",
3864 => x"6c5fb17f",
3865 => x"70810541",
3866 => x"34628105",
3867 => x"430b0b0b",
3868 => x"fad33966",
3869 => x"5260510b",
3870 => x"0b80c8dd",
3871 => x"3f800880",
3872 => x"250b0b0b",
3873 => x"ff943862",
3874 => x"ff054380",
3875 => x"548a5360",
3876 => x"527f510b",
3877 => x"0b0bbbfc",
3878 => x"3f800841",
3879 => x"6f0b0b0b",
3880 => x"81b038a3",
3881 => x"3d08460b",
3882 => x"0b0bfeee",
3883 => x"39669005",
3884 => x"08101067",
3885 => x"05901108",
3886 => x"52560b0b",
3887 => x"0bbec93f",
3888 => x"63800831",
3889 => x"9f065c0b",
3890 => x"0b0bfdf4",
3891 => x"39b93d08",
3892 => x"782e0981",
3893 => x"060b0b0b",
3894 => x"fdd938b8",
3895 => x"3d0870bf",
3896 => x"ffff0657",
3897 => x"5775782e",
3898 => x"0981060b",
3899 => x"0b0bfdc3",
3900 => x"38769ffe",
3901 => x"0a065675",
3902 => x"782e0b0b",
3903 => x"0bfdb438",
3904 => x"6a810564",
3905 => x"8105454b",
3906 => x"81648105",
3907 => x"9f065d58",
3908 => x"6e802e0b",
3909 => x"0b0bfda8",
3910 => x"380b0b0b",
3911 => x"ff8f3979",
3912 => x"5360527f",
3913 => x"510b0b80",
3914 => x"c3bf3f80",
3915 => x"08410b0b",
3916 => x"0bfccf39",
3917 => x"6a663159",
3918 => x"806b114c",
3919 => x"64054481",
3920 => x"527f510b",
3921 => x"0b80c08f",
3922 => x"3f80084a",
3923 => x"0b0b0bfb",
3924 => x"ac398054",
3925 => x"8a536952",
3926 => x"7f510b0b",
3927 => x"0bbab53f",
3928 => x"8008a43d",
3929 => x"08474a0b",
3930 => x"0b0bfdae",
3931 => x"39815c6f",
3932 => x"802e0b0b",
3933 => x"0b82bb38",
3934 => x"8079250b",
3935 => x"0b0b0b90",
3936 => x"38785369",
3937 => x"527f510b",
3938 => x"0b80c4db",
3939 => x"3f80084a",
3940 => x"6948770b",
3941 => x"0b0b82e9",
3942 => x"38815c66",
3943 => x"5260510b",
3944 => x"0b0bdce3",
3945 => x"3f8008b0",
3946 => x"05685361",
3947 => x"52570b0b",
3948 => x"80c6a63f",
3949 => x"80086a54",
3950 => x"67536052",
3951 => x"5a0b0b80",
3952 => x"c6fe3f80",
3953 => x"0856815b",
3954 => x"80088c05",
3955 => x"08802e0b",
3956 => x"0b0b8299",
3957 => x"3875527f",
3958 => x"510b0b0b",
3959 => x"b9923f7a",
3960 => x"62075675",
3961 => x"0b0b0b0b",
3962 => x"9038b93d",
3963 => x"08810656",
3964 => x"75802e0b",
3965 => x"0b0b82c8",
3966 => x"38807a24",
3967 => x"0b0b0b82",
3968 => x"da387962",
3969 => x"0756750b",
3970 => x"0b0b0b90",
3971 => x"38b93d08",
3972 => x"81065675",
3973 => x"802e0b0b",
3974 => x"0b82c038",
3975 => x"7a80240b",
3976 => x"0b0b8883",
3977 => x"38767f70",
3978 => x"81054134",
3979 => x"7b662e0b",
3980 => x"0b0b83fd",
3981 => x"3880548a",
3982 => x"5360527f",
3983 => x"510b0b0b",
3984 => x"b8d23f80",
3985 => x"0841676a",
3986 => x"2e0b0b0b",
3987 => x"83ac3880",
3988 => x"548a5367",
3989 => x"527f510b",
3990 => x"0b0bb8b8",
3991 => x"3f800848",
3992 => x"80548a53",
3993 => x"69527f51",
3994 => x"0b0b0bb8",
3995 => x"a73f8008",
3996 => x"811d5d4a",
3997 => x"66526051",
3998 => x"0b0b0bdb",
3999 => x"8a3f8008",
4000 => x"b0056853",
4001 => x"6152570b",
4002 => x"0b80c4cd",
4003 => x"3f80086a",
4004 => x"54675360",
4005 => x"525a0b0b",
4006 => x"80c5a53f",
4007 => x"80085681",
4008 => x"5b80088c",
4009 => x"05080b0b",
4010 => x"0bfeaa38",
4011 => x"0b0b0b0b",
4012 => x"bc396652",
4013 => x"7e7f8105",
4014 => x"62534056",
4015 => x"0b0b0bda",
4016 => x"c63f8008",
4017 => x"b0055776",
4018 => x"76347b66",
4019 => x"250b0b0b",
4020 => x"82df3880",
4021 => x"548a5360",
4022 => x"527f510b",
4023 => x"0b0bb7b4",
4024 => x"3f800881",
4025 => x"1d5d410b",
4026 => x"0b0b0bc6",
4027 => x"39800852",
4028 => x"60510b0b",
4029 => x"80c3e23f",
4030 => x"80085b0b",
4031 => x"0b0bfdd5",
4032 => x"39698405",
4033 => x"08527f51",
4034 => x"0b0b0bb5",
4035 => x"bc3f8008",
4036 => x"68900508",
4037 => x"10108805",
4038 => x"54688c05",
4039 => x"5380088c",
4040 => x"05524a0b",
4041 => x"0bff94e3",
4042 => x"3f815369",
4043 => x"527f510b",
4044 => x"0b80c1b3",
4045 => x"3f80084a",
4046 => x"815c0b0b",
4047 => x"0bfcdc39",
4048 => x"76b92e0b",
4049 => x"0b0b80d0",
4050 => x"38798024",
4051 => x"1757767f",
4052 => x"70810541",
4053 => x"340b0b0b",
4054 => x"f4eb3980",
4055 => x"7b250b0b",
4056 => x"0b0beb38",
4057 => x"81536052",
4058 => x"7f510b0b",
4059 => x"80c0f83f",
4060 => x"80086753",
4061 => x"80085241",
4062 => x"0b0b80c2",
4063 => x"dc3f800b",
4064 => x"8008250b",
4065 => x"0b0b80c8",
4066 => x"38811757",
4067 => x"76ba2e09",
4068 => x"81060b0b",
4069 => x"0bffb738",
4070 => x"b97f7081",
4071 => x"054134ff",
4072 => x"1f703357",
4073 => x"5f75b92e",
4074 => x"0981060b",
4075 => x"0b0b81d0",
4076 => x"387e6d2e",
4077 => x"0981060b",
4078 => x"0b0b0be3",
4079 => x"38628105",
4080 => x"6d4043b1",
4081 => x"7f708105",
4082 => x"41340b0b",
4083 => x"0bf3f639",
4084 => x"80080b0b",
4085 => x"0bfef738",
4086 => x"76810656",
4087 => x"75802e0b",
4088 => x"0b0bfeea",
4089 => x"38811757",
4090 => x"76ba2e09",
4091 => x"81060b0b",
4092 => x"0bfedb38",
4093 => x"0b0b0bff",
4094 => x"9f398054",
4095 => x"8a536952",
4096 => x"7f510b0b",
4097 => x"0bb58d3f",
4098 => x"80088008",
4099 => x"811e5e49",
4100 => x"4a0b0b0b",
4101 => x"fcde397b",
4102 => x"83240b0b",
4103 => x"0bf7c238",
4104 => x"9c1c6b11",
4105 => x"711b5b4c",
4106 => x"6405440b",
4107 => x"0b0bf7b1",
4108 => x"39815360",
4109 => x"527f510b",
4110 => x"0b0bbfab",
4111 => x"3f800867",
4112 => x"53800852",
4113 => x"410b0b80",
4114 => x"c18f3f80",
4115 => x"0880240b",
4116 => x"0b0bfecb",
4117 => x"3880080b",
4118 => x"0b0b0b8c",
4119 => x"38768106",
4120 => x"56750b0b",
4121 => x"0bfeb838",
4122 => x"ff1f7033",
4123 => x"575f75b0",
4124 => x"2e0b0b0b",
4125 => x"0bf23881",
4126 => x"1f5f0b0b",
4127 => x"0bf2c639",
4128 => x"7e7f8105",
4129 => x"71338105",
4130 => x"58405775",
4131 => x"77340b0b",
4132 => x"0bf2b239",
4133 => x"6a633163",
4134 => x"30a73d0c",
4135 => x"4b804f0b",
4136 => x"0b0bdff1",
4137 => x"39a53d08",
4138 => x"5360527f",
4139 => x"510b0b0b",
4140 => x"bcb73f80",
4141 => x"08410b0b",
4142 => x"0bf5c739",
4143 => x"65101010",
4144 => x"0b0b82f2",
4145 => x"d0058411",
4146 => x"08710856",
4147 => x"56b53d08",
4148 => x"b73d0859",
4149 => x"53567653",
4150 => x"64510b0b",
4151 => x"8180be3f",
4152 => x"a83d08aa",
4153 => x"3d0858b5",
4154 => x"3d0c76b6",
4155 => x"3d0c810b",
4156 => x"b93d08bb",
4157 => x"3d085b59",
4158 => x"5c775178",
4159 => x"520b0b81",
4160 => x"bdeb3f80",
4161 => x"08800853",
4162 => x"65525a0b",
4163 => x"0b81bbbd",
4164 => x"3fa83d08",
4165 => x"aa3d0858",
4166 => x"547655b8",
4167 => x"3d08ba3d",
4168 => x"08585276",
4169 => x"536b510b",
4170 => x"0b80febe",
4171 => x"3faa3d08",
4172 => x"ac3d085a",
4173 => x"b93d0c78",
4174 => x"ba3d0cb0",
4175 => x"1a56757f",
4176 => x"70810541",
4177 => x"347b662e",
4178 => x"0b0b0be7",
4179 => x"f038811c",
4180 => x"5c80c882",
4181 => x"0a568076",
4182 => x"5555b83d",
4183 => x"08ba3d08",
4184 => x"58527653",
4185 => x"64510b0b",
4186 => x"80ffb23f",
4187 => x"a83d08aa",
4188 => x"3d0871bb",
4189 => x"3d0c70bc",
4190 => x"3d0c5a58",
4191 => x"0b0b0bfe",
4192 => x"f839ff1f",
4193 => x"7033575f",
4194 => x"75b02e0b",
4195 => x"0b0b0bf2",
4196 => x"38811f5f",
4197 => x"0b0b0bed",
4198 => x"e6396566",
4199 => x"484a80d0",
4200 => x"820a5680",
4201 => x"765555b8",
4202 => x"3d08ba3d",
4203 => x"08585276",
4204 => x"5364510b",
4205 => x"0b80fdb2",
4206 => x"3fa83d08",
4207 => x"aa3d08b6",
4208 => x"3d08b83d",
4209 => x"08715770",
4210 => x"58735572",
4211 => x"565c5a5c",
4212 => x"5a0b0b81",
4213 => x"b3bb3f80",
4214 => x"0b800825",
4215 => x"0b0b0bf1",
4216 => x"8e3879b9",
4217 => x"3d0c7aba",
4218 => x"3d0c6c5f",
4219 => x"b17f7081",
4220 => x"05413462",
4221 => x"8105430b",
4222 => x"0b0befc9",
4223 => x"3988b316",
4224 => x"5c6d0b0b",
4225 => x"0bf1e338",
4226 => x"b60ba83d",
4227 => x"08316b11",
4228 => x"4c640544",
4229 => x"81527f51",
4230 => x"0b0b0bb6",
4231 => x"ba3f8008",
4232 => x"4a0b0b0b",
4233 => x"f1d73976",
4234 => x"b92e0b0b",
4235 => x"0bfae938",
4236 => x"81175675",
4237 => x"7f708105",
4238 => x"41340b0b",
4239 => x"0bef8639",
4240 => x"f83d0d7a",
4241 => x"5877802e",
4242 => x"0b0b0b81",
4243 => x"bd380b0b",
4244 => x"82f4ec08",
4245 => x"54b81408",
4246 => x"802e0b0b",
4247 => x"0b818238",
4248 => x"8c182270",
4249 => x"902b7090",
4250 => x"2c70832a",
4251 => x"81328106",
4252 => x"5c515754",
4253 => x"780b0b0b",
4254 => x"80df3890",
4255 => x"18085776",
4256 => x"802e0b0b",
4257 => x"0b80d238",
4258 => x"77087731",
4259 => x"77790c76",
4260 => x"83067a58",
4261 => x"5555730b",
4262 => x"0b0b0b85",
4263 => x"38941808",
4264 => x"56758819",
4265 => x"0c807525",
4266 => x"0b0b0b0b",
4267 => x"ac387453",
4268 => x"76529c18",
4269 => x"0851a418",
4270 => x"0854732d",
4271 => x"800b8008",
4272 => x"250b0b0b",
4273 => x"80df3880",
4274 => x"08177580",
4275 => x"08315657",
4276 => x"7480240b",
4277 => x"0b0b0bd6",
4278 => x"38800b80",
4279 => x"0c8a3d0d",
4280 => x"0473510b",
4281 => x"0b0b81f7",
4282 => x"3f8c1822",
4283 => x"70902b70",
4284 => x"902c7083",
4285 => x"2a813281",
4286 => x"065c5157",
4287 => x"54780b0b",
4288 => x"0b0bd638",
4289 => x"0b0b0bfe",
4290 => x"f2390b0b",
4291 => x"8184c052",
4292 => x"0b0b82f4",
4293 => x"ec08510b",
4294 => x"0b0b93b4",
4295 => x"3f800880",
4296 => x"0c8a3d0d",
4297 => x"048c1822",
4298 => x"80c00754",
4299 => x"738c1923",
4300 => x"ff0b800c",
4301 => x"8a3d0d04",
4302 => x"70725180",
4303 => x"710c800b",
4304 => x"84120c80",
4305 => x"0b88120c",
4306 => x"028e0522",
4307 => x"8c122302",
4308 => x"9205228e",
4309 => x"1223800b",
4310 => x"90120c80",
4311 => x"0b94120c",
4312 => x"800b9812",
4313 => x"0c709c12",
4314 => x"0c0b0b81",
4315 => x"d7880ba0",
4316 => x"120c0b0b",
4317 => x"81d7dd0b",
4318 => x"a4120c0b",
4319 => x"0b81d8ec",
4320 => x"0ba8120c",
4321 => x"0b0b81d9",
4322 => x"c60bac12",
4323 => x"0c5004fa",
4324 => x"3d0d7970",
4325 => x"80dc298c",
4326 => x"11547a53",
4327 => x"56570b0b",
4328 => x"0b989f3f",
4329 => x"80088008",
4330 => x"55568008",
4331 => x"802e0b0b",
4332 => x"0b0ba538",
4333 => x"80088c05",
4334 => x"54800b80",
4335 => x"080c7680",
4336 => x"0884050c",
4337 => x"73800888",
4338 => x"050c7453",
4339 => x"80527351",
4340 => x"0b0b0baa",
4341 => x"c03f7554",
4342 => x"73800c88",
4343 => x"3d0d04fc",
4344 => x"3d0d760b",
4345 => x"0b818aa8",
4346 => x"0bbc120c",
4347 => x"55810bb8",
4348 => x"160c800b",
4349 => x"84dc160c",
4350 => x"830b84e0",
4351 => x"160c84e8",
4352 => x"1584e416",
4353 => x"0c745480",
4354 => x"53845284",
4355 => x"1508510b",
4356 => x"0b0bfea4",
4357 => x"3f745481",
4358 => x"53895288",
4359 => x"1508510b",
4360 => x"0b0bfe94",
4361 => x"3f745482",
4362 => x"538a528c",
4363 => x"1508510b",
4364 => x"0b0bfe84",
4365 => x"3f863d0d",
4366 => x"04f93d0d",
4367 => x"790b0b82",
4368 => x"f4ec0854",
4369 => x"57b81308",
4370 => x"802e0b0b",
4371 => x"0b80db38",
4372 => x"84dc1356",
4373 => x"88160884",
4374 => x"1708ff05",
4375 => x"55558074",
4376 => x"240b0b0b",
4377 => x"0ba6388c",
4378 => x"15227090",
4379 => x"2b70902c",
4380 => x"51545872",
4381 => x"802e0b0b",
4382 => x"0b80e838",
4383 => x"80dc15ff",
4384 => x"15555573",
4385 => x"80250b0b",
4386 => x"0b0bdc38",
4387 => x"75085372",
4388 => x"802e0b0b",
4389 => x"0b0bab38",
4390 => x"72568816",
4391 => x"08841708",
4392 => x"ff055555",
4393 => x"0b0b0bff",
4394 => x"b5397251",
4395 => x"0b0b0bfe",
4396 => x"ae3f0b0b",
4397 => x"82f4ec08",
4398 => x"84dc0556",
4399 => x"0b0b0bff",
4400 => x"93398452",
4401 => x"76510b0b",
4402 => x"0bfdc43f",
4403 => x"8008760c",
4404 => x"8008802e",
4405 => x"0b0b0b80",
4406 => x"c4388008",
4407 => x"560b0b0b",
4408 => x"ffb83981",
4409 => x"0b8c1623",
4410 => x"72750c72",
4411 => x"88160c72",
4412 => x"84160c72",
4413 => x"90160c72",
4414 => x"94160c72",
4415 => x"98160cff",
4416 => x"0b8e1623",
4417 => x"72b0160c",
4418 => x"72b4160c",
4419 => x"7280c416",
4420 => x"0c7280c8",
4421 => x"160c7480",
4422 => x"0c893d0d",
4423 => x"048c770c",
4424 => x"800b800c",
4425 => x"893d0d04",
4426 => x"70700b0b",
4427 => x"8184c052",
4428 => x"73510b0b",
4429 => x"0b8f993f",
4430 => x"50500470",
4431 => x"0b0b82f4",
4432 => x"ec08510b",
4433 => x"0b0b0be0",
4434 => x"3f5004fb",
4435 => x"3d0d7770",
4436 => x"52560b0b",
4437 => x"0ba8f03f",
4438 => x"0b0b82fc",
4439 => x"c80b8805",
4440 => x"08841108",
4441 => x"fc06707b",
4442 => x"319fef05",
4443 => x"e08006e0",
4444 => x"80055656",
4445 => x"53a08074",
4446 => x"240b0b0b",
4447 => x"0b9d3880",
4448 => x"5275510b",
4449 => x"0b80cbba",
4450 => x"3f0b0b82",
4451 => x"fcd00815",
4452 => x"53728008",
4453 => x"2e0b0b0b",
4454 => x"0b923875",
4455 => x"510b0b0b",
4456 => x"a8a63f80",
4457 => x"5372800c",
4458 => x"873d0d04",
4459 => x"73305275",
4460 => x"510b0b80",
4461 => x"cb8c3f80",
4462 => x"08ff2e0b",
4463 => x"0b0b0bb1",
4464 => x"380b0b82",
4465 => x"fcc80b88",
4466 => x"05087575",
4467 => x"31810784",
4468 => x"120c530b",
4469 => x"0b82fc8c",
4470 => x"0874310b",
4471 => x"0b82fc8c",
4472 => x"0c75510b",
4473 => x"0b0ba7e0",
4474 => x"3f810b80",
4475 => x"0c873d0d",
4476 => x"04805275",
4477 => x"510b0b80",
4478 => x"cac83f0b",
4479 => x"0b82fcc8",
4480 => x"0b880508",
4481 => x"80087131",
4482 => x"56538f75",
4483 => x"250b0b0b",
4484 => x"ff893880",
4485 => x"080b0b82",
4486 => x"fcbc0831",
4487 => x"0b0b82fc",
4488 => x"8c0c7481",
4489 => x"0784140c",
4490 => x"75510b0b",
4491 => x"0ba7993f",
4492 => x"80530b0b",
4493 => x"0bfeee39",
4494 => x"f63d0d7c",
4495 => x"7e545b72",
4496 => x"802e0b0b",
4497 => x"0b82c838",
4498 => x"7a510b0b",
4499 => x"0ba6f83f",
4500 => x"f8138411",
4501 => x"0870fe06",
4502 => x"70138411",
4503 => x"08fc065d",
4504 => x"58595458",
4505 => x"0b0b82fc",
4506 => x"d008752e",
4507 => x"0b0b0b83",
4508 => x"b5387884",
4509 => x"160c8073",
4510 => x"8106545a",
4511 => x"727a2e0b",
4512 => x"0b0b828f",
4513 => x"38781584",
4514 => x"11088106",
4515 => x"5153720b",
4516 => x"0b0b0ba8",
4517 => x"38781757",
4518 => x"790b0b0b",
4519 => x"82a13888",
4520 => x"15085372",
4521 => x"0b0b82fc",
4522 => x"d02e0b0b",
4523 => x"0b83d738",
4524 => x"8c150870",
4525 => x"8c150c73",
4526 => x"88120c56",
4527 => x"76810784",
4528 => x"190c7618",
4529 => x"77710c53",
4530 => x"790b0b0b",
4531 => x"81b93883",
4532 => x"ff77270b",
4533 => x"0b0b81fb",
4534 => x"3876892a",
4535 => x"77832a56",
4536 => x"5372802e",
4537 => x"0b0b0b80",
4538 => x"d3387686",
4539 => x"2ab80555",
4540 => x"8473270b",
4541 => x"0b0b80c4",
4542 => x"3880db13",
4543 => x"55947327",
4544 => x"0b0b0b0b",
4545 => x"b738768c",
4546 => x"2a80ee05",
4547 => x"5580d473",
4548 => x"270b0b0b",
4549 => x"0ba63876",
4550 => x"8f2a80f7",
4551 => x"055582d4",
4552 => x"73270b0b",
4553 => x"0b0b9538",
4554 => x"76922a80",
4555 => x"fc05558a",
4556 => x"d473270b",
4557 => x"0b0b0b84",
4558 => x"3880fe55",
4559 => x"74101010",
4560 => x"0b0b82fc",
4561 => x"c8058811",
4562 => x"08555673",
4563 => x"762e0b0b",
4564 => x"0b82fa38",
4565 => x"841408fc",
4566 => x"06537673",
4567 => x"270b0b0b",
4568 => x"0b913888",
4569 => x"14085473",
4570 => x"762e0981",
4571 => x"060b0b0b",
4572 => x"0be2388c",
4573 => x"1408708c",
4574 => x"1a0c7488",
4575 => x"1a0c7888",
4576 => x"120c5677",
4577 => x"8c150c7a",
4578 => x"510b0b0b",
4579 => x"a4ba3f8c",
4580 => x"3d0d0477",
4581 => x"08787131",
4582 => x"59770588",
4583 => x"19085457",
4584 => x"720b0b82",
4585 => x"fcd02e0b",
4586 => x"0b0b80f2",
4587 => x"388c1808",
4588 => x"708c150c",
4589 => x"7388120c",
4590 => x"560b0b0b",
4591 => x"fdc73988",
4592 => x"15088c16",
4593 => x"08708c13",
4594 => x"0c578817",
4595 => x"0c0b0b0b",
4596 => x"fdea3976",
4597 => x"832a7054",
4598 => x"55807524",
4599 => x"0b0b0b81",
4600 => x"bd387282",
4601 => x"2c81712b",
4602 => x"0b0b82fc",
4603 => x"cc08070b",
4604 => x"0b82fcc8",
4605 => x"0b84050c",
4606 => x"53741010",
4607 => x"100b0b82",
4608 => x"fcc80588",
4609 => x"11085556",
4610 => x"758c190c",
4611 => x"7388190c",
4612 => x"7788170c",
4613 => x"778c150c",
4614 => x"0b0b0bfe",
4615 => x"ea39815a",
4616 => x"0b0b0bfc",
4617 => x"e0397817",
4618 => x"73810654",
4619 => x"57720b0b",
4620 => x"0b0b9838",
4621 => x"77087871",
4622 => x"31597705",
4623 => x"8c190888",
4624 => x"1a08718c",
4625 => x"120c8812",
4626 => x"0c575776",
4627 => x"81078419",
4628 => x"0c770b0b",
4629 => x"82fcc80b",
4630 => x"88050c0b",
4631 => x"0b82fcc4",
4632 => x"0877260b",
4633 => x"0b0bfe9f",
4634 => x"380b0b82",
4635 => x"fcc00852",
4636 => x"7a510b0b",
4637 => x"0bf9d43f",
4638 => x"7a510b0b",
4639 => x"0ba2c93f",
4640 => x"0b0b0bfe",
4641 => x"8a398178",
4642 => x"8c150c78",
4643 => x"88150c73",
4644 => x"8c1a0c73",
4645 => x"881a0c5a",
4646 => x"0b0b0bfc",
4647 => x"9f398315",
4648 => x"70822c81",
4649 => x"712b0b0b",
4650 => x"82fccc08",
4651 => x"070b0b82",
4652 => x"fcc80b84",
4653 => x"050c5153",
4654 => x"74101010",
4655 => x"0b0b82fc",
4656 => x"c8058811",
4657 => x"0855560b",
4658 => x"0b0bfebc",
4659 => x"39745380",
4660 => x"75240b0b",
4661 => x"0b0bae38",
4662 => x"72822c81",
4663 => x"712b0b0b",
4664 => x"82fccc08",
4665 => x"070b0b82",
4666 => x"fcc80b84",
4667 => x"050c5375",
4668 => x"8c190c73",
4669 => x"88190c77",
4670 => x"88170c77",
4671 => x"8c150c0b",
4672 => x"0b0bfd83",
4673 => x"39831570",
4674 => x"822c8171",
4675 => x"2b0b0b82",
4676 => x"fccc0807",
4677 => x"0b0b82fc",
4678 => x"c80b8405",
4679 => x"0c51530b",
4680 => x"0b0b0bcb",
4681 => x"39f23d0d",
4682 => x"60628811",
4683 => x"08705757",
4684 => x"5f5a7480",
4685 => x"2e0b0b0b",
4686 => x"81b3388c",
4687 => x"1a227083",
4688 => x"2a813270",
4689 => x"81065155",
4690 => x"58730b0b",
4691 => x"0b0b8a38",
4692 => x"901a080b",
4693 => x"0b0b0b97",
4694 => x"3879510b",
4695 => x"0b0bc388",
4696 => x"3fff5480",
4697 => x"080b0b0b",
4698 => x"8183388c",
4699 => x"1a22587d",
4700 => x"08578078",
4701 => x"83ffff06",
4702 => x"700a100a",
4703 => x"70810651",
4704 => x"56575573",
4705 => x"752e0b0b",
4706 => x"0b80e938",
4707 => x"740b0b0b",
4708 => x"0b943876",
4709 => x"08841808",
4710 => x"88195956",
4711 => x"5974802e",
4712 => x"0b0b0b0b",
4713 => x"ee387454",
4714 => x"88807527",
4715 => x"0b0b0b0b",
4716 => x"84388880",
4717 => x"54735378",
4718 => x"529c1a08",
4719 => x"51a41a08",
4720 => x"54732d80",
4721 => x"0b800825",
4722 => x"0b0b0b83",
4723 => x"bf388008",
4724 => x"19758008",
4725 => x"317f8805",
4726 => x"08800831",
4727 => x"70618805",
4728 => x"0c565659",
4729 => x"730b0b0b",
4730 => x"ffa23880",
4731 => x"5473800c",
4732 => x"903d0d04",
4733 => x"75813270",
4734 => x"81067641",
4735 => x"51547380",
4736 => x"2e0b0b0b",
4737 => x"81f03874",
4738 => x"0b0b0b0b",
4739 => x"94387608",
4740 => x"84180888",
4741 => x"19595659",
4742 => x"74802e0b",
4743 => x"0b0b0bee",
4744 => x"38881a08",
4745 => x"7883ffff",
4746 => x"0670892a",
4747 => x"70810651",
4748 => x"56595673",
4749 => x"802e0b0b",
4750 => x"0b83e338",
4751 => x"7575270b",
4752 => x"0b0b0b90",
4753 => x"3877872a",
4754 => x"70810651",
4755 => x"54730b0b",
4756 => x"0b838c38",
4757 => x"7476270b",
4758 => x"0b0b0b83",
4759 => x"38745675",
4760 => x"53785279",
4761 => x"08510b0b",
4762 => x"0b9bb83f",
4763 => x"881a0876",
4764 => x"31881b0c",
4765 => x"7908167a",
4766 => x"0c745675",
4767 => x"19757731",
4768 => x"7f880508",
4769 => x"78317061",
4770 => x"88050c56",
4771 => x"56597380",
4772 => x"2e0b0b0b",
4773 => x"fed5388c",
4774 => x"1a22580b",
4775 => x"0b0bfee7",
4776 => x"39777854",
4777 => x"79537b52",
4778 => x"560b0b0b",
4779 => x"9af53f88",
4780 => x"1a087831",
4781 => x"881b0c79",
4782 => x"08187a0c",
4783 => x"7c76315d",
4784 => x"7c0b0b0b",
4785 => x"0b943879",
4786 => x"510b0b0b",
4787 => x"eef23f80",
4788 => x"080b0b0b",
4789 => x"81b63880",
4790 => x"085f7519",
4791 => x"7577317f",
4792 => x"88050878",
4793 => x"31706188",
4794 => x"050c5656",
4795 => x"5973802e",
4796 => x"0b0b0bfd",
4797 => x"f638740b",
4798 => x"0b0b81a4",
4799 => x"38760884",
4800 => x"18088819",
4801 => x"59565974",
4802 => x"802e0b0b",
4803 => x"0b0bee38",
4804 => x"74538a52",
4805 => x"78510b0b",
4806 => x"0b98bb3f",
4807 => x"80087931",
4808 => x"81055d80",
4809 => x"080b0b0b",
4810 => x"0b843881",
4811 => x"155d815f",
4812 => x"7c58747d",
4813 => x"270b0b0b",
4814 => x"0b833874",
4815 => x"58941a08",
4816 => x"881b0811",
4817 => x"575c807a",
4818 => x"085c5490",
4819 => x"1a087b27",
4820 => x"0b0b0b0b",
4821 => x"83388154",
4822 => x"7578250b",
4823 => x"0b0b0b88",
4824 => x"38730b0b",
4825 => x"0b80c638",
4826 => x"7b78240b",
4827 => x"0b0bfeb1",
4828 => x"387b5378",
4829 => x"529c1a08",
4830 => x"51a41a08",
4831 => x"54732d80",
4832 => x"08568008",
4833 => x"80240b0b",
4834 => x"0bfeb138",
4835 => x"8c1a2280",
4836 => x"c0075473",
4837 => x"8c1b23ff",
4838 => x"5473800c",
4839 => x"903d0d04",
4840 => x"7e0b0b0b",
4841 => x"ff8a380b",
4842 => x"0b0bfee4",
4843 => x"39755378",
4844 => x"527a510b",
4845 => x"0b0b98eb",
4846 => x"3f790816",
4847 => x"7a0c7951",
4848 => x"0b0b0bec",
4849 => x"fb3f8008",
4850 => x"0b0b0bff",
4851 => x"bf387c76",
4852 => x"315d7c0b",
4853 => x"0b0bfe82",
4854 => x"380b0b0b",
4855 => x"fde93990",
4856 => x"1a087a08",
4857 => x"71317611",
4858 => x"70565a57",
4859 => x"520b0b82",
4860 => x"f4ec0851",
4861 => x"0b0b0bb4",
4862 => x"ad3f8008",
4863 => x"802e0b0b",
4864 => x"0bff8938",
4865 => x"8008901b",
4866 => x"0c800816",
4867 => x"7a0c7794",
4868 => x"1b0c7488",
4869 => x"1b0c7456",
4870 => x"0b0b0bfc",
4871 => x"b7397908",
4872 => x"58901a08",
4873 => x"78270b0b",
4874 => x"0b0b8338",
4875 => x"81547575",
4876 => x"270b0b0b",
4877 => x"0b883873",
4878 => x"0b0b0b0b",
4879 => x"bc38941a",
4880 => x"08567575",
4881 => x"260b0b0b",
4882 => x"80e53875",
4883 => x"5378529c",
4884 => x"1a0851a4",
4885 => x"1a085473",
4886 => x"2d800856",
4887 => x"80088024",
4888 => x"0b0b0bfc",
4889 => x"96388c1a",
4890 => x"2280c007",
4891 => x"54738c1b",
4892 => x"23ff540b",
4893 => x"0b0bfea1",
4894 => x"39755378",
4895 => x"5277510b",
4896 => x"0b0b979f",
4897 => x"3f790816",
4898 => x"7a0c7951",
4899 => x"0b0b0beb",
4900 => x"af3f8008",
4901 => x"802e0b0b",
4902 => x"0bfbe038",
4903 => x"8c1a2280",
4904 => x"c0075473",
4905 => x"8c1b23ff",
4906 => x"540b0b0b",
4907 => x"fdeb3974",
4908 => x"75547953",
4909 => x"7852560b",
4910 => x"0b0b96e7",
4911 => x"3f881a08",
4912 => x"7531881b",
4913 => x"0c790815",
4914 => x"7a0c0b0b",
4915 => x"0bfbac39",
4916 => x"f93d0d79",
4917 => x"7b585380",
4918 => x"0b0b0b82",
4919 => x"f4ec0853",
4920 => x"5672722e",
4921 => x"0b0b0b80",
4922 => x"d53884dc",
4923 => x"13557476",
4924 => x"2e0b0b0b",
4925 => x"80c83888",
4926 => x"15088416",
4927 => x"08ff0554",
4928 => x"54807324",
4929 => x"0b0b0b0b",
4930 => x"a4388c14",
4931 => x"2270902b",
4932 => x"70902c51",
4933 => x"5358710b",
4934 => x"0b0b80f6",
4935 => x"3880dc14",
4936 => x"ff145454",
4937 => x"7280250b",
4938 => x"0b0b0bde",
4939 => x"38740855",
4940 => x"740b0b0b",
4941 => x"0bc1380b",
4942 => x"0b82f4ec",
4943 => x"085284dc",
4944 => x"12557480",
4945 => x"2e0b0b0b",
4946 => x"80c13888",
4947 => x"15088416",
4948 => x"08ff0554",
4949 => x"54807324",
4950 => x"0b0b0b0b",
4951 => x"a4388c14",
4952 => x"2270902b",
4953 => x"70902c51",
4954 => x"5358710b",
4955 => x"0b0b0bb8",
4956 => x"3880dc14",
4957 => x"ff145454",
4958 => x"7280250b",
4959 => x"0b0b0bde",
4960 => x"38740855",
4961 => x"740b0b0b",
4962 => x"0bc13875",
4963 => x"800c893d",
4964 => x"0d047351",
4965 => x"762d7580",
4966 => x"080780dc",
4967 => x"15ff1555",
4968 => x"55560b0b",
4969 => x"0bfefd39",
4970 => x"7351762d",
4971 => x"75800807",
4972 => x"80dc15ff",
4973 => x"15555556",
4974 => x"0b0b0bff",
4975 => x"bb39fc3d",
4976 => x"0d767955",
4977 => x"5573802e",
4978 => x"0b0b0b0b",
4979 => x"9f380b0b",
4980 => x"82f1c852",
4981 => x"73510b0b",
4982 => x"0bbe8d3f",
4983 => x"80080b0b",
4984 => x"0b0b9638",
4985 => x"77b0160c",
4986 => x"73b4160c",
4987 => x"0b0b82f1",
4988 => x"c8537280",
4989 => x"0c863d0d",
4990 => x"040b0b82",
4991 => x"f0ec5273",
4992 => x"510b0b0b",
4993 => x"bde23f80",
4994 => x"53800873",
4995 => x"2e098106",
4996 => x"0b0b0b0b",
4997 => x"dd3877b0",
4998 => x"160c73b4",
4999 => x"160c0b0b",
5000 => x"0b0bc939",
5001 => x"0b0b82fc",
5002 => x"8808800c",
5003 => x"040b0b82",
5004 => x"f1d80b80",
5005 => x"0c047070",
5006 => x"70755374",
5007 => x"520b0b82",
5008 => x"f4ec0851",
5009 => x"0b0b0bfe",
5010 => x"f53f5050",
5011 => x"5004700b",
5012 => x"0b82f4ec",
5013 => x"08510b0b",
5014 => x"0b0bd23f",
5015 => x"5004ea3d",
5016 => x"0d688c11",
5017 => x"22700a10",
5018 => x"0a810657",
5019 => x"5856740b",
5020 => x"0b0b8180",
5021 => x"388e1622",
5022 => x"70902b70",
5023 => x"902c5155",
5024 => x"58807424",
5025 => x"0b0b0b80",
5026 => x"c038983d",
5027 => x"c4055373",
5028 => x"520b0b82",
5029 => x"f4ec0851",
5030 => x"0b0b80c1",
5031 => x"ac3f800b",
5032 => x"8008240b",
5033 => x"0b0b0b9d",
5034 => x"387983e0",
5035 => x"80065473",
5036 => x"80c0802e",
5037 => x"0b0b0b81",
5038 => x"aa387382",
5039 => x"80802e0b",
5040 => x"0b0b81ac",
5041 => x"388c1622",
5042 => x"57769080",
5043 => x"0754738c",
5044 => x"17238880",
5045 => x"520b0b82",
5046 => x"f4ec0851",
5047 => x"0b0b0b81",
5048 => x"e13f8008",
5049 => x"0b0b0b0b",
5050 => x"9d388c16",
5051 => x"22820754",
5052 => x"738c1723",
5053 => x"80c31670",
5054 => x"770c9017",
5055 => x"0c810b94",
5056 => x"170c983d",
5057 => x"0d040b0b",
5058 => x"82f4ec08",
5059 => x"0b0b818a",
5060 => x"a80bbc12",
5061 => x"0c548c16",
5062 => x"22818007",
5063 => x"54738c17",
5064 => x"23800876",
5065 => x"0c800890",
5066 => x"170c8880",
5067 => x"0b94170c",
5068 => x"74802e0b",
5069 => x"0b0b0bca",
5070 => x"388e1622",
5071 => x"70902b70",
5072 => x"902c5355",
5073 => x"580b0b80",
5074 => x"ced33f80",
5075 => x"08802e0b",
5076 => x"0b0bffae",
5077 => x"388c1622",
5078 => x"81075473",
5079 => x"8c172398",
5080 => x"3d0d0481",
5081 => x"0b8c1722",
5082 => x"58550b0b",
5083 => x"0bfeda39",
5084 => x"a816080b",
5085 => x"0b81d8ec",
5086 => x"2e098106",
5087 => x"0b0b0bfe",
5088 => x"c4388c16",
5089 => x"22888007",
5090 => x"54738c17",
5091 => x"2388800b",
5092 => x"80cc170c",
5093 => x"0b0b0bfe",
5094 => x"b9397070",
5095 => x"73520b0b",
5096 => x"82f4ec08",
5097 => x"510b0b0b",
5098 => x"0b983f50",
5099 => x"50047070",
5100 => x"73520b0b",
5101 => x"82f4ec08",
5102 => x"510b0b0b",
5103 => x"ecfa3f50",
5104 => x"5004f33d",
5105 => x"0d7f618b",
5106 => x"1170f806",
5107 => x"5c55555e",
5108 => x"7296260b",
5109 => x"0b0b0b83",
5110 => x"38905980",
5111 => x"7924747a",
5112 => x"26075380",
5113 => x"5472742e",
5114 => x"0981060b",
5115 => x"0b0b80d9",
5116 => x"387d510b",
5117 => x"0b0b93cf",
5118 => x"3f7883f7",
5119 => x"260b0b0b",
5120 => x"80ce3878",
5121 => x"832a7010",
5122 => x"10100b0b",
5123 => x"82fcc805",
5124 => x"8c110859",
5125 => x"595a7678",
5126 => x"2e0b0b0b",
5127 => x"84aa3884",
5128 => x"1708fc06",
5129 => x"568c1708",
5130 => x"88180871",
5131 => x"8c120c88",
5132 => x"120c5875",
5133 => x"17841108",
5134 => x"81078412",
5135 => x"0c537d51",
5136 => x"0b0b0b93",
5137 => x"833f8817",
5138 => x"5473800c",
5139 => x"8f3d0d04",
5140 => x"78892a79",
5141 => x"832a5b53",
5142 => x"72802e0b",
5143 => x"0b0b80d3",
5144 => x"3878862a",
5145 => x"b8055a84",
5146 => x"73270b0b",
5147 => x"0b80c438",
5148 => x"80db135a",
5149 => x"9473270b",
5150 => x"0b0b0bb7",
5151 => x"38788c2a",
5152 => x"80ee055a",
5153 => x"80d47327",
5154 => x"0b0b0b0b",
5155 => x"a638788f",
5156 => x"2a80f705",
5157 => x"5a82d473",
5158 => x"270b0b0b",
5159 => x"0b953878",
5160 => x"922a80fc",
5161 => x"055a8ad4",
5162 => x"73270b0b",
5163 => x"0b0b8438",
5164 => x"80fe5a79",
5165 => x"1010100b",
5166 => x"0b82fcc8",
5167 => x"058c1108",
5168 => x"58557675",
5169 => x"2e0b0b0b",
5170 => x"0bad3884",
5171 => x"1708fc06",
5172 => x"707a3155",
5173 => x"56738f24",
5174 => x"0b0b0b8b",
5175 => x"94387380",
5176 => x"250b0b0b",
5177 => x"febf388c",
5178 => x"17085776",
5179 => x"752e0981",
5180 => x"060b0b0b",
5181 => x"0bd53881",
5182 => x"1a5a0b0b",
5183 => x"82fcd808",
5184 => x"57760b0b",
5185 => x"82fcd02e",
5186 => x"0b0b0b83",
5187 => x"9a388417",
5188 => x"08fc0670",
5189 => x"7a315556",
5190 => x"738f240b",
5191 => x"0b0b82c4",
5192 => x"380b0b82",
5193 => x"fcd00b0b",
5194 => x"0b82fcdc",
5195 => x"0c0b0b82",
5196 => x"fcd00b0b",
5197 => x"0b82fcd8",
5198 => x"0c738025",
5199 => x"0b0b0bfd",
5200 => x"f23883ff",
5201 => x"76270b0b",
5202 => x"0b84e238",
5203 => x"75892a76",
5204 => x"832a5553",
5205 => x"72802e0b",
5206 => x"0b0b80d3",
5207 => x"3875862a",
5208 => x"b8055484",
5209 => x"73270b0b",
5210 => x"0b80c438",
5211 => x"80db1354",
5212 => x"9473270b",
5213 => x"0b0b0bb7",
5214 => x"38758c2a",
5215 => x"80ee0554",
5216 => x"80d47327",
5217 => x"0b0b0b0b",
5218 => x"a638758f",
5219 => x"2a80f705",
5220 => x"5482d473",
5221 => x"270b0b0b",
5222 => x"0b953875",
5223 => x"922a80fc",
5224 => x"05548ad4",
5225 => x"73270b0b",
5226 => x"0b0b8438",
5227 => x"80fe5473",
5228 => x"1010100b",
5229 => x"0b82fcc8",
5230 => x"05881108",
5231 => x"56587478",
5232 => x"2e0b0b0b",
5233 => x"88b83884",
5234 => x"1508fc06",
5235 => x"53757327",
5236 => x"0b0b0b0b",
5237 => x"91388815",
5238 => x"08557478",
5239 => x"2e098106",
5240 => x"0b0b0b0b",
5241 => x"e2388c15",
5242 => x"080b0b82",
5243 => x"fcc80b84",
5244 => x"0508718c",
5245 => x"1a0c7688",
5246 => x"1a0c7888",
5247 => x"130c788c",
5248 => x"180c5d58",
5249 => x"7953807a",
5250 => x"240b0b0b",
5251 => x"84e93872",
5252 => x"822c8171",
5253 => x"2b5c537a",
5254 => x"7c260b0b",
5255 => x"0b81c538",
5256 => x"7b7b0653",
5257 => x"720b0b0b",
5258 => x"83d03879",
5259 => x"fc068405",
5260 => x"5a7a1070",
5261 => x"7d06545b",
5262 => x"720b0b0b",
5263 => x"83bc3884",
5264 => x"1a5a0b0b",
5265 => x"0b0bea39",
5266 => x"88178c11",
5267 => x"08585876",
5268 => x"782e0981",
5269 => x"060b0b0b",
5270 => x"fbc53882",
5271 => x"1a5a0b0b",
5272 => x"0bfd9739",
5273 => x"78177981",
5274 => x"0784190c",
5275 => x"700b0b82",
5276 => x"fcdc0c70",
5277 => x"0b0b82fc",
5278 => x"d80c0b0b",
5279 => x"82fcd00b",
5280 => x"8c120c8c",
5281 => x"11088812",
5282 => x"0c748107",
5283 => x"84120c74",
5284 => x"1175710c",
5285 => x"51537d51",
5286 => x"0b0b0b8e",
5287 => x"ab3f8817",
5288 => x"540b0b0b",
5289 => x"fba3390b",
5290 => x"0b82fcc8",
5291 => x"0b840508",
5292 => x"7a545c79",
5293 => x"80250b0b",
5294 => x"0bfed438",
5295 => x"0b0b0b83",
5296 => x"b6397a09",
5297 => x"7c06700b",
5298 => x"0b82fcc8",
5299 => x"0b84050c",
5300 => x"5c7a105b",
5301 => x"7a7c260b",
5302 => x"0b0b0b88",
5303 => x"387a0b0b",
5304 => x"0b86f738",
5305 => x"0b0b82fc",
5306 => x"c80b8805",
5307 => x"08708412",
5308 => x"08fc0670",
5309 => x"7c317c72",
5310 => x"268f7225",
5311 => x"0757575c",
5312 => x"5d557280",
5313 => x"2e0b0b0b",
5314 => x"80f73879",
5315 => x"7a160b0b",
5316 => x"82fcc008",
5317 => x"1b90115a",
5318 => x"55575b0b",
5319 => x"0b82fcbc",
5320 => x"08ff2e0b",
5321 => x"0b0b0b88",
5322 => x"38a08f13",
5323 => x"e0800657",
5324 => x"76527d51",
5325 => x"0b0b0bb0",
5326 => x"893f8008",
5327 => x"548008ff",
5328 => x"2e0b0b0b",
5329 => x"0b983880",
5330 => x"0876270b",
5331 => x"0b0b82e1",
5332 => x"38740b0b",
5333 => x"82fcc82e",
5334 => x"0b0b0b82",
5335 => x"d4380b0b",
5336 => x"82fcc80b",
5337 => x"88050855",
5338 => x"841508fc",
5339 => x"06707a31",
5340 => x"7a72268f",
5341 => x"72250752",
5342 => x"5553720b",
5343 => x"0b0b84ee",
5344 => x"38747981",
5345 => x"0784170c",
5346 => x"7916700b",
5347 => x"0b82fcc8",
5348 => x"0b88050c",
5349 => x"75810784",
5350 => x"120c547e",
5351 => x"52570b0b",
5352 => x"0b8ca53f",
5353 => x"8817540b",
5354 => x"0b0bf99d",
5355 => x"3975832a",
5356 => x"70545480",
5357 => x"74240b0b",
5358 => x"0b81c538",
5359 => x"72822c81",
5360 => x"712b0b0b",
5361 => x"82fccc08",
5362 => x"07700b0b",
5363 => x"82fcc80b",
5364 => x"84050c75",
5365 => x"1010100b",
5366 => x"0b82fcc8",
5367 => x"05881108",
5368 => x"585a5d53",
5369 => x"778c180c",
5370 => x"7488180c",
5371 => x"7688190c",
5372 => x"768c160c",
5373 => x"0b0b0bfc",
5374 => x"8b39797a",
5375 => x"1010100b",
5376 => x"0b82fcc8",
5377 => x"05705759",
5378 => x"5d8c1508",
5379 => x"5776752e",
5380 => x"0b0b0b0b",
5381 => x"ad388417",
5382 => x"08fc0670",
5383 => x"7a315556",
5384 => x"738f240b",
5385 => x"0b0b84d5",
5386 => x"38738025",
5387 => x"0b0b0b85",
5388 => x"92388c17",
5389 => x"08577675",
5390 => x"2e098106",
5391 => x"0b0b0b0b",
5392 => x"d5388815",
5393 => x"811b7083",
5394 => x"06555b55",
5395 => x"720b0b0b",
5396 => x"ffb7387c",
5397 => x"83065372",
5398 => x"802e0b0b",
5399 => x"0bfce338",
5400 => x"ff1df819",
5401 => x"595d8818",
5402 => x"08782e0b",
5403 => x"0b0b0be3",
5404 => x"380b0b0b",
5405 => x"fcdb3983",
5406 => x"1a530b0b",
5407 => x"0bfb9039",
5408 => x"83147082",
5409 => x"2c81712b",
5410 => x"0b0b82fc",
5411 => x"cc080770",
5412 => x"0b0b82fc",
5413 => x"c80b8405",
5414 => x"0c761010",
5415 => x"100b0b82",
5416 => x"fcc80588",
5417 => x"1108595b",
5418 => x"5e51530b",
5419 => x"0b0bfeb4",
5420 => x"390b0b82",
5421 => x"fc8c0817",
5422 => x"58800876",
5423 => x"2e0b0b0b",
5424 => x"81b2380b",
5425 => x"0b82fcbc",
5426 => x"08ff2e0b",
5427 => x"0b0b84e8",
5428 => x"38737631",
5429 => x"180b0b82",
5430 => x"fc8c0c73",
5431 => x"87067057",
5432 => x"5372802e",
5433 => x"0b0b0b0b",
5434 => x"88388873",
5435 => x"31701555",
5436 => x"5676149f",
5437 => x"ff06a080",
5438 => x"71311770",
5439 => x"547f5357",
5440 => x"530b0b0b",
5441 => x"acbc3f80",
5442 => x"08538008",
5443 => x"ff2e0b0b",
5444 => x"0b81d138",
5445 => x"0b0b82fc",
5446 => x"8c081670",
5447 => x"0b0b82fc",
5448 => x"8c0c7475",
5449 => x"0b0b82fc",
5450 => x"c80b8805",
5451 => x"0c747631",
5452 => x"18708107",
5453 => x"51555658",
5454 => x"7b0b0b82",
5455 => x"fcc82e0b",
5456 => x"0b0b8488",
5457 => x"38798f26",
5458 => x"0b0b0b83",
5459 => x"a038810b",
5460 => x"84150c84",
5461 => x"1508fc06",
5462 => x"707a317a",
5463 => x"72268f72",
5464 => x"25075255",
5465 => x"5372802e",
5466 => x"0b0b0bfc",
5467 => x"94380b0b",
5468 => x"0b80fb39",
5469 => x"80089fff",
5470 => x"0653720b",
5471 => x"0b0bfec3",
5472 => x"38770b0b",
5473 => x"82fc8c0c",
5474 => x"0b0b82fc",
5475 => x"c80b8805",
5476 => x"087b1881",
5477 => x"0784120c",
5478 => x"550b0b82",
5479 => x"fcb80878",
5480 => x"270b0b0b",
5481 => x"0b883877",
5482 => x"0b0b82fc",
5483 => x"b80c0b0b",
5484 => x"82fcb408",
5485 => x"78270b0b",
5486 => x"0bfbad38",
5487 => x"770b0b82",
5488 => x"fcb40c84",
5489 => x"1508fc06",
5490 => x"707a317a",
5491 => x"72268f72",
5492 => x"25075255",
5493 => x"5372802e",
5494 => x"0b0b0bfb",
5495 => x"a4380b0b",
5496 => x"0b0b8b39",
5497 => x"80745456",
5498 => x"0b0b0bfe",
5499 => x"a7397d51",
5500 => x"0b0b0b87",
5501 => x"d33f800b",
5502 => x"800c8f3d",
5503 => x"0d047353",
5504 => x"8074240b",
5505 => x"0b0b0bb0",
5506 => x"3872822c",
5507 => x"81712b0b",
5508 => x"0b82fccc",
5509 => x"0807700b",
5510 => x"0b82fcc8",
5511 => x"0b84050c",
5512 => x"5d53778c",
5513 => x"180c7488",
5514 => x"180c7688",
5515 => x"190c768c",
5516 => x"160c0b0b",
5517 => x"0bf7cd39",
5518 => x"83147082",
5519 => x"2c81712b",
5520 => x"0b0b82fc",
5521 => x"cc080770",
5522 => x"0b0b82fc",
5523 => x"c80b8405",
5524 => x"0c5e5153",
5525 => x"0b0b0b0b",
5526 => x"c9397b7b",
5527 => x"0653720b",
5528 => x"0b0bfb96",
5529 => x"38841a7b",
5530 => x"105c5a0b",
5531 => x"0b0b0bea",
5532 => x"39ff1a81",
5533 => x"11515a0b",
5534 => x"0b0bf4fe",
5535 => x"39781779",
5536 => x"81078419",
5537 => x"0c8c1808",
5538 => x"88190871",
5539 => x"8c120c88",
5540 => x"120c5970",
5541 => x"0b0b82fc",
5542 => x"dc0c700b",
5543 => x"0b82fcd8",
5544 => x"0c0b0b82",
5545 => x"fcd00b8c",
5546 => x"120c8c11",
5547 => x"0888120c",
5548 => x"74810784",
5549 => x"120c7411",
5550 => x"75710c51",
5551 => x"530b0b0b",
5552 => x"f7d43975",
5553 => x"17841108",
5554 => x"81078412",
5555 => x"0c538c17",
5556 => x"08881808",
5557 => x"718c120c",
5558 => x"88120c58",
5559 => x"7d510b0b",
5560 => x"0b85e53f",
5561 => x"8817540b",
5562 => x"0b0bf2dd",
5563 => x"39728415",
5564 => x"0cf41af8",
5565 => x"0670841e",
5566 => x"08810607",
5567 => x"841e0c70",
5568 => x"1d545b85",
5569 => x"0b84140c",
5570 => x"850b8814",
5571 => x"0c8f7b27",
5572 => x"0b0b0bfd",
5573 => x"8438881c",
5574 => x"527d510b",
5575 => x"0b0bde98",
5576 => x"3f0b0b82",
5577 => x"fcc80b88",
5578 => x"05080b0b",
5579 => x"82fc8c08",
5580 => x"59550b0b",
5581 => x"0bfce239",
5582 => x"770b0b82",
5583 => x"fc8c0c73",
5584 => x"0b0b82fc",
5585 => x"bc0c0b0b",
5586 => x"0bfb9039",
5587 => x"7284150c",
5588 => x"0b0b0bfc",
5589 => x"c439fa3d",
5590 => x"0d7a7902",
5591 => x"8805a705",
5592 => x"33565253",
5593 => x"8373270b",
5594 => x"0b0b0b8e",
5595 => x"38708306",
5596 => x"5271802e",
5597 => x"0b0b0b0b",
5598 => x"b438ff13",
5599 => x"5372ff2e",
5600 => x"0b0b0b0b",
5601 => x"9f387033",
5602 => x"5273722e",
5603 => x"0b0b0b0b",
5604 => x"95388111",
5605 => x"ff145451",
5606 => x"72ff2e09",
5607 => x"81060b0b",
5608 => x"0b0be338",
5609 => x"80517080",
5610 => x"0c883d0d",
5611 => x"04707257",
5612 => x"55835175",
5613 => x"82802914",
5614 => x"ff125256",
5615 => x"7080250b",
5616 => x"0b0b0bef",
5617 => x"38837327",
5618 => x"0b0b0b80",
5619 => x"ce387408",
5620 => x"76327009",
5621 => x"f7fbfdff",
5622 => x"120670f8",
5623 => x"84828180",
5624 => x"06515151",
5625 => x"70802e0b",
5626 => x"0b0b0ba0",
5627 => x"38745180",
5628 => x"52703357",
5629 => x"73772e0b",
5630 => x"0b0bffaa",
5631 => x"38811181",
5632 => x"13535183",
5633 => x"72270b0b",
5634 => x"0b0be638",
5635 => x"fc138416",
5636 => x"56537283",
5637 => x"260b0b0b",
5638 => x"ffb43874",
5639 => x"510b0b0b",
5640 => x"fed839fa",
5641 => x"3d0d787a",
5642 => x"7c727272",
5643 => x"57575759",
5644 => x"56567476",
5645 => x"270b0b0b",
5646 => x"0bbe3876",
5647 => x"15517571",
5648 => x"270b0b0b",
5649 => x"0bb23870",
5650 => x"7717ff14",
5651 => x"54555371",
5652 => x"ff2e0b0b",
5653 => x"0b0b9a38",
5654 => x"ff14ff14",
5655 => x"54547233",
5656 => x"7434ff12",
5657 => x"5271ff2e",
5658 => x"0981060b",
5659 => x"0b0b0be8",
5660 => x"3875800c",
5661 => x"883d0d04",
5662 => x"768f260b",
5663 => x"0b0b0b9f",
5664 => x"38ff1252",
5665 => x"71ff2e0b",
5666 => x"0b0b0be5",
5667 => x"38727081",
5668 => x"05543374",
5669 => x"70810556",
5670 => x"340b0b0b",
5671 => x"0be33974",
5672 => x"76078306",
5673 => x"51700b0b",
5674 => x"0b0bd638",
5675 => x"75755451",
5676 => x"72708405",
5677 => x"54087170",
5678 => x"8405530c",
5679 => x"72708405",
5680 => x"54087170",
5681 => x"8405530c",
5682 => x"72708405",
5683 => x"54087170",
5684 => x"8405530c",
5685 => x"72708405",
5686 => x"54087170",
5687 => x"8405530c",
5688 => x"f0125271",
5689 => x"8f260b0b",
5690 => x"0b0bc538",
5691 => x"8372270b",
5692 => x"0b0b0b99",
5693 => x"38727084",
5694 => x"05540871",
5695 => x"70840553",
5696 => x"0cfc1252",
5697 => x"7183260b",
5698 => x"0b0b0be9",
5699 => x"3870540b",
5700 => x"0b0bfeed",
5701 => x"39fc3d0d",
5702 => x"76797102",
5703 => x"8c059f05",
5704 => x"33575553",
5705 => x"55837227",
5706 => x"0b0b0b0b",
5707 => x"8e387483",
5708 => x"06517080",
5709 => x"2e0b0b0b",
5710 => x"0baa38ff",
5711 => x"125271ff",
5712 => x"2e0b0b0b",
5713 => x"0b973873",
5714 => x"73708105",
5715 => x"5534ff12",
5716 => x"5271ff2e",
5717 => x"0981060b",
5718 => x"0b0b0beb",
5719 => x"3874800c",
5720 => x"863d0d04",
5721 => x"7474882b",
5722 => x"75077071",
5723 => x"902b0751",
5724 => x"54518f72",
5725 => x"270b0b0b",
5726 => x"0ba93872",
5727 => x"71708405",
5728 => x"530c7271",
5729 => x"70840553",
5730 => x"0c727170",
5731 => x"8405530c",
5732 => x"72717084",
5733 => x"05530cf0",
5734 => x"1252718f",
5735 => x"260b0b0b",
5736 => x"0bd93883",
5737 => x"72270b0b",
5738 => x"0b0b9438",
5739 => x"72717084",
5740 => x"05530cfc",
5741 => x"12527183",
5742 => x"260b0b0b",
5743 => x"0bee3870",
5744 => x"530b0b0b",
5745 => x"fef53904",
5746 => x"04f93d0d",
5747 => x"797b80cc",
5748 => x"12085658",
5749 => x"5673802e",
5750 => x"0b0b0b0b",
5751 => x"a9387610",
5752 => x"10147008",
5753 => x"55557380",
5754 => x"2e0b0b0b",
5755 => x"80c03873",
5756 => x"08750c80",
5757 => x"0b90150c",
5758 => x"800b8c15",
5759 => x"0c735574",
5760 => x"800c893d",
5761 => x"0d049053",
5762 => x"84527551",
5763 => x"0b0b0ba8",
5764 => x"c63f8008",
5765 => x"80cc170c",
5766 => x"80085580",
5767 => x"08802e0b",
5768 => x"0b0b0bdb",
5769 => x"38800854",
5770 => x"0b0b0bff",
5771 => x"b1398177",
5772 => x"2b701010",
5773 => x"94055458",
5774 => x"81527551",
5775 => x"0b0b0ba8",
5776 => x"963f8008",
5777 => x"80085654",
5778 => x"8008802e",
5779 => x"0b0b0bff",
5780 => x"ae387680",
5781 => x"0884050c",
5782 => x"77800888",
5783 => x"050c800b",
5784 => x"90150c80",
5785 => x"0b8c150c",
5786 => x"73550b0b",
5787 => x"0bff9039",
5788 => x"70707452",
5789 => x"71802e0b",
5790 => x"0b0b0b95",
5791 => x"38738413",
5792 => x"08101080",
5793 => x"cc120805",
5794 => x"7008740c",
5795 => x"73710c51",
5796 => x"51505004",
5797 => x"f53d0d7d",
5798 => x"7f616390",
5799 => x"13089414",
5800 => x"5b5d5b5c",
5801 => x"5c5c8057",
5802 => x"8216227a",
5803 => x"71291977",
5804 => x"227c7129",
5805 => x"72902a05",
5806 => x"70902a73",
5807 => x"83ffff06",
5808 => x"72848080",
5809 => x"29057b70",
5810 => x"84055d0c",
5811 => x"811c5c52",
5812 => x"535a5555",
5813 => x"7877240b",
5814 => x"0b0b0bcc",
5815 => x"3877802e",
5816 => x"0b0b0b0b",
5817 => x"9a387888",
5818 => x"1c08250b",
5819 => x"0b0b0b96",
5820 => x"38781010",
5821 => x"1b789412",
5822 => x"0c548119",
5823 => x"901c0c7a",
5824 => x"800c8d3d",
5825 => x"0d04841b",
5826 => x"08810552",
5827 => x"7b510b0b",
5828 => x"0bfdb63f",
5829 => x"8008901c",
5830 => x"08101088",
5831 => x"05548c1c",
5832 => x"5380088c",
5833 => x"0552540b",
5834 => x"0bfedcdf",
5835 => x"3f7a527b",
5836 => x"510b0b0b",
5837 => x"feba3f73",
5838 => x"79101011",
5839 => x"7994120c",
5840 => x"55811a90",
5841 => x"120c5b0b",
5842 => x"0b0bffb3",
5843 => x"39f63d0d",
5844 => x"7c7e6062",
5845 => x"890b8812",
5846 => x"355b5e5c",
5847 => x"59598056",
5848 => x"81557477",
5849 => x"250b0b0b",
5850 => x"0b903874",
5851 => x"10811757",
5852 => x"55767524",
5853 => x"0b0b0b0b",
5854 => x"f2387552",
5855 => x"78510b0b",
5856 => x"0bfcc63f",
5857 => x"80086180",
5858 => x"0894050c",
5859 => x"56810b80",
5860 => x"0890050c",
5861 => x"8957767a",
5862 => x"250b0b0b",
5863 => x"80e13876",
5864 => x"18587770",
5865 => x"81055933",
5866 => x"d005548a",
5867 => x"53755278",
5868 => x"510b0b0b",
5869 => x"fdde3f80",
5870 => x"08811858",
5871 => x"56797724",
5872 => x"0b0b0b0b",
5873 => x"dd388118",
5874 => x"58767b25",
5875 => x"0b0b0b0b",
5876 => x"a7387a77",
5877 => x"31577770",
5878 => x"81055933",
5879 => x"d005548a",
5880 => x"53755278",
5881 => x"510b0b0b",
5882 => x"fdaa3f80",
5883 => x"08ff1858",
5884 => x"56760b0b",
5885 => x"0b0bdf38",
5886 => x"75800c8c",
5887 => x"3d0d048a",
5888 => x"18580b0b",
5889 => x"0b0bc239",
5890 => x"70707074",
5891 => x"528072fc",
5892 => x"80800652",
5893 => x"5370732e",
5894 => x"0981060b",
5895 => x"0b0b0b87",
5896 => x"38907271",
5897 => x"2b535371",
5898 => x"81ff0a06",
5899 => x"51700b0b",
5900 => x"0b0b8838",
5901 => x"88137288",
5902 => x"2b535371",
5903 => x"8f0a0651",
5904 => x"700b0b0b",
5905 => x"0b883884",
5906 => x"1372842b",
5907 => x"53537183",
5908 => x"0a065170",
5909 => x"0b0b0b0b",
5910 => x"88388213",
5911 => x"72822b53",
5912 => x"53807224",
5913 => x"0b0b0b0b",
5914 => x"97388113",
5915 => x"729e2a70",
5916 => x"81065152",
5917 => x"53a05270",
5918 => x"802e0b0b",
5919 => x"0b0b8338",
5920 => x"72527180",
5921 => x"0c505050",
5922 => x"04fc3d0d",
5923 => x"76700870",
5924 => x"87065353",
5925 => x"5570802e",
5926 => x"0b0b0b0b",
5927 => x"b1387181",
5928 => x"06518053",
5929 => x"70732e09",
5930 => x"81060b0b",
5931 => x"0b0b9838",
5932 => x"710a100a",
5933 => x"70810652",
5934 => x"5370802e",
5935 => x"0b0b0b81",
5936 => x"89387275",
5937 => x"0c815372",
5938 => x"800c863d",
5939 => x"0d047072",
5940 => x"83ffff06",
5941 => x"52547080",
5942 => x"2e0b0b0b",
5943 => x"80e03871",
5944 => x"81ff0651",
5945 => x"700b0b0b",
5946 => x"0b883888",
5947 => x"1472882a",
5948 => x"5354718f",
5949 => x"0651700b",
5950 => x"0b0b0b88",
5951 => x"38841472",
5952 => x"842a5354",
5953 => x"71830651",
5954 => x"700b0b0b",
5955 => x"0b883882",
5956 => x"1472822a",
5957 => x"53547181",
5958 => x"0651700b",
5959 => x"0b0b0b94",
5960 => x"38811472",
5961 => x"0a100a53",
5962 => x"54a05371",
5963 => x"802e0b0b",
5964 => x"0bff9438",
5965 => x"71750c73",
5966 => x"800c863d",
5967 => x"0d049072",
5968 => x"712a5354",
5969 => x"0b0b0bff",
5970 => x"96397182",
5971 => x"2a750c82",
5972 => x"0b800c86",
5973 => x"3d0d0470",
5974 => x"70815273",
5975 => x"510b0b0b",
5976 => x"f8e73f74",
5977 => x"80089405",
5978 => x"0c810b80",
5979 => x"0890050c",
5980 => x"505004ee",
5981 => x"3d0d6567",
5982 => x"90120890",
5983 => x"12085856",
5984 => x"57537375",
5985 => x"250b0b0b",
5986 => x"0b8d3872",
5987 => x"76717790",
5988 => x"14085957",
5989 => x"58544274",
5990 => x"14708815",
5991 => x"08248415",
5992 => x"08055365",
5993 => x"525e0b0b",
5994 => x"0bf89e3f",
5995 => x"80088008",
5996 => x"94057060",
5997 => x"822b7211",
5998 => x"43465941",
5999 => x"427f7f27",
6000 => x"0b0b0b0b",
6001 => x"91388077",
6002 => x"70840559",
6003 => x"0c7e7726",
6004 => x"0b0b0b0b",
6005 => x"f1389413",
6006 => x"74101011",
6007 => x"94187710",
6008 => x"10116341",
6009 => x"445d5d5f",
6010 => x"7a61270b",
6011 => x"0b0b81c9",
6012 => x"387a0870",
6013 => x"83ffff06",
6014 => x"59537780",
6015 => x"2e0b0b0b",
6016 => x"80cb387e",
6017 => x"7d575780",
6018 => x"5a767084",
6019 => x"05580870",
6020 => x"83ffff06",
6021 => x"82182271",
6022 => x"7b29057c",
6023 => x"1173902a",
6024 => x"7c297a22",
6025 => x"5e7d0571",
6026 => x"902a0570",
6027 => x"902a5f59",
6028 => x"51515454",
6029 => x"74762372",
6030 => x"82172384",
6031 => x"16567b77",
6032 => x"260b0b0b",
6033 => x"0bc33879",
6034 => x"760c7a08",
6035 => x"5372902a",
6036 => x"5877802e",
6037 => x"0b0b0b80",
6038 => x"d1387e7d",
6039 => x"5757807d",
6040 => x"08705b56",
6041 => x"5a767084",
6042 => x"05580870",
6043 => x"83ffff06",
6044 => x"707a297b",
6045 => x"902a057c",
6046 => x"11515154",
6047 => x"54727623",
6048 => x"74821723",
6049 => x"84167490",
6050 => x"2a792971",
6051 => x"08821322",
6052 => x"5d5b7b05",
6053 => x"74902a05",
6054 => x"70902a5c",
6055 => x"56567b77",
6056 => x"260b0b0b",
6057 => x"ffbf3874",
6058 => x"760c841b",
6059 => x"841e5e5b",
6060 => x"607b260b",
6061 => x"0b0bfeb9",
6062 => x"38626005",
6063 => x"56807e25",
6064 => x"0b0b0b0b",
6065 => x"9838fc16",
6066 => x"5675080b",
6067 => x"0b0b0b8d",
6068 => x"38ff1e5e",
6069 => x"7d80240b",
6070 => x"0b0b0bea",
6071 => x"387d6290",
6072 => x"050c6180",
6073 => x"0c943d0d",
6074 => x"04f73d0d",
6075 => x"7b7d7f70",
6076 => x"83065858",
6077 => x"5a5a740b",
6078 => x"0b0b8181",
6079 => x"3875822c",
6080 => x"5675802e",
6081 => x"0b0b0b80",
6082 => x"cc3880c8",
6083 => x"1a087056",
6084 => x"5776802e",
6085 => x"0b0b0b81",
6086 => x"a3387581",
6087 => x"0655740b",
6088 => x"0b0b0bb8",
6089 => x"3875812c",
6090 => x"5675802e",
6091 => x"0b0b0b0b",
6092 => x"a4387608",
6093 => x"70595574",
6094 => x"802e0b0b",
6095 => x"0b80e038",
6096 => x"74577581",
6097 => x"06557480",
6098 => x"2e0b0b0b",
6099 => x"0bd7380b",
6100 => x"0b0b0b88",
6101 => x"3978800c",
6102 => x"8b3d0d04",
6103 => x"76537852",
6104 => x"79510b0b",
6105 => x"0bfc8c3f",
6106 => x"80087953",
6107 => x"7a52550b",
6108 => x"0b0bf5fc",
6109 => x"3f74590b",
6110 => x"0b0bffa9",
6111 => x"39805474",
6112 => x"10100b0b",
6113 => x"82f49c05",
6114 => x"70085455",
6115 => x"78527951",
6116 => x"0b0b0bf5",
6117 => x"ff3f8008",
6118 => x"590b0b0b",
6119 => x"fedf3976",
6120 => x"53765279",
6121 => x"510b0b0b",
6122 => x"fbc93f80",
6123 => x"08770c80",
6124 => x"08788008",
6125 => x"0c570b0b",
6126 => x"0bff8739",
6127 => x"84f15279",
6128 => x"510b0b0b",
6129 => x"fb913f80",
6130 => x"0880c81b",
6131 => x"0c800875",
6132 => x"80080c76",
6133 => x"81065657",
6134 => x"74802e0b",
6135 => x"0b0bfec5",
6136 => x"380b0b0b",
6137 => x"fef639f5",
6138 => x"3d0d7d7f",
6139 => x"6170852c",
6140 => x"84130890",
6141 => x"14081281",
6142 => x"05881508",
6143 => x"595e5959",
6144 => x"5a5c5c72",
6145 => x"79250b0b",
6146 => x"0b0b9038",
6147 => x"81157310",
6148 => x"54557873",
6149 => x"240b0b0b",
6150 => x"0bf23874",
6151 => x"527b510b",
6152 => x"0b0bf3a5",
6153 => x"3f800880",
6154 => x"08940555",
6155 => x"5a807625",
6156 => x"0b0b0b0b",
6157 => x"94387553",
6158 => x"80747084",
6159 => x"05560cff",
6160 => x"1353720b",
6161 => x"0b0b0bf0",
6162 => x"38941b90",
6163 => x"1c081010",
6164 => x"11799f06",
6165 => x"5a585377",
6166 => x"802e0b0b",
6167 => x"0b80ca38",
6168 => x"a0783155",
6169 => x"80567208",
6170 => x"782b7607",
6171 => x"74708405",
6172 => x"560c7270",
6173 => x"84055408",
6174 => x"752a5676",
6175 => x"73260b0b",
6176 => x"0b0be338",
6177 => x"75740c75",
6178 => x"802e0b0b",
6179 => x"0b0b8438",
6180 => x"811959ff",
6181 => x"19901b0c",
6182 => x"7a527b51",
6183 => x"0b0b0bf3",
6184 => x"cf3f7980",
6185 => x"0c8d3d0d",
6186 => x"04727084",
6187 => x"05540874",
6188 => x"70840556",
6189 => x"0c727727",
6190 => x"0b0b0b0b",
6191 => x"d6387270",
6192 => x"84055408",
6193 => x"74708405",
6194 => x"560c7673",
6195 => x"260b0b0b",
6196 => x"0bd7380b",
6197 => x"0b0bffbb",
6198 => x"39fb3d0d",
6199 => x"77799011",
6200 => x"08901308",
6201 => x"71317056",
6202 => x"54555754",
6203 => x"700b0b0b",
6204 => x"0bb33894",
6205 => x"1473822b",
6206 => x"71117119",
6207 => x"94055254",
6208 => x"5255fc12",
6209 => x"fc127108",
6210 => x"71085656",
6211 => x"52527373",
6212 => x"2e098106",
6213 => x"0b0b0b0b",
6214 => x"93387175",
6215 => x"260b0b0b",
6216 => x"0be03880",
6217 => x"5271800c",
6218 => x"873d0d04",
6219 => x"ff517274",
6220 => x"260b0b0b",
6221 => x"0b833881",
6222 => x"5170800c",
6223 => x"873d0d04",
6224 => x"f33d0d7f",
6225 => x"61637055",
6226 => x"71545754",
6227 => x"560b0b0b",
6228 => x"ff873f80",
6229 => x"08548008",
6230 => x"802e0b0b",
6231 => x"0b81e038",
6232 => x"80547380",
6233 => x"08240b0b",
6234 => x"0b81f638",
6235 => x"84130852",
6236 => x"75510b0b",
6237 => x"0bf0d23f",
6238 => x"80087480",
6239 => x"088c050c",
6240 => x"90140894",
6241 => x"15711010",
6242 => x"11941990",
6243 => x"1a081010",
6244 => x"11800894",
6245 => x"055d415d",
6246 => x"415a5c5d",
6247 => x"805a7770",
6248 => x"84055908",
6249 => x"7083ffff",
6250 => x"067a7084",
6251 => x"055c0870",
6252 => x"83ffff06",
6253 => x"7271311e",
6254 => x"74902a73",
6255 => x"902a3171",
6256 => x"902c1170",
6257 => x"902c4151",
6258 => x"55515657",
6259 => x"57547377",
6260 => x"23728218",
6261 => x"23841757",
6262 => x"7b79260b",
6263 => x"0b0bffbe",
6264 => x"38777e27",
6265 => x"0b0b0b0b",
6266 => x"b0387770",
6267 => x"84055908",
6268 => x"7083ffff",
6269 => x"067b1170",
6270 => x"902c7390",
6271 => x"2a057090",
6272 => x"2c5e5351",
6273 => x"54547377",
6274 => x"23728218",
6275 => x"23841757",
6276 => x"7d78260b",
6277 => x"0b0b0bd2",
6278 => x"38fc1757",
6279 => x"76080b0b",
6280 => x"0b0b9138",
6281 => x"ff1bfc18",
6282 => x"585b7608",
6283 => x"802e0b0b",
6284 => x"0b0bf138",
6285 => x"7a901e0c",
6286 => x"7c800c8f",
6287 => x"3d0d0480",
6288 => x"08527551",
6289 => x"0b0b0bef",
6290 => x"803f8008",
6291 => x"5d810b80",
6292 => x"0890050c",
6293 => x"73800894",
6294 => x"050c7c80",
6295 => x"0c8f3d0d",
6296 => x"04727554",
6297 => x"55810b84",
6298 => x"14085376",
6299 => x"52540b0b",
6300 => x"0beed63f",
6301 => x"80087480",
6302 => x"088c050c",
6303 => x"90140894",
6304 => x"15711010",
6305 => x"11941990",
6306 => x"1a081010",
6307 => x"11800894",
6308 => x"055d415d",
6309 => x"415a5c5d",
6310 => x"805a0b0b",
6311 => x"0bfdff39",
6312 => x"fa3d0d78",
6313 => x"7a7c5457",
6314 => x"7258769f",
6315 => x"fe0a0686",
6316 => x"bf0a0553",
6317 => x"53807225",
6318 => x"0b0b0b0b",
6319 => x"95387154",
6320 => x"80557375",
6321 => x"53730c71",
6322 => x"84140c72",
6323 => x"800c883d",
6324 => x"0d047130",
6325 => x"70942c53",
6326 => x"51937225",
6327 => x"0b0b0b0b",
6328 => x"ab388054",
6329 => x"ec129f71",
6330 => x"3181712b",
6331 => x"5152529e",
6332 => x"72250b0b",
6333 => x"0b0b8338",
6334 => x"81517055",
6335 => x"73755373",
6336 => x"0c718414",
6337 => x"0c72800c",
6338 => x"883d0d04",
6339 => x"a0808072",
6340 => x"2c548055",
6341 => x"0b0b0bff",
6342 => x"a939f63d",
6343 => x"0d7c7e94",
6344 => x"11901208",
6345 => x"101011fc",
6346 => x"11700870",
6347 => x"575a5157",
6348 => x"5853590b",
6349 => x"0b0bf1d0",
6350 => x"3f80087f",
6351 => x"a00b8008",
6352 => x"31710c53",
6353 => x"538a0b80",
6354 => x"08250b0b",
6355 => x"0b80f738",
6356 => x"80577376",
6357 => x"260b0b0b",
6358 => x"80c438f5",
6359 => x"13537280",
6360 => x"2e0b0b0b",
6361 => x"80c838a0",
6362 => x"73317574",
6363 => x"2b78722a",
6364 => x"079ffc0a",
6365 => x"075b5880",
6366 => x"55757427",
6367 => x"0b0b0b0b",
6368 => x"8538fc14",
6369 => x"08557673",
6370 => x"2b75792a",
6371 => x"075b797b",
6372 => x"54790c72",
6373 => x"841a0c78",
6374 => x"800c8c3d",
6375 => x"0d04fc14",
6376 => x"7008f515",
6377 => x"55585472",
6378 => x"0b0b0bff",
6379 => x"ba38749f",
6380 => x"fc0a075a",
6381 => x"765b797b",
6382 => x"54790c72",
6383 => x"841a0c78",
6384 => x"800c8c3d",
6385 => x"0d048b0b",
6386 => x"80083175",
6387 => x"712a9ffc",
6388 => x"0a075b57",
6389 => x"80587574",
6390 => x"270b0b0b",
6391 => x"0b8538fc",
6392 => x"14085895",
6393 => x"1375712b",
6394 => x"79792a07",
6395 => x"5c52797b",
6396 => x"54790c72",
6397 => x"841a0c78",
6398 => x"800c8c3d",
6399 => x"0d04f33d",
6400 => x"0d626462",
6401 => x"64575f75",
6402 => x"405b5981",
6403 => x"527f510b",
6404 => x"0b0bebb5",
6405 => x"3f800880",
6406 => x"0894057e",
6407 => x"70bfffff",
6408 => x"06705f71",
6409 => x"fe0a0670",
6410 => x"4270942a",
6411 => x"5b525755",
6412 => x"59577580",
6413 => x"2e0b0b0b",
6414 => x"0b873873",
6415 => x"90800a07",
6416 => x"5b7d5372",
6417 => x"802e0b0b",
6418 => x"0b80e038",
6419 => x"725c8f3d",
6420 => x"f405510b",
6421 => x"0b0bf0b1",
6422 => x"3f800855",
6423 => x"8008802e",
6424 => x"0b0b0b81",
6425 => x"8d38a00b",
6426 => x"8008317b",
6427 => x"712b7d07",
6428 => x"790c537a",
6429 => x"80082a5b",
6430 => x"7a70841a",
6431 => x"0c703070",
6432 => x"72078025",
6433 => x"82713170",
6434 => x"901c0c51",
6435 => x"51545475",
6436 => x"802e0b0b",
6437 => x"0b0bb638",
6438 => x"7416f7cd",
6439 => x"05790cb5",
6440 => x"75317a0c",
6441 => x"76800c8f",
6442 => x"3d0d048f",
6443 => x"3df00551",
6444 => x"0b0b0bef",
6445 => x"d43f7a78",
6446 => x"0c810b90",
6447 => x"180c810b",
6448 => x"8008a005",
6449 => x"5653750b",
6450 => x"0b0b0bcc",
6451 => x"38f7ce15",
6452 => x"790c7285",
6453 => x"2b731010",
6454 => x"19fc1108",
6455 => x"5354540b",
6456 => x"0b0beea4",
6457 => x"3f738008",
6458 => x"317a0c76",
6459 => x"800c8f3d",
6460 => x"0d047b78",
6461 => x"0c7a7084",
6462 => x"1a0c7030",
6463 => x"70720780",
6464 => x"25827131",
6465 => x"70901c0c",
6466 => x"51515454",
6467 => x"0b0b0bfe",
6468 => x"fe39f03d",
6469 => x"0d626466",
6470 => x"953de411",
6471 => x"577256f8",
6472 => x"05545858",
6473 => x"580b0b0b",
6474 => x"fbf03f92",
6475 => x"3de01154",
6476 => x"7653f005",
6477 => x"510b0b0b",
6478 => x"fbe03f90",
6479 => x"17089017",
6480 => x"0831852b",
6481 => x"7b7b3111",
6482 => x"51568076",
6483 => x"250b0b0b",
6484 => x"0bb03875",
6485 => x"90800a29",
6486 => x"6005407d",
6487 => x"7f585476",
6488 => x"557f6158",
6489 => x"52765392",
6490 => x"3de80551",
6491 => x"0b0b80d6",
6492 => x"ac3f7b7d",
6493 => x"58780c76",
6494 => x"84190c77",
6495 => x"800c923d",
6496 => x"0d047530",
6497 => x"7090800a",
6498 => x"291f5f56",
6499 => x"7d7f5854",
6500 => x"76557f61",
6501 => x"58527653",
6502 => x"923de805",
6503 => x"510b0b80",
6504 => x"d5fb3f7b",
6505 => x"7d58780c",
6506 => x"7684190c",
6507 => x"77800c92",
6508 => x"3d0d04f3",
6509 => x"3d0d7f61",
6510 => x"575c9ffc",
6511 => x"0a578058",
6512 => x"7597240b",
6513 => x"0b0b0b9d",
6514 => x"38751010",
6515 => x"100b0b82",
6516 => x"f2d80584",
6517 => x"11087108",
6518 => x"7e0c841e",
6519 => x"0c7c800c",
6520 => x"568f3d0d",
6521 => x"04807625",
6522 => x"0b0b0b0b",
6523 => x"ab388d3d",
6524 => x"5b80c882",
6525 => x"0a59805a",
6526 => x"78547955",
6527 => x"76527753",
6528 => x"7a510b0b",
6529 => x"0bb6963f",
6530 => x"7c7eff18",
6531 => x"58595775",
6532 => x"80240b0b",
6533 => x"0b0be138",
6534 => x"767c0c77",
6535 => x"841d0c7b",
6536 => x"800c8f3d",
6537 => x"0d04ef3d",
6538 => x"0d636567",
6539 => x"405d427b",
6540 => x"802e0b0b",
6541 => x"0b85ea38",
6542 => x"61510b0b",
6543 => x"0be7883f",
6544 => x"f81c7084",
6545 => x"120870fc",
6546 => x"0670628b",
6547 => x"0570f806",
6548 => x"4159455b",
6549 => x"5c415796",
6550 => x"74270b0b",
6551 => x"0b82fe38",
6552 => x"807b247e",
6553 => x"7c260759",
6554 => x"80547874",
6555 => x"2e098106",
6556 => x"0b0b0b82",
6557 => x"e138777b",
6558 => x"250b0b0b",
6559 => x"82ab3877",
6560 => x"170b0b82",
6561 => x"fcc80b88",
6562 => x"05085e56",
6563 => x"7c762e0b",
6564 => x"0b0b859f",
6565 => x"38841608",
6566 => x"70fe0617",
6567 => x"84110881",
6568 => x"06515555",
6569 => x"730b0b0b",
6570 => x"82bb3874",
6571 => x"fc06597c",
6572 => x"762e0b0b",
6573 => x"0b85c938",
6574 => x"77195f7e",
6575 => x"7b250b0b",
6576 => x"0b82aa38",
6577 => x"79810654",
6578 => x"730b0b0b",
6579 => x"82f53876",
6580 => x"77083184",
6581 => x"1108fc06",
6582 => x"565a7580",
6583 => x"2e0b0b0b",
6584 => x"0b97387c",
6585 => x"762e0b0b",
6586 => x"0b85d438",
6587 => x"74191859",
6588 => x"787b250b",
6589 => x"0b0b84e2",
6590 => x"3879802e",
6591 => x"0b0b0b82",
6592 => x"c2387715",
6593 => x"567a7624",
6594 => x"0b0b0b82",
6595 => x"b6388c1a",
6596 => x"08881b08",
6597 => x"718c120c",
6598 => x"88120c55",
6599 => x"79765957",
6600 => x"881761fc",
6601 => x"05575975",
6602 => x"a4260b0b",
6603 => x"0b86e638",
6604 => x"7b795555",
6605 => x"9376270b",
6606 => x"0b0b80d1",
6607 => x"387b7084",
6608 => x"055d087c",
6609 => x"56790c74",
6610 => x"70840556",
6611 => x"088c180c",
6612 => x"9017549b",
6613 => x"76270b0b",
6614 => x"0b0bb238",
6615 => x"74708405",
6616 => x"5608740c",
6617 => x"74708405",
6618 => x"56089418",
6619 => x"0c981754",
6620 => x"a376270b",
6621 => x"0b0b0b95",
6622 => x"38747084",
6623 => x"05560874",
6624 => x"0c747084",
6625 => x"0556089c",
6626 => x"180ca017",
6627 => x"54747084",
6628 => x"05560874",
6629 => x"70840556",
6630 => x"0c747084",
6631 => x"05560874",
6632 => x"70840556",
6633 => x"0c740874",
6634 => x"0c777b31",
6635 => x"56758f26",
6636 => x"0b0b0b80",
6637 => x"d5388417",
6638 => x"08810678",
6639 => x"0784180c",
6640 => x"77178411",
6641 => x"08810784",
6642 => x"120c5461",
6643 => x"510b0b0b",
6644 => x"e3f63f88",
6645 => x"17547380",
6646 => x"0c933d0d",
6647 => x"04905b0b",
6648 => x"0b0bfcfc",
6649 => x"3978560b",
6650 => x"0b0bfdd8",
6651 => x"398c1608",
6652 => x"88170871",
6653 => x"8c120c88",
6654 => x"120c557e",
6655 => x"707c3157",
6656 => x"588f7627",
6657 => x"0b0b0bff",
6658 => x"ad387a17",
6659 => x"84180881",
6660 => x"067c0784",
6661 => x"190c7681",
6662 => x"0784120c",
6663 => x"76118411",
6664 => x"08810784",
6665 => x"120c5588",
6666 => x"05526151",
6667 => x"0b0bffbc",
6668 => x"873f6151",
6669 => x"0b0b0be3",
6670 => x"8f3f8817",
6671 => x"540b0b0b",
6672 => x"ff94397d",
6673 => x"5261510b",
6674 => x"0b0bcef6",
6675 => x"3f800859",
6676 => x"8008802e",
6677 => x"0b0b0b81",
6678 => x"b7388008",
6679 => x"f8056084",
6680 => x"0508fe06",
6681 => x"61055557",
6682 => x"76742e0b",
6683 => x"0b0b84b7",
6684 => x"38fc1856",
6685 => x"75a4260b",
6686 => x"0b0b81c1",
6687 => x"387b8008",
6688 => x"55559376",
6689 => x"270b0b0b",
6690 => x"80e03874",
6691 => x"70840556",
6692 => x"08800870",
6693 => x"8405800c",
6694 => x"0c800875",
6695 => x"70840557",
6696 => x"08717084",
6697 => x"05530c54",
6698 => x"9b76270b",
6699 => x"0b0b0bba",
6700 => x"38747084",
6701 => x"05560874",
6702 => x"70840556",
6703 => x"0c747084",
6704 => x"05560874",
6705 => x"70840556",
6706 => x"0ca37627",
6707 => x"0b0b0b0b",
6708 => x"99387470",
6709 => x"84055608",
6710 => x"74708405",
6711 => x"560c7470",
6712 => x"84055608",
6713 => x"74708405",
6714 => x"560c7470",
6715 => x"84055608",
6716 => x"74708405",
6717 => x"560c7470",
6718 => x"84055608",
6719 => x"74708405",
6720 => x"560c7408",
6721 => x"740c7b52",
6722 => x"61510b0b",
6723 => x"ffbaa93f",
6724 => x"61510b0b",
6725 => x"0be1b13f",
6726 => x"78547380",
6727 => x"0c933d0d",
6728 => x"047d5261",
6729 => x"510b0b0b",
6730 => x"cd983f80",
6731 => x"08800c93",
6732 => x"3d0d0484",
6733 => x"1608550b",
6734 => x"0b0bfaef",
6735 => x"3975537b",
6736 => x"52800851",
6737 => x"0b0bfec0",
6738 => x"c23f7b52",
6739 => x"61510b0b",
6740 => x"ffb9e53f",
6741 => x"0b0b0bff",
6742 => x"b7398c16",
6743 => x"08881708",
6744 => x"718c120c",
6745 => x"88120c55",
6746 => x"8c1a0888",
6747 => x"1b08718c",
6748 => x"120c8812",
6749 => x"0c557979",
6750 => x"59570b0b",
6751 => x"0bfba139",
6752 => x"7719901c",
6753 => x"55557375",
6754 => x"240b0b0b",
6755 => x"fab6387a",
6756 => x"17700b0b",
6757 => x"82fcc80b",
6758 => x"88050c75",
6759 => x"7c318107",
6760 => x"84120c5d",
6761 => x"84170881",
6762 => x"067b0784",
6763 => x"180c6151",
6764 => x"0b0b0be0",
6765 => x"933f8817",
6766 => x"540b0b0b",
6767 => x"fc983974",
6768 => x"1918901c",
6769 => x"555d737d",
6770 => x"240b0b0b",
6771 => x"faab388c",
6772 => x"1a08881b",
6773 => x"08718c12",
6774 => x"0c88120c",
6775 => x"55881a61",
6776 => x"fc055759",
6777 => x"75a4260b",
6778 => x"0b0b81ca",
6779 => x"387b7955",
6780 => x"55937627",
6781 => x"0b0b0b80",
6782 => x"d1387b70",
6783 => x"84055d08",
6784 => x"7c56790c",
6785 => x"74708405",
6786 => x"56088c1b",
6787 => x"0c901a54",
6788 => x"9b76270b",
6789 => x"0b0b0bb2",
6790 => x"38747084",
6791 => x"05560874",
6792 => x"0c747084",
6793 => x"05560894",
6794 => x"1b0c981a",
6795 => x"54a37627",
6796 => x"0b0b0b0b",
6797 => x"95387470",
6798 => x"84055608",
6799 => x"740c7470",
6800 => x"84055608",
6801 => x"9c1b0ca0",
6802 => x"1a547470",
6803 => x"84055608",
6804 => x"74708405",
6805 => x"560c7470",
6806 => x"84055608",
6807 => x"74708405",
6808 => x"560c7408",
6809 => x"740c7a1a",
6810 => x"700b0b82",
6811 => x"fcc80b88",
6812 => x"050c7d7c",
6813 => x"31810784",
6814 => x"120c5484",
6815 => x"1a088106",
6816 => x"7b07841b",
6817 => x"0c61510b",
6818 => x"0b0bdebc",
6819 => x"3f78540b",
6820 => x"0b0bfd86",
6821 => x"3975537b",
6822 => x"5278510b",
6823 => x"0bfebdeb",
6824 => x"3f0b0b0b",
6825 => x"fa833984",
6826 => x"1708fc06",
6827 => x"18605858",
6828 => x"0b0b0bf9",
6829 => x"f4397553",
6830 => x"7b527851",
6831 => x"0b0bfebd",
6832 => x"ca3f7a1a",
6833 => x"700b0b82",
6834 => x"fcc80b88",
6835 => x"050c7d7c",
6836 => x"31810784",
6837 => x"120c5484",
6838 => x"1a088106",
6839 => x"7b07841b",
6840 => x"0c0b0b0b",
6841 => x"ff9f3970",
6842 => x"70707075",
6843 => x"77535371",
6844 => x"54733070",
6845 => x"75079f2a",
6846 => x"7075fe0a",
6847 => x"06079081",
6848 => x"0a119ffe",
6849 => x"0a723107",
6850 => x"709f2a81",
6851 => x"7131800c",
6852 => x"51515151",
6853 => x"51505050",
6854 => x"50047070",
6855 => x"70707577",
6856 => x"53537154",
6857 => x"73307075",
6858 => x"079f2a70",
6859 => x"75fe0a06",
6860 => x"079ffe0a",
6861 => x"71319f2a",
6862 => x"800c5151",
6863 => x"51505050",
6864 => x"50047070",
6865 => x"7070800b",
6866 => x"0b0b8385",
6867 => x"840c7651",
6868 => x"0b0b0b8c",
6869 => x"f33f8008",
6870 => x"538008ff",
6871 => x"2e0b0b0b",
6872 => x"0b893872",
6873 => x"800c5050",
6874 => x"5050040b",
6875 => x"0b838584",
6876 => x"08547380",
6877 => x"2e0b0b0b",
6878 => x"0be93875",
6879 => x"74710c52",
6880 => x"72800c50",
6881 => x"50505004",
6882 => x"f93d0d79",
6883 => x"7c557b54",
6884 => x"8e112270",
6885 => x"902b7090",
6886 => x"2c55570b",
6887 => x"0b82f4ec",
6888 => x"08535856",
6889 => x"0b0b0b88",
6890 => x"ac3f8008",
6891 => x"57800b80",
6892 => x"08240b0b",
6893 => x"0b0b9338",
6894 => x"80d01608",
6895 => x"80080580",
6896 => x"d0170c76",
6897 => x"800c893d",
6898 => x"0d048c16",
6899 => x"2283dfff",
6900 => x"0655748c",
6901 => x"17237680",
6902 => x"0c893d0d",
6903 => x"04fa3d0d",
6904 => x"788c1122",
6905 => x"70882a70",
6906 => x"81065157",
6907 => x"5856740b",
6908 => x"0b0b0bae",
6909 => x"388c1622",
6910 => x"83dfff06",
6911 => x"55748c17",
6912 => x"237a5479",
6913 => x"538e1622",
6914 => x"70902b70",
6915 => x"902c5456",
6916 => x"0b0b82f4",
6917 => x"ec085256",
6918 => x"0b0b0b83",
6919 => x"f33f883d",
6920 => x"0d048254",
6921 => x"80538e16",
6922 => x"2270902b",
6923 => x"70902c54",
6924 => x"560b0b82",
6925 => x"f4ec0852",
6926 => x"570b0b0b",
6927 => x"86d03f8c",
6928 => x"162283df",
6929 => x"ff065574",
6930 => x"8c17237a",
6931 => x"5479538e",
6932 => x"16227090",
6933 => x"2b70902c",
6934 => x"54560b0b",
6935 => x"82f4ec08",
6936 => x"52560b0b",
6937 => x"0b83a93f",
6938 => x"883d0d04",
6939 => x"f93d0d79",
6940 => x"7c557b54",
6941 => x"8e112270",
6942 => x"902b7090",
6943 => x"2c55570b",
6944 => x"0b82f4ec",
6945 => x"08535856",
6946 => x"0b0b0b86",
6947 => x"813f8008",
6948 => x"578008ff",
6949 => x"2e0b0b0b",
6950 => x"0b99388c",
6951 => x"1622a080",
6952 => x"0755748c",
6953 => x"17238008",
6954 => x"80d0170c",
6955 => x"76800c89",
6956 => x"3d0d048c",
6957 => x"162283df",
6958 => x"ff065574",
6959 => x"8c172376",
6960 => x"800c893d",
6961 => x"0d047070",
6962 => x"70748e11",
6963 => x"2270902b",
6964 => x"70902c55",
6965 => x"5151530b",
6966 => x"0b82f4ec",
6967 => x"08510b0b",
6968 => x"0b84a03f",
6969 => x"50505004",
6970 => x"fb3d0d77",
6971 => x"79707207",
6972 => x"83065354",
6973 => x"52700b0b",
6974 => x"0b0b9638",
6975 => x"71737308",
6976 => x"54565471",
6977 => x"73082e0b",
6978 => x"0b0b80d0",
6979 => x"38737554",
6980 => x"52713370",
6981 => x"81ff0652",
6982 => x"5470802e",
6983 => x"0b0b0b0b",
6984 => x"a5387233",
6985 => x"5570752e",
6986 => x"0981060b",
6987 => x"0b0b0b99",
6988 => x"38811281",
6989 => x"14713370",
6990 => x"81ff0654",
6991 => x"56545270",
6992 => x"0b0b0b0b",
6993 => x"dd387233",
6994 => x"557381ff",
6995 => x"067581ff",
6996 => x"06717131",
6997 => x"800c5252",
6998 => x"873d0d04",
6999 => x"710970f7",
7000 => x"fbfdff14",
7001 => x"0670f884",
7002 => x"82818006",
7003 => x"51515170",
7004 => x"0b0b0b0b",
7005 => x"9e388414",
7006 => x"84167108",
7007 => x"54565471",
7008 => x"75082e0b",
7009 => x"0b0b0bd4",
7010 => x"38737554",
7011 => x"520b0b0b",
7012 => x"feff3980",
7013 => x"0b800c87",
7014 => x"3d0d0470",
7015 => x"70707075",
7016 => x"70718306",
7017 => x"53555270",
7018 => x"0b0b0b80",
7019 => x"c0387170",
7020 => x"087009f7",
7021 => x"fbfdff12",
7022 => x"0670f884",
7023 => x"82818006",
7024 => x"51515253",
7025 => x"700b0b0b",
7026 => x"0ba13884",
7027 => x"13700870",
7028 => x"09f7fbfd",
7029 => x"ff120670",
7030 => x"f8848281",
7031 => x"80065151",
7032 => x"52537080",
7033 => x"2e0b0b0b",
7034 => x"0be13872",
7035 => x"52713351",
7036 => x"70802e0b",
7037 => x"0b0b0b8e",
7038 => x"38811270",
7039 => x"33525270",
7040 => x"0b0b0b0b",
7041 => x"f4387174",
7042 => x"31800c50",
7043 => x"50505004",
7044 => x"fb3d0d80",
7045 => x"0b0b0b83",
7046 => x"85840c7a",
7047 => x"53795278",
7048 => x"510b0b0b",
7049 => x"88de3f80",
7050 => x"08558008",
7051 => x"ff2e0b0b",
7052 => x"0b0b8838",
7053 => x"74800c87",
7054 => x"3d0d040b",
7055 => x"0b838584",
7056 => x"08567580",
7057 => x"2e0b0b0b",
7058 => x"0bea3877",
7059 => x"76710c54",
7060 => x"74800c87",
7061 => x"3d0d04fb",
7062 => x"3d0d787a",
7063 => x"29527751",
7064 => x"0b0b0bc2",
7065 => x"dd3f8008",
7066 => x"80085556",
7067 => x"8008802e",
7068 => x"0b0b0b80",
7069 => x"f2388008",
7070 => x"fc0508fc",
7071 => x"06fc0555",
7072 => x"74a4260b",
7073 => x"0b0b80e6",
7074 => x"38937527",
7075 => x"0b0b0b80",
7076 => x"c338800b",
7077 => x"80087084",
7078 => x"05800c0c",
7079 => x"80085480",
7080 => x"74708405",
7081 => x"560c9b75",
7082 => x"270b0b0b",
7083 => x"0ba63880",
7084 => x"74708405",
7085 => x"560c8074",
7086 => x"70840556",
7087 => x"0ca37527",
7088 => x"0b0b0b0b",
7089 => x"8f388074",
7090 => x"70840556",
7091 => x"0c807470",
7092 => x"8405560c",
7093 => x"80747084",
7094 => x"05560c80",
7095 => x"74708405",
7096 => x"560c8074",
7097 => x"0c755473",
7098 => x"800c873d",
7099 => x"0d047453",
7100 => x"80528008",
7101 => x"510b0b0b",
7102 => x"d49b3f75",
7103 => x"540b0b0b",
7104 => x"0be53970",
7105 => x"70707080",
7106 => x"0b0b0b83",
7107 => x"85840c76",
7108 => x"510b0b0b",
7109 => x"8a943f80",
7110 => x"08538008",
7111 => x"ff2e0b0b",
7112 => x"0b0b8938",
7113 => x"72800c50",
7114 => x"50505004",
7115 => x"0b0b8385",
7116 => x"84085473",
7117 => x"802e0b0b",
7118 => x"0b0be938",
7119 => x"7574710c",
7120 => x"5272800c",
7121 => x"50505050",
7122 => x"04fc3d0d",
7123 => x"800b0b0b",
7124 => x"8385840c",
7125 => x"78527751",
7126 => x"0b0b0b8d",
7127 => x"823f8008",
7128 => x"548008ff",
7129 => x"2e0b0b0b",
7130 => x"0b883873",
7131 => x"800c863d",
7132 => x"0d040b0b",
7133 => x"83858408",
7134 => x"5574802e",
7135 => x"0b0b0b0b",
7136 => x"ea387675",
7137 => x"710c5373",
7138 => x"800c863d",
7139 => x"0d04fb3d",
7140 => x"0d800b0b",
7141 => x"0b838584",
7142 => x"0c7a5379",
7143 => x"5278510b",
7144 => x"0b0b8a9e",
7145 => x"3f800855",
7146 => x"8008ff2e",
7147 => x"0b0b0b0b",
7148 => x"88387480",
7149 => x"0c873d0d",
7150 => x"040b0b83",
7151 => x"85840856",
7152 => x"75802e0b",
7153 => x"0b0b0bea",
7154 => x"38777671",
7155 => x"0c547480",
7156 => x"0c873d0d",
7157 => x"04fb3d0d",
7158 => x"800b0b0b",
7159 => x"8385840c",
7160 => x"7a537952",
7161 => x"78510b0b",
7162 => x"0b86b13f",
7163 => x"80085580",
7164 => x"08ff2e0b",
7165 => x"0b0b0b88",
7166 => x"3874800c",
7167 => x"873d0d04",
7168 => x"0b0b8385",
7169 => x"84085675",
7170 => x"802e0b0b",
7171 => x"0b0bea38",
7172 => x"7776710c",
7173 => x"5474800c",
7174 => x"873d0d04",
7175 => x"fc3d0d76",
7176 => x"78700855",
7177 => x"5555720b",
7178 => x"0b0b0b8f",
7179 => x"38735274",
7180 => x"510b0bff",
7181 => x"ac823f86",
7182 => x"3d0d0472",
7183 => x"5274510b",
7184 => x"0b0b0bd8",
7185 => x"3f735274",
7186 => x"510b0bff",
7187 => x"abea3f86",
7188 => x"3d0d04fb",
7189 => x"3d0d7755",
7190 => x"740b0b82",
7191 => x"f4ec082e",
7192 => x"0b0b0b80",
7193 => x"fe3880cc",
7194 => x"15085380",
7195 => x"5672762e",
7196 => x"0981060b",
7197 => x"0b0b8180",
7198 => x"3882c815",
7199 => x"08537280",
7200 => x"2e0b0b0b",
7201 => x"0bb23882",
7202 => x"cc155672",
7203 => x"762e0b0b",
7204 => x"0b0ba538",
7205 => x"72547574",
7206 => x"2e0b0b0b",
7207 => x"0b9a3873",
7208 => x"74085552",
7209 => x"74510b0b",
7210 => x"ffab8d3f",
7211 => x"75742e09",
7212 => x"81060b0b",
7213 => x"0b0be838",
7214 => x"80d41508",
7215 => x"53720b0b",
7216 => x"0b80d938",
7217 => x"b8150880",
7218 => x"2e0b0b0b",
7219 => x"0b953874",
7220 => x"51bc1508",
7221 => x"53722d84",
7222 => x"dc150853",
7223 => x"720b0b0b",
7224 => x"80ca3887",
7225 => x"3d0d0481",
7226 => x"1656758e",
7227 => x"240b0b0b",
7228 => x"80c83880",
7229 => x"cc150853",
7230 => x"75101013",
7231 => x"70085553",
7232 => x"73802e0b",
7233 => x"0b0b0bdf",
7234 => x"38737408",
7235 => x"55527451",
7236 => x"0b0bffaa",
7237 => x"a33f0b0b",
7238 => x"0b0be539",
7239 => x"72527451",
7240 => x"0b0bffaa",
7241 => x"933f0b0b",
7242 => x"0bff9939",
7243 => x"72527451",
7244 => x"0b0b0bfd",
7245 => x"e73f873d",
7246 => x"0d0480cc",
7247 => x"15085274",
7248 => x"510b0bff",
7249 => x"a9f23f0b",
7250 => x"0b0bfead",
7251 => x"39fb3d0d",
7252 => x"77567580",
7253 => x"2e0b0b0b",
7254 => x"80dc3882",
7255 => x"c8160855",
7256 => x"74802e0b",
7257 => x"0b0b0bb5",
7258 => x"38841508",
7259 => x"ff055480",
7260 => x"74240b0b",
7261 => x"0b0b9c38",
7262 => x"73101015",
7263 => x"88055372",
7264 => x"08fc1454",
7265 => x"52712dff",
7266 => x"14547380",
7267 => x"250b0b0b",
7268 => x"0bed3874",
7269 => x"0855740b",
7270 => x"0b0b0bcd",
7271 => x"38bc1608",
7272 => x"0b0b0b0b",
7273 => x"8538873d",
7274 => x"0d047551",
7275 => x"bc160852",
7276 => x"712d873d",
7277 => x"0d040b0b",
7278 => x"82f4ec08",
7279 => x"82c81108",
7280 => x"56560b0b",
7281 => x"0bff9939",
7282 => x"7070700b",
7283 => x"0b8384fc",
7284 => x"080b0b0b",
7285 => x"0b8d380b",
7286 => x"0b838588",
7287 => x"0b0b0b83",
7288 => x"84fc0c0b",
7289 => x"0b8384fc",
7290 => x"08751152",
7291 => x"52ff5370",
7292 => x"0b87fb80",
7293 => x"80260b0b",
7294 => x"0b0b8a38",
7295 => x"700b0b83",
7296 => x"84fc0c71",
7297 => x"5372800c",
7298 => x"50505004",
7299 => x"fd3d0d80",
7300 => x"0b0b0b82",
7301 => x"f4e00854",
7302 => x"5472812e",
7303 => x"0b0b0b0b",
7304 => x"ab38730b",
7305 => x"0b838580",
7306 => x"0c0b0bfe",
7307 => x"a5853f0b",
7308 => x"0bfea3cc",
7309 => x"3f0b0b83",
7310 => x"84d05281",
7311 => x"510b0bfe",
7312 => x"a7dd3f80",
7313 => x"08510b0b",
7314 => x"0b89973f",
7315 => x"720b0b83",
7316 => x"85800c0b",
7317 => x"0bfea4db",
7318 => x"3f0b0bfe",
7319 => x"a3a23f0b",
7320 => x"0b8384d0",
7321 => x"5281510b",
7322 => x"0bfea7b3",
7323 => x"3f800851",
7324 => x"0b0b0b88",
7325 => x"ed3f000b",
7326 => x"0b0b0bfb",
7327 => x"39000b0b",
7328 => x"0b0bfb39",
7329 => x"f53d0d7e",
7330 => x"600b0b83",
7331 => x"85800870",
7332 => x"5b585b5b",
7333 => x"750b0b0b",
7334 => x"80db3877",
7335 => x"7a250b0b",
7336 => x"0b0bac38",
7337 => x"771b7033",
7338 => x"7081ff06",
7339 => x"58585975",
7340 => x"8a2e0b0b",
7341 => x"0b0b9f38",
7342 => x"7681ff06",
7343 => x"510b0bfe",
7344 => x"a3cc3f81",
7345 => x"18587978",
7346 => x"240b0b0b",
7347 => x"0bd63879",
7348 => x"800c8d3d",
7349 => x"0d048d51",
7350 => x"0b0bfea3",
7351 => x"b13f7833",
7352 => x"7081ff06",
7353 => x"52570b0b",
7354 => x"fea3a33f",
7355 => x"8118580b",
7356 => x"0b0b0bd2",
7357 => x"3979557a",
7358 => x"547d5385",
7359 => x"528d3dfc",
7360 => x"05510b0b",
7361 => x"fea2c03f",
7362 => x"8008560b",
7363 => x"0b0b87c9",
7364 => x"3f7b8008",
7365 => x"0c75800c",
7366 => x"8d3d0d04",
7367 => x"f63d0d7d",
7368 => x"7f0b0b83",
7369 => x"85800870",
7370 => x"5b585a5a",
7371 => x"750b0b0b",
7372 => x"80d63877",
7373 => x"79250b0b",
7374 => x"0b80c438",
7375 => x"0b0bfea2",
7376 => x"a43f8008",
7377 => x"81ff0670",
7378 => x"8d327030",
7379 => x"709f2a51",
7380 => x"51575776",
7381 => x"8a2e0b0b",
7382 => x"0b80d438",
7383 => x"75802e0b",
7384 => x"0b0b80cb",
7385 => x"38771a56",
7386 => x"76763476",
7387 => x"510b0bfe",
7388 => x"a29c3f81",
7389 => x"18587878",
7390 => x"240b0b0b",
7391 => x"ffbe3877",
7392 => x"5675800c",
7393 => x"8c3d0d04",
7394 => x"78557954",
7395 => x"7c538452",
7396 => x"8c3dfc05",
7397 => x"510b0bfe",
7398 => x"a1ad3f80",
7399 => x"08560b0b",
7400 => x"0b86b63f",
7401 => x"7a80080c",
7402 => x"75800c8c",
7403 => x"3d0d0477",
7404 => x"1a568a76",
7405 => x"34811858",
7406 => x"8d510b0b",
7407 => x"fea1cf3f",
7408 => x"8a510b0b",
7409 => x"fea1c73f",
7410 => x"77560b0b",
7411 => x"0bffb239",
7412 => x"f93d0d79",
7413 => x"570b0b83",
7414 => x"85800880",
7415 => x"2e0b0b0b",
7416 => x"0bb53876",
7417 => x"510b0b0b",
7418 => x"f3b13f7b",
7419 => x"567a5580",
7420 => x"08810554",
7421 => x"76538252",
7422 => x"893dfc05",
7423 => x"510b0bfe",
7424 => x"a0c53f80",
7425 => x"08570b0b",
7426 => x"0b85ce3f",
7427 => x"7780080c",
7428 => x"76800c89",
7429 => x"3d0d040b",
7430 => x"0b0b85bd",
7431 => x"3f850b80",
7432 => x"080cff0b",
7433 => x"800c893d",
7434 => x"0d04fb3d",
7435 => x"0d0b0b83",
7436 => x"85800870",
7437 => x"5654730b",
7438 => x"0b0b0b88",
7439 => x"3874800c",
7440 => x"873d0d04",
7441 => x"77538352",
7442 => x"873dfc05",
7443 => x"510b0bfe",
7444 => x"9ff53f80",
7445 => x"08540b0b",
7446 => x"0b84fe3f",
7447 => x"7580080c",
7448 => x"73800c87",
7449 => x"3d0d04ff",
7450 => x"0b800c04",
7451 => x"fb3d0d77",
7452 => x"550b0b83",
7453 => x"85800880",
7454 => x"2e0b0b0b",
7455 => x"0bb13874",
7456 => x"510b0b0b",
7457 => x"f2953f80",
7458 => x"08810554",
7459 => x"74538752",
7460 => x"873dfc05",
7461 => x"510b0bfe",
7462 => x"9fad3f80",
7463 => x"08550b0b",
7464 => x"0b84b63f",
7465 => x"7580080c",
7466 => x"74800c87",
7467 => x"3d0d040b",
7468 => x"0b0b84a5",
7469 => x"3f850b80",
7470 => x"080cff0b",
7471 => x"800c873d",
7472 => x"0d04fa3d",
7473 => x"0d0b0b83",
7474 => x"85800880",
7475 => x"2e0b0b0b",
7476 => x"0ba8387a",
7477 => x"55795478",
7478 => x"53865288",
7479 => x"3dfc0551",
7480 => x"0b0bfe9e",
7481 => x"e23f8008",
7482 => x"560b0b0b",
7483 => x"83eb3f76",
7484 => x"80080c75",
7485 => x"800c883d",
7486 => x"0d040b0b",
7487 => x"0b83da3f",
7488 => x"9d0b8008",
7489 => x"0cff0b80",
7490 => x"0c883d0d",
7491 => x"04fb3d0d",
7492 => x"77795656",
7493 => x"80705454",
7494 => x"7375250b",
7495 => x"0b0b0ba3",
7496 => x"38741010",
7497 => x"10f80552",
7498 => x"72167033",
7499 => x"70742b76",
7500 => x"078116f8",
7501 => x"16565656",
7502 => x"51517473",
7503 => x"240b0b0b",
7504 => x"0be63873",
7505 => x"800c873d",
7506 => x"0d04fc3d",
7507 => x"0d767855",
7508 => x"55bc5380",
7509 => x"5273510b",
7510 => x"0b0bc7b9",
7511 => x"3f845274",
7512 => x"510b0b0b",
7513 => x"ffa73f80",
7514 => x"08742384",
7515 => x"52841551",
7516 => x"0b0b0bff",
7517 => x"983f8008",
7518 => x"82152384",
7519 => x"52881551",
7520 => x"0b0b0bff",
7521 => x"883f8008",
7522 => x"84150c84",
7523 => x"528c1551",
7524 => x"0b0b0bfe",
7525 => x"f83f8008",
7526 => x"88152384",
7527 => x"52901551",
7528 => x"0b0b0bfe",
7529 => x"e83f8008",
7530 => x"8a152384",
7531 => x"52941551",
7532 => x"0b0b0bfe",
7533 => x"d83f8008",
7534 => x"8c152384",
7535 => x"52981551",
7536 => x"0b0b0bfe",
7537 => x"c83f8008",
7538 => x"8e152388",
7539 => x"529c1551",
7540 => x"0b0b0bfe",
7541 => x"b83f8008",
7542 => x"90150c86",
7543 => x"3d0d04e9",
7544 => x"3d0d6a0b",
7545 => x"0b838580",
7546 => x"08575775",
7547 => x"0b0b0b0b",
7548 => x"933880c0",
7549 => x"800b8418",
7550 => x"0c75ac18",
7551 => x"0c75800c",
7552 => x"993d0d04",
7553 => x"893d7055",
7554 => x"6a54558a",
7555 => x"52993dff",
7556 => x"bc05510b",
7557 => x"0bfe9caf",
7558 => x"3f800877",
7559 => x"53755256",
7560 => x"0b0b0bfe",
7561 => x"a53f0b0b",
7562 => x"0b81ae3f",
7563 => x"7780080c",
7564 => x"75800c99",
7565 => x"3d0d04e9",
7566 => x"3d0d6957",
7567 => x"0b0b8385",
7568 => x"8008802e",
7569 => x"0b0b0b80",
7570 => x"c1387651",
7571 => x"0b0b0bee",
7572 => x"ca3f893d",
7573 => x"70568008",
7574 => x"81055577",
7575 => x"54568f52",
7576 => x"993dffbc",
7577 => x"05510b0b",
7578 => x"fe9bdc3f",
7579 => x"80086b53",
7580 => x"7652570b",
7581 => x"0b0bfdd2",
7582 => x"3f0b0b0b",
7583 => x"80db3f77",
7584 => x"80080c76",
7585 => x"800c993d",
7586 => x"0d040b0b",
7587 => x"0b80ca3f",
7588 => x"850b8008",
7589 => x"0cff0b80",
7590 => x"0c993d0d",
7591 => x"04fc3d0d",
7592 => x"81540b0b",
7593 => x"83858008",
7594 => x"0b0b0b0b",
7595 => x"88387380",
7596 => x"0c863d0d",
7597 => x"04765397",
7598 => x"b952863d",
7599 => x"fc05510b",
7600 => x"0bfe9b83",
7601 => x"3f800854",
7602 => x"0b0b0b0b",
7603 => x"8c3f7480",
7604 => x"080c7380",
7605 => x"0c863d0d",
7606 => x"040b0b82",
7607 => x"f4ec0880",
7608 => x"0c04f73d",
7609 => x"0d7b0b0b",
7610 => x"82f4ec08",
7611 => x"82c81108",
7612 => x"5a545a77",
7613 => x"802e0b0b",
7614 => x"0b80ee38",
7615 => x"81881884",
7616 => x"1908ff05",
7617 => x"81712b59",
7618 => x"55598074",
7619 => x"240b0b0b",
7620 => x"81893880",
7621 => x"74240b0b",
7622 => x"0b0bbd38",
7623 => x"73822b78",
7624 => x"11880556",
7625 => x"56818019",
7626 => x"08770653",
7627 => x"72802e0b",
7628 => x"0b0b80c6",
7629 => x"38781670",
7630 => x"08535379",
7631 => x"51740853",
7632 => x"722dff14",
7633 => x"fc17fc17",
7634 => x"79812c5a",
7635 => x"57575473",
7636 => x"80250b0b",
7637 => x"0b0bce38",
7638 => x"77085877",
7639 => x"0b0b0bff",
7640 => x"9b380b0b",
7641 => x"82f4ec08",
7642 => x"53bc1308",
7643 => x"0b0b0b0b",
7644 => x"b2387951",
7645 => x"0b0b0bf5",
7646 => x"fd3f7408",
7647 => x"53722dff",
7648 => x"14fc17fc",
7649 => x"1779812c",
7650 => x"5a575754",
7651 => x"7380250b",
7652 => x"0b0bff91",
7653 => x"380b0b0b",
7654 => x"ffbe3980",
7655 => x"570b0b0b",
7656 => x"fef13972",
7657 => x"51bc1308",
7658 => x"53722d79",
7659 => x"510b0b0b",
7660 => x"f5c43f8c",
7661 => x"08028c0c",
7662 => x"d43d0d8c",
7663 => x"08880508",
7664 => x"510b0b0b",
7665 => x"8fb43f80",
7666 => x"08547380",
7667 => x"2e0b0b0b",
7668 => x"0b93388c",
7669 => x"08880508",
7670 => x"708c08d0",
7671 => x"050c540b",
7672 => x"0b0b8e8a",
7673 => x"398c088c",
7674 => x"0508510b",
7675 => x"0b0b8f8a",
7676 => x"3f800854",
7677 => x"73802e0b",
7678 => x"0b0b0b93",
7679 => x"388c088c",
7680 => x"0508708c",
7681 => x"08d0050c",
7682 => x"540b0b0b",
7683 => x"8de0398c",
7684 => x"08880508",
7685 => x"510b0b0b",
7686 => x"8eaa3f80",
7687 => x"08547380",
7688 => x"2e0b0b0b",
7689 => x"80d9388c",
7690 => x"088c0508",
7691 => x"510b0b0b",
7692 => x"8e923f80",
7693 => x"08547380",
7694 => x"2e0b0b0b",
7695 => x"0baf388c",
7696 => x"08880508",
7697 => x"8c088c05",
7698 => x"08555584",
7699 => x"15088415",
7700 => x"082e0b0b",
7701 => x"0b0b9638",
7702 => x"0b0b0b8d",
7703 => x"d43f8008",
7704 => x"708c08d0",
7705 => x"050c540b",
7706 => x"0b0b8d82",
7707 => x"398c0888",
7708 => x"0508708c",
7709 => x"08d0050c",
7710 => x"540b0b0b",
7711 => x"8cf0398c",
7712 => x"088c0508",
7713 => x"510b0b0b",
7714 => x"8dba3f80",
7715 => x"08547380",
7716 => x"2e0b0b0b",
7717 => x"0b93388c",
7718 => x"088c0508",
7719 => x"708c08d0",
7720 => x"050c540b",
7721 => x"0b0b8cc6",
7722 => x"398c088c",
7723 => x"0508510b",
7724 => x"0b0b8cc7",
7725 => x"3f800854",
7726 => x"73802e0b",
7727 => x"0b0b80f5",
7728 => x"388c0888",
7729 => x"0508510b",
7730 => x"0b0b8caf",
7731 => x"3f800854",
7732 => x"73802e0b",
7733 => x"0b0b80cb",
7734 => x"388c0890",
7735 => x"05088c08",
7736 => x"88050871",
7737 => x"58565494",
7738 => x"70547553",
7739 => x"7652540b",
7740 => x"0bfea197",
7741 => x"3f8c0890",
7742 => x"05088c08",
7743 => x"8805088c",
7744 => x"088c0508",
7745 => x"84120884",
7746 => x"12080684",
7747 => x"140c8c08",
7748 => x"90050870",
7749 => x"8c08d005",
7750 => x"0c515656",
7751 => x"560b0b0b",
7752 => x"8bcc398c",
7753 => x"08880508",
7754 => x"708c08d0",
7755 => x"050c540b",
7756 => x"0b0b8bba",
7757 => x"398c0888",
7758 => x"0508510b",
7759 => x"0b0b8bbb",
7760 => x"3f800854",
7761 => x"73802e0b",
7762 => x"0b0b0b93",
7763 => x"388c088c",
7764 => x"0508708c",
7765 => x"08d0050c",
7766 => x"540b0b0b",
7767 => x"8b90398c",
7768 => x"08880508",
7769 => x"8811088c",
7770 => x"08f4050c",
7771 => x"8c088c05",
7772 => x"08881108",
7773 => x"8c08f005",
7774 => x"0c8c0888",
7775 => x"05085151",
7776 => x"54901408",
7777 => x"8c150855",
7778 => x"55738c08",
7779 => x"e8050c74",
7780 => x"8c08ec05",
7781 => x"0c8c088c",
7782 => x"05085490",
7783 => x"14088c15",
7784 => x"08555573",
7785 => x"8c08e005",
7786 => x"0c748c08",
7787 => x"e4050c8c",
7788 => x"08f40508",
7789 => x"8c08f005",
7790 => x"08318c08",
7791 => x"dc050c8c",
7792 => x"08dc0508",
7793 => x"80250b0b",
7794 => x"0b0b8c38",
7795 => x"8c08dc05",
7796 => x"08308c08",
7797 => x"dc050c8c",
7798 => x"08dc0508",
7799 => x"bf240b0b",
7800 => x"0b81bf38",
7801 => x"8c08f005",
7802 => x"088c08f4",
7803 => x"0508250b",
7804 => x"0b0b80cf",
7805 => x"388c08f0",
7806 => x"05088105",
7807 => x"8c08f005",
7808 => x"0c8c08e0",
7809 => x"05088006",
7810 => x"8c08e405",
7811 => x"0881068c",
7812 => x"08e00508",
7813 => x"9f2b8c08",
7814 => x"e4050881",
7815 => x"2a707207",
7816 => x"8c08e005",
7817 => x"08812a70",
7818 => x"76078c08",
7819 => x"e0050c74",
7820 => x"72078c08",
7821 => x"e4050c59",
7822 => x"595b5b58",
7823 => x"560b0b0b",
7824 => x"ffa2398c",
7825 => x"08f40508",
7826 => x"8c08f005",
7827 => x"08250b0b",
7828 => x"0b819a38",
7829 => x"8c08f405",
7830 => x"0881058c",
7831 => x"08f4050c",
7832 => x"8c08e805",
7833 => x"0880068c",
7834 => x"08ec0508",
7835 => x"81068c08",
7836 => x"e805089f",
7837 => x"2b8c08ec",
7838 => x"0508812a",
7839 => x"7072078c",
7840 => x"08e80508",
7841 => x"812a7076",
7842 => x"078c08e8",
7843 => x"050c7472",
7844 => x"078c08ec",
7845 => x"050c5959",
7846 => x"5b5b5856",
7847 => x"0b0b0bff",
7848 => x"a2398c08",
7849 => x"f005088c",
7850 => x"08f40508",
7851 => x"250b0b0b",
7852 => x"0ba1388c",
7853 => x"08f40508",
7854 => x"8c08f005",
7855 => x"0c805480",
7856 => x"55738c08",
7857 => x"e0050c74",
7858 => x"8c08e405",
7859 => x"0c0b0b0b",
7860 => x"0b9b398c",
7861 => x"08f00508",
7862 => x"8c08f405",
7863 => x"0c805480",
7864 => x"55738c08",
7865 => x"e8050c74",
7866 => x"8c08ec05",
7867 => x"0c8c0888",
7868 => x"05088c08",
7869 => x"8c050855",
7870 => x"55841508",
7871 => x"8415082e",
7872 => x"0b0b0b85",
7873 => x"85388c08",
7874 => x"88050854",
7875 => x"84140880",
7876 => x"2e0b0b0b",
7877 => x"81bc388c",
7878 => x"08e00508",
7879 => x"8c08e405",
7880 => x"08565473",
7881 => x"8c08c805",
7882 => x"0c748c08",
7883 => x"cc050c8c",
7884 => x"08e80508",
7885 => x"8c08ec05",
7886 => x"08575574",
7887 => x"8c08c005",
7888 => x"0c758c08",
7889 => x"c4050c8c",
7890 => x"08cc0508",
7891 => x"8c08c405",
7892 => x"08717131",
7893 => x"708c08ff",
7894 => x"bc050c52",
7895 => x"5556810b",
7896 => x"8c08ffb4",
7897 => x"050c8c08",
7898 => x"ffbc0508",
7899 => x"8c08cc05",
7900 => x"08575574",
7901 => x"76260b0b",
7902 => x"0b0b8938",
7903 => x"800b8c08",
7904 => x"ffb4050c",
7905 => x"8c08c805",
7906 => x"088c08c0",
7907 => x"05087171",
7908 => x"31708c08",
7909 => x"ffb8050c",
7910 => x"8c08ffb8",
7911 => x"0508708c",
7912 => x"08ffb405",
7913 => x"0831708c",
7914 => x"08ffb805",
7915 => x"0c525952",
7916 => x"56548c08",
7917 => x"ffb80508",
7918 => x"8c08ffbc",
7919 => x"05085654",
7920 => x"738c08f8",
7921 => x"050c748c",
7922 => x"08fc050c",
7923 => x"0b0b0b81",
7924 => x"bf398c08",
7925 => x"e805088c",
7926 => x"08ec0508",
7927 => x"5755748c",
7928 => x"08ffac05",
7929 => x"0c758c08",
7930 => x"ffb0050c",
7931 => x"8c08e005",
7932 => x"088c08e4",
7933 => x"05085654",
7934 => x"738c08ff",
7935 => x"a4050c74",
7936 => x"8c08ffa8",
7937 => x"050c8c08",
7938 => x"ffb00508",
7939 => x"8c08ffa8",
7940 => x"05087171",
7941 => x"31708c08",
7942 => x"ffa0050c",
7943 => x"52575581",
7944 => x"0b8c08ff",
7945 => x"98050c8c",
7946 => x"08ffa005",
7947 => x"088c08ff",
7948 => x"b0050856",
7949 => x"54737526",
7950 => x"0b0b0b0b",
7951 => x"8938800b",
7952 => x"8c08ff98",
7953 => x"050c8c08",
7954 => x"ffac0508",
7955 => x"8c08ffa4",
7956 => x"05087171",
7957 => x"31708c08",
7958 => x"ff9c050c",
7959 => x"8c08ff9c",
7960 => x"0508708c",
7961 => x"08ff9805",
7962 => x"0831708c",
7963 => x"08ff9c05",
7964 => x"0c535852",
7965 => x"55568c08",
7966 => x"ff9c0508",
7967 => x"8c08ffa0",
7968 => x"05085654",
7969 => x"738c08f8",
7970 => x"050c748c",
7971 => x"08fc050c",
7972 => x"800b8c08",
7973 => x"f8050824",
7974 => x"0b0b0b0b",
7975 => x"ba388c08",
7976 => x"90050854",
7977 => x"800b8415",
7978 => x"0c8c0890",
7979 => x"05088c08",
7980 => x"f4050888",
7981 => x"120c8c08",
7982 => x"90050857",
7983 => x"548c08f8",
7984 => x"05088c08",
7985 => x"fc050856",
7986 => x"54738c17",
7987 => x"0c749017",
7988 => x"0c0b0b0b",
7989 => x"80d1398c",
7990 => x"08900508",
7991 => x"54810b84",
7992 => x"150c8c08",
7993 => x"9005088c",
7994 => x"08f40508",
7995 => x"88120c8c",
7996 => x"08900508",
7997 => x"8c08d405",
7998 => x"5858548c",
7999 => x"08f80508",
8000 => x"8c08fc05",
8001 => x"08565473",
8002 => x"52745375",
8003 => x"510b0b80",
8004 => x"cfcb3f8c",
8005 => x"08d40508",
8006 => x"8c08d805",
8007 => x"08565473",
8008 => x"8c180c74",
8009 => x"90180c8c",
8010 => x"08900508",
8011 => x"548c1408",
8012 => x"f00a260b",
8013 => x"0b0b82bb",
8014 => x"388c0890",
8015 => x"05088c11",
8016 => x"08709013",
8017 => x"08075155",
8018 => x"5573802e",
8019 => x"0b0b0b82",
8020 => x"a2388c08",
8021 => x"9005088c",
8022 => x"08900508",
8023 => x"9011089f",
8024 => x"2a8c1208",
8025 => x"10707207",
8026 => x"8c150c90",
8027 => x"13081090",
8028 => x"150c8c08",
8029 => x"90050888",
8030 => x"1108ff05",
8031 => x"88120c53",
8032 => x"58585557",
8033 => x"0b0b0bff",
8034 => x"9e398c08",
8035 => x"9005088c",
8036 => x"08880508",
8037 => x"84110884",
8038 => x"130c8c08",
8039 => x"9005088c",
8040 => x"08f40508",
8041 => x"88120c8c",
8042 => x"08900508",
8043 => x"8c08ff94",
8044 => x"050c5256",
8045 => x"548c08e8",
8046 => x"05088c08",
8047 => x"ec050857",
8048 => x"55748c08",
8049 => x"ff8c050c",
8050 => x"758c08ff",
8051 => x"90050c8c",
8052 => x"08e00508",
8053 => x"8c08e405",
8054 => x"08565473",
8055 => x"8c08ff84",
8056 => x"050c748c",
8057 => x"08ff8805",
8058 => x"0c8c08ff",
8059 => x"9005088c",
8060 => x"08ff8805",
8061 => x"08701270",
8062 => x"8c08ff80",
8063 => x"050c5257",
8064 => x"55810b8c",
8065 => x"08fef805",
8066 => x"0c8c08ff",
8067 => x"8005088c",
8068 => x"08ff9005",
8069 => x"08565474",
8070 => x"74260b0b",
8071 => x"0b0b8938",
8072 => x"800b8c08",
8073 => x"fef8050c",
8074 => x"8c08ff8c",
8075 => x"05088c08",
8076 => x"ff840508",
8077 => x"7012708c",
8078 => x"08fefc05",
8079 => x"0c8c08fe",
8080 => x"fc05088c",
8081 => x"08fef805",
8082 => x"0811708c",
8083 => x"08fefc05",
8084 => x"0c535852",
8085 => x"55568c08",
8086 => x"fefc0508",
8087 => x"8c08ff80",
8088 => x"05088c08",
8089 => x"ff940508",
8090 => x"58565473",
8091 => x"8c170c74",
8092 => x"90170c8c",
8093 => x"08900508",
8094 => x"5483740c",
8095 => x"8c089005",
8096 => x"08548c14",
8097 => x"08f80a26",
8098 => x"0b0b0b0b",
8099 => x"87380b0b",
8100 => x"0b80cf39",
8101 => x"8c089005",
8102 => x"088c0890",
8103 => x"05088c11",
8104 => x"08800690",
8105 => x"12088106",
8106 => x"8c089005",
8107 => x"088c1108",
8108 => x"9f2b9012",
8109 => x"08812a70",
8110 => x"72078c14",
8111 => x"08812a70",
8112 => x"77078c1a",
8113 => x"0c757207",
8114 => x"901a0c8c",
8115 => x"08900508",
8116 => x"88110881",
8117 => x"0588120c",
8118 => x"51575c5f",
8119 => x"5f5c5a58",
8120 => x"555b8c08",
8121 => x"90050870",
8122 => x"8c08d005",
8123 => x"0c548c08",
8124 => x"d0050880",
8125 => x"0cae3d0d",
8126 => x"8c0c048c",
8127 => x"08028c0c",
8128 => x"7070800b",
8129 => x"8c08fc05",
8130 => x"0c8c0888",
8131 => x"05085170",
8132 => x"08822e09",
8133 => x"81060b0b",
8134 => x"0b0b8838",
8135 => x"810b8c08",
8136 => x"fc050c8c",
8137 => x"08fc0508",
8138 => x"70800c51",
8139 => x"50508c0c",
8140 => x"048c0802",
8141 => x"8c0c700b",
8142 => x"0b82f4b8",
8143 => x"70800c51",
8144 => x"508c0c04",
8145 => x"8c08028c",
8146 => x"0c707080",
8147 => x"0b8c08fc",
8148 => x"050c8c08",
8149 => x"88050851",
8150 => x"7008842e",
8151 => x"0981060b",
8152 => x"0b0b0b88",
8153 => x"38810b8c",
8154 => x"08fc050c",
8155 => x"8c08fc05",
8156 => x"0870800c",
8157 => x"5150508c",
8158 => x"0c048c08",
8159 => x"028c0c70",
8160 => x"70800b8c",
8161 => x"08fc050c",
8162 => x"8c088805",
8163 => x"08517008",
8164 => x"802e0b0b",
8165 => x"0b0b9738",
8166 => x"8c088805",
8167 => x"08517008",
8168 => x"812e0b0b",
8169 => x"0b0b8738",
8170 => x"0b0b0b0b",
8171 => x"8839810b",
8172 => x"8c08fc05",
8173 => x"0c8c08fc",
8174 => x"05087080",
8175 => x"0c515050",
8176 => x"8c0c048c",
8177 => x"08028c0c",
8178 => x"e73d0d8c",
8179 => x"08880508",
8180 => x"568c088c",
8181 => x"05088c08",
8182 => x"90050856",
8183 => x"54738c08",
8184 => x"ffb8050c",
8185 => x"748c08ff",
8186 => x"bc050c8c",
8187 => x"08940508",
8188 => x"8c089805",
8189 => x"08565473",
8190 => x"8c08ffb0",
8191 => x"050c748c",
8192 => x"08ffb405",
8193 => x"0c8c08ec",
8194 => x"0570538c",
8195 => x"08ffb805",
8196 => x"70535154",
8197 => x"0b0b80de",
8198 => x"c13f8c08",
8199 => x"d8057053",
8200 => x"8c08ffb0",
8201 => x"05705351",
8202 => x"540b0b80",
8203 => x"deac3f8c",
8204 => x"08c40570",
8205 => x"548c08d8",
8206 => x"0570548c",
8207 => x"08ec0570",
8208 => x"54515154",
8209 => x"0b0b0bee",
8210 => x"ea3f8008",
8211 => x"708c08c0",
8212 => x"050c8c08",
8213 => x"c0050853",
8214 => x"7652540b",
8215 => x"0b80ccb8",
8216 => x"3f75800c",
8217 => x"9b3d0d8c",
8218 => x"0c048c08",
8219 => x"028c0ce7",
8220 => x"3d0d8c08",
8221 => x"88050856",
8222 => x"8c088c05",
8223 => x"088c0890",
8224 => x"05085654",
8225 => x"738c08ff",
8226 => x"b8050c74",
8227 => x"8c08ffbc",
8228 => x"050c8c08",
8229 => x"9405088c",
8230 => x"08980508",
8231 => x"5654738c",
8232 => x"08ffb005",
8233 => x"0c748c08",
8234 => x"ffb4050c",
8235 => x"8c08ec05",
8236 => x"70538c08",
8237 => x"ffb80570",
8238 => x"5351540b",
8239 => x"0b80dd9a",
8240 => x"3f8c08d8",
8241 => x"0570538c",
8242 => x"08ffb005",
8243 => x"70535154",
8244 => x"0b0b80dd",
8245 => x"853f8c08",
8246 => x"dc050881",
8247 => x"328c08dc",
8248 => x"050c8c08",
8249 => x"c4057054",
8250 => x"8c08d805",
8251 => x"70548c08",
8252 => x"ec057054",
8253 => x"5151540b",
8254 => x"0b0bedb7",
8255 => x"3f800870",
8256 => x"8c08c005",
8257 => x"0c8c08c0",
8258 => x"05085376",
8259 => x"52540b0b",
8260 => x"80cb853f",
8261 => x"75800c9b",
8262 => x"3d0d8c0c",
8263 => x"048c0802",
8264 => x"8c0cff83",
8265 => x"3d0d8c08",
8266 => x"8c05088c",
8267 => x"08900508",
8268 => x"5856758c",
8269 => x"08ffb805",
8270 => x"0c768c08",
8271 => x"ffbc050c",
8272 => x"8c089405",
8273 => x"088c0898",
8274 => x"05085856",
8275 => x"758c08ff",
8276 => x"b0050c76",
8277 => x"8c08ffb4",
8278 => x"050c8c08",
8279 => x"ec057053",
8280 => x"8c08ffb8",
8281 => x"05705351",
8282 => x"560b0b80",
8283 => x"dbec3f8c",
8284 => x"08d80570",
8285 => x"538c08ff",
8286 => x"b0057053",
8287 => x"51560b0b",
8288 => x"80dbd73f",
8289 => x"8c08ec05",
8290 => x"8c08ffac",
8291 => x"050c8c08",
8292 => x"d8058c08",
8293 => x"ffa8050c",
8294 => x"8c08c405",
8295 => x"8c08ffa4",
8296 => x"050c8056",
8297 => x"8057758c",
8298 => x"08ff9805",
8299 => x"0c768c08",
8300 => x"ff9c050c",
8301 => x"80568057",
8302 => x"758c08ff",
8303 => x"90050c76",
8304 => x"8c08ff94",
8305 => x"050c8c08",
8306 => x"ffac0508",
8307 => x"510b0b0b",
8308 => x"9d823f80",
8309 => x"08567580",
8310 => x"2e0b0b0b",
8311 => x"80da388c",
8312 => x"08ffac05",
8313 => x"088c08fe",
8314 => x"c4050c80",
8315 => x"0b8c08fe",
8316 => x"c0050c8c",
8317 => x"08ffac05",
8318 => x"088c08ff",
8319 => x"a8050857",
8320 => x"57841708",
8321 => x"8417082e",
8322 => x"0b0b0b0b",
8323 => x"8938810b",
8324 => x"8c08fec0",
8325 => x"050c8c08",
8326 => x"fec40508",
8327 => x"8c08fec0",
8328 => x"05088412",
8329 => x"0c8c08ff",
8330 => x"ac05088c",
8331 => x"08ffa005",
8332 => x"0c560b0b",
8333 => x"0b9af139",
8334 => x"8c08ffa8",
8335 => x"0508510b",
8336 => x"0b0b9c90",
8337 => x"3f800856",
8338 => x"75802e0b",
8339 => x"0b0b80da",
8340 => x"388c08ff",
8341 => x"a805088c",
8342 => x"08febc05",
8343 => x"0c800b8c",
8344 => x"08feb805",
8345 => x"0c8c08ff",
8346 => x"ac05088c",
8347 => x"08ffa805",
8348 => x"08575784",
8349 => x"17088417",
8350 => x"082e0b0b",
8351 => x"0b0b8938",
8352 => x"810b8c08",
8353 => x"feb8050c",
8354 => x"8c08febc",
8355 => x"05088c08",
8356 => x"feb80508",
8357 => x"84120c8c",
8358 => x"08ffa805",
8359 => x"088c08ff",
8360 => x"a0050c57",
8361 => x"0b0b0b99",
8362 => x"ff398c08",
8363 => x"ffac0508",
8364 => x"510b0b0b",
8365 => x"9ae83f80",
8366 => x"08567580",
8367 => x"2e0b0b0b",
8368 => x"8189388c",
8369 => x"08ffa805",
8370 => x"08510b0b",
8371 => x"0b9a993f",
8372 => x"80085675",
8373 => x"802e0b0b",
8374 => x"0b0b9738",
8375 => x"0b0b0b99",
8376 => x"f43f8008",
8377 => x"708c08ff",
8378 => x"a0050c56",
8379 => x"0b0b0b99",
8380 => x"b7398c08",
8381 => x"ffac0508",
8382 => x"8c08feb4",
8383 => x"050c800b",
8384 => x"8c08feb0",
8385 => x"050c8c08",
8386 => x"ffac0508",
8387 => x"8c08ffa8",
8388 => x"05085757",
8389 => x"84170884",
8390 => x"17082e0b",
8391 => x"0b0b0b89",
8392 => x"38810b8c",
8393 => x"08feb005",
8394 => x"0c8c08fe",
8395 => x"b405088c",
8396 => x"08feb005",
8397 => x"0884120c",
8398 => x"8c08ffac",
8399 => x"05088c08",
8400 => x"ffa0050c",
8401 => x"560b0b0b",
8402 => x"98de398c",
8403 => x"08ffa805",
8404 => x"08510b0b",
8405 => x"0b99c73f",
8406 => x"80085675",
8407 => x"802e0b0b",
8408 => x"0b818938",
8409 => x"8c08ffac",
8410 => x"0508510b",
8411 => x"0b0b98f8",
8412 => x"3f800856",
8413 => x"75802e0b",
8414 => x"0b0b0b97",
8415 => x"380b0b0b",
8416 => x"98d33f80",
8417 => x"08708c08",
8418 => x"ffa0050c",
8419 => x"560b0b0b",
8420 => x"9896398c",
8421 => x"08ffa805",
8422 => x"088c08fe",
8423 => x"ac050c80",
8424 => x"0b8c08fe",
8425 => x"a8050c8c",
8426 => x"08ffac05",
8427 => x"088c08ff",
8428 => x"a8050857",
8429 => x"57841708",
8430 => x"8417082e",
8431 => x"0b0b0b0b",
8432 => x"8938810b",
8433 => x"8c08fea8",
8434 => x"050c8c08",
8435 => x"feac0508",
8436 => x"8c08fea8",
8437 => x"05088412",
8438 => x"0c8c08ff",
8439 => x"a805088c",
8440 => x"08ffa005",
8441 => x"0c570b0b",
8442 => x"0b97bd39",
8443 => x"8c08ffac",
8444 => x"0508510b",
8445 => x"0b0b97f0",
8446 => x"3f800856",
8447 => x"75802e0b",
8448 => x"0b0b80da",
8449 => x"388c08ff",
8450 => x"ac05088c",
8451 => x"08fea405",
8452 => x"0c800b8c",
8453 => x"08fea005",
8454 => x"0c8c08ff",
8455 => x"ac05088c",
8456 => x"08ffa805",
8457 => x"08575784",
8458 => x"17088417",
8459 => x"082e0b0b",
8460 => x"0b0b8938",
8461 => x"810b8c08",
8462 => x"fea0050c",
8463 => x"8c08fea4",
8464 => x"05088c08",
8465 => x"fea00508",
8466 => x"84120c8c",
8467 => x"08ffac05",
8468 => x"088c08ff",
8469 => x"a0050c56",
8470 => x"0b0b0b96",
8471 => x"cb398c08",
8472 => x"ffa80508",
8473 => x"510b0b0b",
8474 => x"96fe3f80",
8475 => x"08567580",
8476 => x"2e0b0b0b",
8477 => x"80da388c",
8478 => x"08ffa805",
8479 => x"088c08fe",
8480 => x"9c050c80",
8481 => x"0b8c08fe",
8482 => x"98050c8c",
8483 => x"08ffac05",
8484 => x"088c08ff",
8485 => x"a8050857",
8486 => x"57841708",
8487 => x"8417082e",
8488 => x"0b0b0b0b",
8489 => x"8938810b",
8490 => x"8c08fe98",
8491 => x"050c8c08",
8492 => x"fe9c0508",
8493 => x"8c08fe98",
8494 => x"05088412",
8495 => x"0c8c08ff",
8496 => x"a805088c",
8497 => x"08ffa005",
8498 => x"0c570b0b",
8499 => x"0b95d939",
8500 => x"8c08ffac",
8501 => x"05089011",
8502 => x"088c08ff",
8503 => x"8c050c8c",
8504 => x"08ffac05",
8505 => x"088c1108",
8506 => x"802a5959",
8507 => x"5680778c",
8508 => x"08ff8805",
8509 => x"0c8c08ff",
8510 => x"a8050890",
8511 => x"11088c08",
8512 => x"ff84050c",
8513 => x"8c08ffa8",
8514 => x"05088c11",
8515 => x"08802a5a",
8516 => x"5a515680",
8517 => x"778c08ff",
8518 => x"80050c8c",
8519 => x"08ff8405",
8520 => x"085a5680",
8521 => x"0b8c08ff",
8522 => x"8c050858",
8523 => x"58800b8c",
8524 => x"08fef005",
8525 => x"5b567554",
8526 => x"76557752",
8527 => x"78537951",
8528 => x"0b0b0bbb",
8529 => x"b23f8c08",
8530 => x"fef00508",
8531 => x"8c08fef4",
8532 => x"05085856",
8533 => x"758c08fe",
8534 => x"f8050c76",
8535 => x"8c08fefc",
8536 => x"050c8c08",
8537 => x"ff800508",
8538 => x"59800b8c",
8539 => x"08ff8c05",
8540 => x"08585880",
8541 => x"0b8c08fe",
8542 => x"e8055b56",
8543 => x"75547655",
8544 => x"77527853",
8545 => x"79510b0b",
8546 => x"0bbaec3f",
8547 => x"8c08fee8",
8548 => x"05088c08",
8549 => x"feec0508",
8550 => x"5856758c",
8551 => x"08fef005",
8552 => x"0c768c08",
8553 => x"fef4050c",
8554 => x"8c08ff84",
8555 => x"05085980",
8556 => x"0b8c08ff",
8557 => x"88050858",
8558 => x"58800b8c",
8559 => x"08fee005",
8560 => x"5b567554",
8561 => x"76557752",
8562 => x"78537951",
8563 => x"0b0b0bba",
8564 => x"a63f8c08",
8565 => x"fee00508",
8566 => x"8c08fee4",
8567 => x"05085856",
8568 => x"758c08fe",
8569 => x"e8050c76",
8570 => x"8c08feec",
8571 => x"050c8c08",
8572 => x"ff800508",
8573 => x"59800b8c",
8574 => x"08ff8805",
8575 => x"08585880",
8576 => x"0b8c08fe",
8577 => x"d8055b56",
8578 => x"75547655",
8579 => x"77527853",
8580 => x"79510b0b",
8581 => x"0bb9e03f",
8582 => x"8c08fed8",
8583 => x"05088c08",
8584 => x"fedc0508",
8585 => x"5856758c",
8586 => x"08fee005",
8587 => x"0c768c08",
8588 => x"fee4050c",
8589 => x"80568057",
8590 => x"758c08fe",
8591 => x"d8050c76",
8592 => x"8c08fedc",
8593 => x"050c8056",
8594 => x"8057758c",
8595 => x"08fed005",
8596 => x"0c768c08",
8597 => x"fed4050c",
8598 => x"8c08fef0",
8599 => x"05088c08",
8600 => x"fef40508",
8601 => x"5856758c",
8602 => x"08fe9005",
8603 => x"0c768c08",
8604 => x"fe94050c",
8605 => x"8c08fee8",
8606 => x"05088c08",
8607 => x"feec0508",
8608 => x"5856758c",
8609 => x"08fe8805",
8610 => x"0c768c08",
8611 => x"fe8c050c",
8612 => x"8c08fe94",
8613 => x"05088c08",
8614 => x"fe8c0508",
8615 => x"7012708c",
8616 => x"08fe8405",
8617 => x"0c525757",
8618 => x"810b8c08",
8619 => x"fdfc050c",
8620 => x"8c08fe84",
8621 => x"05088c08",
8622 => x"fe940508",
8623 => x"57577577",
8624 => x"260b0b0b",
8625 => x"0b893880",
8626 => x"0b8c08fd",
8627 => x"fc050c8c",
8628 => x"08fe9005",
8629 => x"088c08fe",
8630 => x"88050870",
8631 => x"12708c08",
8632 => x"fe80050c",
8633 => x"8c08fe80",
8634 => x"05088c08",
8635 => x"fdfc0508",
8636 => x"11708c08",
8637 => x"fe80050c",
8638 => x"53515257",
8639 => x"578c08fe",
8640 => x"8005088c",
8641 => x"08fe8405",
8642 => x"08585675",
8643 => x"8c08fec8",
8644 => x"050c768c",
8645 => x"08fecc05",
8646 => x"0c8c08fe",
8647 => x"f005088c",
8648 => x"08fec805",
8649 => x"08260b0b",
8650 => x"0b0bb038",
8651 => x"8c08fef0",
8652 => x"05088c08",
8653 => x"fec80508",
8654 => x"2e098106",
8655 => x"0b0b0b81",
8656 => x"d1388c08",
8657 => x"fef40508",
8658 => x"8c08fecc",
8659 => x"0508260b",
8660 => x"0b0b0b87",
8661 => x"380b0b0b",
8662 => x"81b8398c",
8663 => x"08fed805",
8664 => x"088c08fe",
8665 => x"dc050858",
8666 => x"56758c08",
8667 => x"fdf4050c",
8668 => x"768c08fd",
8669 => x"f8050c81",
8670 => x"56805775",
8671 => x"8c08fdec",
8672 => x"050c768c",
8673 => x"08fdf005",
8674 => x"0c8c08fd",
8675 => x"f805088c",
8676 => x"08fdf005",
8677 => x"08701270",
8678 => x"8c08fde8",
8679 => x"050c5257",
8680 => x"57810b8c",
8681 => x"08fde005",
8682 => x"0c8c08fd",
8683 => x"e805088c",
8684 => x"08fdf805",
8685 => x"08575775",
8686 => x"77260b0b",
8687 => x"0b0b8938",
8688 => x"800b8c08",
8689 => x"fde0050c",
8690 => x"8c08fdf4",
8691 => x"05088c08",
8692 => x"fdec0508",
8693 => x"7012708c",
8694 => x"08fde405",
8695 => x"0c8c08fd",
8696 => x"e405088c",
8697 => x"08fde005",
8698 => x"0811708c",
8699 => x"08fde405",
8700 => x"0c535152",
8701 => x"57578c08",
8702 => x"fde40508",
8703 => x"8c08fde8",
8704 => x"05085856",
8705 => x"758c08fe",
8706 => x"d8050c76",
8707 => x"8c08fedc",
8708 => x"050c8c08",
8709 => x"fecc0508",
8710 => x"57807780",
8711 => x"2b8c08fe",
8712 => x"f0050c56",
8713 => x"800b8c08",
8714 => x"fef4050c",
8715 => x"8c08fef8",
8716 => x"05088c08",
8717 => x"fefc0508",
8718 => x"5856758c",
8719 => x"08fdd805",
8720 => x"0c768c08",
8721 => x"fddc050c",
8722 => x"8c08fef0",
8723 => x"05088c08",
8724 => x"fef40508",
8725 => x"5856758c",
8726 => x"08fdd005",
8727 => x"0c768c08",
8728 => x"fdd4050c",
8729 => x"8c08fddc",
8730 => x"05088c08",
8731 => x"fdd40508",
8732 => x"7012708c",
8733 => x"08fdcc05",
8734 => x"0c525757",
8735 => x"810b8c08",
8736 => x"fdc4050c",
8737 => x"8c08fdcc",
8738 => x"05088c08",
8739 => x"fddc0508",
8740 => x"57577577",
8741 => x"260b0b0b",
8742 => x"0b893880",
8743 => x"0b8c08fd",
8744 => x"c4050c8c",
8745 => x"08fdd805",
8746 => x"088c08fd",
8747 => x"d0050870",
8748 => x"12708c08",
8749 => x"fdc8050c",
8750 => x"8c08fdc8",
8751 => x"05088c08",
8752 => x"fdc40508",
8753 => x"11708c08",
8754 => x"fdc8050c",
8755 => x"53515257",
8756 => x"578c08fd",
8757 => x"c805088c",
8758 => x"08fdcc05",
8759 => x"08585675",
8760 => x"8c08fed0",
8761 => x"050c768c",
8762 => x"08fed405",
8763 => x"0c8c08fe",
8764 => x"f805088c",
8765 => x"08fed005",
8766 => x"08260b0b",
8767 => x"0b0bb038",
8768 => x"8c08fef8",
8769 => x"05088c08",
8770 => x"fed00508",
8771 => x"2e098106",
8772 => x"0b0b0b81",
8773 => x"d1388c08",
8774 => x"fefc0508",
8775 => x"8c08fed4",
8776 => x"0508260b",
8777 => x"0b0b0b87",
8778 => x"380b0b0b",
8779 => x"81b8398c",
8780 => x"08fed805",
8781 => x"088c08fe",
8782 => x"dc050858",
8783 => x"56758c08",
8784 => x"fdbc050c",
8785 => x"768c08fd",
8786 => x"c0050c80",
8787 => x"56815775",
8788 => x"8c08fdb4",
8789 => x"050c768c",
8790 => x"08fdb805",
8791 => x"0c8c08fd",
8792 => x"c005088c",
8793 => x"08fdb805",
8794 => x"08701270",
8795 => x"8c08fdb0",
8796 => x"050c5257",
8797 => x"57810b8c",
8798 => x"08fda805",
8799 => x"0c8c08fd",
8800 => x"b005088c",
8801 => x"08fdc005",
8802 => x"08575775",
8803 => x"77260b0b",
8804 => x"0b0b8938",
8805 => x"800b8c08",
8806 => x"fda8050c",
8807 => x"8c08fdbc",
8808 => x"05088c08",
8809 => x"fdb40508",
8810 => x"7012708c",
8811 => x"08fdac05",
8812 => x"0c8c08fd",
8813 => x"ac05088c",
8814 => x"08fda805",
8815 => x"0811708c",
8816 => x"08fdac05",
8817 => x"0c535152",
8818 => x"57578c08",
8819 => x"fdac0508",
8820 => x"8c08fdb0",
8821 => x"05085856",
8822 => x"758c08fe",
8823 => x"d8050c76",
8824 => x"8c08fedc",
8825 => x"050c8c08",
8826 => x"fec80508",
8827 => x"802a708c",
8828 => x"08fda405",
8829 => x"0c578070",
8830 => x"8c08fda0",
8831 => x"050c568c",
8832 => x"08fda005",
8833 => x"088c08fd",
8834 => x"a4050858",
8835 => x"56758c08",
8836 => x"fda0050c",
8837 => x"768c08fd",
8838 => x"a4050c8c",
8839 => x"08fee005",
8840 => x"088c08fe",
8841 => x"e4050858",
8842 => x"56758c08",
8843 => x"fd98050c",
8844 => x"768c08fd",
8845 => x"9c050c8c",
8846 => x"08fda405",
8847 => x"088c08fd",
8848 => x"9c050870",
8849 => x"12708c08",
8850 => x"fd94050c",
8851 => x"52575781",
8852 => x"0b8c08fd",
8853 => x"8c050c8c",
8854 => x"08fd9405",
8855 => x"088c08fd",
8856 => x"a4050857",
8857 => x"57757726",
8858 => x"0b0b0b0b",
8859 => x"8938800b",
8860 => x"8c08fd8c",
8861 => x"050c8c08",
8862 => x"fda00508",
8863 => x"8c08fd98",
8864 => x"05087012",
8865 => x"708c08fd",
8866 => x"90050c8c",
8867 => x"08fd9005",
8868 => x"088c08fd",
8869 => x"8c050811",
8870 => x"708c08fd",
8871 => x"90050c53",
8872 => x"51525757",
8873 => x"8c08fed8",
8874 => x"05088c08",
8875 => x"fedc0508",
8876 => x"5856758c",
8877 => x"08fd8405",
8878 => x"0c768c08",
8879 => x"fd88050c",
8880 => x"8c08fd88",
8881 => x"05088c08",
8882 => x"fd940508",
8883 => x"7012708c",
8884 => x"08fd8005",
8885 => x"0c525757",
8886 => x"810b8c08",
8887 => x"fcf8050c",
8888 => x"8c08fd80",
8889 => x"05088c08",
8890 => x"fd880508",
8891 => x"57577577",
8892 => x"260b0b0b",
8893 => x"0b893880",
8894 => x"0b8c08fc",
8895 => x"f8050c8c",
8896 => x"08fd8405",
8897 => x"088c08fd",
8898 => x"90050870",
8899 => x"12708c08",
8900 => x"fcfc050c",
8901 => x"8c08fcfc",
8902 => x"05088c08",
8903 => x"fcf80508",
8904 => x"11708c08",
8905 => x"fcfc050c",
8906 => x"53515257",
8907 => x"578c08fc",
8908 => x"fc05088c",
8909 => x"08fd8005",
8910 => x"08585675",
8911 => x"8c08fed8",
8912 => x"050c768c",
8913 => x"08fedc05",
8914 => x"0c8c08fe",
8915 => x"d805088c",
8916 => x"08fedc05",
8917 => x"08585675",
8918 => x"8c08ff90",
8919 => x"050c768c",
8920 => x"08ff9405",
8921 => x"0c8c08fe",
8922 => x"d005088c",
8923 => x"08fed405",
8924 => x"08585675",
8925 => x"8c08ff98",
8926 => x"050c768c",
8927 => x"08ff9c05",
8928 => x"0c8c08ff",
8929 => x"a405088c",
8930 => x"08ffac05",
8931 => x"088c08ff",
8932 => x"a8050888",
8933 => x"12088812",
8934 => x"08058411",
8935 => x"88150c8c",
8936 => x"08ffa405",
8937 => x"088c08fc",
8938 => x"f4050c51",
8939 => x"58585880",
8940 => x"0b8c08fc",
8941 => x"f0050c8c",
8942 => x"08ffac05",
8943 => x"088c08ff",
8944 => x"a8050857",
8945 => x"57841708",
8946 => x"8417082e",
8947 => x"0b0b0b0b",
8948 => x"8938810b",
8949 => x"8c08fcf0",
8950 => x"050c8c08",
8951 => x"fcf40508",
8952 => x"8c08fcf0",
8953 => x"05088412",
8954 => x"0c578c08",
8955 => x"ff900508",
8956 => x"f80a260b",
8957 => x"0b0b0b87",
8958 => x"380b0b0b",
8959 => x"81ae398c",
8960 => x"08ffa405",
8961 => x"08881108",
8962 => x"81058812",
8963 => x"0c8c08ff",
8964 => x"90050880",
8965 => x"068c08ff",
8966 => x"94050881",
8967 => x"06705259",
8968 => x"51567580",
8969 => x"2e0b0b0b",
8970 => x"80cf388c",
8971 => x"08ff9805",
8972 => x"089f2b8c",
8973 => x"08ff9c05",
8974 => x"08812a70",
8975 => x"72078c08",
8976 => x"ff980508",
8977 => x"812a5959",
8978 => x"5959758c",
8979 => x"08ff9805",
8980 => x"0c768c08",
8981 => x"ff9c050c",
8982 => x"8c08ff98",
8983 => x"0508810a",
8984 => x"078c08ff",
8985 => x"9c050880",
8986 => x"07585675",
8987 => x"8c08ff98",
8988 => x"050c768c",
8989 => x"08ff9c05",
8990 => x"0c8c08ff",
8991 => x"9005089f",
8992 => x"2b8c08ff",
8993 => x"94050881",
8994 => x"2a707207",
8995 => x"8c08ff90",
8996 => x"0508812a",
8997 => x"59595959",
8998 => x"758c08ff",
8999 => x"90050c76",
9000 => x"8c08ff94",
9001 => x"050c0b0b",
9002 => x"0bfebf39",
9003 => x"8c08ff90",
9004 => x"0508f00a",
9005 => x"260b0b0b",
9006 => x"81a1388c",
9007 => x"08ffa405",
9008 => x"08881108",
9009 => x"ff058812",
9010 => x"0c8c08ff",
9011 => x"9405089f",
9012 => x"2a8c08ff",
9013 => x"90050810",
9014 => x"7072078c",
9015 => x"08ff9405",
9016 => x"08105b53",
9017 => x"5a5a5675",
9018 => x"8c08ff90",
9019 => x"050c768c",
9020 => x"08ff9405",
9021 => x"0c800b8c",
9022 => x"08ff9805",
9023 => x"08240b0b",
9024 => x"0b0b8738",
9025 => x"0b0b0b0b",
9026 => x"a1398c08",
9027 => x"ff900508",
9028 => x"80078c08",
9029 => x"ff940508",
9030 => x"81075856",
9031 => x"758c08ff",
9032 => x"90050c76",
9033 => x"8c08ff94",
9034 => x"050c8c08",
9035 => x"ff9c0508",
9036 => x"9f2a8c08",
9037 => x"ff980508",
9038 => x"10707207",
9039 => x"8c08ff9c",
9040 => x"0508105a",
9041 => x"58595975",
9042 => x"8c08ff98",
9043 => x"050c768c",
9044 => x"08ff9c05",
9045 => x"0c0b0b0b",
9046 => x"fed2398c",
9047 => x"08ff9005",
9048 => x"08800670",
9049 => x"8c08fce8",
9050 => x"050c8c08",
9051 => x"ff940508",
9052 => x"81ff0670",
9053 => x"8c08fcec",
9054 => x"050c5856",
9055 => x"8c08fce8",
9056 => x"05088c08",
9057 => x"fcec0508",
9058 => x"5856758c",
9059 => x"08fce805",
9060 => x"0c768c08",
9061 => x"fcec050c",
9062 => x"8c08fce8",
9063 => x"05085776",
9064 => x"0b0b0b83",
9065 => x"d0388c08",
9066 => x"fcec0508",
9067 => x"56758180",
9068 => x"2e098106",
9069 => x"0b0b0b83",
9070 => x"bc388c08",
9071 => x"ff900508",
9072 => x"982b8c08",
9073 => x"ff940508",
9074 => x"882a7072",
9075 => x"078c08ff",
9076 => x"90050888",
9077 => x"2a718106",
9078 => x"51595959",
9079 => x"5975802e",
9080 => x"0b0b0b81",
9081 => x"bf388c08",
9082 => x"ff900508",
9083 => x"8c08ff94",
9084 => x"05085856",
9085 => x"758c08fc",
9086 => x"e0050c76",
9087 => x"8c08fce4",
9088 => x"050c8056",
9089 => x"81805775",
9090 => x"8c08fcd8",
9091 => x"050c768c",
9092 => x"08fcdc05",
9093 => x"0c8c08fc",
9094 => x"e405088c",
9095 => x"08fcdc05",
9096 => x"08701270",
9097 => x"8c08fcd4",
9098 => x"050c5257",
9099 => x"57810b8c",
9100 => x"08fccc05",
9101 => x"0c8c08fc",
9102 => x"d405088c",
9103 => x"08fce405",
9104 => x"08575775",
9105 => x"77260b0b",
9106 => x"0b0b8938",
9107 => x"800b8c08",
9108 => x"fccc050c",
9109 => x"8c08fce0",
9110 => x"05088c08",
9111 => x"fcd80508",
9112 => x"7012708c",
9113 => x"08fcd005",
9114 => x"0c8c08fc",
9115 => x"d005088c",
9116 => x"08fccc05",
9117 => x"0811708c",
9118 => x"08fcd005",
9119 => x"0c535152",
9120 => x"57578c08",
9121 => x"fcd00508",
9122 => x"8c08fcd4",
9123 => x"05085856",
9124 => x"758c08ff",
9125 => x"90050c76",
9126 => x"8c08ff94",
9127 => x"050c0b0b",
9128 => x"0b81d239",
9129 => x"8c08ff98",
9130 => x"0508708c",
9131 => x"08ff9c05",
9132 => x"08075156",
9133 => x"75802e0b",
9134 => x"0b0b81b9",
9135 => x"388c08ff",
9136 => x"9005088c",
9137 => x"08ff9405",
9138 => x"08585675",
9139 => x"8c08fcc4",
9140 => x"050c768c",
9141 => x"08fcc805",
9142 => x"0c805681",
9143 => x"8057758c",
9144 => x"08fcbc05",
9145 => x"0c768c08",
9146 => x"fcc0050c",
9147 => x"8c08fcc8",
9148 => x"05088c08",
9149 => x"fcc00508",
9150 => x"7012708c",
9151 => x"08fcb805",
9152 => x"0c525757",
9153 => x"810b8c08",
9154 => x"fcb0050c",
9155 => x"8c08fcb8",
9156 => x"05088c08",
9157 => x"fcc80508",
9158 => x"57577577",
9159 => x"260b0b0b",
9160 => x"0b893880",
9161 => x"0b8c08fc",
9162 => x"b0050c8c",
9163 => x"08fcc405",
9164 => x"088c08fc",
9165 => x"bc050870",
9166 => x"12708c08",
9167 => x"fcb4050c",
9168 => x"8c08fcb4",
9169 => x"05088c08",
9170 => x"fcb00508",
9171 => x"11708c08",
9172 => x"fcb4050c",
9173 => x"53515257",
9174 => x"578c08fc",
9175 => x"b405088c",
9176 => x"08fcb805",
9177 => x"08585675",
9178 => x"8c08ff90",
9179 => x"050c768c",
9180 => x"08ff9405",
9181 => x"0c8c08ff",
9182 => x"a4050856",
9183 => x"8c08ff90",
9184 => x"05088c08",
9185 => x"ff940508",
9186 => x"5957768c",
9187 => x"170c7790",
9188 => x"170c8c08",
9189 => x"ffa40508",
9190 => x"5683760c",
9191 => x"8c08ffa4",
9192 => x"05088c08",
9193 => x"ffa0050c",
9194 => x"8c08ffa0",
9195 => x"0508708c",
9196 => x"08c0050c",
9197 => x"8c08c005",
9198 => x"08538c08",
9199 => x"88050852",
9200 => x"560b0b0b",
9201 => x"add23f8c",
9202 => x"08880508",
9203 => x"800c80ff",
9204 => x"3d0d8c0c",
9205 => x"048c0802",
9206 => x"8c0c700b",
9207 => x"0b82f4b8",
9208 => x"70800c51",
9209 => x"508c0c04",
9210 => x"8c08028c",
9211 => x"0c707080",
9212 => x"0b8c08fc",
9213 => x"050c8c08",
9214 => x"88050851",
9215 => x"7008822e",
9216 => x"0981060b",
9217 => x"0b0b0b88",
9218 => x"38810b8c",
9219 => x"08fc050c",
9220 => x"8c08fc05",
9221 => x"0870800c",
9222 => x"5150508c",
9223 => x"0c048c08",
9224 => x"028c0c70",
9225 => x"70800b8c",
9226 => x"08fc050c",
9227 => x"8c088805",
9228 => x"08517008",
9229 => x"842e0981",
9230 => x"060b0b0b",
9231 => x"0b883881",
9232 => x"0b8c08fc",
9233 => x"050c8c08",
9234 => x"fc050870",
9235 => x"800c5150",
9236 => x"508c0c04",
9237 => x"8c08028c",
9238 => x"0c707080",
9239 => x"0b8c08fc",
9240 => x"050c8c08",
9241 => x"88050851",
9242 => x"7008802e",
9243 => x"0b0b0b0b",
9244 => x"97388c08",
9245 => x"88050851",
9246 => x"7008812e",
9247 => x"0b0b0b0b",
9248 => x"87380b0b",
9249 => x"0b0b8839",
9250 => x"810b8c08",
9251 => x"fc050c8c",
9252 => x"08fc0508",
9253 => x"70800c51",
9254 => x"50508c0c",
9255 => x"048c0802",
9256 => x"8c0cffbc",
9257 => x"3d0d8c08",
9258 => x"8c05088c",
9259 => x"08900508",
9260 => x"5553728c",
9261 => x"08cc050c",
9262 => x"738c08d0",
9263 => x"050c8c08",
9264 => x"9405088c",
9265 => x"08980508",
9266 => x"5553728c",
9267 => x"08c4050c",
9268 => x"738c08c8",
9269 => x"050c8c08",
9270 => x"ec057053",
9271 => x"8c08cc05",
9272 => x"70535153",
9273 => x"0b0b0bbc",
9274 => x"f13f8c08",
9275 => x"d8057053",
9276 => x"8c08c405",
9277 => x"70535153",
9278 => x"0b0b0bbc",
9279 => x"dd3f8c08",
9280 => x"ec058c08",
9281 => x"c0050c8c",
9282 => x"08d8058c",
9283 => x"08ffbc05",
9284 => x"0c8c08c0",
9285 => x"0508510b",
9286 => x"0b0b9084",
9287 => x"3f800853",
9288 => x"72802e0b",
9289 => x"0b0b0b92",
9290 => x"388c08c0",
9291 => x"05088c08",
9292 => x"ffb8050c",
9293 => x"0b0b0b8e",
9294 => x"bb398c08",
9295 => x"ffbc0508",
9296 => x"510b0b0b",
9297 => x"8fda3f80",
9298 => x"08537280",
9299 => x"2e0b0b0b",
9300 => x"0b93388c",
9301 => x"08ffbc05",
9302 => x"088c08ff",
9303 => x"b8050c0b",
9304 => x"0b0b8e90",
9305 => x"398c08c0",
9306 => x"05088c08",
9307 => x"c005088c",
9308 => x"08ffbc05",
9309 => x"08841208",
9310 => x"84120832",
9311 => x"84140c8c",
9312 => x"08c00508",
9313 => x"54555555",
9314 => x"0b0b0b8e",
9315 => x"dd3f8008",
9316 => x"53720b0b",
9317 => x"0b0b9d38",
9318 => x"8c08c005",
9319 => x"08510b0b",
9320 => x"0b8e913f",
9321 => x"80085372",
9322 => x"0b0b0b0b",
9323 => x"87380b0b",
9324 => x"0b80c339",
9325 => x"8c08c005",
9326 => x"088c08ff",
9327 => x"bc050854",
9328 => x"54730873",
9329 => x"082e0981",
9330 => x"060b0b0b",
9331 => x"0b97380b",
9332 => x"0b0b8dcd",
9333 => x"3f800870",
9334 => x"8c08ffb8",
9335 => x"050c530b",
9336 => x"0b0b8d90",
9337 => x"398c08c0",
9338 => x"05088c08",
9339 => x"ffb8050c",
9340 => x"0b0b0b8c",
9341 => x"ff398c08",
9342 => x"ffbc0508",
9343 => x"510b0b0b",
9344 => x"8de83f80",
9345 => x"08537280",
9346 => x"2e0b0b0b",
9347 => x"0baf388c",
9348 => x"08c00508",
9349 => x"53805480",
9350 => x"55738c14",
9351 => x"0c749014",
9352 => x"0c8c08c0",
9353 => x"05085380",
9354 => x"0b88140c",
9355 => x"8c08c005",
9356 => x"088c08ff",
9357 => x"b8050c0b",
9358 => x"0b0b8cb8",
9359 => x"398c08ff",
9360 => x"bc050851",
9361 => x"0b0b0b8c",
9362 => x"eb3f8008",
9363 => x"5372802e",
9364 => x"0b0b0b0b",
9365 => x"9b388c08",
9366 => x"c0050853",
9367 => x"84730c8c",
9368 => x"08c00508",
9369 => x"8c08ffb8",
9370 => x"050c0b0b",
9371 => x"0b8c8539",
9372 => x"8c08c005",
9373 => x"088c08c0",
9374 => x"05088c08",
9375 => x"ffbc0508",
9376 => x"88120888",
9377 => x"12083188",
9378 => x"140c8c08",
9379 => x"c0050851",
9380 => x"55555590",
9381 => x"13088c14",
9382 => x"08545472",
9383 => x"8c08ffa8",
9384 => x"050c738c",
9385 => x"08ffac05",
9386 => x"0c8c08ff",
9387 => x"bc050853",
9388 => x"9013088c",
9389 => x"14085454",
9390 => x"728c08ff",
9391 => x"a0050c73",
9392 => x"8c08ffa4",
9393 => x"050c8c08",
9394 => x"ffa00508",
9395 => x"8c08ffa8",
9396 => x"0508260b",
9397 => x"0b0b0bb0",
9398 => x"388c08ff",
9399 => x"a005088c",
9400 => x"08ffa805",
9401 => x"082e0981",
9402 => x"060b0b0b",
9403 => x"81e9388c",
9404 => x"08ffa405",
9405 => x"088c08ff",
9406 => x"ac050826",
9407 => x"0b0b0b0b",
9408 => x"87380b0b",
9409 => x"0b81d039",
9410 => x"8c08ffa8",
9411 => x"05088c08",
9412 => x"ffac0508",
9413 => x"5553728c",
9414 => x"08ff9005",
9415 => x"0c738c08",
9416 => x"ff94050c",
9417 => x"8c08ff90",
9418 => x"05088c08",
9419 => x"ff940508",
9420 => x"5553728c",
9421 => x"08ff8805",
9422 => x"0c738c08",
9423 => x"ff8c050c",
9424 => x"8c08ff8c",
9425 => x"05088c08",
9426 => x"ff940508",
9427 => x"7012708c",
9428 => x"08ff8405",
9429 => x"0c525454",
9430 => x"810b8c08",
9431 => x"fefc050c",
9432 => x"8c08ff84",
9433 => x"05088c08",
9434 => x"ff8c0508",
9435 => x"54547274",
9436 => x"260b0b0b",
9437 => x"0b893880",
9438 => x"0b8c08fe",
9439 => x"fc050c8c",
9440 => x"08ff8805",
9441 => x"088c08ff",
9442 => x"90050870",
9443 => x"12708c08",
9444 => x"ff80050c",
9445 => x"8c08ff80",
9446 => x"05088c08",
9447 => x"fefc0508",
9448 => x"11708c08",
9449 => x"ff80050c",
9450 => x"53515254",
9451 => x"548c08ff",
9452 => x"8005088c",
9453 => x"08ff8405",
9454 => x"08555372",
9455 => x"8c08ffa8",
9456 => x"050c738c",
9457 => x"08ffac05",
9458 => x"0c8c08c0",
9459 => x"05088811",
9460 => x"08ff0588",
9461 => x"120c5388",
9462 => x"0a538054",
9463 => x"728c08ff",
9464 => x"b0050c73",
9465 => x"8c08ffb4",
9466 => x"050c8053",
9467 => x"8054728c",
9468 => x"08ff9805",
9469 => x"0c738c08",
9470 => x"ff9c050c",
9471 => x"8c08ffb0",
9472 => x"0508708c",
9473 => x"08ffb405",
9474 => x"08075153",
9475 => x"72802e0b",
9476 => x"0b0b849f",
9477 => x"388c08ff",
9478 => x"a005088c",
9479 => x"08ffa805",
9480 => x"08260b0b",
9481 => x"0b829838",
9482 => x"8c08ffa0",
9483 => x"05088c08",
9484 => x"ffa80508",
9485 => x"2e098106",
9486 => x"0b0b0b0b",
9487 => x"94388c08",
9488 => x"ffa40508",
9489 => x"8c08ffac",
9490 => x"0508260b",
9491 => x"0b0b81ef",
9492 => x"388c08ff",
9493 => x"9805088c",
9494 => x"08ffb005",
9495 => x"08078c08",
9496 => x"ff9c0508",
9497 => x"8c08ffb4",
9498 => x"05080755",
9499 => x"53728c08",
9500 => x"ff98050c",
9501 => x"738c08ff",
9502 => x"9c050c8c",
9503 => x"08ffa805",
9504 => x"088c08ff",
9505 => x"ac050855",
9506 => x"53728c08",
9507 => x"fef4050c",
9508 => x"738c08fe",
9509 => x"f8050c8c",
9510 => x"08ffa005",
9511 => x"088c08ff",
9512 => x"a4050855",
9513 => x"53728c08",
9514 => x"feec050c",
9515 => x"738c08fe",
9516 => x"f0050c8c",
9517 => x"08fef805",
9518 => x"088c08fe",
9519 => x"f0050871",
9520 => x"7131708c",
9521 => x"08fee805",
9522 => x"0c525454",
9523 => x"810b8c08",
9524 => x"fee0050c",
9525 => x"8c08fee8",
9526 => x"05088c08",
9527 => x"fef80508",
9528 => x"54547373",
9529 => x"260b0b0b",
9530 => x"0b893880",
9531 => x"0b8c08fe",
9532 => x"e0050c8c",
9533 => x"08fef405",
9534 => x"088c08fe",
9535 => x"ec050871",
9536 => x"7131708c",
9537 => x"08fee405",
9538 => x"0c8c08fe",
9539 => x"e4050870",
9540 => x"8c08fee0",
9541 => x"05083170",
9542 => x"8c08fee4",
9543 => x"050c5351",
9544 => x"5254548c",
9545 => x"08fee405",
9546 => x"088c08fe",
9547 => x"e8050855",
9548 => x"53728c08",
9549 => x"ffa8050c",
9550 => x"738c08ff",
9551 => x"ac050c8c",
9552 => x"08ffb005",
9553 => x"089f2b8c",
9554 => x"08ffb405",
9555 => x"08812a70",
9556 => x"72078c08",
9557 => x"ffb00508",
9558 => x"812a5656",
9559 => x"5656728c",
9560 => x"08ffb005",
9561 => x"0c738c08",
9562 => x"ffb4050c",
9563 => x"8c08ffa8",
9564 => x"05088c08",
9565 => x"ffac0508",
9566 => x"5553728c",
9567 => x"08fed805",
9568 => x"0c738c08",
9569 => x"fedc050c",
9570 => x"8c08fed8",
9571 => x"05088c08",
9572 => x"fedc0508",
9573 => x"5553728c",
9574 => x"08fed005",
9575 => x"0c738c08",
9576 => x"fed4050c",
9577 => x"8c08fed4",
9578 => x"05088c08",
9579 => x"fedc0508",
9580 => x"7012708c",
9581 => x"08fecc05",
9582 => x"0c525454",
9583 => x"810b8c08",
9584 => x"fec4050c",
9585 => x"8c08fecc",
9586 => x"05088c08",
9587 => x"fed40508",
9588 => x"54547274",
9589 => x"260b0b0b",
9590 => x"0b893880",
9591 => x"0b8c08fe",
9592 => x"c4050c8c",
9593 => x"08fed005",
9594 => x"088c08fe",
9595 => x"d8050870",
9596 => x"12708c08",
9597 => x"fec8050c",
9598 => x"8c08fec8",
9599 => x"05088c08",
9600 => x"fec40508",
9601 => x"11708c08",
9602 => x"fec8050c",
9603 => x"53515254",
9604 => x"548c08fe",
9605 => x"c805088c",
9606 => x"08fecc05",
9607 => x"08555372",
9608 => x"8c08ffa8",
9609 => x"050c738c",
9610 => x"08ffac05",
9611 => x"0c0b0b0b",
9612 => x"fbca398c",
9613 => x"08ff9805",
9614 => x"08800670",
9615 => x"8c08febc",
9616 => x"050c8c08",
9617 => x"ff9c0508",
9618 => x"81ff0670",
9619 => x"8c08fec0",
9620 => x"050c5454",
9621 => x"8c08febc",
9622 => x"05088c08",
9623 => x"fec00508",
9624 => x"5553728c",
9625 => x"08febc05",
9626 => x"0c738c08",
9627 => x"fec0050c",
9628 => x"8c08febc",
9629 => x"05085473",
9630 => x"0b0b0b83",
9631 => x"d0388c08",
9632 => x"fec00508",
9633 => x"53728180",
9634 => x"2e098106",
9635 => x"0b0b0b83",
9636 => x"bc388c08",
9637 => x"ff980508",
9638 => x"982b8c08",
9639 => x"ff9c0508",
9640 => x"882a7072",
9641 => x"078c08ff",
9642 => x"98050888",
9643 => x"2a718106",
9644 => x"51565656",
9645 => x"5672802e",
9646 => x"0b0b0b81",
9647 => x"bf388c08",
9648 => x"ff980508",
9649 => x"8c08ff9c",
9650 => x"05085553",
9651 => x"728c08fe",
9652 => x"b4050c73",
9653 => x"8c08feb8",
9654 => x"050c8053",
9655 => x"81805472",
9656 => x"8c08feac",
9657 => x"050c738c",
9658 => x"08feb005",
9659 => x"0c8c08fe",
9660 => x"b805088c",
9661 => x"08feb005",
9662 => x"08701270",
9663 => x"8c08fea8",
9664 => x"050c5254",
9665 => x"54810b8c",
9666 => x"08fea005",
9667 => x"0c8c08fe",
9668 => x"a805088c",
9669 => x"08feb805",
9670 => x"08545472",
9671 => x"74260b0b",
9672 => x"0b0b8938",
9673 => x"800b8c08",
9674 => x"fea0050c",
9675 => x"8c08feb4",
9676 => x"05088c08",
9677 => x"feac0508",
9678 => x"7012708c",
9679 => x"08fea405",
9680 => x"0c8c08fe",
9681 => x"a405088c",
9682 => x"08fea005",
9683 => x"0811708c",
9684 => x"08fea405",
9685 => x"0c535152",
9686 => x"54548c08",
9687 => x"fea40508",
9688 => x"8c08fea8",
9689 => x"05085553",
9690 => x"728c08ff",
9691 => x"98050c73",
9692 => x"8c08ff9c",
9693 => x"050c0b0b",
9694 => x"0b81d239",
9695 => x"8c08ffa8",
9696 => x"0508708c",
9697 => x"08ffac05",
9698 => x"08075153",
9699 => x"72802e0b",
9700 => x"0b0b81b9",
9701 => x"388c08ff",
9702 => x"9805088c",
9703 => x"08ff9c05",
9704 => x"08555372",
9705 => x"8c08fe98",
9706 => x"050c738c",
9707 => x"08fe9c05",
9708 => x"0c805381",
9709 => x"8054728c",
9710 => x"08fe9005",
9711 => x"0c738c08",
9712 => x"fe94050c",
9713 => x"8c08fe9c",
9714 => x"05088c08",
9715 => x"fe940508",
9716 => x"7012708c",
9717 => x"08fe8c05",
9718 => x"0c525454",
9719 => x"810b8c08",
9720 => x"fe84050c",
9721 => x"8c08fe8c",
9722 => x"05088c08",
9723 => x"fe9c0508",
9724 => x"54547274",
9725 => x"260b0b0b",
9726 => x"0b893880",
9727 => x"0b8c08fe",
9728 => x"84050c8c",
9729 => x"08fe9805",
9730 => x"088c08fe",
9731 => x"90050870",
9732 => x"12708c08",
9733 => x"fe88050c",
9734 => x"8c08fe88",
9735 => x"05088c08",
9736 => x"fe840508",
9737 => x"11708c08",
9738 => x"fe88050c",
9739 => x"53515254",
9740 => x"548c08fe",
9741 => x"8805088c",
9742 => x"08fe8c05",
9743 => x"08555372",
9744 => x"8c08ff98",
9745 => x"050c738c",
9746 => x"08ff9c05",
9747 => x"0c8c08c0",
9748 => x"0508558c",
9749 => x"08ff9805",
9750 => x"088c08ff",
9751 => x"9c050855",
9752 => x"53728c16",
9753 => x"0c739016",
9754 => x"0c8c08c0",
9755 => x"05088c08",
9756 => x"ffb8050c",
9757 => x"8c08ffb8",
9758 => x"0508708c",
9759 => x"08d4050c",
9760 => x"8c08d405",
9761 => x"08538c08",
9762 => x"88050852",
9763 => x"530b0b0b",
9764 => x"9c863f8c",
9765 => x"08880508",
9766 => x"800c80c6",
9767 => x"3d0d8c0c",
9768 => x"048c0802",
9769 => x"8c0c700b",
9770 => x"0b82f4b8",
9771 => x"70800c51",
9772 => x"508c0c04",
9773 => x"8c08028c",
9774 => x"0c707080",
9775 => x"0b8c08fc",
9776 => x"050c8c08",
9777 => x"88050851",
9778 => x"7008822e",
9779 => x"0981060b",
9780 => x"0b0b0b88",
9781 => x"38810b8c",
9782 => x"08fc050c",
9783 => x"8c08fc05",
9784 => x"0870800c",
9785 => x"5150508c",
9786 => x"0c048c08",
9787 => x"028c0c70",
9788 => x"70800b8c",
9789 => x"08fc050c",
9790 => x"8c088805",
9791 => x"08517008",
9792 => x"842e0981",
9793 => x"060b0b0b",
9794 => x"0b883881",
9795 => x"0b8c08fc",
9796 => x"050c8c08",
9797 => x"fc050870",
9798 => x"800c5150",
9799 => x"508c0c04",
9800 => x"8c08028c",
9801 => x"0c707080",
9802 => x"0b8c08fc",
9803 => x"050c8c08",
9804 => x"88050851",
9805 => x"7008802e",
9806 => x"0b0b0b0b",
9807 => x"97388c08",
9808 => x"88050851",
9809 => x"7008812e",
9810 => x"0b0b0b0b",
9811 => x"87380b0b",
9812 => x"0b0b8839",
9813 => x"810b8c08",
9814 => x"fc050c8c",
9815 => x"08fc0508",
9816 => x"70800c51",
9817 => x"50508c0c",
9818 => x"048c0802",
9819 => x"8c0cee3d",
9820 => x"0d8c0888",
9821 => x"05088c08",
9822 => x"8c050855",
9823 => x"53728c08",
9824 => x"d0050c73",
9825 => x"8c08d405",
9826 => x"0c8c0890",
9827 => x"05088c08",
9828 => x"94050855",
9829 => x"53728c08",
9830 => x"c8050c73",
9831 => x"8c08cc05",
9832 => x"0c8c08ec",
9833 => x"0570538c",
9834 => x"08d00570",
9835 => x"5351530b",
9836 => x"0b0baba6",
9837 => x"3f8c08d8",
9838 => x"0570538c",
9839 => x"08c80570",
9840 => x"5351530b",
9841 => x"0b0bab92",
9842 => x"3f8c08ec",
9843 => x"05705253",
9844 => x"0b0b0b80",
9845 => x"df3f8008",
9846 => x"53720b0b",
9847 => x"0b0b9e38",
9848 => x"8c08d805",
9849 => x"7052530b",
9850 => x"0b0b80c8",
9851 => x"3f800853",
9852 => x"720b0b0b",
9853 => x"0b87380b",
9854 => x"0b0b0b8e",
9855 => x"39810b8c",
9856 => x"08c4050c",
9857 => x"0b0b0b0b",
9858 => x"9e398c08",
9859 => x"d8057053",
9860 => x"8c08ec05",
9861 => x"70535153",
9862 => x"0b0b0bae",
9863 => x"c53f8008",
9864 => x"708c08c4",
9865 => x"050c538c",
9866 => x"08c40508",
9867 => x"800c943d",
9868 => x"0d8c0c04",
9869 => x"8c08028c",
9870 => x"0c707080",
9871 => x"0b8c08fc",
9872 => x"050c8c08",
9873 => x"88050851",
9874 => x"7008802e",
9875 => x"0b0b0b0b",
9876 => x"97388c08",
9877 => x"88050851",
9878 => x"7008812e",
9879 => x"0b0b0b0b",
9880 => x"87380b0b",
9881 => x"0b0b8839",
9882 => x"810b8c08",
9883 => x"fc050c8c",
9884 => x"08fc0508",
9885 => x"70800c51",
9886 => x"50508c0c",
9887 => x"048c0802",
9888 => x"8c0cee3d",
9889 => x"0d8c0888",
9890 => x"05088c08",
9891 => x"8c050855",
9892 => x"53728c08",
9893 => x"d0050c73",
9894 => x"8c08d405",
9895 => x"0c8c0890",
9896 => x"05088c08",
9897 => x"94050855",
9898 => x"53728c08",
9899 => x"c8050c73",
9900 => x"8c08cc05",
9901 => x"0c8c08ec",
9902 => x"0570538c",
9903 => x"08d00570",
9904 => x"5351530b",
9905 => x"0b0ba992",
9906 => x"3f8c08d8",
9907 => x"0570538c",
9908 => x"08c80570",
9909 => x"5351530b",
9910 => x"0b0ba8fe",
9911 => x"3f8c08ec",
9912 => x"05705253",
9913 => x"0b0b0b80",
9914 => x"df3f8008",
9915 => x"53720b0b",
9916 => x"0b0b9e38",
9917 => x"8c08d805",
9918 => x"7052530b",
9919 => x"0b0b80c8",
9920 => x"3f800853",
9921 => x"720b0b0b",
9922 => x"0b87380b",
9923 => x"0b0b0b8e",
9924 => x"39810b8c",
9925 => x"08c4050c",
9926 => x"0b0b0b0b",
9927 => x"9e398c08",
9928 => x"d8057053",
9929 => x"8c08ec05",
9930 => x"70535153",
9931 => x"0b0b0bac",
9932 => x"b13f8008",
9933 => x"708c08c4",
9934 => x"050c538c",
9935 => x"08c40508",
9936 => x"800c943d",
9937 => x"0d8c0c04",
9938 => x"8c08028c",
9939 => x"0c707080",
9940 => x"0b8c08fc",
9941 => x"050c8c08",
9942 => x"88050851",
9943 => x"7008802e",
9944 => x"0b0b0b0b",
9945 => x"97388c08",
9946 => x"88050851",
9947 => x"7008812e",
9948 => x"0b0b0b0b",
9949 => x"87380b0b",
9950 => x"0b0b8839",
9951 => x"810b8c08",
9952 => x"fc050c8c",
9953 => x"08fc0508",
9954 => x"70800c51",
9955 => x"50508c0c",
9956 => x"048c0802",
9957 => x"8c0cee3d",
9958 => x"0d8c0888",
9959 => x"05088c08",
9960 => x"8c050855",
9961 => x"53728c08",
9962 => x"d0050c73",
9963 => x"8c08d405",
9964 => x"0c8c0890",
9965 => x"05088c08",
9966 => x"94050855",
9967 => x"53728c08",
9968 => x"c8050c73",
9969 => x"8c08cc05",
9970 => x"0c8c08ec",
9971 => x"0570538c",
9972 => x"08d00570",
9973 => x"5351530b",
9974 => x"0b0ba6fe",
9975 => x"3f8c08d8",
9976 => x"0570538c",
9977 => x"08c80570",
9978 => x"5351530b",
9979 => x"0b0ba6ea",
9980 => x"3f8c08ec",
9981 => x"05705253",
9982 => x"0b0b0b80",
9983 => x"df3f8008",
9984 => x"53720b0b",
9985 => x"0b0b9e38",
9986 => x"8c08d805",
9987 => x"7052530b",
9988 => x"0b0b80c8",
9989 => x"3f800853",
9990 => x"720b0b0b",
9991 => x"0b87380b",
9992 => x"0b0b0b8e",
9993 => x"39ff0b8c",
9994 => x"08c4050c",
9995 => x"0b0b0b0b",
9996 => x"9e398c08",
9997 => x"d8057053",
9998 => x"8c08ec05",
9999 => x"70535153",
10000 => x"0b0b0baa",
10001 => x"9d3f8008",
10002 => x"708c08c4",
10003 => x"050c538c",
10004 => x"08c40508",
10005 => x"800c943d",
10006 => x"0d8c0c04",
10007 => x"8c08028c",
10008 => x"0c707080",
10009 => x"0b8c08fc",
10010 => x"050c8c08",
10011 => x"88050851",
10012 => x"7008802e",
10013 => x"0b0b0b0b",
10014 => x"97388c08",
10015 => x"88050851",
10016 => x"7008812e",
10017 => x"0b0b0b0b",
10018 => x"87380b0b",
10019 => x"0b0b8839",
10020 => x"810b8c08",
10021 => x"fc050c8c",
10022 => x"08fc0508",
10023 => x"70800c51",
10024 => x"50508c0c",
10025 => x"048c0802",
10026 => x"8c0cee3d",
10027 => x"0d8c0888",
10028 => x"05088c08",
10029 => x"8c050855",
10030 => x"53728c08",
10031 => x"d0050c73",
10032 => x"8c08d405",
10033 => x"0c8c0890",
10034 => x"05088c08",
10035 => x"94050855",
10036 => x"53728c08",
10037 => x"c8050c73",
10038 => x"8c08cc05",
10039 => x"0c8c08ec",
10040 => x"0570538c",
10041 => x"08d00570",
10042 => x"5351530b",
10043 => x"0b0ba4ea",
10044 => x"3f8c08d8",
10045 => x"0570538c",
10046 => x"08c80570",
10047 => x"5351530b",
10048 => x"0b0ba4d6",
10049 => x"3f8c08ec",
10050 => x"05705253",
10051 => x"0b0b0b80",
10052 => x"df3f8008",
10053 => x"53720b0b",
10054 => x"0b0b9e38",
10055 => x"8c08d805",
10056 => x"7052530b",
10057 => x"0b0b80c8",
10058 => x"3f800853",
10059 => x"720b0b0b",
10060 => x"0b87380b",
10061 => x"0b0b0b8e",
10062 => x"39810b8c",
10063 => x"08c4050c",
10064 => x"0b0b0b0b",
10065 => x"9e398c08",
10066 => x"d8057053",
10067 => x"8c08ec05",
10068 => x"70535153",
10069 => x"0b0b0ba8",
10070 => x"893f8008",
10071 => x"708c08c4",
10072 => x"050c538c",
10073 => x"08c40508",
10074 => x"800c943d",
10075 => x"0d8c0c04",
10076 => x"8c08028c",
10077 => x"0c707080",
10078 => x"0b8c08fc",
10079 => x"050c8c08",
10080 => x"88050851",
10081 => x"7008802e",
10082 => x"0b0b0b0b",
10083 => x"97388c08",
10084 => x"88050851",
10085 => x"7008812e",
10086 => x"0b0b0b0b",
10087 => x"87380b0b",
10088 => x"0b0b8839",
10089 => x"810b8c08",
10090 => x"fc050c8c",
10091 => x"08fc0508",
10092 => x"70800c51",
10093 => x"50508c0c",
10094 => x"048c0802",
10095 => x"8c0cee3d",
10096 => x"0d8c0888",
10097 => x"05088c08",
10098 => x"8c050855",
10099 => x"53728c08",
10100 => x"d0050c73",
10101 => x"8c08d405",
10102 => x"0c8c0890",
10103 => x"05088c08",
10104 => x"94050855",
10105 => x"53728c08",
10106 => x"c8050c73",
10107 => x"8c08cc05",
10108 => x"0c8c08ec",
10109 => x"0570538c",
10110 => x"08d00570",
10111 => x"5351530b",
10112 => x"0b0ba2d6",
10113 => x"3f8c08d8",
10114 => x"0570538c",
10115 => x"08c80570",
10116 => x"5351530b",
10117 => x"0b0ba2c2",
10118 => x"3f8c08ec",
10119 => x"05705253",
10120 => x"0b0b0b80",
10121 => x"df3f8008",
10122 => x"53720b0b",
10123 => x"0b0b9e38",
10124 => x"8c08d805",
10125 => x"7052530b",
10126 => x"0b0b80c8",
10127 => x"3f800853",
10128 => x"720b0b0b",
10129 => x"0b87380b",
10130 => x"0b0b0b8e",
10131 => x"39810b8c",
10132 => x"08c4050c",
10133 => x"0b0b0b0b",
10134 => x"9e398c08",
10135 => x"d8057053",
10136 => x"8c08ec05",
10137 => x"70535153",
10138 => x"0b0b0ba5",
10139 => x"f53f8008",
10140 => x"708c08c4",
10141 => x"050c538c",
10142 => x"08c40508",
10143 => x"800c943d",
10144 => x"0d8c0c04",
10145 => x"8c08028c",
10146 => x"0c707080",
10147 => x"0b8c08fc",
10148 => x"050c8c08",
10149 => x"88050851",
10150 => x"7008802e",
10151 => x"0b0b0b0b",
10152 => x"97388c08",
10153 => x"88050851",
10154 => x"7008812e",
10155 => x"0b0b0b0b",
10156 => x"87380b0b",
10157 => x"0b0b8839",
10158 => x"810b8c08",
10159 => x"fc050c8c",
10160 => x"08fc0508",
10161 => x"70800c51",
10162 => x"50508c0c",
10163 => x"048c0802",
10164 => x"8c0cf63d",
10165 => x"0d830b8c",
10166 => x"08ec050c",
10167 => x"800b8c08",
10168 => x"e8050c8c",
10169 => x"088c0508",
10170 => x"80250b0b",
10171 => x"0b0b8838",
10172 => x"810b8c08",
10173 => x"e8050c8c",
10174 => x"08e80508",
10175 => x"8c08f005",
10176 => x"0c8c088c",
10177 => x"05080b0b",
10178 => x"0b0b8e38",
10179 => x"820b8c08",
10180 => x"ec050c0b",
10181 => x"0b0b81b5",
10182 => x"39bc0b8c",
10183 => x"08f4050c",
10184 => x"8c08f005",
10185 => x"08802e0b",
10186 => x"0b0b80c9",
10187 => x"388c088c",
10188 => x"0508810a",
10189 => x"2e098106",
10190 => x"0b0b0b0b",
10191 => x"9b388f83",
10192 => x"0a53800b",
10193 => x"8c088805",
10194 => x"08565472",
10195 => x"750c7384",
10196 => x"160c0b0b",
10197 => x"0b818939",
10198 => x"8c088c05",
10199 => x"0830708c",
10200 => x"08fc050c",
10201 => x"709f2c70",
10202 => x"8c08f805",
10203 => x"0c51530b",
10204 => x"0b0b0b97",
10205 => x"398c088c",
10206 => x"0508708c",
10207 => x"08fc050c",
10208 => x"709f2c70",
10209 => x"8c08f805",
10210 => x"0c51538c",
10211 => x"08f80508",
10212 => x"f00a260b",
10213 => x"0b0b0bb5",
10214 => x"388c08fc",
10215 => x"05089f2a",
10216 => x"8c08f805",
10217 => x"08107072",
10218 => x"078c08f8",
10219 => x"050c8c08",
10220 => x"fc050810",
10221 => x"8c08fc05",
10222 => x"0c8c08f4",
10223 => x"0508ff05",
10224 => x"8c08f405",
10225 => x"0c54540b",
10226 => x"0b0bffbf",
10227 => x"398c08ec",
10228 => x"0570538c",
10229 => x"08880508",
10230 => x"52530b0b",
10231 => x"0b8db93f",
10232 => x"8c088805",
10233 => x"08800c8c",
10234 => x"3d0d8c0c",
10235 => x"048c0802",
10236 => x"8c0cec3d",
10237 => x"0d8c0888",
10238 => x"05088c08",
10239 => x"8c050857",
10240 => x"55748c08",
10241 => x"e0050c75",
10242 => x"8c08e405",
10243 => x"0c8c08ec",
10244 => x"0570538c",
10245 => x"08e00570",
10246 => x"5351550b",
10247 => x"0b0b9eba",
10248 => x"3f8c08ec",
10249 => x"05705255",
10250 => x"0b0b0b83",
10251 => x"d93f8008",
10252 => x"5574802e",
10253 => x"0b0b0b0b",
10254 => x"8e38800b",
10255 => x"8c08d405",
10256 => x"0c0b0b0b",
10257 => x"82b4398c",
10258 => x"08ec0570",
10259 => x"52550b0b",
10260 => x"0b82ea3f",
10261 => x"80085574",
10262 => x"802e0b0b",
10263 => x"0b0b8e38",
10264 => x"800b8c08",
10265 => x"d4050c0b",
10266 => x"0b0b828e",
10267 => x"398c08ec",
10268 => x"05705255",
10269 => x"0b0b0b82",
10270 => x"8e3f8008",
10271 => x"5574802e",
10272 => x"0b0b0b0b",
10273 => x"b4388c08",
10274 => x"f0050880",
10275 => x"2e0b0b0b",
10276 => x"0b8f3881",
10277 => x"0a0b8c08",
10278 => x"d0050c0b",
10279 => x"0b0b0b89",
10280 => x"39fe0a0b",
10281 => x"8c08d005",
10282 => x"0c8c08d0",
10283 => x"05088c08",
10284 => x"d4050c0b",
10285 => x"0b0b81c2",
10286 => x"398c08f4",
10287 => x"05088025",
10288 => x"0b0b0b0b",
10289 => x"8e38800b",
10290 => x"8c08d405",
10291 => x"0c0b0b0b",
10292 => x"81a8399e",
10293 => x"0b8c08f4",
10294 => x"0508250b",
10295 => x"0b0b0bb4",
10296 => x"388c08f0",
10297 => x"0508802e",
10298 => x"0b0b0b0b",
10299 => x"8f38810a",
10300 => x"0b8c08cc",
10301 => x"050c0b0b",
10302 => x"0b0b8939",
10303 => x"fe0a0b8c",
10304 => x"08cc050c",
10305 => x"8c08cc05",
10306 => x"088c08d4",
10307 => x"050c0b0b",
10308 => x"0b80e739",
10309 => x"bc0b8c08",
10310 => x"f4050831",
10311 => x"8c08d805",
10312 => x"71565855",
10313 => x"8c08f805",
10314 => x"088c08fc",
10315 => x"05085755",
10316 => x"74527553",
10317 => x"76510b0b",
10318 => x"0b88d53f",
10319 => x"8c08d805",
10320 => x"088c08dc",
10321 => x"0508708c",
10322 => x"08e8050c",
10323 => x"8c08e805",
10324 => x"088c08c8",
10325 => x"050c5755",
10326 => x"8c08f005",
10327 => x"08802e0b",
10328 => x"0b0b0b8c",
10329 => x"388c08c8",
10330 => x"0508308c",
10331 => x"08c8050c",
10332 => x"8c08c805",
10333 => x"088c08d4",
10334 => x"050c8c08",
10335 => x"d4050880",
10336 => x"0c963d0d",
10337 => x"8c0c048c",
10338 => x"08028c0c",
10339 => x"7070800b",
10340 => x"8c08fc05",
10341 => x"0c8c0888",
10342 => x"05085170",
10343 => x"08842e09",
10344 => x"81060b0b",
10345 => x"0b0b8838",
10346 => x"810b8c08",
10347 => x"fc050c8c",
10348 => x"08fc0508",
10349 => x"70800c51",
10350 => x"50508c0c",
10351 => x"048c0802",
10352 => x"8c0c7070",
10353 => x"800b8c08",
10354 => x"fc050c8c",
10355 => x"08880508",
10356 => x"51700880",
10357 => x"2e0b0b0b",
10358 => x"0b97388c",
10359 => x"08880508",
10360 => x"51700881",
10361 => x"2e0b0b0b",
10362 => x"0b87380b",
10363 => x"0b0b0b88",
10364 => x"39810b8c",
10365 => x"08fc050c",
10366 => x"8c08fc05",
10367 => x"0870800c",
10368 => x"5150508c",
10369 => x"0c048c08",
10370 => x"028c0c70",
10371 => x"70800b8c",
10372 => x"08fc050c",
10373 => x"8c088805",
10374 => x"08517008",
10375 => x"822e0981",
10376 => x"060b0b0b",
10377 => x"0b883881",
10378 => x"0b8c08fc",
10379 => x"050c8c08",
10380 => x"fc050870",
10381 => x"800c5150",
10382 => x"508c0c04",
10383 => x"8c08028c",
10384 => x"0c707070",
10385 => x"7080538c",
10386 => x"088c0508",
10387 => x"528c0888",
10388 => x"0508510b",
10389 => x"0bfdccbf",
10390 => x"3f800870",
10391 => x"800c5450",
10392 => x"5050508c",
10393 => x"0c048c08",
10394 => x"028c0c70",
10395 => x"70707081",
10396 => x"538c088c",
10397 => x"0508528c",
10398 => x"08880508",
10399 => x"510b0bfd",
10400 => x"cc953f80",
10401 => x"0870800c",
10402 => x"54505050",
10403 => x"508c0c04",
10404 => x"8c08028c",
10405 => x"0c707080",
10406 => x"0b8c08fc",
10407 => x"050c8c08",
10408 => x"88050881",
10409 => x"06ff1170",
10410 => x"09708c08",
10411 => x"8c050806",
10412 => x"8c08fc05",
10413 => x"08118c08",
10414 => x"fc050c8c",
10415 => x"08880508",
10416 => x"812a8c08",
10417 => x"88050c8c",
10418 => x"088c0508",
10419 => x"108c088c",
10420 => x"050c5151",
10421 => x"51518c08",
10422 => x"88050880",
10423 => x"2e0b0b0b",
10424 => x"0b87380b",
10425 => x"0b0bffb6",
10426 => x"398c08fc",
10427 => x"05087080",
10428 => x"0c515050",
10429 => x"8c0c048c",
10430 => x"08028c0c",
10431 => x"eb3d0d80",
10432 => x"0b8c08f0",
10433 => x"050c800b",
10434 => x"8c08f405",
10435 => x"0c8c088c",
10436 => x"05088c08",
10437 => x"90050856",
10438 => x"54738c08",
10439 => x"f0050c74",
10440 => x"8c08f405",
10441 => x"0c8c08f8",
10442 => x"058c08f0",
10443 => x"05565688",
10444 => x"70547553",
10445 => x"7652540b",
10446 => x"0bfdcccf",
10447 => x"3f800b8c",
10448 => x"08e8050c",
10449 => x"800b8c08",
10450 => x"ec050c8c",
10451 => x"08940508",
10452 => x"8c089805",
10453 => x"08565473",
10454 => x"8c08e805",
10455 => x"0c748c08",
10456 => x"ec050c8c",
10457 => x"08f0058c",
10458 => x"08e80556",
10459 => x"56887054",
10460 => x"75537652",
10461 => x"540b0bfd",
10462 => x"cc913f80",
10463 => x"0b8c08e8",
10464 => x"050c800b",
10465 => x"8c08ec05",
10466 => x"0c8c08fc",
10467 => x"050883ff",
10468 => x"ff068c08",
10469 => x"cc050c8c",
10470 => x"08fc0508",
10471 => x"902a8c08",
10472 => x"c4050c8c",
10473 => x"08f40508",
10474 => x"83ffff06",
10475 => x"8c08c805",
10476 => x"0c8c08f4",
10477 => x"0508902a",
10478 => x"8c08c005",
10479 => x"0c8c08cc",
10480 => x"05088c08",
10481 => x"c8050829",
10482 => x"708c08dc",
10483 => x"050c8c08",
10484 => x"cc05088c",
10485 => x"08c00508",
10486 => x"29708c08",
10487 => x"d8050c8c",
10488 => x"08c40508",
10489 => x"8c08c805",
10490 => x"0829708c",
10491 => x"08d4050c",
10492 => x"8c08c405",
10493 => x"088c08c0",
10494 => x"05082970",
10495 => x"8c08d005",
10496 => x"0c8c08dc",
10497 => x"0508902a",
10498 => x"8c08d805",
10499 => x"08118c08",
10500 => x"d8050c8c",
10501 => x"08d80508",
10502 => x"8c08d405",
10503 => x"08058c08",
10504 => x"d8050c51",
10505 => x"51515154",
10506 => x"8c08d805",
10507 => x"088c08d4",
10508 => x"0508270b",
10509 => x"0b0b0b8f",
10510 => x"388c08d0",
10511 => x"05088480",
10512 => x"80058c08",
10513 => x"d0050c8c",
10514 => x"08d80508",
10515 => x"902a8c08",
10516 => x"d0050811",
10517 => x"8c08e005",
10518 => x"0c8c08d8",
10519 => x"050883ff",
10520 => x"ff067090",
10521 => x"2b8c08dc",
10522 => x"050883ff",
10523 => x"ff067012",
10524 => x"8c08e405",
10525 => x"0c525751",
10526 => x"548c08e0",
10527 => x"05088c08",
10528 => x"e4050856",
10529 => x"54738c08",
10530 => x"e8050c74",
10531 => x"8c08ec05",
10532 => x"0c8c08fc",
10533 => x"05088c08",
10534 => x"f0050829",
10535 => x"8c08f805",
10536 => x"088c08f4",
10537 => x"05082970",
10538 => x"128c08e8",
10539 => x"0508118c",
10540 => x"08e8050c",
10541 => x"5155558c",
10542 => x"08e80508",
10543 => x"8c08ec05",
10544 => x"088c0888",
10545 => x"05085856",
10546 => x"5473760c",
10547 => x"7484170c",
10548 => x"8c088805",
10549 => x"08800c97",
10550 => x"3d0d8c0c",
10551 => x"048c0802",
10552 => x"8c0cf63d",
10553 => x"0d800b8c",
10554 => x"08f0050c",
10555 => x"800b8c08",
10556 => x"f4050c8c",
10557 => x"088c0508",
10558 => x"8c089005",
10559 => x"08565473",
10560 => x"8c08f005",
10561 => x"0c748c08",
10562 => x"f4050c8c",
10563 => x"08f8058c",
10564 => x"08f00556",
10565 => x"56887054",
10566 => x"75537652",
10567 => x"540b0bfd",
10568 => x"c8e93f80",
10569 => x"0b8c08f0",
10570 => x"050c800b",
10571 => x"8c08f405",
10572 => x"0c8c08f8",
10573 => x"0508308c",
10574 => x"08ec050c",
10575 => x"8c08fc05",
10576 => x"08802e0b",
10577 => x"0b0b0b8d",
10578 => x"388c08ec",
10579 => x"0508ff05",
10580 => x"8c08ec05",
10581 => x"0c8c08ec",
10582 => x"05088c08",
10583 => x"f0050c8c",
10584 => x"08fc0508",
10585 => x"308c08f4",
10586 => x"050c8c08",
10587 => x"f005088c",
10588 => x"08f40508",
10589 => x"8c088805",
10590 => x"08585654",
10591 => x"73760c74",
10592 => x"84170c8c",
10593 => x"08880508",
10594 => x"800c8c3d",
10595 => x"0d8c0c04",
10596 => x"8c08028c",
10597 => x"0cf53d0d",
10598 => x"8c089405",
10599 => x"080b0b0b",
10600 => x"0ba0388c",
10601 => x"088c0508",
10602 => x"8c089005",
10603 => x"088c0888",
10604 => x"05085856",
10605 => x"5473760c",
10606 => x"7484170c",
10607 => x"0b0b0b81",
10608 => x"ca39800b",
10609 => x"8c08f005",
10610 => x"0c800b8c",
10611 => x"08f4050c",
10612 => x"8c088c05",
10613 => x"088c0890",
10614 => x"05085654",
10615 => x"738c08f0",
10616 => x"050c748c",
10617 => x"08f4050c",
10618 => x"8c08f805",
10619 => x"8c08f005",
10620 => x"56568870",
10621 => x"54755376",
10622 => x"52540b0b",
10623 => x"fdc78c3f",
10624 => x"a00b8c08",
10625 => x"94050831",
10626 => x"8c08ec05",
10627 => x"0c8c08ec",
10628 => x"05088024",
10629 => x"0b0b0b0b",
10630 => x"a138800b",
10631 => x"8c08f005",
10632 => x"0c8c08ec",
10633 => x"0508308c",
10634 => x"08f80508",
10635 => x"712a8c08",
10636 => x"f4050c54",
10637 => x"0b0b0b0b",
10638 => x"b9398c08",
10639 => x"f805088c",
10640 => x"08ec0508",
10641 => x"2b8c08e8",
10642 => x"050c8c08",
10643 => x"f805088c",
10644 => x"08940508",
10645 => x"2a8c08f0",
10646 => x"050c8c08",
10647 => x"fc05088c",
10648 => x"08940508",
10649 => x"2a708c08",
10650 => x"e8050807",
10651 => x"8c08f405",
10652 => x"0c548c08",
10653 => x"f005088c",
10654 => x"08f40508",
10655 => x"8c088805",
10656 => x"08585654",
10657 => x"73760c74",
10658 => x"84170c8c",
10659 => x"08880508",
10660 => x"800c8d3d",
10661 => x"0d8c0c04",
10662 => x"8c08028c",
10663 => x"0cc73d0d",
10664 => x"8c088c05",
10665 => x"08559015",
10666 => x"088c1608",
10667 => x"5656748c",
10668 => x"08f0050c",
10669 => x"758c08f4",
10670 => x"050c8c08",
10671 => x"8c050884",
10672 => x"11088c08",
10673 => x"ec050c55",
10674 => x"800b8c08",
10675 => x"e8050c8c",
10676 => x"088c0508",
10677 => x"510b0b0b",
10678 => x"90b73f80",
10679 => x"08557480",
10680 => x"2e0b0b0b",
10681 => x"0bad388f",
10682 => x"ff0b8c08",
10683 => x"e8050c8c",
10684 => x"08f00508",
10685 => x"a0808007",
10686 => x"8c08f405",
10687 => x"08800757",
10688 => x"55748c08",
10689 => x"f0050c75",
10690 => x"8c08f405",
10691 => x"0c0b0b0b",
10692 => x"8df4398c",
10693 => x"088c0508",
10694 => x"510b0b0b",
10695 => x"8fbd3f80",
10696 => x"08557480",
10697 => x"2e0b0b0b",
10698 => x"0b9f388f",
10699 => x"ff0b8c08",
10700 => x"e8050c80",
10701 => x"55805674",
10702 => x"8c08f005",
10703 => x"0c758c08",
10704 => x"f4050c0b",
10705 => x"0b0b8dbe",
10706 => x"398c088c",
10707 => x"0508510b",
10708 => x"0b0b8ed1",
10709 => x"3f800855",
10710 => x"74802e0b",
10711 => x"0b0b0b9e",
10712 => x"38800b8c",
10713 => x"08e8050c",
10714 => x"80558056",
10715 => x"748c08f0",
10716 => x"050c758c",
10717 => x"08f4050c",
10718 => x"0b0b0b8d",
10719 => x"89398c08",
10720 => x"f0050870",
10721 => x"8c08f405",
10722 => x"08075155",
10723 => x"740b0b0b",
10724 => x"0b8e3880",
10725 => x"0b8c08e8",
10726 => x"050c0b0b",
10727 => x"0b8ce739",
10728 => x"8c088c05",
10729 => x"08558815",
10730 => x"08f88225",
10731 => x"0b0b0b87",
10732 => x"af388c08",
10733 => x"8c0508f8",
10734 => x"820b8812",
10735 => x"08318c08",
10736 => x"e4050c55",
10737 => x"800b8c08",
10738 => x"e8050cb8",
10739 => x"0b8c08e4",
10740 => x"0508250b",
10741 => x"0b0b0b97",
10742 => x"38805580",
10743 => x"56748c08",
10744 => x"f0050c75",
10745 => x"8c08f405",
10746 => x"0c0b0b0b",
10747 => x"82b03980",
10748 => x"0b8c08e0",
10749 => x"050c8c08",
10750 => x"d8055780",
10751 => x"55810b8c",
10752 => x"08e40508",
10753 => x"55567452",
10754 => x"75537651",
10755 => x"0b0bfdbc",
10756 => x"ab3f8c08",
10757 => x"d805088c",
10758 => x"08dc0508",
10759 => x"5755748c",
10760 => x"08d0050c",
10761 => x"758c08d4",
10762 => x"050cff56",
10763 => x"ff57758c",
10764 => x"08c8050c",
10765 => x"768c08cc",
10766 => x"050c8c08",
10767 => x"d405088c",
10768 => x"08cc0508",
10769 => x"7012708c",
10770 => x"08c4050c",
10771 => x"52565781",
10772 => x"0b8c08ff",
10773 => x"bc050c8c",
10774 => x"08c40508",
10775 => x"8c08d405",
10776 => x"08585676",
10777 => x"76260b0b",
10778 => x"0b0b8938",
10779 => x"800b8c08",
10780 => x"ffbc050c",
10781 => x"8c08d005",
10782 => x"088c08c8",
10783 => x"05087012",
10784 => x"708c08c0",
10785 => x"050c8c08",
10786 => x"c005088c",
10787 => x"08ffbc05",
10788 => x"0811708c",
10789 => x"08c0050c",
10790 => x"8c08c005",
10791 => x"08708c08",
10792 => x"f0050806",
10793 => x"8c08c405",
10794 => x"08708c08",
10795 => x"f4050806",
10796 => x"72707207",
10797 => x"51525752",
10798 => x"5252525a",
10799 => x"52575576",
10800 => x"802e0b0b",
10801 => x"0b0b8838",
10802 => x"810b8c08",
10803 => x"e0050c8c",
10804 => x"08d8058c",
10805 => x"08e40508",
10806 => x"55578c08",
10807 => x"f005088c",
10808 => x"08f40508",
10809 => x"57557452",
10810 => x"75537651",
10811 => x"0b0b0bf9",
10812 => x"9f3f8c08",
10813 => x"d805088c",
10814 => x"08dc0508",
10815 => x"8c08e005",
10816 => x"089f2c8c",
10817 => x"08e00508",
10818 => x"71707507",
10819 => x"8c08f005",
10820 => x"0c737207",
10821 => x"8c08f405",
10822 => x"0c59595b",
10823 => x"59578c08",
10824 => x"f0050880",
10825 => x"06708c08",
10826 => x"ffb4050c",
10827 => x"8c08f405",
10828 => x"0881ff06",
10829 => x"708c08ff",
10830 => x"b8050c57",
10831 => x"558c08ff",
10832 => x"b405088c",
10833 => x"08ffb805",
10834 => x"08575574",
10835 => x"8c08ffb4",
10836 => x"050c758c",
10837 => x"08ffb805",
10838 => x"0c8c08ff",
10839 => x"b4050856",
10840 => x"750b0b0b",
10841 => x"81f8388c",
10842 => x"08ffb805",
10843 => x"08577681",
10844 => x"802e0981",
10845 => x"060b0b0b",
10846 => x"81e4388c",
10847 => x"08f00508",
10848 => x"982b8c08",
10849 => x"f4050888",
10850 => x"2a707207",
10851 => x"8c08f005",
10852 => x"08882a71",
10853 => x"81065158",
10854 => x"58585874",
10855 => x"802e0b0b",
10856 => x"0b82ef38",
10857 => x"8c08f005",
10858 => x"088c08f4",
10859 => x"05085755",
10860 => x"748c08ff",
10861 => x"ac050c75",
10862 => x"8c08ffb0",
10863 => x"050c8056",
10864 => x"81805775",
10865 => x"8c08ffa4",
10866 => x"050c768c",
10867 => x"08ffa805",
10868 => x"0c8c08ff",
10869 => x"b005088c",
10870 => x"08ffa805",
10871 => x"08701270",
10872 => x"8c08ffa0",
10873 => x"050c5256",
10874 => x"57810b8c",
10875 => x"08ff9805",
10876 => x"0c8c08ff",
10877 => x"a005088c",
10878 => x"08ffb005",
10879 => x"08585676",
10880 => x"76260b0b",
10881 => x"0b0b8938",
10882 => x"800b8c08",
10883 => x"ff98050c",
10884 => x"8c08ffac",
10885 => x"05088c08",
10886 => x"ffa40508",
10887 => x"7012708c",
10888 => x"08ff9c05",
10889 => x"0c8c08ff",
10890 => x"9c05088c",
10891 => x"08ff9805",
10892 => x"0811708c",
10893 => x"08ff9c05",
10894 => x"0c525a52",
10895 => x"57558c08",
10896 => x"ff9c0508",
10897 => x"8c08ffa0",
10898 => x"05085755",
10899 => x"748c08f0",
10900 => x"050c758c",
10901 => x"08f4050c",
10902 => x"0b0b0b81",
10903 => x"b5398c08",
10904 => x"f005088c",
10905 => x"08f40508",
10906 => x"5856758c",
10907 => x"08ff9005",
10908 => x"0c768c08",
10909 => x"ff94050c",
10910 => x"805580ff",
10911 => x"56748c08",
10912 => x"ff88050c",
10913 => x"758c08ff",
10914 => x"8c050c8c",
10915 => x"08ff9405",
10916 => x"088c08ff",
10917 => x"8c050870",
10918 => x"12708c08",
10919 => x"ff84050c",
10920 => x"52585681",
10921 => x"0b8c08fe",
10922 => x"fc050c8c",
10923 => x"08ff8405",
10924 => x"088c08ff",
10925 => x"94050857",
10926 => x"55757526",
10927 => x"0b0b0b0b",
10928 => x"8938800b",
10929 => x"8c08fefc",
10930 => x"050c8c08",
10931 => x"ff900508",
10932 => x"8c08ff88",
10933 => x"05087012",
10934 => x"708c08ff",
10935 => x"80050c8c",
10936 => x"08ff8005",
10937 => x"088c08fe",
10938 => x"fc050811",
10939 => x"708c08ff",
10940 => x"80050c53",
10941 => x"59525657",
10942 => x"8c08ff80",
10943 => x"05088c08",
10944 => x"ff840508",
10945 => x"5755748c",
10946 => x"08f0050c",
10947 => x"758c08f4",
10948 => x"050c8c08",
10949 => x"f00508f0",
10950 => x"0a260b0b",
10951 => x"0b0b8738",
10952 => x"0b0b0b0b",
10953 => x"8d398c08",
10954 => x"e8050881",
10955 => x"058c08e8",
10956 => x"050c8c08",
10957 => x"f0050898",
10958 => x"2b8c08f4",
10959 => x"0508882a",
10960 => x"7072078c",
10961 => x"08f00508",
10962 => x"882a5858",
10963 => x"5858748c",
10964 => x"08f0050c",
10965 => x"758c08f4",
10966 => x"050c0b0b",
10967 => x"0b85a739",
10968 => x"8c088c05",
10969 => x"085587ff",
10970 => x"0b881608",
10971 => x"250b0b0b",
10972 => x"0b9f388f",
10973 => x"ff0b8c08",
10974 => x"e8050c80",
10975 => x"55805674",
10976 => x"8c08f005",
10977 => x"0c758c08",
10978 => x"f4050c0b",
10979 => x"0b0b84f6",
10980 => x"398c088c",
10981 => x"05088811",
10982 => x"0887ff05",
10983 => x"8c08e805",
10984 => x"0c8c08f0",
10985 => x"05088006",
10986 => x"708c08fe",
10987 => x"f4050c8c",
10988 => x"08f40508",
10989 => x"81ff0670",
10990 => x"8c08fef8",
10991 => x"050c5957",
10992 => x"558c08fe",
10993 => x"f405088c",
10994 => x"08fef805",
10995 => x"08575574",
10996 => x"8c08fef4",
10997 => x"050c758c",
10998 => x"08fef805",
10999 => x"0c8c08fe",
11000 => x"f4050856",
11001 => x"750b0b0b",
11002 => x"81f8388c",
11003 => x"08fef805",
11004 => x"08577681",
11005 => x"802e0981",
11006 => x"060b0b0b",
11007 => x"81e4388c",
11008 => x"08f00508",
11009 => x"982b8c08",
11010 => x"f4050888",
11011 => x"2a707207",
11012 => x"8c08f005",
11013 => x"08882a71",
11014 => x"81065158",
11015 => x"58585874",
11016 => x"802e0b0b",
11017 => x"0b82ef38",
11018 => x"8c08f005",
11019 => x"088c08f4",
11020 => x"05085755",
11021 => x"748c08fe",
11022 => x"ec050c75",
11023 => x"8c08fef0",
11024 => x"050c8056",
11025 => x"81805775",
11026 => x"8c08fee4",
11027 => x"050c768c",
11028 => x"08fee805",
11029 => x"0c8c08fe",
11030 => x"f005088c",
11031 => x"08fee805",
11032 => x"08701270",
11033 => x"8c08fee0",
11034 => x"050c5256",
11035 => x"57810b8c",
11036 => x"08fed805",
11037 => x"0c8c08fe",
11038 => x"e005088c",
11039 => x"08fef005",
11040 => x"08585676",
11041 => x"76260b0b",
11042 => x"0b0b8938",
11043 => x"800b8c08",
11044 => x"fed8050c",
11045 => x"8c08feec",
11046 => x"05088c08",
11047 => x"fee40508",
11048 => x"7012708c",
11049 => x"08fedc05",
11050 => x"0c8c08fe",
11051 => x"dc05088c",
11052 => x"08fed805",
11053 => x"0811708c",
11054 => x"08fedc05",
11055 => x"0c525a52",
11056 => x"57558c08",
11057 => x"fedc0508",
11058 => x"8c08fee0",
11059 => x"05085755",
11060 => x"748c08f0",
11061 => x"050c758c",
11062 => x"08f4050c",
11063 => x"0b0b0b81",
11064 => x"b5398c08",
11065 => x"f005088c",
11066 => x"08f40508",
11067 => x"5856758c",
11068 => x"08fed005",
11069 => x"0c768c08",
11070 => x"fed4050c",
11071 => x"805580ff",
11072 => x"56748c08",
11073 => x"fec8050c",
11074 => x"758c08fe",
11075 => x"cc050c8c",
11076 => x"08fed405",
11077 => x"088c08fe",
11078 => x"cc050870",
11079 => x"12708c08",
11080 => x"fec4050c",
11081 => x"52585681",
11082 => x"0b8c08fe",
11083 => x"bc050c8c",
11084 => x"08fec405",
11085 => x"088c08fe",
11086 => x"d4050857",
11087 => x"55757526",
11088 => x"0b0b0b0b",
11089 => x"8938800b",
11090 => x"8c08febc",
11091 => x"050c8c08",
11092 => x"fed00508",
11093 => x"8c08fec8",
11094 => x"05087012",
11095 => x"708c08fe",
11096 => x"c0050c8c",
11097 => x"08fec005",
11098 => x"088c08fe",
11099 => x"bc050811",
11100 => x"708c08fe",
11101 => x"c0050c53",
11102 => x"59525657",
11103 => x"8c08fec0",
11104 => x"05088c08",
11105 => x"fec40508",
11106 => x"5755748c",
11107 => x"08f0050c",
11108 => x"758c08f4",
11109 => x"050c8c08",
11110 => x"f00508f8",
11111 => x"0a260b0b",
11112 => x"0b0b8738",
11113 => x"0b0b0b0b",
11114 => x"b5398c08",
11115 => x"f005089f",
11116 => x"2b8c08f4",
11117 => x"0508812a",
11118 => x"7072078c",
11119 => x"08f00508",
11120 => x"812a5858",
11121 => x"5858748c",
11122 => x"08f0050c",
11123 => x"758c08f4",
11124 => x"050c8c08",
11125 => x"e8050881",
11126 => x"058c08e8",
11127 => x"050c8c08",
11128 => x"f0050898",
11129 => x"2b8c08f4",
11130 => x"0508882a",
11131 => x"7072078c",
11132 => x"08f00508",
11133 => x"882a5858",
11134 => x"5858748c",
11135 => x"08f0050c",
11136 => x"758c08f4",
11137 => x"050c8c08",
11138 => x"f00508bf",
11139 => x"ffff068c",
11140 => x"08f8050c",
11141 => x"8c08f405",
11142 => x"08ff068c",
11143 => x"08fc050c",
11144 => x"8c08e805",
11145 => x"08568070",
11146 => x"8006778f",
11147 => x"ff067094",
11148 => x"2b535a58",
11149 => x"55800b8c",
11150 => x"08f80508",
11151 => x"76078c08",
11152 => x"f8050c70",
11153 => x"8c08fc05",
11154 => x"08078c08",
11155 => x"fc050c8c",
11156 => x"08ec0508",
11157 => x"51568070",
11158 => x"80067781",
11159 => x"06709f2b",
11160 => x"535a5855",
11161 => x"800b8c08",
11162 => x"f8050876",
11163 => x"078c08f8",
11164 => x"050c708c",
11165 => x"08fc0508",
11166 => x"078c08fc",
11167 => x"050c568c",
11168 => x"08f80508",
11169 => x"8c08fc05",
11170 => x"088c0888",
11171 => x"05085957",
11172 => x"5574770c",
11173 => x"7584180c",
11174 => x"8c088805",
11175 => x"08800cbb",
11176 => x"3d0d8c0c",
11177 => x"048c0802",
11178 => x"8c0c7070",
11179 => x"800b8c08",
11180 => x"fc050c8c",
11181 => x"08880508",
11182 => x"51700882",
11183 => x"2e098106",
11184 => x"0b0b0b0b",
11185 => x"8838810b",
11186 => x"8c08fc05",
11187 => x"0c8c08fc",
11188 => x"05087080",
11189 => x"0c515050",
11190 => x"8c0c048c",
11191 => x"08028c0c",
11192 => x"7070800b",
11193 => x"8c08fc05",
11194 => x"0c8c0888",
11195 => x"05085170",
11196 => x"08842e09",
11197 => x"81060b0b",
11198 => x"0b0b8838",
11199 => x"810b8c08",
11200 => x"fc050c8c",
11201 => x"08fc0508",
11202 => x"70800c51",
11203 => x"50508c0c",
11204 => x"048c0802",
11205 => x"8c0c7070",
11206 => x"800b8c08",
11207 => x"fc050c8c",
11208 => x"08880508",
11209 => x"51700880",
11210 => x"2e0b0b0b",
11211 => x"0b97388c",
11212 => x"08880508",
11213 => x"51700881",
11214 => x"2e0b0b0b",
11215 => x"0b87380b",
11216 => x"0b0b0b88",
11217 => x"39810b8c",
11218 => x"08fc050c",
11219 => x"8c08fc05",
11220 => x"0870800c",
11221 => x"5150508c",
11222 => x"0c048c08",
11223 => x"028c0cf8",
11224 => x"3d0d8c08",
11225 => x"88050870",
11226 => x"08bfffff",
11227 => x"068c08f8",
11228 => x"050c8411",
11229 => x"08ff068c",
11230 => x"08fc050c",
11231 => x"8c088805",
11232 => x"08700894",
11233 => x"2a545451",
11234 => x"80728fff",
11235 => x"068c08f4",
11236 => x"050c8c08",
11237 => x"88050870",
11238 => x"089f2a54",
11239 => x"54518072",
11240 => x"81068c08",
11241 => x"f0050c8c",
11242 => x"088c0508",
11243 => x"8c08f005",
11244 => x"0884120c",
11245 => x"51518c08",
11246 => x"f405080b",
11247 => x"0b0b81cf",
11248 => x"388c08f8",
11249 => x"0508708c",
11250 => x"08fc0508",
11251 => x"07515170",
11252 => x"0b0b0b0b",
11253 => x"90388c08",
11254 => x"8c050851",
11255 => x"82710c0b",
11256 => x"0b0b82f8",
11257 => x"398c088c",
11258 => x"05088c08",
11259 => x"f40508f8",
11260 => x"82058812",
11261 => x"0c8c08fc",
11262 => x"0508982a",
11263 => x"8c08f805",
11264 => x"08882b70",
11265 => x"72078c08",
11266 => x"fc050888",
11267 => x"2b565355",
11268 => x"5551708c",
11269 => x"08f8050c",
11270 => x"718c08fc",
11271 => x"050c8c08",
11272 => x"8c050851",
11273 => x"83710c8c",
11274 => x"08f80508",
11275 => x"f00a260b",
11276 => x"0b0b0bbb",
11277 => x"388c08fc",
11278 => x"05089f2a",
11279 => x"8c08f805",
11280 => x"08107072",
11281 => x"078c08fc",
11282 => x"05081055",
11283 => x"53545470",
11284 => x"8c08f805",
11285 => x"0c718c08",
11286 => x"fc050c8c",
11287 => x"088c0508",
11288 => x"881108ff",
11289 => x"0588120c",
11290 => x"510b0b0b",
11291 => x"ffb9398c",
11292 => x"088c0508",
11293 => x"538c08f8",
11294 => x"05088c08",
11295 => x"fc050853",
11296 => x"51708c14",
11297 => x"0c719014",
11298 => x"0c0b0b0b",
11299 => x"81ce398c",
11300 => x"08f40508",
11301 => x"8fff2e09",
11302 => x"81060b0b",
11303 => x"0b80f438",
11304 => x"8c08f805",
11305 => x"08708c08",
11306 => x"fc050807",
11307 => x"5151700b",
11308 => x"0b0b0b90",
11309 => x"388c088c",
11310 => x"05085184",
11311 => x"710c0b0b",
11312 => x"0b819939",
11313 => x"8c08f805",
11314 => x"08932a52",
11315 => x"80728106",
11316 => x"51517080",
11317 => x"2e0b0b0b",
11318 => x"0b90388c",
11319 => x"088c0508",
11320 => x"5181710c",
11321 => x"0b0b0b0b",
11322 => x"8a398c08",
11323 => x"8c050851",
11324 => x"80710c8c",
11325 => x"088c0508",
11326 => x"538c08f8",
11327 => x"05088c08",
11328 => x"fc050853",
11329 => x"51708c14",
11330 => x"0c719014",
11331 => x"0c0b0b0b",
11332 => x"80ca398c",
11333 => x"088c0508",
11334 => x"8c08f405",
11335 => x"08f88105",
11336 => x"88120c8c",
11337 => x"088c0508",
11338 => x"51518371",
11339 => x"0c8c088c",
11340 => x"05088c08",
11341 => x"fc050898",
11342 => x"2a8c08f8",
11343 => x"0508882b",
11344 => x"7072078c",
11345 => x"08fc0508",
11346 => x"882b7188",
11347 => x"0a078c16",
11348 => x"0c708007",
11349 => x"90160c56",
11350 => x"54555555",
11351 => x"8a3d0d8c",
11352 => x"0c048c08",
11353 => x"028c0cf0",
11354 => x"3d0d8c08",
11355 => x"88050851",
11356 => x"0b0b0b89",
11357 => x"993f8008",
11358 => x"52710b0b",
11359 => x"0b0b9d38",
11360 => x"8c088c05",
11361 => x"08510b0b",
11362 => x"0b89833f",
11363 => x"80085271",
11364 => x"0b0b0b0b",
11365 => x"87380b0b",
11366 => x"0b0b8e39",
11367 => x"810b8c08",
11368 => x"fc050c0b",
11369 => x"0b0b87ed",
11370 => x"398c0888",
11371 => x"0508510b",
11372 => x"0b0b88a4",
11373 => x"3f800852",
11374 => x"71802e0b",
11375 => x"0b0b0bb9",
11376 => x"388c088c",
11377 => x"0508510b",
11378 => x"0b0b888c",
11379 => x"3f800852",
11380 => x"71802e0b",
11381 => x"0b0b0ba1",
11382 => x"388c088c",
11383 => x"05088c08",
11384 => x"88050884",
11385 => x"12088412",
11386 => x"0831708c",
11387 => x"08fc050c",
11388 => x"5254520b",
11389 => x"0b0b879d",
11390 => x"398c0888",
11391 => x"0508510b",
11392 => x"0b0b87d4",
11393 => x"3f800852",
11394 => x"71802e0b",
11395 => x"0b0b0bb6",
11396 => x"388c0888",
11397 => x"05085284",
11398 => x"1208802e",
11399 => x"0b0b0b0b",
11400 => x"8e38ff0b",
11401 => x"8c08f805",
11402 => x"0c0b0b0b",
11403 => x"0b883981",
11404 => x"0b8c08f8",
11405 => x"050c8c08",
11406 => x"f805088c",
11407 => x"08fc050c",
11408 => x"0b0b0b86",
11409 => x"d0398c08",
11410 => x"8c050851",
11411 => x"0b0b0b87",
11412 => x"873f8008",
11413 => x"5271802e",
11414 => x"0b0b0b0b",
11415 => x"b6388c08",
11416 => x"8c050852",
11417 => x"84120880",
11418 => x"2e0b0b0b",
11419 => x"0b8e3881",
11420 => x"0b8c08f4",
11421 => x"050c0b0b",
11422 => x"0b0b8839",
11423 => x"ff0b8c08",
11424 => x"f4050c8c",
11425 => x"08f40508",
11426 => x"8c08fc05",
11427 => x"0c0b0b0b",
11428 => x"8683398c",
11429 => x"08880508",
11430 => x"510b0b0b",
11431 => x"86843f80",
11432 => x"08527180",
11433 => x"2e0b0b0b",
11434 => x"0ba6388c",
11435 => x"088c0508",
11436 => x"510b0b0b",
11437 => x"85ec3f80",
11438 => x"08527180",
11439 => x"2e0b0b0b",
11440 => x"0b8e3880",
11441 => x"0b8c08fc",
11442 => x"050c0b0b",
11443 => x"0b85c639",
11444 => x"8c088805",
11445 => x"08510b0b",
11446 => x"0b85c73f",
11447 => x"80085271",
11448 => x"802e0b0b",
11449 => x"0b0bb638",
11450 => x"8c088c05",
11451 => x"08528412",
11452 => x"08802e0b",
11453 => x"0b0b0b8e",
11454 => x"38810b8c",
11455 => x"08f0050c",
11456 => x"0b0b0b0b",
11457 => x"8839ff0b",
11458 => x"8c08f005",
11459 => x"0c8c08f0",
11460 => x"05088c08",
11461 => x"fc050c0b",
11462 => x"0b0b84f9",
11463 => x"398c088c",
11464 => x"0508510b",
11465 => x"0b0b84fa",
11466 => x"3f800852",
11467 => x"71802e0b",
11468 => x"0b0b0bb6",
11469 => x"388c0888",
11470 => x"05085284",
11471 => x"1208802e",
11472 => x"0b0b0b0b",
11473 => x"8e38ff0b",
11474 => x"8c08ec05",
11475 => x"0c0b0b0b",
11476 => x"0b883981",
11477 => x"0b8c08ec",
11478 => x"050c8c08",
11479 => x"ec05088c",
11480 => x"08fc050c",
11481 => x"0b0b0b84",
11482 => x"ac398c08",
11483 => x"8805088c",
11484 => x"088c0508",
11485 => x"53538413",
11486 => x"08841308",
11487 => x"2e0b0b0b",
11488 => x"0bb6388c",
11489 => x"08880508",
11490 => x"52841208",
11491 => x"802e0b0b",
11492 => x"0b0b8e38",
11493 => x"ff0b8c08",
11494 => x"e8050c0b",
11495 => x"0b0b0b88",
11496 => x"39810b8c",
11497 => x"08e8050c",
11498 => x"8c08e805",
11499 => x"088c08fc",
11500 => x"050c0b0b",
11501 => x"0b83de39",
11502 => x"8c088805",
11503 => x"088c088c",
11504 => x"05085353",
11505 => x"88120888",
11506 => x"1408250b",
11507 => x"0b0b0bb6",
11508 => x"388c0888",
11509 => x"05085284",
11510 => x"1208802e",
11511 => x"0b0b0b0b",
11512 => x"8e38ff0b",
11513 => x"8c08e405",
11514 => x"0c0b0b0b",
11515 => x"0b883981",
11516 => x"0b8c08e4",
11517 => x"050c8c08",
11518 => x"e405088c",
11519 => x"08fc050c",
11520 => x"0b0b0b83",
11521 => x"90398c08",
11522 => x"8805088c",
11523 => x"088c0508",
11524 => x"53538813",
11525 => x"08881308",
11526 => x"250b0b0b",
11527 => x"0bb6388c",
11528 => x"08880508",
11529 => x"52841208",
11530 => x"802e0b0b",
11531 => x"0b0b8e38",
11532 => x"810b8c08",
11533 => x"e0050c0b",
11534 => x"0b0b0b88",
11535 => x"39ff0b8c",
11536 => x"08e0050c",
11537 => x"8c08e005",
11538 => x"088c08fc",
11539 => x"050c0b0b",
11540 => x"0b82c239",
11541 => x"8c088805",
11542 => x"088c08dc",
11543 => x"050c8c08",
11544 => x"8c05088c",
11545 => x"08d8050c",
11546 => x"8c08dc05",
11547 => x"088c08d8",
11548 => x"05085452",
11549 => x"8c12088c",
11550 => x"1408260b",
11551 => x"0b0b0bbc",
11552 => x"388c08dc",
11553 => x"05088c08",
11554 => x"d8050854",
11555 => x"528c1208",
11556 => x"8c14082e",
11557 => x"0981060b",
11558 => x"0b0b80d5",
11559 => x"388c08dc",
11560 => x"05088c08",
11561 => x"d8050854",
11562 => x"52901208",
11563 => x"90140826",
11564 => x"0b0b0b0b",
11565 => x"87380b0b",
11566 => x"0b0bb639",
11567 => x"8c088805",
11568 => x"08528412",
11569 => x"08802e0b",
11570 => x"0b0b0b8e",
11571 => x"38ff0b8c",
11572 => x"08d4050c",
11573 => x"0b0b0b0b",
11574 => x"8839810b",
11575 => x"8c08d405",
11576 => x"0c8c08d4",
11577 => x"05088c08",
11578 => x"fc050c0b",
11579 => x"0b0b81a5",
11580 => x"398c088c",
11581 => x"05088c08",
11582 => x"d0050c8c",
11583 => x"08880508",
11584 => x"8c08cc05",
11585 => x"0c8c08d0",
11586 => x"05088c08",
11587 => x"cc050854",
11588 => x"528c1208",
11589 => x"8c140826",
11590 => x"0b0b0b0b",
11591 => x"bc388c08",
11592 => x"d005088c",
11593 => x"08cc0508",
11594 => x"54528c12",
11595 => x"088c1408",
11596 => x"2e098106",
11597 => x"0b0b0b80",
11598 => x"d5388c08",
11599 => x"d005088c",
11600 => x"08cc0508",
11601 => x"54529012",
11602 => x"08901408",
11603 => x"260b0b0b",
11604 => x"0b87380b",
11605 => x"0b0b0bb6",
11606 => x"398c0888",
11607 => x"05085284",
11608 => x"1208802e",
11609 => x"0b0b0b0b",
11610 => x"8e38810b",
11611 => x"8c08c805",
11612 => x"0c0b0b0b",
11613 => x"0b8839ff",
11614 => x"0b8c08c8",
11615 => x"050c8c08",
11616 => x"c805088c",
11617 => x"08fc050c",
11618 => x"0b0b0b0b",
11619 => x"8839800b",
11620 => x"8c08fc05",
11621 => x"0c8c08fc",
11622 => x"0508800c",
11623 => x"923d0d8c",
11624 => x"0c048c08",
11625 => x"028c0c70",
11626 => x"70800b8c",
11627 => x"08fc050c",
11628 => x"8c088805",
11629 => x"08517008",
11630 => x"822e0981",
11631 => x"060b0b0b",
11632 => x"0b883881",
11633 => x"0b8c08fc",
11634 => x"050c8c08",
11635 => x"fc050870",
11636 => x"800c5150",
11637 => x"508c0c04",
11638 => x"8c08028c",
11639 => x"0c707080",
11640 => x"0b8c08fc",
11641 => x"050c8c08",
11642 => x"88050851",
11643 => x"7008842e",
11644 => x"0981060b",
11645 => x"0b0b0b88",
11646 => x"38810b8c",
11647 => x"08fc050c",
11648 => x"8c08fc05",
11649 => x"0870800c",
11650 => x"5150508c",
11651 => x"0c048c08",
11652 => x"028c0c70",
11653 => x"70800b8c",
11654 => x"08fc050c",
11655 => x"8c088805",
11656 => x"08517008",
11657 => x"802e0b0b",
11658 => x"0b0b9738",
11659 => x"8c088805",
11660 => x"08517008",
11661 => x"812e0b0b",
11662 => x"0b0b8738",
11663 => x"0b0b0b0b",
11664 => x"8839810b",
11665 => x"8c08fc05",
11666 => x"0c8c08fc",
11667 => x"05087080",
11668 => x"0c515050",
11669 => x"8c0c0470",
11670 => x"700b0b83",
11671 => x"84d80bfc",
11672 => x"05700852",
11673 => x"5270ff2e",
11674 => x"0b0b0b0b",
11675 => x"9538702d",
11676 => x"fc127008",
11677 => x"525270ff",
11678 => x"2e098106",
11679 => x"0b0b0b0b",
11680 => x"ed385050",
11681 => x"04040b0b",
11682 => x"fd9e993f",
11683 => x"04000000",
11684 => x"00000040",
11685 => x"48656c6c",
11686 => x"6f20776f",
11687 => x"726c6421",
11688 => x"0a000000",
11689 => x"20202020",
11690 => x"20202020",
11691 => x"20202020",
11692 => x"20202020",
11693 => x"30303030",
11694 => x"30303030",
11695 => x"30303030",
11696 => x"30303030",
11697 => x"0000164c",
11698 => x"000010d6",
11699 => x"000010d6",
11700 => x"0000163f",
11701 => x"000010d6",
11702 => x"000010d6",
11703 => x"000010d6",
11704 => x"000010d6",
11705 => x"000010d6",
11706 => x"000010d6",
11707 => x"000010a4",
11708 => x"000015c6",
11709 => x"000010d6",
11710 => x"000010b9",
11711 => x"000012d9",
11712 => x"000010d6",
11713 => x"000015fe",
11714 => x"000015d5",
11715 => x"000015d5",
11716 => x"000015d5",
11717 => x"000015d5",
11718 => x"000015d5",
11719 => x"000015d5",
11720 => x"000015d5",
11721 => x"000015d5",
11722 => x"000015d5",
11723 => x"000010d6",
11724 => x"000010d6",
11725 => x"000010d6",
11726 => x"000010d6",
11727 => x"000010d6",
11728 => x"000010d6",
11729 => x"000010d6",
11730 => x"000010d6",
11731 => x"000010d6",
11732 => x"00001476",
11733 => x"00001060",
11734 => x"000013e5",
11735 => x"000010d6",
11736 => x"000013e5",
11737 => x"000010d6",
11738 => x"000010d6",
11739 => x"000010d6",
11740 => x"000010d6",
11741 => x"0000160c",
11742 => x"000010d6",
11743 => x"000010d6",
11744 => x"00001024",
11745 => x"000010d6",
11746 => x"000010d6",
11747 => x"000010d6",
11748 => x"0000152a",
11749 => x"000010d6",
11750 => x"00000ce0",
11751 => x"000010d6",
11752 => x"000010d6",
11753 => x"000014d2",
11754 => x"000010d6",
11755 => x"000010d6",
11756 => x"000010d6",
11757 => x"000010d6",
11758 => x"000010d6",
11759 => x"000010d6",
11760 => x"000010d6",
11761 => x"000010d6",
11762 => x"000010d6",
11763 => x"000010d6",
11764 => x"00001476",
11765 => x"00001064",
11766 => x"000013e5",
11767 => x"000013e5",
11768 => x"000013e5",
11769 => x"000013d7",
11770 => x"00001064",
11771 => x"000010d6",
11772 => x"000010d6",
11773 => x"000012b5",
11774 => x"000010d6",
11775 => x"00001592",
11776 => x"00001028",
11777 => x"0000132c",
11778 => x"000010c9",
11779 => x"000010d6",
11780 => x"0000152a",
11781 => x"000010d6",
11782 => x"00000ce4",
11783 => x"000010d6",
11784 => x"000010d6",
11785 => x"00001619",
11786 => x"62756720",
11787 => x"696e2076",
11788 => x"66707269",
11789 => x"6e74663a",
11790 => x"20626164",
11791 => x"20626173",
11792 => x"65000000",
11793 => x"30313233",
11794 => x"34353637",
11795 => x"38396162",
11796 => x"63646566",
11797 => x"00000000",
11798 => x"496e6600",
11799 => x"30313233",
11800 => x"34353637",
11801 => x"38394142",
11802 => x"43444546",
11803 => x"00000000",
11804 => x"30000000",
11805 => x"2e000000",
11806 => x"4e614e00",
11807 => x"286e756c",
11808 => x"6c290000",
11809 => x"432d5554",
11810 => x"462d3800",
11811 => x"432d534a",
11812 => x"49530000",
11813 => x"432d4555",
11814 => x"434a5000",
11815 => x"432d4a49",
11816 => x"53000000",
11817 => x"496e6669",
11818 => x"6e697479",
11819 => x"00000000",
11820 => x"000037a9",
11821 => x"000037a9",
11822 => x"0000378d",
11823 => x"000031e6",
11824 => x"00003792",
11825 => x"000031eb",
11826 => x"43000000",
11827 => x"49534f2d",
11828 => x"38383539",
11829 => x"2d310000",
11830 => x"0000b874",
11831 => x"0000b86c",
11832 => x"0000b86c",
11833 => x"0000b86c",
11834 => x"0000b86c",
11835 => x"0000b86c",
11836 => x"0000b86c",
11837 => x"0000b86c",
11838 => x"0000b86c",
11839 => x"0000b86c",
11840 => x"ffffffff",
11841 => x"ffffffff",
11842 => x"3c9cd2b2",
11843 => x"97d889bc",
11844 => x"3949f623",
11845 => x"d5a8a733",
11846 => x"32a50ffd",
11847 => x"44f4a73d",
11848 => x"255bba08",
11849 => x"cf8c979d",
11850 => x"0ac80628",
11851 => x"64ac6f43",
11852 => x"4341c379",
11853 => x"37e08000",
11854 => x"4693b8b5",
11855 => x"b5056e17",
11856 => x"4d384f03",
11857 => x"e93ff9f5",
11858 => x"5a827748",
11859 => x"f9301d32",
11860 => x"75154fdd",
11861 => x"7f73bf3c",
11862 => x"3ff00000",
11863 => x"00000000",
11864 => x"40240000",
11865 => x"00000000",
11866 => x"40590000",
11867 => x"00000000",
11868 => x"408f4000",
11869 => x"00000000",
11870 => x"40c38800",
11871 => x"00000000",
11872 => x"40f86a00",
11873 => x"00000000",
11874 => x"412e8480",
11875 => x"00000000",
11876 => x"416312d0",
11877 => x"00000000",
11878 => x"4197d784",
11879 => x"00000000",
11880 => x"41cdcd65",
11881 => x"00000000",
11882 => x"4202a05f",
11883 => x"20000000",
11884 => x"42374876",
11885 => x"e8000000",
11886 => x"426d1a94",
11887 => x"a2000000",
11888 => x"42a2309c",
11889 => x"e5400000",
11890 => x"42d6bcc4",
11891 => x"1e900000",
11892 => x"430c6bf5",
11893 => x"26340000",
11894 => x"4341c379",
11895 => x"37e08000",
11896 => x"43763457",
11897 => x"85d8a000",
11898 => x"43abc16d",
11899 => x"674ec800",
11900 => x"43e158e4",
11901 => x"60913d00",
11902 => x"4415af1d",
11903 => x"78b58c40",
11904 => x"444b1ae4",
11905 => x"d6e2ef50",
11906 => x"4480f0cf",
11907 => x"064dd592",
11908 => x"44b52d02",
11909 => x"c7e14af6",
11910 => x"44ea7843",
11911 => x"79d99db4",
11912 => x"00000005",
11913 => x"00000019",
11914 => x"0000007d",
11915 => x"64756d6d",
11916 => x"792e6578",
11917 => x"65000000",
11918 => x"00000000",
11919 => x"00000000",
11920 => x"00000000",
11921 => x"00000000",
11922 => x"00000000",
11923 => x"00ffffff",
11924 => x"ff00ffff",
11925 => x"ffff00ff",
11926 => x"ffffff00",
11927 => x"00000000",
11928 => x"00000000",
11929 => x"00000000",
11930 => x"0000c260",
11931 => x"0000ba70",
11932 => x"00000000",
11933 => x"0000bcd8",
11934 => x"0000bd34",
11935 => x"0000bd90",
11936 => x"00000000",
11937 => x"00000000",
11938 => x"00000000",
11939 => x"00000000",
11940 => x"00000000",
11941 => x"00000000",
11942 => x"00000000",
11943 => x"00000000",
11944 => x"00000000",
11945 => x"0000b8c8",
11946 => x"00000000",
11947 => x"00000000",
11948 => x"00000000",
11949 => x"00000000",
11950 => x"00000000",
11951 => x"00000000",
11952 => x"00000000",
11953 => x"00000000",
11954 => x"00000000",
11955 => x"00000000",
11956 => x"00000000",
11957 => x"00000000",
11958 => x"00000000",
11959 => x"00000000",
11960 => x"00000000",
11961 => x"00000000",
11962 => x"00000000",
11963 => x"00000000",
11964 => x"00000000",
11965 => x"00000000",
11966 => x"00000000",
11967 => x"00000000",
11968 => x"00000000",
11969 => x"00000000",
11970 => x"00000000",
11971 => x"00000000",
11972 => x"00000000",
11973 => x"00000000",
11974 => x"00000001",
11975 => x"330eabcd",
11976 => x"1234e66d",
11977 => x"deec0005",
11978 => x"000b0000",
11979 => x"00000000",
11980 => x"00000000",
11981 => x"00000000",
11982 => x"00000000",
11983 => x"00000000",
11984 => x"00000000",
11985 => x"00000000",
11986 => x"00000000",
11987 => x"00000000",
11988 => x"00000000",
11989 => x"00000000",
11990 => x"00000000",
11991 => x"00000000",
11992 => x"00000000",
11993 => x"00000000",
11994 => x"00000000",
11995 => x"00000000",
11996 => x"00000000",
11997 => x"00000000",
11998 => x"00000000",
11999 => x"00000000",
12000 => x"00000000",
12001 => x"00000000",
12002 => x"00000000",
12003 => x"00000000",
12004 => x"00000000",
12005 => x"00000000",
12006 => x"00000000",
12007 => x"00000000",
12008 => x"00000000",
12009 => x"00000000",
12010 => x"00000000",
12011 => x"00000000",
12012 => x"00000000",
12013 => x"00000000",
12014 => x"00000000",
12015 => x"00000000",
12016 => x"00000000",
12017 => x"00000000",
12018 => x"00000000",
12019 => x"00000000",
12020 => x"00000000",
12021 => x"00000000",
12022 => x"00000000",
12023 => x"00000000",
12024 => x"00000000",
12025 => x"00000000",
12026 => x"00000000",
12027 => x"00000000",
12028 => x"00000000",
12029 => x"00000000",
12030 => x"00000000",
12031 => x"00000000",
12032 => x"00000000",
12033 => x"00000000",
12034 => x"00000000",
12035 => x"00000000",
12036 => x"00000000",
12037 => x"00000000",
12038 => x"00000000",
12039 => x"00000000",
12040 => x"00000000",
12041 => x"00000000",
12042 => x"00000000",
12043 => x"00000000",
12044 => x"00000000",
12045 => x"00000000",
12046 => x"00000000",
12047 => x"00000000",
12048 => x"00000000",
12049 => x"00000000",
12050 => x"00000000",
12051 => x"00000000",
12052 => x"00000000",
12053 => x"00000000",
12054 => x"00000000",
12055 => x"00000000",
12056 => x"00000000",
12057 => x"00000000",
12058 => x"00000000",
12059 => x"00000000",
12060 => x"00000000",
12061 => x"00000000",
12062 => x"00000000",
12063 => x"00000000",
12064 => x"00000000",
12065 => x"00000000",
12066 => x"00000000",
12067 => x"00000000",
12068 => x"00000000",
12069 => x"00000000",
12070 => x"00000000",
12071 => x"00000000",
12072 => x"00000000",
12073 => x"00000000",
12074 => x"00000000",
12075 => x"00000000",
12076 => x"00000000",
12077 => x"00000000",
12078 => x"00000000",
12079 => x"00000000",
12080 => x"00000000",
12081 => x"00000000",
12082 => x"00000000",
12083 => x"00000000",
12084 => x"00000000",
12085 => x"00000000",
12086 => x"00000000",
12087 => x"00000000",
12088 => x"00000000",
12089 => x"00000000",
12090 => x"00000000",
12091 => x"00000000",
12092 => x"00000000",
12093 => x"00000000",
12094 => x"00000000",
12095 => x"00000000",
12096 => x"00000000",
12097 => x"00000000",
12098 => x"00000000",
12099 => x"00000000",
12100 => x"00000000",
12101 => x"00000000",
12102 => x"00000000",
12103 => x"00000000",
12104 => x"00000000",
12105 => x"00000000",
12106 => x"00000000",
12107 => x"00000000",
12108 => x"00000000",
12109 => x"00000000",
12110 => x"00000000",
12111 => x"00000000",
12112 => x"00000000",
12113 => x"00000000",
12114 => x"00000000",
12115 => x"00000000",
12116 => x"00000000",
12117 => x"00000000",
12118 => x"00000000",
12119 => x"00000000",
12120 => x"00000000",
12121 => x"00000000",
12122 => x"00000000",
12123 => x"00000000",
12124 => x"00000000",
12125 => x"00000000",
12126 => x"00000000",
12127 => x"00000000",
12128 => x"00000000",
12129 => x"00000000",
12130 => x"00000000",
12131 => x"00000000",
12132 => x"00000000",
12133 => x"00000000",
12134 => x"00000000",
12135 => x"00000000",
12136 => x"00000000",
12137 => x"00000000",
12138 => x"00000000",
12139 => x"00000000",
12140 => x"00000000",
12141 => x"00000000",
12142 => x"00000000",
12143 => x"00000000",
12144 => x"00000000",
12145 => x"00000000",
12146 => x"00000000",
12147 => x"00000000",
12148 => x"00000000",
12149 => x"00000000",
12150 => x"00000000",
12151 => x"00000000",
12152 => x"00000000",
12153 => x"00000000",
12154 => x"00000000",
12155 => x"43000000",
12156 => x"00000000",
12157 => x"00000000",
12158 => x"00000000",
12159 => x"00000000",
12160 => x"00000000",
12161 => x"00000001",
12162 => x"0000b8cc",
12163 => x"00000000",
12164 => x"00000000",
12165 => x"00000000",
12166 => x"00000000",
12167 => x"00000000",
12168 => x"00000000",
12169 => x"00000000",
12170 => x"00000000",
12171 => x"00000000",
12172 => x"00000000",
12173 => x"00000000",
12174 => x"00000000",
12175 => x"ffffffff",
12176 => x"00000000",
12177 => x"00020000",
12178 => x"00000000",
12179 => x"00000000",
12180 => x"0000be48",
12181 => x"0000be48",
12182 => x"0000be50",
12183 => x"0000be50",
12184 => x"0000be58",
12185 => x"0000be58",
12186 => x"0000be60",
12187 => x"0000be60",
12188 => x"0000be68",
12189 => x"0000be68",
12190 => x"0000be70",
12191 => x"0000be70",
12192 => x"0000be78",
12193 => x"0000be78",
12194 => x"0000be80",
12195 => x"0000be80",
12196 => x"0000be88",
12197 => x"0000be88",
12198 => x"0000be90",
12199 => x"0000be90",
12200 => x"0000be98",
12201 => x"0000be98",
12202 => x"0000bea0",
12203 => x"0000bea0",
12204 => x"0000bea8",
12205 => x"0000bea8",
12206 => x"0000beb0",
12207 => x"0000beb0",
12208 => x"0000beb8",
12209 => x"0000beb8",
12210 => x"0000bec0",
12211 => x"0000bec0",
12212 => x"0000bec8",
12213 => x"0000bec8",
12214 => x"0000bed0",
12215 => x"0000bed0",
12216 => x"0000bed8",
12217 => x"0000bed8",
12218 => x"0000bee0",
12219 => x"0000bee0",
12220 => x"0000bee8",
12221 => x"0000bee8",
12222 => x"0000bef0",
12223 => x"0000bef0",
12224 => x"0000bef8",
12225 => x"0000bef8",
12226 => x"0000bf00",
12227 => x"0000bf00",
12228 => x"0000bf08",
12229 => x"0000bf08",
12230 => x"0000bf10",
12231 => x"0000bf10",
12232 => x"0000bf18",
12233 => x"0000bf18",
12234 => x"0000bf20",
12235 => x"0000bf20",
12236 => x"0000bf28",
12237 => x"0000bf28",
12238 => x"0000bf30",
12239 => x"0000bf30",
12240 => x"0000bf38",
12241 => x"0000bf38",
12242 => x"0000bf40",
12243 => x"0000bf40",
12244 => x"0000bf48",
12245 => x"0000bf48",
12246 => x"0000bf50",
12247 => x"0000bf50",
12248 => x"0000bf58",
12249 => x"0000bf58",
12250 => x"0000bf60",
12251 => x"0000bf60",
12252 => x"0000bf68",
12253 => x"0000bf68",
12254 => x"0000bf70",
12255 => x"0000bf70",
12256 => x"0000bf78",
12257 => x"0000bf78",
12258 => x"0000bf80",
12259 => x"0000bf80",
12260 => x"0000bf88",
12261 => x"0000bf88",
12262 => x"0000bf90",
12263 => x"0000bf90",
12264 => x"0000bf98",
12265 => x"0000bf98",
12266 => x"0000bfa0",
12267 => x"0000bfa0",
12268 => x"0000bfa8",
12269 => x"0000bfa8",
12270 => x"0000bfb0",
12271 => x"0000bfb0",
12272 => x"0000bfb8",
12273 => x"0000bfb8",
12274 => x"0000bfc0",
12275 => x"0000bfc0",
12276 => x"0000bfc8",
12277 => x"0000bfc8",
12278 => x"0000bfd0",
12279 => x"0000bfd0",
12280 => x"0000bfd8",
12281 => x"0000bfd8",
12282 => x"0000bfe0",
12283 => x"0000bfe0",
12284 => x"0000bfe8",
12285 => x"0000bfe8",
12286 => x"0000bff0",
12287 => x"0000bff0",
12288 => x"0000bff8",
12289 => x"0000bff8",
12290 => x"0000c000",
12291 => x"0000c000",
12292 => x"0000c008",
12293 => x"0000c008",
12294 => x"0000c010",
12295 => x"0000c010",
12296 => x"0000c018",
12297 => x"0000c018",
12298 => x"0000c020",
12299 => x"0000c020",
12300 => x"0000c028",
12301 => x"0000c028",
12302 => x"0000c030",
12303 => x"0000c030",
12304 => x"0000c038",
12305 => x"0000c038",
12306 => x"0000c040",
12307 => x"0000c040",
12308 => x"0000c048",
12309 => x"0000c048",
12310 => x"0000c050",
12311 => x"0000c050",
12312 => x"0000c058",
12313 => x"0000c058",
12314 => x"0000c060",
12315 => x"0000c060",
12316 => x"0000c068",
12317 => x"0000c068",
12318 => x"0000c070",
12319 => x"0000c070",
12320 => x"0000c078",
12321 => x"0000c078",
12322 => x"0000c080",
12323 => x"0000c080",
12324 => x"0000c088",
12325 => x"0000c088",
12326 => x"0000c090",
12327 => x"0000c090",
12328 => x"0000c098",
12329 => x"0000c098",
12330 => x"0000c0a0",
12331 => x"0000c0a0",
12332 => x"0000c0a8",
12333 => x"0000c0a8",
12334 => x"0000c0b0",
12335 => x"0000c0b0",
12336 => x"0000c0b8",
12337 => x"0000c0b8",
12338 => x"0000c0c0",
12339 => x"0000c0c0",
12340 => x"0000c0c8",
12341 => x"0000c0c8",
12342 => x"0000c0d0",
12343 => x"0000c0d0",
12344 => x"0000c0d8",
12345 => x"0000c0d8",
12346 => x"0000c0e0",
12347 => x"0000c0e0",
12348 => x"0000c0e8",
12349 => x"0000c0e8",
12350 => x"0000c0f0",
12351 => x"0000c0f0",
12352 => x"0000c0f8",
12353 => x"0000c0f8",
12354 => x"0000c100",
12355 => x"0000c100",
12356 => x"0000c108",
12357 => x"0000c108",
12358 => x"0000c110",
12359 => x"0000c110",
12360 => x"0000c118",
12361 => x"0000c118",
12362 => x"0000c120",
12363 => x"0000c120",
12364 => x"0000c128",
12365 => x"0000c128",
12366 => x"0000c130",
12367 => x"0000c130",
12368 => x"0000c138",
12369 => x"0000c138",
12370 => x"0000c140",
12371 => x"0000c140",
12372 => x"0000c148",
12373 => x"0000c148",
12374 => x"0000c150",
12375 => x"0000c150",
12376 => x"0000c158",
12377 => x"0000c158",
12378 => x"0000c160",
12379 => x"0000c160",
12380 => x"0000c168",
12381 => x"0000c168",
12382 => x"0000c170",
12383 => x"0000c170",
12384 => x"0000c178",
12385 => x"0000c178",
12386 => x"0000c180",
12387 => x"0000c180",
12388 => x"0000c188",
12389 => x"0000c188",
12390 => x"0000c190",
12391 => x"0000c190",
12392 => x"0000c198",
12393 => x"0000c198",
12394 => x"0000c1a0",
12395 => x"0000c1a0",
12396 => x"0000c1a8",
12397 => x"0000c1a8",
12398 => x"0000c1b0",
12399 => x"0000c1b0",
12400 => x"0000c1b8",
12401 => x"0000c1b8",
12402 => x"0000c1c0",
12403 => x"0000c1c0",
12404 => x"0000c1c8",
12405 => x"0000c1c8",
12406 => x"0000c1d0",
12407 => x"0000c1d0",
12408 => x"0000c1d8",
12409 => x"0000c1d8",
12410 => x"0000c1e0",
12411 => x"0000c1e0",
12412 => x"0000c1e8",
12413 => x"0000c1e8",
12414 => x"0000c1f0",
12415 => x"0000c1f0",
12416 => x"0000c1f8",
12417 => x"0000c1f8",
12418 => x"0000c200",
12419 => x"0000c200",
12420 => x"0000c208",
12421 => x"0000c208",
12422 => x"0000c210",
12423 => x"0000c210",
12424 => x"0000c218",
12425 => x"0000c218",
12426 => x"0000c220",
12427 => x"0000c220",
12428 => x"0000c228",
12429 => x"0000c228",
12430 => x"0000c230",
12431 => x"0000c230",
12432 => x"0000c238",
12433 => x"0000c238",
12434 => x"0000c240",
12435 => x"0000c240",
12436 => x"0000ba2c",
12437 => x"ffffffff",
12438 => x"00000000",
12439 => x"ffffffff",
12440 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(conv_integer(memAAddr)) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(conv_integer(memAAddr));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(conv_integer(memBAddr)) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(conv_integer(memBAddr));
		end if;
	end if;
end process;




end dualport_ram_arch;
