-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b80ea",
     1 => x"ec040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b80ed",
     9 => x"d3040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b80ed",
    73 => x"85040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b80ece8",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b81bf",
   162 => x"c0738306",
   163 => x"10100508",
   164 => x"060b0b80",
   165 => x"eceb0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b80ed",
   169 => x"ba040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b80ed",
   177 => x"a1040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"81bfd00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053370",
   258 => x"525280ea",
   259 => x"ae3f7151",
   260 => x"80eaf83f",
   261 => x"71b00c83",
   262 => x"3d0d04ff",
   263 => x"3d0d81bf",
   264 => x"ac08b811",
   265 => x"08535180",
   266 => x"0bb8120c",
   267 => x"71b00c83",
   268 => x"3d0d0480",
   269 => x"0b81e2e0",
   270 => x"34800bb0",
   271 => x"0c04fb3d",
   272 => x"0d815180",
   273 => x"c6ef3fb0",
   274 => x"08538251",
   275 => x"80c6e63f",
   276 => x"b00856b0",
   277 => x"08833890",
   278 => x"5672fc06",
   279 => x"5575812e",
   280 => x"80fb3880",
   281 => x"54737627",
   282 => x"ad387383",
   283 => x"06537280",
   284 => x"2eb23881",
   285 => x"9cb45180",
   286 => x"e59a3f74",
   287 => x"70840556",
   288 => x"0852a051",
   289 => x"80e5b03f",
   290 => x"a05180e4",
   291 => x"ed3f8114",
   292 => x"54757426",
   293 => x"d5388a51",
   294 => x"80e4df3f",
   295 => x"800bb00c",
   296 => x"873d0d04",
   297 => x"819cb851",
   298 => x"80e4e93f",
   299 => x"7452a051",
   300 => x"80e5843f",
   301 => x"81a9a451",
   302 => x"80e4d93f",
   303 => x"819cb451",
   304 => x"80e4d13f",
   305 => x"74708405",
   306 => x"560852a0",
   307 => x"5180e4e7",
   308 => x"3fa05180",
   309 => x"e4a43f81",
   310 => x"1454ffb5",
   311 => x"39819cb4",
   312 => x"5180e4b0",
   313 => x"3f740852",
   314 => x"a05180e4",
   315 => x"ca3f8a51",
   316 => x"80e4873f",
   317 => x"800bb00c",
   318 => x"873d0d04",
   319 => x"fc3d0d81",
   320 => x"5180c5b1",
   321 => x"3fb00852",
   322 => x"825180c3",
   323 => x"f63fb008",
   324 => x"81ff0672",
   325 => x"56538354",
   326 => x"72802ea2",
   327 => x"38735180",
   328 => x"c5933f81",
   329 => x"147081ff",
   330 => x"06ff1570",
   331 => x"81ff06b0",
   332 => x"08797084",
   333 => x"055b0c56",
   334 => x"52555272",
   335 => x"e03872b0",
   336 => x"0c863d0d",
   337 => x"04803d0d",
   338 => x"8c5180e3",
   339 => x"ad3f800b",
   340 => x"b00c823d",
   341 => x"0d04fb3d",
   342 => x"0d800b81",
   343 => x"9cbc5256",
   344 => x"80e3b13f",
   345 => x"75557410",
   346 => x"81fe0653",
   347 => x"81d05281",
   348 => x"bfd80851",
   349 => x"80c9d33f",
   350 => x"b008982b",
   351 => x"54807424",
   352 => x"a238819c",
   353 => x"c85180e3",
   354 => x"8b3f7452",
   355 => x"885180e3",
   356 => x"a63f819c",
   357 => x"d45180e2",
   358 => x"fb3f8116",
   359 => x"7083ffff",
   360 => x"06575481",
   361 => x"157081ff",
   362 => x"0670982b",
   363 => x"52565473",
   364 => x"8025ffb2",
   365 => x"3875b00c",
   366 => x"873d0d04",
   367 => x"f33d0d7f",
   368 => x"02840580",
   369 => x"c3053302",
   370 => x"880580c6",
   371 => x"0522819c",
   372 => x"e4545b55",
   373 => x"5880e2bc",
   374 => x"3f785180",
   375 => x"e4803f81",
   376 => x"9cf05180",
   377 => x"e2ae3f73",
   378 => x"52885180",
   379 => x"e2c93f81",
   380 => x"9d8c5180",
   381 => x"e29e3f80",
   382 => x"57767927",
   383 => x"81a13873",
   384 => x"108e3d5d",
   385 => x"5a7981ff",
   386 => x"06538190",
   387 => x"52775180",
   388 => x"c8b83f76",
   389 => x"882a5390",
   390 => x"52775180",
   391 => x"c8ac3f76",
   392 => x"81ff0653",
   393 => x"90527751",
   394 => x"80c89f3f",
   395 => x"811a7081",
   396 => x"ff065455",
   397 => x"81905277",
   398 => x"5180c88e",
   399 => x"3f805380",
   400 => x"e0527751",
   401 => x"80c8833f",
   402 => x"b008982b",
   403 => x"54807424",
   404 => x"8a388818",
   405 => x"087081ff",
   406 => x"065c567a",
   407 => x"81ff0681",
   408 => x"9cb45256",
   409 => x"80e1ad3f",
   410 => x"75528851",
   411 => x"80e1c83f",
   412 => x"81a78051",
   413 => x"80e19d3f",
   414 => x"e0165480",
   415 => x"df7427b6",
   416 => x"38768706",
   417 => x"701d5755",
   418 => x"a0763474",
   419 => x"872eb938",
   420 => x"81177083",
   421 => x"ffff0658",
   422 => x"55787726",
   423 => x"fee73880",
   424 => x"e00b8c19",
   425 => x"0c8c1808",
   426 => x"70812a81",
   427 => x"06585a76",
   428 => x"f4388f3d",
   429 => x"0d047687",
   430 => x"06701d55",
   431 => x"55757434",
   432 => x"74872e09",
   433 => x"8106c938",
   434 => x"7b5180e0",
   435 => x"c73f8a51",
   436 => x"80e0a73f",
   437 => x"81177083",
   438 => x"ffff0658",
   439 => x"55787726",
   440 => x"fea338ff",
   441 => x"ba39fb3d",
   442 => x"0d815180",
   443 => x"c0953fb0",
   444 => x"0881ff06",
   445 => x"54825180",
   446 => x"c1bb3fb0",
   447 => x"0881ff06",
   448 => x"568351bf",
   449 => x"fe3fb008",
   450 => x"83ffff06",
   451 => x"55739c38",
   452 => x"81bfd808",
   453 => x"54748438",
   454 => x"81805574",
   455 => x"53755273",
   456 => x"51fd993f",
   457 => x"74b00c87",
   458 => x"3d0d0481",
   459 => x"bfdc0854",
   460 => x"e439f83d",
   461 => x"0d02aa05",
   462 => x"2281bfb4",
   463 => x"3381f706",
   464 => x"58587681",
   465 => x"bfb43481",
   466 => x"bfd80855",
   467 => x"80c05381",
   468 => x"90527451",
   469 => x"80c5f33f",
   470 => x"745180c6",
   471 => x"9f3fb008",
   472 => x"81ff0654",
   473 => x"73802e84",
   474 => x"90387653",
   475 => x"80d05274",
   476 => x"5180c5d6",
   477 => x"3f80598f",
   478 => x"5781bfb4",
   479 => x"3381fe06",
   480 => x"547381bf",
   481 => x"b43481bf",
   482 => x"d8087457",
   483 => x"5580c053",
   484 => x"81905274",
   485 => x"5180c5b2",
   486 => x"3f745180",
   487 => x"c5de3fb0",
   488 => x"0881ff06",
   489 => x"5473802e",
   490 => x"83c43875",
   491 => x"5380d052",
   492 => x"745180c5",
   493 => x"953f7777",
   494 => x"2c810655",
   495 => x"74802e83",
   496 => x"a23881bf",
   497 => x"b4338207",
   498 => x"547381bf",
   499 => x"b43481bf",
   500 => x"d8087457",
   501 => x"5580c053",
   502 => x"81905274",
   503 => x"5180c4ea",
   504 => x"3f745180",
   505 => x"c5963fb0",
   506 => x"0881ff06",
   507 => x"5473802e",
   508 => x"82e63875",
   509 => x"5380d052",
   510 => x"745180c4",
   511 => x"cd3f81bf",
   512 => x"d8085580",
   513 => x"c1538190",
   514 => x"52745180",
   515 => x"c4bc3f74",
   516 => x"5180c4e8",
   517 => x"3fb00881",
   518 => x"ff065675",
   519 => x"802e828c",
   520 => x"38805380",
   521 => x"e0527451",
   522 => x"80c49f3f",
   523 => x"745180c4",
   524 => x"cb3fb008",
   525 => x"81ff0654",
   526 => x"73802e81",
   527 => x"ef388815",
   528 => x"0870902b",
   529 => x"70902c56",
   530 => x"56567382",
   531 => x"2a810654",
   532 => x"73802e8d",
   533 => x"3881772b",
   534 => x"79077083",
   535 => x"ffff065a",
   536 => x"5681bfb4",
   537 => x"33810754",
   538 => x"7381bfb4",
   539 => x"3481bfd8",
   540 => x"08745755",
   541 => x"80c05381",
   542 => x"90527451",
   543 => x"80c3cb3f",
   544 => x"745180c3",
   545 => x"f73fb008",
   546 => x"81ff0654",
   547 => x"73802e81",
   548 => x"a8387553",
   549 => x"80d05274",
   550 => x"5180c3ae",
   551 => x"3f768180",
   552 => x"0a2981ff",
   553 => x"0a057098",
   554 => x"2c585676",
   555 => x"8025fdc9",
   556 => x"3881bfb4",
   557 => x"33820757",
   558 => x"7681bfb4",
   559 => x"3481bfd8",
   560 => x"085580c0",
   561 => x"53819052",
   562 => x"745180c2",
   563 => x"fd3f7451",
   564 => x"80c3a93f",
   565 => x"b00881ff",
   566 => x"06587780",
   567 => x"2e81b838",
   568 => x"765380d0",
   569 => x"52745180",
   570 => x"c2e03f81",
   571 => x"bfb43388",
   572 => x"07577681",
   573 => x"bfb43481",
   574 => x"bfd80855",
   575 => x"80c05381",
   576 => x"90527451",
   577 => x"80c2c33f",
   578 => x"745180c2",
   579 => x"ef3fb008",
   580 => x"81ff0658",
   581 => x"77802e80",
   582 => x"ef387653",
   583 => x"80d05274",
   584 => x"5180c2a6",
   585 => x"3f78b00c",
   586 => x"8a3d0d04",
   587 => x"819d9051",
   588 => x"80dbe13f",
   589 => x"ff54fe92",
   590 => x"39819d90",
   591 => x"5180dbd4",
   592 => x"3f768180",
   593 => x"0a2981ff",
   594 => x"0a057098",
   595 => x"2c585676",
   596 => x"8025fca5",
   597 => x"38feda39",
   598 => x"819d9051",
   599 => x"80dbb53f",
   600 => x"fd9c3981",
   601 => x"bfb43381",
   602 => x"fd0654fc",
   603 => x"dc39819d",
   604 => x"905180db",
   605 => x"9f3ffcbe",
   606 => x"39819d90",
   607 => x"5180db94",
   608 => x"3f80598f",
   609 => x"57fbf239",
   610 => x"819d9051",
   611 => x"80db853f",
   612 => x"78b00c8a",
   613 => x"3d0d0481",
   614 => x"9d905180",
   615 => x"daf63ffe",
   616 => x"ca39ff3d",
   617 => x"0d8151ba",
   618 => x"da3fb008",
   619 => x"81ff0652",
   620 => x"818051fa",
   621 => x"fd3f8280",
   622 => x"51faf73f",
   623 => x"848351fa",
   624 => x"f13f86f1",
   625 => x"51faeb3f",
   626 => x"71832b88",
   627 => x"830751fa",
   628 => x"e13f71b0",
   629 => x"0c833d0d",
   630 => x"04fe3d0d",
   631 => x"74708106",
   632 => x"53537185",
   633 => x"d0387281",
   634 => x"2a708106",
   635 => x"51527185",
   636 => x"ac387282",
   637 => x"2a708106",
   638 => x"51527185",
   639 => x"88387283",
   640 => x"2a708106",
   641 => x"51527184",
   642 => x"e4387284",
   643 => x"2a708106",
   644 => x"51527184",
   645 => x"c0387285",
   646 => x"2a708106",
   647 => x"51527184",
   648 => x"9c387286",
   649 => x"2a708106",
   650 => x"51527183",
   651 => x"f8387287",
   652 => x"2a708106",
   653 => x"51527183",
   654 => x"d4387288",
   655 => x"2a708106",
   656 => x"51527183",
   657 => x"b0387289",
   658 => x"2a708106",
   659 => x"51527183",
   660 => x"8c38728a",
   661 => x"2a708106",
   662 => x"51527182",
   663 => x"e838728b",
   664 => x"2a708106",
   665 => x"51527182",
   666 => x"c438728c",
   667 => x"2a708106",
   668 => x"51527182",
   669 => x"a038728d",
   670 => x"2a708106",
   671 => x"51527181",
   672 => x"fc38728e",
   673 => x"2a708106",
   674 => x"51527181",
   675 => x"d838728f",
   676 => x"2a708106",
   677 => x"51527181",
   678 => x"b4387290",
   679 => x"2a708106",
   680 => x"51527181",
   681 => x"90387291",
   682 => x"2a708106",
   683 => x"51527180",
   684 => x"ec387292",
   685 => x"2a708106",
   686 => x"51527180",
   687 => x"c8387293",
   688 => x"2a708106",
   689 => x"515271a6",
   690 => x"3872942a",
   691 => x"70810651",
   692 => x"52718b38",
   693 => x"80732483",
   694 => x"f438843d",
   695 => x"0d04819d",
   696 => x"c85180d8",
   697 => x"af3f7280",
   698 => x"25f03883",
   699 => x"e039819d",
   700 => x"e45180d8",
   701 => x"9f3f7294",
   702 => x"2a708106",
   703 => x"51527180",
   704 => x"2ed238da",
   705 => x"39819e80",
   706 => x"5180d888",
   707 => x"3f72932a",
   708 => x"70810651",
   709 => x"5271802e",
   710 => x"ffaf38d2",
   711 => x"39819e9c",
   712 => x"5180d7f0",
   713 => x"3f72922a",
   714 => x"70810651",
   715 => x"5271802e",
   716 => x"ff8c38d1",
   717 => x"39819eb8",
   718 => x"5180d7d8",
   719 => x"3f72912a",
   720 => x"70810651",
   721 => x"5271802e",
   722 => x"fee838d1",
   723 => x"39819ed8",
   724 => x"5180d7c0",
   725 => x"3f72902a",
   726 => x"70810651",
   727 => x"5271802e",
   728 => x"fec438d1",
   729 => x"39819ef8",
   730 => x"5180d7a8",
   731 => x"3f728f2a",
   732 => x"70810651",
   733 => x"5271802e",
   734 => x"fea038d1",
   735 => x"39819f98",
   736 => x"5180d790",
   737 => x"3f728e2a",
   738 => x"70810651",
   739 => x"5271802e",
   740 => x"fdfc38d1",
   741 => x"39819fb8",
   742 => x"5180d6f8",
   743 => x"3f728d2a",
   744 => x"70810651",
   745 => x"5271802e",
   746 => x"fdd838d1",
   747 => x"39819fcc",
   748 => x"5180d6e0",
   749 => x"3f728c2a",
   750 => x"70810651",
   751 => x"5271802e",
   752 => x"fdb438d1",
   753 => x"39819fec",
   754 => x"5180d6c8",
   755 => x"3f728b2a",
   756 => x"70810651",
   757 => x"5271802e",
   758 => x"fd9038d1",
   759 => x"3981a094",
   760 => x"5180d6b0",
   761 => x"3f728a2a",
   762 => x"70810651",
   763 => x"5271802e",
   764 => x"fcec38d1",
   765 => x"3981a0b4",
   766 => x"5180d698",
   767 => x"3f72892a",
   768 => x"70810651",
   769 => x"5271802e",
   770 => x"fcc838d1",
   771 => x"3981a0d4",
   772 => x"5180d680",
   773 => x"3f72882a",
   774 => x"70810651",
   775 => x"5271802e",
   776 => x"fca438d1",
   777 => x"3981a0fc",
   778 => x"5180d5e8",
   779 => x"3f72872a",
   780 => x"70810651",
   781 => x"5271802e",
   782 => x"fc8038d1",
   783 => x"3981a19c",
   784 => x"5180d5d0",
   785 => x"3f72862a",
   786 => x"70810651",
   787 => x"5271802e",
   788 => x"fbdc38d1",
   789 => x"3981a1bc",
   790 => x"5180d5b8",
   791 => x"3f72852a",
   792 => x"70810651",
   793 => x"5271802e",
   794 => x"fbb838d1",
   795 => x"3981a1e4",
   796 => x"5180d5a0",
   797 => x"3f72842a",
   798 => x"70810651",
   799 => x"5271802e",
   800 => x"fb9438d1",
   801 => x"3981a284",
   802 => x"5180d588",
   803 => x"3f72832a",
   804 => x"70810651",
   805 => x"5271802e",
   806 => x"faf038d1",
   807 => x"3981a2a4",
   808 => x"5180d4f0",
   809 => x"3f72822a",
   810 => x"70810651",
   811 => x"5271802e",
   812 => x"facc38d1",
   813 => x"3981a2cc",
   814 => x"5180d4d8",
   815 => x"3f72812a",
   816 => x"70810651",
   817 => x"5271802e",
   818 => x"faa838d1",
   819 => x"3981a2ec",
   820 => x"5180d4c0",
   821 => x"3f843d0d",
   822 => x"04fd3d0d",
   823 => x"81a38051",
   824 => x"80d4b13f",
   825 => x"81bfe408",
   826 => x"7008709e",
   827 => x"2a708106",
   828 => x"51525553",
   829 => x"81547283",
   830 => x"38725473",
   831 => x"802e88c4",
   832 => x"3881a39c",
   833 => x"5180d48c",
   834 => x"3f81a3a4",
   835 => x"5180d484",
   836 => x"3f81bfe4",
   837 => x"08841108",
   838 => x"709d2a81",
   839 => x"06515553",
   840 => x"73802e87",
   841 => x"b03881a3",
   842 => x"c05180d3",
   843 => x"e73f81a3",
   844 => x"cc5180d3",
   845 => x"df3f81bf",
   846 => x"ac0880d4",
   847 => x"11085254",
   848 => x"80d59b3f",
   849 => x"81a3e851",
   850 => x"80d3c93f",
   851 => x"81bfac08",
   852 => x"80d01108",
   853 => x"525380d5",
   854 => x"853f8a51",
   855 => x"80d39b3f",
   856 => x"81a48451",
   857 => x"80d3ad3f",
   858 => x"81a4a851",
   859 => x"80d3a53f",
   860 => x"81a4f051",
   861 => x"80d39d3f",
   862 => x"81a5b851",
   863 => x"80d3953f",
   864 => x"81bfac08",
   865 => x"70085254",
   866 => x"80d4d33f",
   867 => x"b00881ff",
   868 => x"0653728c",
   869 => x"279438a0",
   870 => x"5180d2de",
   871 => x"3f811370",
   872 => x"81ff0651",
   873 => x"538c7326",
   874 => x"ee3881bf",
   875 => x"ac088411",
   876 => x"08525480",
   877 => x"d4a83fb0",
   878 => x"0881ff06",
   879 => x"53728c27",
   880 => x"9438a051",
   881 => x"80d2b33f",
   882 => x"81137081",
   883 => x"ff065153",
   884 => x"8c7326ee",
   885 => x"3881bfac",
   886 => x"08881108",
   887 => x"525480d3",
   888 => x"fd3fb008",
   889 => x"81ff0653",
   890 => x"728c2794",
   891 => x"38a05180",
   892 => x"d2883f81",
   893 => x"137081ff",
   894 => x"0651538c",
   895 => x"7326ee38",
   896 => x"81bfac08",
   897 => x"8c110852",
   898 => x"5480d3d2",
   899 => x"3fb00881",
   900 => x"ff065372",
   901 => x"8c279438",
   902 => x"a05180d1",
   903 => x"dd3f8113",
   904 => x"7081ff06",
   905 => x"51538c73",
   906 => x"26ee3881",
   907 => x"a5d45180",
   908 => x"d1e23f81",
   909 => x"bfac0890",
   910 => x"11085254",
   911 => x"80d39f3f",
   912 => x"b00881ff",
   913 => x"0653728c",
   914 => x"279438a0",
   915 => x"5180d1aa",
   916 => x"3f811370",
   917 => x"81ff0651",
   918 => x"538c7326",
   919 => x"ee3881bf",
   920 => x"ac089411",
   921 => x"08525480",
   922 => x"d2f43fb0",
   923 => x"0881ff06",
   924 => x"53728c27",
   925 => x"9438a051",
   926 => x"80d0ff3f",
   927 => x"81137081",
   928 => x"ff065153",
   929 => x"8c7326ee",
   930 => x"3881bfac",
   931 => x"08981108",
   932 => x"525480d2",
   933 => x"c93fb008",
   934 => x"81ff0653",
   935 => x"728c2794",
   936 => x"38a05180",
   937 => x"d0d43f81",
   938 => x"137081ff",
   939 => x"0651538c",
   940 => x"7326ee38",
   941 => x"81bfac08",
   942 => x"9c110852",
   943 => x"5480d29e",
   944 => x"3fb00881",
   945 => x"ff065372",
   946 => x"8c279438",
   947 => x"a05180d0",
   948 => x"a93f8113",
   949 => x"7081ff06",
   950 => x"51538c73",
   951 => x"26ee3881",
   952 => x"a5f05180",
   953 => x"d0ae3f81",
   954 => x"bfac0854",
   955 => x"810bb015",
   956 => x"0cb01408",
   957 => x"53728025",
   958 => x"f838a014",
   959 => x"085180d1",
   960 => x"dd3fb008",
   961 => x"81ff0653",
   962 => x"728c2794",
   963 => x"38a05180",
   964 => x"cfe83f81",
   965 => x"137081ff",
   966 => x"0654548c",
   967 => x"7326ee38",
   968 => x"81bfac08",
   969 => x"a4110852",
   970 => x"5380d1b2",
   971 => x"3fb00881",
   972 => x"ff065372",
   973 => x"8c279438",
   974 => x"a05180cf",
   975 => x"bd3f8113",
   976 => x"7081ff06",
   977 => x"54548c73",
   978 => x"26ee3881",
   979 => x"bfac08a8",
   980 => x"11085253",
   981 => x"80d1873f",
   982 => x"b00881ff",
   983 => x"0653728c",
   984 => x"279438a0",
   985 => x"5180cf92",
   986 => x"3f811370",
   987 => x"81ff0654",
   988 => x"548c7326",
   989 => x"ee3881bf",
   990 => x"ac08ac11",
   991 => x"08525380",
   992 => x"d0dc3fb0",
   993 => x"0881ff06",
   994 => x"53728c27",
   995 => x"9438a051",
   996 => x"80cee73f",
   997 => x"81137081",
   998 => x"ff065454",
   999 => x"8c7326ee",
  1000 => x"3881a68c",
  1001 => x"5180ceec",
  1002 => x"3f81bfac",
  1003 => x"0880e011",
  1004 => x"08525380",
  1005 => x"d0a83f81",
  1006 => x"a6a05180",
  1007 => x"ced63f81",
  1008 => x"bfac08b0",
  1009 => x"1108fe0a",
  1010 => x"06525480",
  1011 => x"d0903f81",
  1012 => x"bfac0854",
  1013 => x"800bb015",
  1014 => x"0c81a6b4",
  1015 => x"5180ceb4",
  1016 => x"3f81a6cc",
  1017 => x"5180ceac",
  1018 => x"3f81bfac",
  1019 => x"0880c011",
  1020 => x"08525380",
  1021 => x"cfe83fb0",
  1022 => x"0881ff06",
  1023 => x"53729827",
  1024 => x"9438a051",
  1025 => x"80cdf33f",
  1026 => x"81137081",
  1027 => x"ff065454",
  1028 => x"987326ee",
  1029 => x"3881bfac",
  1030 => x"0880c811",
  1031 => x"08525380",
  1032 => x"cfbc3fb0",
  1033 => x"0881ff06",
  1034 => x"53729827",
  1035 => x"9438a051",
  1036 => x"80cdc73f",
  1037 => x"81137081",
  1038 => x"ff065454",
  1039 => x"987326ee",
  1040 => x"3881a6e8",
  1041 => x"5180cdcc",
  1042 => x"3f81bfac",
  1043 => x"0880c411",
  1044 => x"08525380",
  1045 => x"cf883fb0",
  1046 => x"0881ff06",
  1047 => x"53729827",
  1048 => x"9438a051",
  1049 => x"80cd933f",
  1050 => x"81137081",
  1051 => x"ff065454",
  1052 => x"987326ee",
  1053 => x"3881bfac",
  1054 => x"0880cc11",
  1055 => x"08525380",
  1056 => x"cedc3fb0",
  1057 => x"0881ff06",
  1058 => x"53729827",
  1059 => x"9438a051",
  1060 => x"80cce73f",
  1061 => x"81137081",
  1062 => x"ff065454",
  1063 => x"987326ee",
  1064 => x"388a5180",
  1065 => x"ccd43f81",
  1066 => x"bfac08b4",
  1067 => x"110881a7",
  1068 => x"84535153",
  1069 => x"80ccdd3f",
  1070 => x"725180ce",
  1071 => x"a13fa051",
  1072 => x"80ccb73f",
  1073 => x"72862681",
  1074 => x"8e387210",
  1075 => x"1081b394",
  1076 => x"05547308",
  1077 => x"0481a798",
  1078 => x"5180ccb8",
  1079 => x"3f81a3cc",
  1080 => x"5180ccb0",
  1081 => x"3f81bfac",
  1082 => x"0880d411",
  1083 => x"08525480",
  1084 => x"cdec3f81",
  1085 => x"a3e85180",
  1086 => x"cc9a3f81",
  1087 => x"bfac0880",
  1088 => x"d0110852",
  1089 => x"5380cdd6",
  1090 => x"3f8a5180",
  1091 => x"cbec3f81",
  1092 => x"a4845180",
  1093 => x"cbfe3f81",
  1094 => x"a4a85180",
  1095 => x"cbf63f81",
  1096 => x"a4f05180",
  1097 => x"cbee3f81",
  1098 => x"a5b85180",
  1099 => x"cbe63f81",
  1100 => x"bfac0870",
  1101 => x"08525480",
  1102 => x"cda43fb0",
  1103 => x"0881ff06",
  1104 => x"53f8cf39",
  1105 => x"81a7a051",
  1106 => x"80cbc93f",
  1107 => x"f7b33981",
  1108 => x"a7a85180",
  1109 => x"cbbe3f81",
  1110 => x"bfac08b8",
  1111 => x"110881a7",
  1112 => x"b4535454",
  1113 => x"80cbad3f",
  1114 => x"7252a051",
  1115 => x"80cbc83f",
  1116 => x"7251f0e5",
  1117 => x"3f8a5180",
  1118 => x"cb803f80",
  1119 => x"0bb00c85",
  1120 => x"3d0d0481",
  1121 => x"a7c85180",
  1122 => x"cb8a3fcb",
  1123 => x"3981a7d4",
  1124 => x"5180cb80",
  1125 => x"3fc13981",
  1126 => x"a7e05180",
  1127 => x"caf63fff",
  1128 => x"b63981a7",
  1129 => x"e45180ca",
  1130 => x"eb3fffab",
  1131 => x"3981a7f0",
  1132 => x"5180cae0",
  1133 => x"3fffa039",
  1134 => x"81a7fc51",
  1135 => x"80cad53f",
  1136 => x"ff9539fe",
  1137 => x"3d0d8151",
  1138 => x"aab93fb0",
  1139 => x"0881ff06",
  1140 => x"81bfac08",
  1141 => x"71b4120c",
  1142 => x"53b00c84",
  1143 => x"3d0d04fe",
  1144 => x"3d0d880a",
  1145 => x"53840a0b",
  1146 => x"81bfa808",
  1147 => x"8c110851",
  1148 => x"52528071",
  1149 => x"27953880",
  1150 => x"73708405",
  1151 => x"550c8072",
  1152 => x"70840554",
  1153 => x"0cff1151",
  1154 => x"70ed3880",
  1155 => x"0bb00c84",
  1156 => x"3d0d04fa",
  1157 => x"3d0d880a",
  1158 => x"57840a56",
  1159 => x"8151a9e3",
  1160 => x"3fb00883",
  1161 => x"ffff0654",
  1162 => x"73833890",
  1163 => x"54805574",
  1164 => x"742781c2",
  1165 => x"38750870",
  1166 => x"902c5253",
  1167 => x"80cb9f3f",
  1168 => x"b00881ff",
  1169 => x"0652718a",
  1170 => x"279438a0",
  1171 => x"5180c9aa",
  1172 => x"3f811270",
  1173 => x"81ff0651",
  1174 => x"528a7226",
  1175 => x"ee387290",
  1176 => x"2b70902c",
  1177 => x"525280ca",
  1178 => x"f53fb008",
  1179 => x"81ff0652",
  1180 => x"718a2794",
  1181 => x"38a05180",
  1182 => x"c9803f81",
  1183 => x"127081ff",
  1184 => x"0653538a",
  1185 => x"7226ee38",
  1186 => x"76087090",
  1187 => x"2c525380",
  1188 => x"cacc3fb0",
  1189 => x"0881ff06",
  1190 => x"52718a27",
  1191 => x"9438a051",
  1192 => x"80c8d73f",
  1193 => x"81127081",
  1194 => x"ff065152",
  1195 => x"8a7226ee",
  1196 => x"3872902b",
  1197 => x"70902c52",
  1198 => x"5280caa2",
  1199 => x"3fb00881",
  1200 => x"ff065271",
  1201 => x"8a279438",
  1202 => x"a05180c8",
  1203 => x"ad3f8112",
  1204 => x"7081ff06",
  1205 => x"53538a72",
  1206 => x"26ee388a",
  1207 => x"5180c89a",
  1208 => x"3f841784",
  1209 => x"17811770",
  1210 => x"83ffff06",
  1211 => x"58545757",
  1212 => x"737526fe",
  1213 => x"c03873b0",
  1214 => x"0c883d0d",
  1215 => x"04fd3d0d",
  1216 => x"8151a7ff",
  1217 => x"3fb00881",
  1218 => x"ff065473",
  1219 => x"802ea438",
  1220 => x"73842690",
  1221 => x"3881bfa8",
  1222 => x"0874710c",
  1223 => x"5373b00c",
  1224 => x"853d0d04",
  1225 => x"81bfa808",
  1226 => x"5380730c",
  1227 => x"73b00c85",
  1228 => x"3d0d0481",
  1229 => x"a9885180",
  1230 => x"c7da3f81",
  1231 => x"a9985180",
  1232 => x"c7d23f81",
  1233 => x"bfa80870",
  1234 => x"08525380",
  1235 => x"c9903f81",
  1236 => x"a9a85180",
  1237 => x"c7be3f81",
  1238 => x"bfa80884",
  1239 => x"11085353",
  1240 => x"a05180c7",
  1241 => x"d23f81a9",
  1242 => x"bc5180c7",
  1243 => x"a73f81bf",
  1244 => x"a8088811",
  1245 => x"085353a0",
  1246 => x"5180c7bb",
  1247 => x"3f81a9d0",
  1248 => x"5180c790",
  1249 => x"3f81bfa8",
  1250 => x"088c1108",
  1251 => x"525380c8",
  1252 => x"cd3f8a51",
  1253 => x"80c6e33f",
  1254 => x"73b00c85",
  1255 => x"3d0d04bc",
  1256 => x"0802bc0c",
  1257 => x"f93d0d02",
  1258 => x"bc08fc05",
  1259 => x"0c880a0b",
  1260 => x"bc08f405",
  1261 => x"0cfc3d0d",
  1262 => x"823dbc08",
  1263 => x"f0050c81",
  1264 => x"51a6c03f",
  1265 => x"b00881ff",
  1266 => x"06bc08f8",
  1267 => x"050c8251",
  1268 => x"a6b13fb0",
  1269 => x"08bc08f0",
  1270 => x"05082383",
  1271 => x"51a6a43f",
  1272 => x"b008bc08",
  1273 => x"f0050882",
  1274 => x"05238451",
  1275 => x"a6953fb0",
  1276 => x"08bc08f0",
  1277 => x"05088405",
  1278 => x"238551a6",
  1279 => x"863fb008",
  1280 => x"bc08f005",
  1281 => x"08860523",
  1282 => x"8651a5f7",
  1283 => x"3fb008bc",
  1284 => x"08f00508",
  1285 => x"88052387",
  1286 => x"51a5e83f",
  1287 => x"b008bc08",
  1288 => x"f005088a",
  1289 => x"05238851",
  1290 => x"a5d93fb0",
  1291 => x"08bc08f0",
  1292 => x"05088c05",
  1293 => x"238951a5",
  1294 => x"ca3fb008",
  1295 => x"bc08f005",
  1296 => x"088e0523",
  1297 => x"800b81bf",
  1298 => x"a808708c",
  1299 => x"050851bc",
  1300 => x"08e4050c",
  1301 => x"bc08ec05",
  1302 => x"0cbc08ec",
  1303 => x"0508bc08",
  1304 => x"e4050827",
  1305 => x"818f38bc",
  1306 => x"08e40508",
  1307 => x"bc08e805",
  1308 => x"0cbc08f8",
  1309 => x"0508802e",
  1310 => x"81b638bc",
  1311 => x"08ec0508",
  1312 => x"10bc08f0",
  1313 => x"05080570",
  1314 => x"22bc08f4",
  1315 => x"05088205",
  1316 => x"2271902b",
  1317 => x"07bc08f4",
  1318 => x"05080cbc",
  1319 => x"08e4050c",
  1320 => x"bc08f805",
  1321 => x"0cbc08ec",
  1322 => x"05088105",
  1323 => x"7081ff06",
  1324 => x"bc08e405",
  1325 => x"0cbc08f8",
  1326 => x"050c860b",
  1327 => x"bc08ec05",
  1328 => x"08278838",
  1329 => x"800bbc08",
  1330 => x"e4050cbc",
  1331 => x"08e40508",
  1332 => x"bc08f405",
  1333 => x"088405bc",
  1334 => x"08e80508",
  1335 => x"ff05bc08",
  1336 => x"e8050cbc",
  1337 => x"08f4050c",
  1338 => x"bc08ec05",
  1339 => x"0cbc08e8",
  1340 => x"0508ff87",
  1341 => x"38bc08fc",
  1342 => x"05080d80",
  1343 => x"0bb00c89",
  1344 => x"3d0dbc0c",
  1345 => x"04bc08e4",
  1346 => x"0508bc08",
  1347 => x"f4050884",
  1348 => x"05bc08e8",
  1349 => x"0508ff05",
  1350 => x"bc08e805",
  1351 => x"0cbc08f4",
  1352 => x"050cbc08",
  1353 => x"ec050cbc",
  1354 => x"08e80508",
  1355 => x"802ec638",
  1356 => x"bc08ec05",
  1357 => x"0810bc08",
  1358 => x"f0050805",
  1359 => x"70227090",
  1360 => x"2bbc08f4",
  1361 => x"050808fc",
  1362 => x"80800671",
  1363 => x"902c07bc",
  1364 => x"08f40508",
  1365 => x"0c52bc08",
  1366 => x"e4050cbc",
  1367 => x"08f8050c",
  1368 => x"800bbc08",
  1369 => x"e4050cbc",
  1370 => x"08ec0508",
  1371 => x"8626ff95",
  1372 => x"38bc08ec",
  1373 => x"05088105",
  1374 => x"7081ff06",
  1375 => x"bc08f405",
  1376 => x"088405bc",
  1377 => x"08e80508",
  1378 => x"ff05bc08",
  1379 => x"e8050cbc",
  1380 => x"08f4050c",
  1381 => x"bc08ec05",
  1382 => x"0cbc08e4",
  1383 => x"050cbc08",
  1384 => x"e80508ff",
  1385 => x"8b38fecd",
  1386 => x"39fb3d0d",
  1387 => x"029f0533",
  1388 => x"79982b70",
  1389 => x"982c5154",
  1390 => x"55810a54",
  1391 => x"805672e8",
  1392 => x"25bd38e8",
  1393 => x"53751081",
  1394 => x"07738180",
  1395 => x"0a298180",
  1396 => x"0a057098",
  1397 => x"2c515456",
  1398 => x"807324e9",
  1399 => x"38807325",
  1400 => x"80c73873",
  1401 => x"812a810a",
  1402 => x"07738180",
  1403 => x"0a2981ff",
  1404 => x"0a057098",
  1405 => x"2c515454",
  1406 => x"728024e7",
  1407 => x"38ab3997",
  1408 => x"73259a38",
  1409 => x"9774812a",
  1410 => x"810a0771",
  1411 => x"81800a29",
  1412 => x"81ff0a05",
  1413 => x"70982c51",
  1414 => x"525553dc",
  1415 => x"39807324",
  1416 => x"ffa33872",
  1417 => x"8024ffbb",
  1418 => x"38745280",
  1419 => x"51a8e33f",
  1420 => x"7381ff06",
  1421 => x"51a9e13f",
  1422 => x"74528151",
  1423 => x"a8d43f73",
  1424 => x"882a7081",
  1425 => x"ff065253",
  1426 => x"a9ce3f74",
  1427 => x"528251a8",
  1428 => x"c13f7390",
  1429 => x"2a7081ff",
  1430 => x"065253a9",
  1431 => x"bb3f7452",
  1432 => x"8351a8ae",
  1433 => x"3f73982a",
  1434 => x"51a9ad3f",
  1435 => x"74528451",
  1436 => x"a8a03f75",
  1437 => x"81ff0651",
  1438 => x"a99e3f74",
  1439 => x"528551a8",
  1440 => x"913f7588",
  1441 => x"2a7081ff",
  1442 => x"065253a9",
  1443 => x"8b3f7452",
  1444 => x"8651a7fe",
  1445 => x"3f75902a",
  1446 => x"7081ff06",
  1447 => x"5254a8f8",
  1448 => x"3f745287",
  1449 => x"51a7eb3f",
  1450 => x"75982a51",
  1451 => x"a8ea3f87",
  1452 => x"3d0d04f2",
  1453 => x"3d0d0280",
  1454 => x"c3053302",
  1455 => x"840580c7",
  1456 => x"05338180",
  1457 => x"0a712b98",
  1458 => x"2a81bfa8",
  1459 => x"088c1108",
  1460 => x"71084453",
  1461 => x"565c5557",
  1462 => x"80730c80",
  1463 => x"7071725c",
  1464 => x"5a5e5b80",
  1465 => x"56757a27",
  1466 => x"80d73881",
  1467 => x"772783c6",
  1468 => x"387783ff",
  1469 => x"ff068119",
  1470 => x"71101084",
  1471 => x"0a057930",
  1472 => x"7a823270",
  1473 => x"30728025",
  1474 => x"71802507",
  1475 => x"56585841",
  1476 => x"57595c7b",
  1477 => x"802e83cd",
  1478 => x"38821522",
  1479 => x"5372902b",
  1480 => x"70902c54",
  1481 => x"55727b25",
  1482 => x"8338725b",
  1483 => x"7c732583",
  1484 => x"38725d81",
  1485 => x"167081ff",
  1486 => x"06575e79",
  1487 => x"7626ffb1",
  1488 => x"38811970",
  1489 => x"81ff065a",
  1490 => x"5680e579",
  1491 => x"27ff9438",
  1492 => x"987d3590",
  1493 => x"2b70902c",
  1494 => x"7c309871",
  1495 => x"35902b70",
  1496 => x"902c5c5c",
  1497 => x"55565477",
  1498 => x"54777525",
  1499 => x"83387454",
  1500 => x"73902b70",
  1501 => x"902c5d55",
  1502 => x"7b54807c",
  1503 => x"2583cf38",
  1504 => x"73902b70",
  1505 => x"902c5f56",
  1506 => x"80705d58",
  1507 => x"80705a56",
  1508 => x"757a2780",
  1509 => x"e4388177",
  1510 => x"27838438",
  1511 => x"7783ffff",
  1512 => x"06811971",
  1513 => x"1010840a",
  1514 => x"0579307a",
  1515 => x"82327030",
  1516 => x"72802571",
  1517 => x"80250753",
  1518 => x"51575357",
  1519 => x"59547380",
  1520 => x"2e839c38",
  1521 => x"82152254",
  1522 => x"73902b70",
  1523 => x"902c719f",
  1524 => x"2c707232",
  1525 => x"7131799f",
  1526 => x"2c707b32",
  1527 => x"71315154",
  1528 => x"51565653",
  1529 => x"72742583",
  1530 => x"38745681",
  1531 => x"197081ff",
  1532 => x"065a5579",
  1533 => x"7926ffa4",
  1534 => x"387d7635",
  1535 => x"982b7098",
  1536 => x"2c53547b",
  1537 => x"51fba23f",
  1538 => x"811c7081",
  1539 => x"ff065d59",
  1540 => x"80e57c27",
  1541 => x"fef63881",
  1542 => x"bfa8087f",
  1543 => x"710c5880",
  1544 => x"5281b484",
  1545 => x"51a8e13f",
  1546 => x"81e3c408",
  1547 => x"80eacc0b",
  1548 => x"81e3c40c",
  1549 => x"5f805280",
  1550 => x"51a4d73f",
  1551 => x"81a9e051",
  1552 => x"bdd23f7c",
  1553 => x"51bf973f",
  1554 => x"80528751",
  1555 => x"a4c43f81",
  1556 => x"a9e851bd",
  1557 => x"bf3f7a51",
  1558 => x"bf843f80",
  1559 => x"d2528051",
  1560 => x"a4b03f81",
  1561 => x"a9f051bd",
  1562 => x"ab3f7651",
  1563 => x"bef03f80",
  1564 => x"c0528751",
  1565 => x"a49c3f81",
  1566 => x"a9f851bd",
  1567 => x"973f7980",
  1568 => x"e62951be",
  1569 => x"d93f7e81",
  1570 => x"e3c40c90",
  1571 => x"3d0d0474",
  1572 => x"22537290",
  1573 => x"2b70902c",
  1574 => x"545c727b",
  1575 => x"25833872",
  1576 => x"5b7c7325",
  1577 => x"8338725d",
  1578 => x"81167081",
  1579 => x"ff06575e",
  1580 => x"757a27fd",
  1581 => x"8c387783",
  1582 => x"ffff0681",
  1583 => x"19711010",
  1584 => x"880a0579",
  1585 => x"307a8232",
  1586 => x"70307280",
  1587 => x"25718025",
  1588 => x"07565840",
  1589 => x"41575954",
  1590 => x"73802eff",
  1591 => x"b2388215",
  1592 => x"2253ffae",
  1593 => x"39742253",
  1594 => x"fcb33974",
  1595 => x"22547390",
  1596 => x"2b70902c",
  1597 => x"719f2c70",
  1598 => x"72327131",
  1599 => x"799f2c70",
  1600 => x"7b327131",
  1601 => x"51545156",
  1602 => x"56537274",
  1603 => x"25833874",
  1604 => x"56811970",
  1605 => x"81ff065a",
  1606 => x"55787a27",
  1607 => x"fddb3877",
  1608 => x"83ffff06",
  1609 => x"81197110",
  1610 => x"10880a05",
  1611 => x"79307a82",
  1612 => x"32703072",
  1613 => x"80257180",
  1614 => x"25075351",
  1615 => x"57535759",
  1616 => x"5473802e",
  1617 => x"ffa53882",
  1618 => x"152254ff",
  1619 => x"a1398170",
  1620 => x"902b7090",
  1621 => x"2c405754",
  1622 => x"80705d58",
  1623 => x"fcae3974",
  1624 => x"2254fce4",
  1625 => x"39fa3d0d",
  1626 => x"8a51bb8e",
  1627 => x"3f978f3f",
  1628 => x"99d95381",
  1629 => x"aa805281",
  1630 => x"aa945197",
  1631 => x"943fa3c3",
  1632 => x"5381aa98",
  1633 => x"5281aac0",
  1634 => x"5197863f",
  1635 => x"bb895381",
  1636 => x"aac85281",
  1637 => x"aad85196",
  1638 => x"f83fa5fd",
  1639 => x"5381aae0",
  1640 => x"5281ab84",
  1641 => x"5196ea3f",
  1642 => x"bdcc5381",
  1643 => x"ab8c5281",
  1644 => x"abac5196",
  1645 => x"dc3fbeea",
  1646 => x"5381abb0",
  1647 => x"5281abd4",
  1648 => x"5196ce3f",
  1649 => x"bba05381",
  1650 => x"abdc5281",
  1651 => x"a7985196",
  1652 => x"c03fbbe1",
  1653 => x"5381ac80",
  1654 => x"5281aca8",
  1655 => x"5196b23f",
  1656 => x"bd895381",
  1657 => x"acb05281",
  1658 => x"acd05196",
  1659 => x"a43f889b",
  1660 => x"5381acd8",
  1661 => x"5281acf4",
  1662 => x"5196963f",
  1663 => x"a4935381",
  1664 => x"acfc5281",
  1665 => x"acc85196",
  1666 => x"883fa3df",
  1667 => x"5381ad98",
  1668 => x"5281adac",
  1669 => x"5195fa3f",
  1670 => x"b8c85381",
  1671 => x"adb45281",
  1672 => x"add05195",
  1673 => x"ec3fb8ee",
  1674 => x"5381add8",
  1675 => x"5281adec",
  1676 => x"5195de3f",
  1677 => x"a79f5381",
  1678 => x"adf45281",
  1679 => x"ae985195",
  1680 => x"d03fbfc8",
  1681 => x"5381aea0",
  1682 => x"5281aeb0",
  1683 => x"5195c23f",
  1684 => x"80c29353",
  1685 => x"81aeb452",
  1686 => x"81aed051",
  1687 => x"95b33fba",
  1688 => x"cf5381ae",
  1689 => x"d85281ae",
  1690 => x"f05195a5",
  1691 => x"3f80c29b",
  1692 => x"5381aef8",
  1693 => x"5281af8c",
  1694 => x"5195963f",
  1695 => x"8ad65381",
  1696 => x"af945281",
  1697 => x"afa85195",
  1698 => x"883f8de6",
  1699 => x"5381afac",
  1700 => x"5281afd4",
  1701 => x"5194fa3f",
  1702 => x"baeb5381",
  1703 => x"afdc5281",
  1704 => x"affc5194",
  1705 => x"ec3f93a2",
  1706 => x"5381b084",
  1707 => x"5281b098",
  1708 => x"5194de3f",
  1709 => x"88be5381",
  1710 => x"b0a05281",
  1711 => x"b0ac5194",
  1712 => x"d03f89fc",
  1713 => x"5381b0b0",
  1714 => x"5281b0d8",
  1715 => x"5194c23f",
  1716 => x"88be5381",
  1717 => x"b0e05281",
  1718 => x"a9b85194",
  1719 => x"b43f8ac5",
  1720 => x"5381b180",
  1721 => x"5281b190",
  1722 => x"5194a63f",
  1723 => x"88b35381",
  1724 => x"9cc45281",
  1725 => x"9ca45194",
  1726 => x"983f80d0",
  1727 => x"e753819c",
  1728 => x"c452819c",
  1729 => x"ac519489",
  1730 => x"3f9adc3f",
  1731 => x"94cf3f81",
  1732 => x"0b81e2e0",
  1733 => x"3481cfc0",
  1734 => x"337081ff",
  1735 => x"06555573",
  1736 => x"b038bbe2",
  1737 => x"3fb00890",
  1738 => x"3894c03f",
  1739 => x"81e2e033",
  1740 => x"5675e238",
  1741 => x"883d0d04",
  1742 => x"bbdf3fb0",
  1743 => x"0881ff06",
  1744 => x"5195963f",
  1745 => x"94a53f81",
  1746 => x"e2e03356",
  1747 => x"75c738e4",
  1748 => x"39800b81",
  1749 => x"cfc0349b",
  1750 => x"ae3f81bf",
  1751 => x"e4087008",
  1752 => x"70872a81",
  1753 => x"06525754",
  1754 => x"73802e8f",
  1755 => x"3876802e",
  1756 => x"81c338ff",
  1757 => x"177081ff",
  1758 => x"06585475",
  1759 => x"862a8106",
  1760 => x"5574802e",
  1761 => x"aa387680",
  1762 => x"f6388196",
  1763 => x"0b81bfe4",
  1764 => x"08841108",
  1765 => x"70efff0a",
  1766 => x"06ae800a",
  1767 => x"0784130c",
  1768 => x"57841108",
  1769 => x"70be800a",
  1770 => x"0784130c",
  1771 => x"57555775",
  1772 => x"852a8106",
  1773 => x"5574802e",
  1774 => x"963876b9",
  1775 => x"3881960b",
  1776 => x"81bfac08",
  1777 => x"b8110857",
  1778 => x"5557800b",
  1779 => x"b8150c75",
  1780 => x"842a8106",
  1781 => x"5675802e",
  1782 => x"fec83876",
  1783 => x"802eab38",
  1784 => x"ff177081",
  1785 => x"ff065855",
  1786 => x"ba9c3fb0",
  1787 => x"08802efe",
  1788 => x"b838fec4",
  1789 => x"39ff1770",
  1790 => x"81ff0658",
  1791 => x"55d139ff",
  1792 => x"177081ff",
  1793 => x"065854ff",
  1794 => x"a6398196",
  1795 => x"0b81bfe4",
  1796 => x"08841108",
  1797 => x"840a0784",
  1798 => x"120c5657",
  1799 => x"9e973f80",
  1800 => x"5281b484",
  1801 => x"51a0e13f",
  1802 => x"b9dc3fb0",
  1803 => x"08802efd",
  1804 => x"f838fe84",
  1805 => x"39819676",
  1806 => x"822a8306",
  1807 => x"53768306",
  1808 => x"5257f4ef",
  1809 => x"3ffeb439",
  1810 => x"fe3d0d81",
  1811 => x"5195b43f",
  1812 => x"b00881ff",
  1813 => x"06538251",
  1814 => x"95a93fb0",
  1815 => x"0881ff06",
  1816 => x"527251f4",
  1817 => x"ce3f800b",
  1818 => x"b00c843d",
  1819 => x"0d04f93d",
  1820 => x"0d815195",
  1821 => x"8e3fb008",
  1822 => x"81ff0681",
  1823 => x"b1985257",
  1824 => x"b5923f81",
  1825 => x"b1ac51b5",
  1826 => x"8b3ff880",
  1827 => x"809a8054",
  1828 => x"80557370",
  1829 => x"84055508",
  1830 => x"74708405",
  1831 => x"56085456",
  1832 => x"72a03881",
  1833 => x"157081ff",
  1834 => x"06565687",
  1835 => x"7527e338",
  1836 => x"76812e80",
  1837 => x"d8388a51",
  1838 => x"b4c03f76",
  1839 => x"b00c893d",
  1840 => x"0d048a51",
  1841 => x"b4b43f72",
  1842 => x"51b6933f",
  1843 => x"b00881ff",
  1844 => x"0653728c",
  1845 => x"279338a0",
  1846 => x"51b49f3f",
  1847 => x"81137081",
  1848 => x"ff065153",
  1849 => x"8c7326ef",
  1850 => x"3881b1c4",
  1851 => x"51b4a53f",
  1852 => x"7552a051",
  1853 => x"b4c13f75",
  1854 => x"51d9de3f",
  1855 => x"81157081",
  1856 => x"ff065656",
  1857 => x"877527ff",
  1858 => x"8938ffa4",
  1859 => x"39f88080",
  1860 => x"9a805480",
  1861 => x"53807470",
  1862 => x"8405560c",
  1863 => x"80747084",
  1864 => x"05560c81",
  1865 => x"137081ff",
  1866 => x"06545572",
  1867 => x"8726ff86",
  1868 => x"38807470",
  1869 => x"8405560c",
  1870 => x"80747084",
  1871 => x"05560c81",
  1872 => x"137081ff",
  1873 => x"06545587",
  1874 => x"7327ca38",
  1875 => x"fee839fe",
  1876 => x"3d0d8151",
  1877 => x"93ad3fb0",
  1878 => x"0881ff06",
  1879 => x"81bfa408",
  1880 => x"7188120c",
  1881 => x"53b00c84",
  1882 => x"3d0d0480",
  1883 => x"3d0d8151",
  1884 => x"94c33fb0",
  1885 => x"0883ffff",
  1886 => x"0651d3b6",
  1887 => x"3fb00883",
  1888 => x"ffff06b0",
  1889 => x"0c823d0d",
  1890 => x"04803d0d",
  1891 => x"81bff008",
  1892 => x"51f8bb95",
  1893 => x"86a1710c",
  1894 => x"810bb00c",
  1895 => x"823d0d04",
  1896 => x"fc3d0d81",
  1897 => x"5192dc3f",
  1898 => x"b00881ff",
  1899 => x"06548251",
  1900 => x"92d13fb0",
  1901 => x"0881ff06",
  1902 => x"81bfe408",
  1903 => x"84110870",
  1904 => x"fe8f0a06",
  1905 => x"77982b07",
  1906 => x"51545653",
  1907 => x"72802e86",
  1908 => x"3871810a",
  1909 => x"07527184",
  1910 => x"160c71b0",
  1911 => x"0c863d0d",
  1912 => x"04fd3d0d",
  1913 => x"81bfe408",
  1914 => x"84110855",
  1915 => x"53815192",
  1916 => x"923fb008",
  1917 => x"81ff0674",
  1918 => x"dfffff06",
  1919 => x"54527180",
  1920 => x"2e873873",
  1921 => x"a0808007",
  1922 => x"53825191",
  1923 => x"f63fb008",
  1924 => x"81ff0673",
  1925 => x"efff0a06",
  1926 => x"55527180",
  1927 => x"2e873872",
  1928 => x"90800a07",
  1929 => x"54835191",
  1930 => x"da3fb008",
  1931 => x"81ff0674",
  1932 => x"f7ff0a06",
  1933 => x"54527180",
  1934 => x"2e873873",
  1935 => x"88800a07",
  1936 => x"53845191",
  1937 => x"be3fb008",
  1938 => x"81ff0673",
  1939 => x"fbff0a06",
  1940 => x"55527180",
  1941 => x"2e873872",
  1942 => x"84800a07",
  1943 => x"54855191",
  1944 => x"a23fb008",
  1945 => x"81ff0674",
  1946 => x"fdff0a06",
  1947 => x"54527180",
  1948 => x"2e873873",
  1949 => x"82800a07",
  1950 => x"5381bfe4",
  1951 => x"08738412",
  1952 => x"0c5472b0",
  1953 => x"0c853d0d",
  1954 => x"04fa3d0d",
  1955 => x"880a0b81",
  1956 => x"bfa8088c",
  1957 => x"11085955",
  1958 => x"56815190",
  1959 => x"e63fb008",
  1960 => x"902b7090",
  1961 => x"2c565380",
  1962 => x"77279938",
  1963 => x"80775454",
  1964 => x"7383ffff",
  1965 => x"06767084",
  1966 => x"05580cff",
  1967 => x"13751555",
  1968 => x"5372ed38",
  1969 => x"800bb00c",
  1970 => x"883d0d04",
  1971 => x"fc3d0d81",
  1972 => x"b1cc51b0",
  1973 => x"bf3f81bf",
  1974 => x"e4087008",
  1975 => x"709e2a70",
  1976 => x"81065154",
  1977 => x"54548153",
  1978 => x"71833871",
  1979 => x"5372802e",
  1980 => x"80d23881",
  1981 => x"b1dc51b0",
  1982 => x"9b3f8151",
  1983 => x"90853fb0",
  1984 => x"0881ff06",
  1985 => x"81b1cc52",
  1986 => x"55b0893f",
  1987 => x"74802eab",
  1988 => x"3881b1e4",
  1989 => x"51affd3f",
  1990 => x"81bfe408",
  1991 => x"84110870",
  1992 => x"fd0a0654",
  1993 => x"54547480",
  1994 => x"2e863872",
  1995 => x"820a0752",
  1996 => x"7184150c",
  1997 => x"71b00c86",
  1998 => x"3d0d0481",
  1999 => x"a7a051af",
  2000 => x"d33fce39",
  2001 => x"81a7a051",
  2002 => x"afca3f81",
  2003 => x"b1dc51af",
  2004 => x"c33f8151",
  2005 => x"8fad3fb0",
  2006 => x"0881ff06",
  2007 => x"81b1cc52",
  2008 => x"55afb13f",
  2009 => x"74ffaa38",
  2010 => x"d239fd3d",
  2011 => x"0d81518f",
  2012 => x"923fb008",
  2013 => x"81ff0681",
  2014 => x"b1f05254",
  2015 => x"af963f73",
  2016 => x"a43881a7",
  2017 => x"9851af8c",
  2018 => x"3f81bfe4",
  2019 => x"08841108",
  2020 => x"70fb0a06",
  2021 => x"84130c53",
  2022 => x"538a51ae",
  2023 => x"dd3f73b0",
  2024 => x"0c853d0d",
  2025 => x"0481a3c0",
  2026 => x"51aee93f",
  2027 => x"81bfe408",
  2028 => x"84110870",
  2029 => x"840a0784",
  2030 => x"130c5353",
  2031 => x"8a51aeba",
  2032 => x"3f73b00c",
  2033 => x"853d0d04",
  2034 => x"fd3d0d81",
  2035 => x"cfbc0852",
  2036 => x"f881c08e",
  2037 => x"800b81bf",
  2038 => x"e4085553",
  2039 => x"71802e80",
  2040 => x"f7387281",
  2041 => x"ff068415",
  2042 => x"0c81bfa0",
  2043 => x"337081ff",
  2044 => x"06515271",
  2045 => x"802e80c2",
  2046 => x"38729f2a",
  2047 => x"73100753",
  2048 => x"81cfc033",
  2049 => x"7081ff06",
  2050 => x"51527180",
  2051 => x"2ed43880",
  2052 => x"0b81cfc0",
  2053 => x"3491f03f",
  2054 => x"81bfb033",
  2055 => x"547380e2",
  2056 => x"3881bfe4",
  2057 => x"087381ff",
  2058 => x"0684120c",
  2059 => x"81bfa033",
  2060 => x"7081ff06",
  2061 => x"51535471",
  2062 => x"c0387281",
  2063 => x"2a739f2b",
  2064 => x"0753ffbc",
  2065 => x"3972812a",
  2066 => x"739f2b07",
  2067 => x"5380fd51",
  2068 => x"b0d53f81",
  2069 => x"bfe40854",
  2070 => x"7281ff06",
  2071 => x"84150c81",
  2072 => x"bfa03370",
  2073 => x"81ff0653",
  2074 => x"5471802e",
  2075 => x"d838729f",
  2076 => x"2a731007",
  2077 => x"5380fd51",
  2078 => x"b0ad3f81",
  2079 => x"bfe40854",
  2080 => x"d739800b",
  2081 => x"b00c853d",
  2082 => x"0d04f73d",
  2083 => x"0d853d54",
  2084 => x"965381b2",
  2085 => x"84527351",
  2086 => x"b3cb3f96",
  2087 => x"893f8151",
  2088 => x"8ce13f80",
  2089 => x"52805193",
  2090 => x"e93f7353",
  2091 => x"805281b4",
  2092 => x"8451a8a8",
  2093 => x"3f805281",
  2094 => x"5193d73f",
  2095 => x"73538252",
  2096 => x"81b48451",
  2097 => x"a8963f80",
  2098 => x"52825193",
  2099 => x"c53f7353",
  2100 => x"815281b4",
  2101 => x"8451a884",
  2102 => x"3f805284",
  2103 => x"5193b33f",
  2104 => x"73538452",
  2105 => x"81b48451",
  2106 => x"a7f23f80",
  2107 => x"52855193",
  2108 => x"a13f7353",
  2109 => x"905281b4",
  2110 => x"8451a7e0",
  2111 => x"3f805286",
  2112 => x"51938f3f",
  2113 => x"73538352",
  2114 => x"81b48451",
  2115 => x"a7ce3f8b",
  2116 => x"3d0d04fe",
  2117 => x"f53f800b",
  2118 => x"b00c04fc",
  2119 => x"3d0d8196",
  2120 => x"bc548055",
  2121 => x"84527451",
  2122 => x"92e83f80",
  2123 => x"53737081",
  2124 => x"05553351",
  2125 => x"93e23f81",
  2126 => x"137081ff",
  2127 => x"06515380",
  2128 => x"dc7327e9",
  2129 => x"38811570",
  2130 => x"81ff0656",
  2131 => x"53877527",
  2132 => x"d338800b",
  2133 => x"b00c863d",
  2134 => x"0d04fd3d",
  2135 => x"0d81bfa0",
  2136 => x"337081ff",
  2137 => x"06545472",
  2138 => x"bf26ac38",
  2139 => x"81bfa033",
  2140 => x"7081ff06",
  2141 => x"81bfa408",
  2142 => x"5288120c",
  2143 => x"5480e452",
  2144 => x"80c2da51",
  2145 => x"8fe13f81",
  2146 => x"bfa03381",
  2147 => x"05537281",
  2148 => x"bfa03485",
  2149 => x"3d0d0480",
  2150 => x"e45280c3",
  2151 => x"b1518fc7",
  2152 => x"3f81bfa0",
  2153 => x"33810553",
  2154 => x"7281bfa0",
  2155 => x"34853d0d",
  2156 => x"04fd3d0d",
  2157 => x"81bfa033",
  2158 => x"7081ff06",
  2159 => x"545472bf",
  2160 => x"2680c938",
  2161 => x"81bfa033",
  2162 => x"7081ff06",
  2163 => x"81bfa408",
  2164 => x"5688160c",
  2165 => x"5381bfa0",
  2166 => x"337081ff",
  2167 => x"06555373",
  2168 => x"bf2e80d1",
  2169 => x"3880e452",
  2170 => x"80c3b151",
  2171 => x"8ef93f81",
  2172 => x"bfa03381",
  2173 => x"05537281",
  2174 => x"bfa03481",
  2175 => x"bfa03380",
  2176 => x"ff065372",
  2177 => x"81bfa034",
  2178 => x"853d0d04",
  2179 => x"81bfa033",
  2180 => x"7081ff06",
  2181 => x"80ff7131",
  2182 => x"81bfa408",
  2183 => x"5288120c",
  2184 => x"555381bf",
  2185 => x"a0337081",
  2186 => x"ff065553",
  2187 => x"73bf2e09",
  2188 => x"8106ffb1",
  2189 => x"3880ce90",
  2190 => x"5280c3b1",
  2191 => x"518ea83f",
  2192 => x"81bfa033",
  2193 => x"81055372",
  2194 => x"81bfa034",
  2195 => x"81bfa033",
  2196 => x"80ff0653",
  2197 => x"7281bfa0",
  2198 => x"34853d0d",
  2199 => x"04810b81",
  2200 => x"bfb03404",
  2201 => x"fe3d0d81",
  2202 => x"bfe80898",
  2203 => x"11087084",
  2204 => x"2a708106",
  2205 => x"51535353",
  2206 => x"70802e8d",
  2207 => x"3871ef06",
  2208 => x"98140c81",
  2209 => x"0b81cfc0",
  2210 => x"34843d0d",
  2211 => x"04fb3d0d",
  2212 => x"81bfe408",
  2213 => x"7008810a",
  2214 => x"0681cfbc",
  2215 => x"0c54acaa",
  2216 => x"3faccd3f",
  2217 => x"8efe3f81",
  2218 => x"bfe80898",
  2219 => x"11088807",
  2220 => x"98120c54",
  2221 => x"81cfbc08",
  2222 => x"80ede455",
  2223 => x"53728438",
  2224 => x"88805473",
  2225 => x"81e3c40c",
  2226 => x"72802e84",
  2227 => x"a338819d",
  2228 => x"8c51a8c0",
  2229 => x"3f8c51a8",
  2230 => x"a13f81b2",
  2231 => x"8451a8b4",
  2232 => x"3f81cfbc",
  2233 => x"08802e81",
  2234 => x"db3881b2",
  2235 => x"9c51a8a4",
  2236 => x"3f81cfbc",
  2237 => x"08547380",
  2238 => x"2e82c638",
  2239 => x"81bfa808",
  2240 => x"5481740c",
  2241 => x"81bfe408",
  2242 => x"84110870",
  2243 => x"56575580",
  2244 => x"5373fe8f",
  2245 => x"0a067398",
  2246 => x"2b077084",
  2247 => x"170c8114",
  2248 => x"7081ff06",
  2249 => x"5154548f",
  2250 => x"7327e638",
  2251 => x"7584160c",
  2252 => x"81bfac08",
  2253 => x"54800bb8",
  2254 => x"150ca080",
  2255 => x"870a0851",
  2256 => x"a99c3f82",
  2257 => x"5280c4dd",
  2258 => x"518c9c3f",
  2259 => x"f881c08e",
  2260 => x"800b81bf",
  2261 => x"e4085654",
  2262 => x"81cfbc08",
  2263 => x"802e81b7",
  2264 => x"387381ff",
  2265 => x"0684160c",
  2266 => x"81bfa033",
  2267 => x"7081ff06",
  2268 => x"54567280",
  2269 => x"2e80c238",
  2270 => x"739f2a74",
  2271 => x"10075481",
  2272 => x"cfc03370",
  2273 => x"81ff0657",
  2274 => x"5375802e",
  2275 => x"d438800b",
  2276 => x"81cfc034",
  2277 => x"8af13f81",
  2278 => x"bfb03355",
  2279 => x"7482dc38",
  2280 => x"81bfe408",
  2281 => x"7481ff06",
  2282 => x"84120c81",
  2283 => x"bfa03370",
  2284 => x"81ff0655",
  2285 => x"575572c0",
  2286 => x"3873812a",
  2287 => x"749f2b07",
  2288 => x"54ffbc39",
  2289 => x"81b2a851",
  2290 => x"a6ca3f81",
  2291 => x"0a51a6c4",
  2292 => x"3f81b2bc",
  2293 => x"51a6bd3f",
  2294 => x"81b2e451",
  2295 => x"a6b63fb4",
  2296 => x"51a7fb3f",
  2297 => x"81b2f851",
  2298 => x"a6aa3f81",
  2299 => x"b38051a6",
  2300 => x"a33f81b3",
  2301 => x"8c51a69c",
  2302 => x"3f81cfbc",
  2303 => x"085473fd",
  2304 => x"fb38be39",
  2305 => x"73812a74",
  2306 => x"9f2b0754",
  2307 => x"80fd51a9",
  2308 => x"963f81bf",
  2309 => x"e4085573",
  2310 => x"81ff0684",
  2311 => x"160c81bf",
  2312 => x"a0337081",
  2313 => x"ff065656",
  2314 => x"74802ed8",
  2315 => x"38739f2a",
  2316 => x"74100754",
  2317 => x"80fd51a8",
  2318 => x"ee3f81bf",
  2319 => x"e40855d7",
  2320 => x"3981bfac",
  2321 => x"0874b412",
  2322 => x"0c568180",
  2323 => x"51c5e33f",
  2324 => x"828051c5",
  2325 => x"dd3f8483",
  2326 => x"51c5d73f",
  2327 => x"86f151c5",
  2328 => x"d13f8883",
  2329 => x"51c5cb3f",
  2330 => x"81bfe408",
  2331 => x"7008709e",
  2332 => x"2a708106",
  2333 => x"51555654",
  2334 => x"81557280",
  2335 => x"2e80f738",
  2336 => x"7481ff06",
  2337 => x"84150870",
  2338 => x"fd0a0658",
  2339 => x"56537280",
  2340 => x"2e863874",
  2341 => x"820a0756",
  2342 => x"7584150c",
  2343 => x"841408be",
  2344 => x"800a0784",
  2345 => x"150c8414",
  2346 => x"08840a07",
  2347 => x"84150c81",
  2348 => x"bfac0855",
  2349 => x"800bb816",
  2350 => x"0c81bfa8",
  2351 => x"08548174",
  2352 => x"0c93c452",
  2353 => x"80c29b51",
  2354 => x"899d3f87",
  2355 => x"e85280c2",
  2356 => x"da518993",
  2357 => x"3fe98e3f",
  2358 => x"81bfa808",
  2359 => x"5481740c",
  2360 => x"81bfe408",
  2361 => x"84110870",
  2362 => x"56575580",
  2363 => x"53fca239",
  2364 => x"8db43ffb",
  2365 => x"d9397255",
  2366 => x"ff8639aa",
  2367 => x"db3f800b",
  2368 => x"81e2d834",
  2369 => x"800b81e2",
  2370 => x"d434800b",
  2371 => x"81e2dc0c",
  2372 => x"04fc3d0d",
  2373 => x"765281e2",
  2374 => x"d4337010",
  2375 => x"10107110",
  2376 => x"0581cfc4",
  2377 => x"055254af",
  2378 => x"ca3f7752",
  2379 => x"81e2d433",
  2380 => x"70902971",
  2381 => x"31701010",
  2382 => x"81d28405",
  2383 => x"535555af",
  2384 => x"b23f81e2",
  2385 => x"d4337010",
  2386 => x"1081e184",
  2387 => x"057a710c",
  2388 => x"54810553",
  2389 => x"7281e2d4",
  2390 => x"34863d0d",
  2391 => x"04803d0d",
  2392 => x"81b3d051",
  2393 => x"a3ae3f82",
  2394 => x"3d0d04fe",
  2395 => x"3d0d81e2",
  2396 => x"dc085372",
  2397 => x"8538843d",
  2398 => x"0d04722d",
  2399 => x"b0085380",
  2400 => x"0b81e2dc",
  2401 => x"0cb0088c",
  2402 => x"3881b3d0",
  2403 => x"51a3853f",
  2404 => x"843d0d04",
  2405 => x"819cb451",
  2406 => x"a2fa3f72",
  2407 => x"83ffff26",
  2408 => x"aa3881ff",
  2409 => x"73279638",
  2410 => x"72529051",
  2411 => x"a3893f8a",
  2412 => x"51a2c73f",
  2413 => x"81b3d051",
  2414 => x"a2da3fd4",
  2415 => x"39725288",
  2416 => x"51a2f43f",
  2417 => x"8a51a2b2",
  2418 => x"3fea3972",
  2419 => x"52a051a2",
  2420 => x"e63f8a51",
  2421 => x"a2a43fdc",
  2422 => x"39fa3d0d",
  2423 => x"02a30533",
  2424 => x"56758d2e",
  2425 => x"80f43875",
  2426 => x"88327030",
  2427 => x"7780ff32",
  2428 => x"70307280",
  2429 => x"25718025",
  2430 => x"07545156",
  2431 => x"58557495",
  2432 => x"389f7627",
  2433 => x"8c3881e2",
  2434 => x"d8335580",
  2435 => x"ce7527ae",
  2436 => x"38883d0d",
  2437 => x"0481e2d8",
  2438 => x"33567580",
  2439 => x"2ef33888",
  2440 => x"51a1d73f",
  2441 => x"a051a1d2",
  2442 => x"3f8851a1",
  2443 => x"cd3f81e2",
  2444 => x"d833ff05",
  2445 => x"577681e2",
  2446 => x"d834883d",
  2447 => x"0d047551",
  2448 => x"a1b83f81",
  2449 => x"e2d83381",
  2450 => x"11555773",
  2451 => x"81e2d834",
  2452 => x"7581e284",
  2453 => x"1834883d",
  2454 => x"0d048a51",
  2455 => x"a19c3f81",
  2456 => x"e2d83381",
  2457 => x"11565474",
  2458 => x"81e2d834",
  2459 => x"800b81e2",
  2460 => x"84153480",
  2461 => x"56800b81",
  2462 => x"e2841733",
  2463 => x"565474a0",
  2464 => x"2e833881",
  2465 => x"5474802e",
  2466 => x"90387380",
  2467 => x"2e8b3881",
  2468 => x"167081ff",
  2469 => x"065757dd",
  2470 => x"3975802e",
  2471 => x"bf38800b",
  2472 => x"81e2d433",
  2473 => x"55557474",
  2474 => x"27ab3873",
  2475 => x"57741010",
  2476 => x"10751005",
  2477 => x"765481e2",
  2478 => x"845381cf",
  2479 => x"c40551ad",
  2480 => x"fe3fb008",
  2481 => x"802ea638",
  2482 => x"81157081",
  2483 => x"ff065654",
  2484 => x"767526d9",
  2485 => x"3881b3d4",
  2486 => x"51a0b93f",
  2487 => x"81b3d051",
  2488 => x"a0b23f80",
  2489 => x"0b81e2d8",
  2490 => x"34883d0d",
  2491 => x"04741010",
  2492 => x"81e18405",
  2493 => x"700881e2",
  2494 => x"dc0c5680",
  2495 => x"0b81e2d8",
  2496 => x"34e739f7",
  2497 => x"3d0d02af",
  2498 => x"05335980",
  2499 => x"0b81e284",
  2500 => x"3381e284",
  2501 => x"59555673",
  2502 => x"a02e0981",
  2503 => x"06963881",
  2504 => x"167081ff",
  2505 => x"0681e284",
  2506 => x"11703353",
  2507 => x"59575473",
  2508 => x"a02eec38",
  2509 => x"80587779",
  2510 => x"2780ea38",
  2511 => x"80773356",
  2512 => x"5474742e",
  2513 => x"83388154",
  2514 => x"74a02e9a",
  2515 => x"387380c5",
  2516 => x"3874a02e",
  2517 => x"91388118",
  2518 => x"7081ff06",
  2519 => x"59557878",
  2520 => x"26da3880",
  2521 => x"c0398116",
  2522 => x"7081ff06",
  2523 => x"81e28411",
  2524 => x"70335752",
  2525 => x"575773a0",
  2526 => x"2e098106",
  2527 => x"d9388116",
  2528 => x"7081ff06",
  2529 => x"81e28411",
  2530 => x"70335752",
  2531 => x"575773a0",
  2532 => x"2ed438c2",
  2533 => x"39811670",
  2534 => x"81ff0681",
  2535 => x"e2841159",
  2536 => x"5755ff98",
  2537 => x"398a538b",
  2538 => x"3dfc0552",
  2539 => x"7651b0d4",
  2540 => x"3f8b3d0d",
  2541 => x"04f73d0d",
  2542 => x"02af0533",
  2543 => x"59800b81",
  2544 => x"e2843381",
  2545 => x"e2845955",
  2546 => x"5673a02e",
  2547 => x"09810696",
  2548 => x"38811670",
  2549 => x"81ff0681",
  2550 => x"e2841170",
  2551 => x"33535957",
  2552 => x"5473a02e",
  2553 => x"ec388058",
  2554 => x"77792780",
  2555 => x"ea388077",
  2556 => x"33565474",
  2557 => x"742e8338",
  2558 => x"815474a0",
  2559 => x"2e9a3873",
  2560 => x"80c53874",
  2561 => x"a02e9138",
  2562 => x"81187081",
  2563 => x"ff065955",
  2564 => x"787826da",
  2565 => x"3880c039",
  2566 => x"81167081",
  2567 => x"ff0681e2",
  2568 => x"84117033",
  2569 => x"57525757",
  2570 => x"73a02e09",
  2571 => x"8106d938",
  2572 => x"81167081",
  2573 => x"ff0681e2",
  2574 => x"84117033",
  2575 => x"57525757",
  2576 => x"73a02ed4",
  2577 => x"38c23981",
  2578 => x"167081ff",
  2579 => x"0681e284",
  2580 => x"11595755",
  2581 => x"ff983990",
  2582 => x"538b3dfc",
  2583 => x"05527651",
  2584 => x"b2bf3f8b",
  2585 => x"3d0d04fc",
  2586 => x"3d0d8a51",
  2587 => x"9d8c3f81",
  2588 => x"b3e8519d",
  2589 => x"9f3f800b",
  2590 => x"81e2d433",
  2591 => x"53537272",
  2592 => x"2780f538",
  2593 => x"72101010",
  2594 => x"73100581",
  2595 => x"cfc40570",
  2596 => x"52549d80",
  2597 => x"3f72842b",
  2598 => x"70743182",
  2599 => x"2b81d284",
  2600 => x"11335153",
  2601 => x"5571802e",
  2602 => x"b7387351",
  2603 => x"a9b23fb0",
  2604 => x"0881ff06",
  2605 => x"52718926",
  2606 => x"9338a051",
  2607 => x"9cbc3f81",
  2608 => x"127081ff",
  2609 => x"06535489",
  2610 => x"7227ef38",
  2611 => x"81b48051",
  2612 => x"9cc23f74",
  2613 => x"7331822b",
  2614 => x"81d28405",
  2615 => x"519cb53f",
  2616 => x"8a519c96",
  2617 => x"3f811370",
  2618 => x"81ff0681",
  2619 => x"e2d43354",
  2620 => x"54557173",
  2621 => x"26ff8d38",
  2622 => x"8a519bfe",
  2623 => x"3f81e2d4",
  2624 => x"33b00c86",
  2625 => x"3d0d04fe",
  2626 => x"3d0d81e3",
  2627 => x"b422ff05",
  2628 => x"517081e3",
  2629 => x"b4237083",
  2630 => x"ffff0651",
  2631 => x"7080c438",
  2632 => x"81e3b833",
  2633 => x"517081ff",
  2634 => x"2eb93870",
  2635 => x"10101081",
  2636 => x"e2e40552",
  2637 => x"713381e3",
  2638 => x"b834fe72",
  2639 => x"3481e3b8",
  2640 => x"33701010",
  2641 => x"1081e2e4",
  2642 => x"05525382",
  2643 => x"112281e3",
  2644 => x"b4238412",
  2645 => x"0853722d",
  2646 => x"81e3b422",
  2647 => x"5170802e",
  2648 => x"ffbe3884",
  2649 => x"3d0d04f9",
  2650 => x"3d0d02aa",
  2651 => x"05225680",
  2652 => x"55741010",
  2653 => x"1081e2e4",
  2654 => x"05703352",
  2655 => x"527081fe",
  2656 => x"2e993881",
  2657 => x"157081ff",
  2658 => x"06565274",
  2659 => x"8a2e0981",
  2660 => x"06df3881",
  2661 => x"0bb00c89",
  2662 => x"3d0d0481",
  2663 => x"e3b83370",
  2664 => x"81ff0681",
  2665 => x"e3b42253",
  2666 => x"54587281",
  2667 => x"ff2eb038",
  2668 => x"72832b54",
  2669 => x"70762780",
  2670 => x"de387571",
  2671 => x"317083ff",
  2672 => x"ff067481",
  2673 => x"e2e41733",
  2674 => x"70832b81",
  2675 => x"e2e61122",
  2676 => x"56585652",
  2677 => x"57577281",
  2678 => x"ff2e0981",
  2679 => x"06d63872",
  2680 => x"72347582",
  2681 => x"13237984",
  2682 => x"130c7781",
  2683 => x"ff065473",
  2684 => x"732e9638",
  2685 => x"76101010",
  2686 => x"81e2e405",
  2687 => x"53747334",
  2688 => x"805170b0",
  2689 => x"0c893d0d",
  2690 => x"047481e3",
  2691 => x"b8347581",
  2692 => x"e3b42380",
  2693 => x"51ec3970",
  2694 => x"76315170",
  2695 => x"81e2e615",
  2696 => x"23ffbc39",
  2697 => x"ff3d0d8a",
  2698 => x"52711010",
  2699 => x"1081e2dc",
  2700 => x"0551fe71",
  2701 => x"34ff1270",
  2702 => x"81ff0653",
  2703 => x"5171ea38",
  2704 => x"ff0b81e3",
  2705 => x"b834833d",
  2706 => x"0d04fe3d",
  2707 => x"0d740284",
  2708 => x"05970533",
  2709 => x"0288059b",
  2710 => x"05338813",
  2711 => x"0c8c120c",
  2712 => x"538c1308",
  2713 => x"70812a81",
  2714 => x"06515271",
  2715 => x"f4388c13",
  2716 => x"087081ff",
  2717 => x"06b00c51",
  2718 => x"843d0d04",
  2719 => x"803d0d72",
  2720 => x"8c110870",
  2721 => x"872a8132",
  2722 => x"8106b00c",
  2723 => x"5151823d",
  2724 => x"0d04fd3d",
  2725 => x"0d029705",
  2726 => x"33028405",
  2727 => x"9b053371",
  2728 => x"81b00781",
  2729 => x"bf065354",
  2730 => x"54f88080",
  2731 => x"98807171",
  2732 => x"0c73842a",
  2733 => x"9007710c",
  2734 => x"738f0671",
  2735 => x"0c527281",
  2736 => x"bfb83473",
  2737 => x"81bfbc34",
  2738 => x"853d0d04",
  2739 => x"fd3d0d02",
  2740 => x"97053381",
  2741 => x"bfbc3354",
  2742 => x"73058706",
  2743 => x"0284059a",
  2744 => x"052281bf",
  2745 => x"b8335473",
  2746 => x"057081ff",
  2747 => x"067281b0",
  2748 => x"07545154",
  2749 => x"54f88080",
  2750 => x"98807171",
  2751 => x"0c73842a",
  2752 => x"9007710c",
  2753 => x"738f0671",
  2754 => x"0c527281",
  2755 => x"bfb83473",
  2756 => x"81bfbc34",
  2757 => x"853d0d04",
  2758 => x"ff3d0d02",
  2759 => x"8f0533f8",
  2760 => x"80809884",
  2761 => x"0c81bfb8",
  2762 => x"33810551",
  2763 => x"7081bfb8",
  2764 => x"34833d0d",
  2765 => x"04ff3d0d",
  2766 => x"80527181",
  2767 => x"b00781bf",
  2768 => x"06f88080",
  2769 => x"98800c90",
  2770 => x"0bf88080",
  2771 => x"98800c80",
  2772 => x"0bf88080",
  2773 => x"98800c80",
  2774 => x"51800bf8",
  2775 => x"80809884",
  2776 => x"0c811170",
  2777 => x"81ff0651",
  2778 => x"5180e571",
  2779 => x"27eb3881",
  2780 => x"127081ff",
  2781 => x"06535187",
  2782 => x"7227ffbe",
  2783 => x"3881b00b",
  2784 => x"f8808098",
  2785 => x"800c900b",
  2786 => x"f8808098",
  2787 => x"800c800b",
  2788 => x"f8808098",
  2789 => x"800c800b",
  2790 => x"81bfb834",
  2791 => x"800b81bf",
  2792 => x"bc34833d",
  2793 => x"0d04ff3d",
  2794 => x"0d80c00b",
  2795 => x"f8808098",
  2796 => x"800c81a1",
  2797 => x"0bf88080",
  2798 => x"98800c81",
  2799 => x"c00bf880",
  2800 => x"8098800c",
  2801 => x"81a40bf8",
  2802 => x"80809880",
  2803 => x"0c81a60b",
  2804 => x"f8808098",
  2805 => x"800c81a2",
  2806 => x"0bf88080",
  2807 => x"98800caf",
  2808 => x"0bf88080",
  2809 => x"98800ca5",
  2810 => x"0bf88080",
  2811 => x"98800c81",
  2812 => x"810bf880",
  2813 => x"8098800c",
  2814 => x"9d0bf880",
  2815 => x"8098800c",
  2816 => x"81fa0bf8",
  2817 => x"80809880",
  2818 => x"0c800bf8",
  2819 => x"80809880",
  2820 => x"0c805271",
  2821 => x"81b00781",
  2822 => x"bf06f880",
  2823 => x"8098800c",
  2824 => x"900bf880",
  2825 => x"8098800c",
  2826 => x"800bf880",
  2827 => x"8098800c",
  2828 => x"8051800b",
  2829 => x"f8808098",
  2830 => x"840c8111",
  2831 => x"7081ff06",
  2832 => x"515180e5",
  2833 => x"7127eb38",
  2834 => x"81127081",
  2835 => x"ff065351",
  2836 => x"877227ff",
  2837 => x"be3881b0",
  2838 => x"0bf88080",
  2839 => x"98800c90",
  2840 => x"0bf88080",
  2841 => x"98800c80",
  2842 => x"0bf88080",
  2843 => x"98800c80",
  2844 => x"0b81bfb8",
  2845 => x"34800b81",
  2846 => x"bfbc3481",
  2847 => x"af0bf880",
  2848 => x"8098800c",
  2849 => x"833d0d04",
  2850 => x"803d0d02",
  2851 => x"8f053373",
  2852 => x"81e3bc0c",
  2853 => x"517081e3",
  2854 => x"c034823d",
  2855 => x"0d04ee3d",
  2856 => x"0d640284",
  2857 => x"0580d705",
  2858 => x"33028805",
  2859 => x"80db0533",
  2860 => x"59575980",
  2861 => x"76810677",
  2862 => x"812a8106",
  2863 => x"78832b81",
  2864 => x"80067982",
  2865 => x"2a810657",
  2866 => x"5e415f5d",
  2867 => x"81ff4272",
  2868 => x"7d2e0981",
  2869 => x"0683387c",
  2870 => x"42768a2e",
  2871 => x"83b93888",
  2872 => x"19085574",
  2873 => x"802e83a4",
  2874 => x"38851933",
  2875 => x"5aff5376",
  2876 => x"7a268e38",
  2877 => x"84193354",
  2878 => x"73772685",
  2879 => x"38767431",
  2880 => x"53741370",
  2881 => x"33545872",
  2882 => x"81ff0683",
  2883 => x"1a337098",
  2884 => x"2b81ff0a",
  2885 => x"119b2a81",
  2886 => x"055b4542",
  2887 => x"40815374",
  2888 => x"83387453",
  2889 => x"7281ff06",
  2890 => x"43807a81",
  2891 => x"ff06545c",
  2892 => x"ff547673",
  2893 => x"268b3884",
  2894 => x"19335376",
  2895 => x"732783f4",
  2896 => x"38737481",
  2897 => x"ff065553",
  2898 => x"805a7973",
  2899 => x"24ab3874",
  2900 => x"7a2e0981",
  2901 => x"0682e138",
  2902 => x"60982b81",
  2903 => x"ff0a119b",
  2904 => x"2a821b33",
  2905 => x"71712911",
  2906 => x"7081ff06",
  2907 => x"7871298c",
  2908 => x"1f080552",
  2909 => x"455d575d",
  2910 => x"537f6305",
  2911 => x"7081ff06",
  2912 => x"70612b70",
  2913 => x"81ff067b",
  2914 => x"622b7081",
  2915 => x"ff067b83",
  2916 => x"2a81065f",
  2917 => x"5358525e",
  2918 => x"42557880",
  2919 => x"2e8f3881",
  2920 => x"bfb83361",
  2921 => x"05567580",
  2922 => x"e62483c5",
  2923 => x"387f7829",
  2924 => x"61304157",
  2925 => x"7c7e2c98",
  2926 => x"2b70982c",
  2927 => x"55557377",
  2928 => x"25818238",
  2929 => x"ff1c7d81",
  2930 => x"065a537c",
  2931 => x"732e83c4",
  2932 => x"387e86a6",
  2933 => x"386184eb",
  2934 => x"387d802e",
  2935 => x"82a43879",
  2936 => x"14703370",
  2937 => x"58545580",
  2938 => x"5578752e",
  2939 => x"85387284",
  2940 => x"2a567583",
  2941 => x"2a708106",
  2942 => x"51537280",
  2943 => x"2e843881",
  2944 => x"c0557582",
  2945 => x"2a708106",
  2946 => x"51537280",
  2947 => x"2e853874",
  2948 => x"b0075575",
  2949 => x"812a7081",
  2950 => x"06515372",
  2951 => x"802e8538",
  2952 => x"748c0755",
  2953 => x"75810653",
  2954 => x"72802e85",
  2955 => x"38748307",
  2956 => x"557451f9",
  2957 => x"e33f7714",
  2958 => x"982b7098",
  2959 => x"2c555676",
  2960 => x"7424ff9b",
  2961 => x"3862802e",
  2962 => x"953861ff",
  2963 => x"1d54547c",
  2964 => x"732e81fb",
  2965 => x"387351f9",
  2966 => x"bf3f7e81",
  2967 => x"ea387f52",
  2968 => x"8151f8e8",
  2969 => x"3f811d70",
  2970 => x"81ff065e",
  2971 => x"547b7d26",
  2972 => x"fec23860",
  2973 => x"527b3070",
  2974 => x"982b7098",
  2975 => x"2c53585b",
  2976 => x"f8ca3f60",
  2977 => x"5372b00c",
  2978 => x"943d0d04",
  2979 => x"82193385",
  2980 => x"1a335b53",
  2981 => x"fcf13981",
  2982 => x"bfbc3353",
  2983 => x"72872681",
  2984 => x"9a388113",
  2985 => x"56805275",
  2986 => x"81ff0651",
  2987 => x"f7e43f80",
  2988 => x"5372b00c",
  2989 => x"943d0d04",
  2990 => x"73802eaf",
  2991 => x"38ff1470",
  2992 => x"81ff0655",
  2993 => x"5a7381ff",
  2994 => x"2ea13874",
  2995 => x"70810556",
  2996 => x"337c0570",
  2997 => x"83ffff06",
  2998 => x"ff167081",
  2999 => x"ff06575c",
  3000 => x"5d537381",
  3001 => x"ff2e0981",
  3002 => x"06e13860",
  3003 => x"982b81ff",
  3004 => x"0a119b2a",
  3005 => x"707e291e",
  3006 => x"8c1c0805",
  3007 => x"5c4255fc",
  3008 => x"f8397914",
  3009 => x"70335259",
  3010 => x"f88e3f77",
  3011 => x"14982b70",
  3012 => x"982c5556",
  3013 => x"737725fe",
  3014 => x"ac387914",
  3015 => x"70335259",
  3016 => x"f7f63f77",
  3017 => x"14982b70",
  3018 => x"982c5556",
  3019 => x"767424d2",
  3020 => x"38fe9239",
  3021 => x"76733154",
  3022 => x"fc873980",
  3023 => x"528051f6",
  3024 => x"d13f8053",
  3025 => x"feeb3973",
  3026 => x"51f7cd3f",
  3027 => x"fe903961",
  3028 => x"7b327081",
  3029 => x"ff065555",
  3030 => x"7d802efd",
  3031 => x"f8387a81",
  3032 => x"2a743270",
  3033 => x"5254f7b0",
  3034 => x"3f7e802e",
  3035 => x"fdf038d7",
  3036 => x"3981bfbc",
  3037 => x"337c0553",
  3038 => x"80527281",
  3039 => x"ff0651f6",
  3040 => x"913f8053",
  3041 => x"76a02efd",
  3042 => x"fc387f78",
  3043 => x"29613041",
  3044 => x"57fca139",
  3045 => x"7e87ad38",
  3046 => x"6185eb38",
  3047 => x"7d802e80",
  3048 => x"ec387914",
  3049 => x"70337c07",
  3050 => x"70525456",
  3051 => x"80557875",
  3052 => x"2e853872",
  3053 => x"842a5675",
  3054 => x"832a7081",
  3055 => x"06515372",
  3056 => x"802e8438",
  3057 => x"81c05575",
  3058 => x"822a7081",
  3059 => x"06515372",
  3060 => x"802e8538",
  3061 => x"74b00755",
  3062 => x"75812a70",
  3063 => x"81065153",
  3064 => x"72802e85",
  3065 => x"38748c07",
  3066 => x"55758106",
  3067 => x"5372802e",
  3068 => x"85387483",
  3069 => x"07557451",
  3070 => x"f69e3f77",
  3071 => x"14982b70",
  3072 => x"982c5553",
  3073 => x"767424ff",
  3074 => x"9938fcb9",
  3075 => x"39791470",
  3076 => x"337c0752",
  3077 => x"56f6813f",
  3078 => x"7714982b",
  3079 => x"70982c55",
  3080 => x"59737725",
  3081 => x"fc9f3879",
  3082 => x"1470337c",
  3083 => x"075256f5",
  3084 => x"e73f7714",
  3085 => x"982b7098",
  3086 => x"2c555976",
  3087 => x"7424ce38",
  3088 => x"fc83397d",
  3089 => x"802e80f0",
  3090 => x"38791470",
  3091 => x"33705854",
  3092 => x"55805578",
  3093 => x"752e8538",
  3094 => x"72842a56",
  3095 => x"75832a70",
  3096 => x"81065153",
  3097 => x"72802e84",
  3098 => x"3881c055",
  3099 => x"75822a70",
  3100 => x"81065153",
  3101 => x"72802e85",
  3102 => x"3874b007",
  3103 => x"5575812a",
  3104 => x"70810651",
  3105 => x"5372802e",
  3106 => x"8538748c",
  3107 => x"07557581",
  3108 => x"06537280",
  3109 => x"2e853874",
  3110 => x"83075574",
  3111 => x"097081ff",
  3112 => x"065253f4",
  3113 => x"f33f7714",
  3114 => x"982b7098",
  3115 => x"2c555676",
  3116 => x"7424ff95",
  3117 => x"38fb8e39",
  3118 => x"79147033",
  3119 => x"70097081",
  3120 => x"ff065458",
  3121 => x"5455f4d0",
  3122 => x"3f771498",
  3123 => x"2b70982c",
  3124 => x"55597377",
  3125 => x"25faee38",
  3126 => x"79147033",
  3127 => x"70097081",
  3128 => x"ff065458",
  3129 => x"5455f4b0",
  3130 => x"3f771498",
  3131 => x"2b70982c",
  3132 => x"55597674",
  3133 => x"24c238fa",
  3134 => x"cc396180",
  3135 => x"2e81ce38",
  3136 => x"7d802e80",
  3137 => x"f7387914",
  3138 => x"70337058",
  3139 => x"54558055",
  3140 => x"78752e85",
  3141 => x"3872842a",
  3142 => x"5675832a",
  3143 => x"70810651",
  3144 => x"5372802e",
  3145 => x"843881c0",
  3146 => x"5575822a",
  3147 => x"70810651",
  3148 => x"5372802e",
  3149 => x"853874b0",
  3150 => x"07557581",
  3151 => x"2a708106",
  3152 => x"51537280",
  3153 => x"2e853874",
  3154 => x"8c075575",
  3155 => x"81065372",
  3156 => x"802e8538",
  3157 => x"74830755",
  3158 => x"74097081",
  3159 => x"ff067053",
  3160 => x"5753f3b4",
  3161 => x"3f7551f3",
  3162 => x"af3f7714",
  3163 => x"982b7098",
  3164 => x"2c555576",
  3165 => x"7424ff8e",
  3166 => x"38f9ca39",
  3167 => x"79147033",
  3168 => x"70097081",
  3169 => x"ff067055",
  3170 => x"59555659",
  3171 => x"f38a3f75",
  3172 => x"51f3853f",
  3173 => x"7714982b",
  3174 => x"70982c55",
  3175 => x"59737725",
  3176 => x"f9a33879",
  3177 => x"14703370",
  3178 => x"097081ff",
  3179 => x"06705559",
  3180 => x"555659f2",
  3181 => x"e33f7551",
  3182 => x"f2de3f77",
  3183 => x"14982b70",
  3184 => x"982c5559",
  3185 => x"767424ff",
  3186 => x"b338f8f9",
  3187 => x"397d802e",
  3188 => x"80f43879",
  3189 => x"14703370",
  3190 => x"58545580",
  3191 => x"5578752e",
  3192 => x"85387284",
  3193 => x"2a567583",
  3194 => x"2a708106",
  3195 => x"51537280",
  3196 => x"2e843881",
  3197 => x"c0557582",
  3198 => x"2a708106",
  3199 => x"51537280",
  3200 => x"2e853874",
  3201 => x"b0075575",
  3202 => x"812a7081",
  3203 => x"06515372",
  3204 => x"802e8538",
  3205 => x"748c0755",
  3206 => x"75810653",
  3207 => x"72802e85",
  3208 => x"38748307",
  3209 => x"557481ff",
  3210 => x"06705256",
  3211 => x"f1ea3f75",
  3212 => x"51f1e53f",
  3213 => x"7714982b",
  3214 => x"70982c55",
  3215 => x"55767424",
  3216 => x"ff9138f8",
  3217 => x"80397914",
  3218 => x"70337053",
  3219 => x"5753f1c8",
  3220 => x"3f7551f1",
  3221 => x"c33f7714",
  3222 => x"982b7098",
  3223 => x"2c555973",
  3224 => x"7725f7e1",
  3225 => x"38791470",
  3226 => x"33705357",
  3227 => x"53f1a93f",
  3228 => x"7551f1a4",
  3229 => x"3f771498",
  3230 => x"2b70982c",
  3231 => x"55597674",
  3232 => x"24c438f7",
  3233 => x"c0397d80",
  3234 => x"2e80f238",
  3235 => x"79147033",
  3236 => x"7c077052",
  3237 => x"54568055",
  3238 => x"78752e85",
  3239 => x"3872842a",
  3240 => x"5675832a",
  3241 => x"70810651",
  3242 => x"5372802e",
  3243 => x"843881c0",
  3244 => x"5575822a",
  3245 => x"70810651",
  3246 => x"5372802e",
  3247 => x"853874b0",
  3248 => x"07557581",
  3249 => x"2a708106",
  3250 => x"51537280",
  3251 => x"2e853874",
  3252 => x"8c075575",
  3253 => x"81065372",
  3254 => x"802e8538",
  3255 => x"74830755",
  3256 => x"74097081",
  3257 => x"ff065256",
  3258 => x"f0ae3f77",
  3259 => x"14982b70",
  3260 => x"982c5553",
  3261 => x"767424ff",
  3262 => x"9338f6c9",
  3263 => x"39791470",
  3264 => x"337c0770",
  3265 => x"097081ff",
  3266 => x"06545556",
  3267 => x"59f0893f",
  3268 => x"7714982b",
  3269 => x"70982c55",
  3270 => x"59737725",
  3271 => x"f6a73879",
  3272 => x"1470337c",
  3273 => x"07700970",
  3274 => x"81ff0654",
  3275 => x"555659ef",
  3276 => x"e73f7714",
  3277 => x"982b7098",
  3278 => x"2c555976",
  3279 => x"7424ffbd",
  3280 => x"38f68239",
  3281 => x"61802e81",
  3282 => x"d4387d80",
  3283 => x"2e80f938",
  3284 => x"79147033",
  3285 => x"7c077052",
  3286 => x"54568055",
  3287 => x"78752e85",
  3288 => x"3872842a",
  3289 => x"5675832a",
  3290 => x"70810651",
  3291 => x"5372802e",
  3292 => x"843881c0",
  3293 => x"5575822a",
  3294 => x"70810651",
  3295 => x"5372802e",
  3296 => x"853874b0",
  3297 => x"07557581",
  3298 => x"2a708106",
  3299 => x"51537280",
  3300 => x"2e853874",
  3301 => x"8c075575",
  3302 => x"81065372",
  3303 => x"802e8538",
  3304 => x"74830755",
  3305 => x"74097081",
  3306 => x"ff067053",
  3307 => x"5456eee8",
  3308 => x"3f7251ee",
  3309 => x"e33f7714",
  3310 => x"982b7098",
  3311 => x"2c555676",
  3312 => x"7424ff8c",
  3313 => x"38f4fe39",
  3314 => x"79147033",
  3315 => x"7c077009",
  3316 => x"7081ff06",
  3317 => x"70555357",
  3318 => x"5753eebc",
  3319 => x"3f7251ee",
  3320 => x"b73f7714",
  3321 => x"982b7098",
  3322 => x"2c555973",
  3323 => x"7725f4d5",
  3324 => x"38791470",
  3325 => x"337c0770",
  3326 => x"097081ff",
  3327 => x"06705553",
  3328 => x"575753ee",
  3329 => x"933f7251",
  3330 => x"ee8e3f77",
  3331 => x"14982b70",
  3332 => x"982c5559",
  3333 => x"767424ff",
  3334 => x"af38f4a9",
  3335 => x"397d802e",
  3336 => x"80f63879",
  3337 => x"1470337c",
  3338 => x"07705254",
  3339 => x"56805578",
  3340 => x"752e8538",
  3341 => x"72842a56",
  3342 => x"75832a70",
  3343 => x"81065153",
  3344 => x"72802e84",
  3345 => x"3881c055",
  3346 => x"75822a70",
  3347 => x"81065153",
  3348 => x"72802e85",
  3349 => x"3874b007",
  3350 => x"5575812a",
  3351 => x"70810651",
  3352 => x"5372802e",
  3353 => x"8538748c",
  3354 => x"07557581",
  3355 => x"06537280",
  3356 => x"2e853874",
  3357 => x"83075574",
  3358 => x"81ff0670",
  3359 => x"5256ed98",
  3360 => x"3f7551ed",
  3361 => x"933f7714",
  3362 => x"982b7098",
  3363 => x"2c555376",
  3364 => x"7424ff8f",
  3365 => x"38f3ae39",
  3366 => x"79147033",
  3367 => x"7c077053",
  3368 => x"5456ecf4",
  3369 => x"3f7251ec",
  3370 => x"ef3f7714",
  3371 => x"982b7098",
  3372 => x"2c555973",
  3373 => x"7725f38d",
  3374 => x"38791470",
  3375 => x"337c0770",
  3376 => x"535456ec",
  3377 => x"d33f7251",
  3378 => x"ecce3f77",
  3379 => x"14982b70",
  3380 => x"982c5559",
  3381 => x"767424c0",
  3382 => x"38f2ea39",
  3383 => x"f83d0d7a",
  3384 => x"7d028805",
  3385 => x"af05335a",
  3386 => x"55598074",
  3387 => x"70810556",
  3388 => x"33755856",
  3389 => x"5774772e",
  3390 => x"09810688",
  3391 => x"3876b00c",
  3392 => x"8a3d0d04",
  3393 => x"74537752",
  3394 => x"7851ef92",
  3395 => x"3fb00881",
  3396 => x"ff067705",
  3397 => x"7083ffff",
  3398 => x"06777081",
  3399 => x"05593352",
  3400 => x"58557480",
  3401 => x"2ed73874",
  3402 => x"53775278",
  3403 => x"51eeef3f",
  3404 => x"b00881ff",
  3405 => x"06770570",
  3406 => x"83ffff06",
  3407 => x"77708105",
  3408 => x"59335258",
  3409 => x"5574ffbc",
  3410 => x"38ffb239",
  3411 => x"fe3d0d02",
  3412 => x"93053353",
  3413 => x"81e3c033",
  3414 => x"5281e3bc",
  3415 => x"0851eebe",
  3416 => x"3fb00881",
  3417 => x"ff06b00c",
  3418 => x"843d0d04",
  3419 => x"da9f3f04",
  3420 => x"fb3d0d77",
  3421 => x"79555580",
  3422 => x"56757524",
  3423 => x"ab388074",
  3424 => x"249d3880",
  3425 => x"53735274",
  3426 => x"5180e13f",
  3427 => x"b0085475",
  3428 => x"802e8538",
  3429 => x"b0083054",
  3430 => x"73b00c87",
  3431 => x"3d0d0473",
  3432 => x"30768132",
  3433 => x"5754dc39",
  3434 => x"74305581",
  3435 => x"56738025",
  3436 => x"d238ec39",
  3437 => x"fa3d0d78",
  3438 => x"7a575580",
  3439 => x"57767524",
  3440 => x"a438759f",
  3441 => x"2c548153",
  3442 => x"75743274",
  3443 => x"31527451",
  3444 => x"9b3fb008",
  3445 => x"5476802e",
  3446 => x"8538b008",
  3447 => x"305473b0",
  3448 => x"0c883d0d",
  3449 => x"04743055",
  3450 => x"8157d739",
  3451 => x"fc3d0d76",
  3452 => x"78535481",
  3453 => x"53807473",
  3454 => x"26525572",
  3455 => x"802e9838",
  3456 => x"70802ea9",
  3457 => x"38807224",
  3458 => x"a4387110",
  3459 => x"73107572",
  3460 => x"26535452",
  3461 => x"72ea3873",
  3462 => x"51788338",
  3463 => x"745170b0",
  3464 => x"0c863d0d",
  3465 => x"0472812a",
  3466 => x"72812a53",
  3467 => x"5372802e",
  3468 => x"e6387174",
  3469 => x"26ef3873",
  3470 => x"72317574",
  3471 => x"0774812a",
  3472 => x"74812a55",
  3473 => x"555654e5",
  3474 => x"39101010",
  3475 => x"10101010",
  3476 => x"10101010",
  3477 => x"10101010",
  3478 => x"10101010",
  3479 => x"10101010",
  3480 => x"10101010",
  3481 => x"10101010",
  3482 => x"53510473",
  3483 => x"81ff0673",
  3484 => x"83060981",
  3485 => x"05830510",
  3486 => x"10102b07",
  3487 => x"72fc060c",
  3488 => x"5151043c",
  3489 => x"04727280",
  3490 => x"728106ff",
  3491 => x"05097206",
  3492 => x"05711052",
  3493 => x"720a100a",
  3494 => x"5372ed38",
  3495 => x"51515351",
  3496 => x"04b008b4",
  3497 => x"08b80875",
  3498 => x"7580ebb4",
  3499 => x"2d5050b0",
  3500 => x"0856b80c",
  3501 => x"b40cb00c",
  3502 => x"5104b008",
  3503 => x"b408b808",
  3504 => x"757580ea",
  3505 => x"f02d5050",
  3506 => x"b00856b8",
  3507 => x"0cb40cb0",
  3508 => x"0c5104b0",
  3509 => x"08b408b8",
  3510 => x"0880c4e4",
  3511 => x"2db80cb4",
  3512 => x"0cb00c04",
  3513 => x"ff3d0d02",
  3514 => x"8f053381",
  3515 => x"bff40852",
  3516 => x"710c800b",
  3517 => x"b00c833d",
  3518 => x"0d04ff3d",
  3519 => x"0d028f05",
  3520 => x"335181e3",
  3521 => x"c4085271",
  3522 => x"2db00881",
  3523 => x"ff06b00c",
  3524 => x"833d0d04",
  3525 => x"fe3d0d74",
  3526 => x"70335353",
  3527 => x"71802e93",
  3528 => x"38811372",
  3529 => x"5281e3c4",
  3530 => x"08535371",
  3531 => x"2d723352",
  3532 => x"71ef3884",
  3533 => x"3d0d04f4",
  3534 => x"3d0d7f02",
  3535 => x"8405bb05",
  3536 => x"33555788",
  3537 => x"0b8c3d5b",
  3538 => x"59895381",
  3539 => x"bd8c5279",
  3540 => x"5186923f",
  3541 => x"73792e80",
  3542 => x"ff387856",
  3543 => x"73902e80",
  3544 => x"ec3802a7",
  3545 => x"0558768f",
  3546 => x"06547389",
  3547 => x"2680c238",
  3548 => x"7518b015",
  3549 => x"55557375",
  3550 => x"3476842a",
  3551 => x"ff177081",
  3552 => x"ff065855",
  3553 => x"5775df38",
  3554 => x"781a5575",
  3555 => x"75347970",
  3556 => x"33555573",
  3557 => x"802e9338",
  3558 => x"81157452",
  3559 => x"81e3c408",
  3560 => x"5755752d",
  3561 => x"74335473",
  3562 => x"ef3878b0",
  3563 => x"0c8e3d0d",
  3564 => x"047518b7",
  3565 => x"15555573",
  3566 => x"75347684",
  3567 => x"2aff1770",
  3568 => x"81ff0658",
  3569 => x"555775ff",
  3570 => x"9d38ffbc",
  3571 => x"39847057",
  3572 => x"5902a705",
  3573 => x"58ff8f39",
  3574 => x"82705759",
  3575 => x"f439f13d",
  3576 => x"0d618d3d",
  3577 => x"705b5c5a",
  3578 => x"807a5657",
  3579 => x"767a2481",
  3580 => x"85387817",
  3581 => x"548a5274",
  3582 => x"5184b83f",
  3583 => x"b008b005",
  3584 => x"53727434",
  3585 => x"8117578a",
  3586 => x"52745184",
  3587 => x"813fb008",
  3588 => x"55b008de",
  3589 => x"38b00877",
  3590 => x"9f2a1870",
  3591 => x"812c5a56",
  3592 => x"56807825",
  3593 => x"9e387817",
  3594 => x"ff055575",
  3595 => x"19703355",
  3596 => x"53743373",
  3597 => x"34737534",
  3598 => x"8116ff16",
  3599 => x"56567776",
  3600 => x"24e93876",
  3601 => x"19588078",
  3602 => x"34807a24",
  3603 => x"177081ff",
  3604 => x"067c7033",
  3605 => x"56575556",
  3606 => x"72802e93",
  3607 => x"38811573",
  3608 => x"5281e3c4",
  3609 => x"08585576",
  3610 => x"2d743353",
  3611 => x"72ef3873",
  3612 => x"b00c913d",
  3613 => x"0d04ad7b",
  3614 => x"3402ad05",
  3615 => x"7a307119",
  3616 => x"5656598a",
  3617 => x"52745183",
  3618 => x"aa3fb008",
  3619 => x"b0055372",
  3620 => x"74348117",
  3621 => x"578a5274",
  3622 => x"5182f33f",
  3623 => x"b00855b0",
  3624 => x"08fecf38",
  3625 => x"feef39fd",
  3626 => x"3d0d81bf",
  3627 => x"e80876b2",
  3628 => x"e4299412",
  3629 => x"0c54850b",
  3630 => x"98150c98",
  3631 => x"14087081",
  3632 => x"06515372",
  3633 => x"f638853d",
  3634 => x"0d04803d",
  3635 => x"0d81bfe8",
  3636 => x"0851870b",
  3637 => x"84120cff",
  3638 => x"0ba4120c",
  3639 => x"a70ba812",
  3640 => x"0cb2e40b",
  3641 => x"94120c87",
  3642 => x"0b98120c",
  3643 => x"823d0d04",
  3644 => x"803d0d81",
  3645 => x"bfec0851",
  3646 => x"b80b8c12",
  3647 => x"0c830b88",
  3648 => x"120c823d",
  3649 => x"0d04803d",
  3650 => x"0d81bfec",
  3651 => x"08841108",
  3652 => x"8106b00c",
  3653 => x"51823d0d",
  3654 => x"04ff3d0d",
  3655 => x"81bfec08",
  3656 => x"52841208",
  3657 => x"70810651",
  3658 => x"5170802e",
  3659 => x"f4387108",
  3660 => x"7081ff06",
  3661 => x"b00c5183",
  3662 => x"3d0d04fe",
  3663 => x"3d0d0293",
  3664 => x"05335372",
  3665 => x"8a2e9c38",
  3666 => x"81bfec08",
  3667 => x"52841208",
  3668 => x"70892a70",
  3669 => x"81065151",
  3670 => x"5170f238",
  3671 => x"72720c84",
  3672 => x"3d0d0481",
  3673 => x"bfec0852",
  3674 => x"84120870",
  3675 => x"892a7081",
  3676 => x"06515151",
  3677 => x"70f2388d",
  3678 => x"720c8412",
  3679 => x"0870892a",
  3680 => x"70810651",
  3681 => x"515170c5",
  3682 => x"38d239fa",
  3683 => x"3d0d02a3",
  3684 => x"053381bf",
  3685 => x"e00881e3",
  3686 => x"c8337081",
  3687 => x"ff067010",
  3688 => x"101181e3",
  3689 => x"cc337081",
  3690 => x"ff067290",
  3691 => x"29117088",
  3692 => x"2b780777",
  3693 => x"0c535b5b",
  3694 => x"55555954",
  3695 => x"54738a2e",
  3696 => x"98387480",
  3697 => x"cf2e9238",
  3698 => x"738c2ea4",
  3699 => x"38811653",
  3700 => x"7281e3cc",
  3701 => x"34883d0d",
  3702 => x"0471a326",
  3703 => x"a3388117",
  3704 => x"527181e3",
  3705 => x"c834800b",
  3706 => x"81e3cc34",
  3707 => x"883d0d04",
  3708 => x"80527188",
  3709 => x"2b730c81",
  3710 => x"12529790",
  3711 => x"7226f338",
  3712 => x"800b81e3",
  3713 => x"c834800b",
  3714 => x"81e3cc34",
  3715 => x"df39bc08",
  3716 => x"02bc0cfd",
  3717 => x"3d0d8053",
  3718 => x"bc088c05",
  3719 => x"0852bc08",
  3720 => x"88050851",
  3721 => x"f7c63fb0",
  3722 => x"0870b00c",
  3723 => x"54853d0d",
  3724 => x"bc0c04bc",
  3725 => x"0802bc0c",
  3726 => x"fd3d0d81",
  3727 => x"53bc088c",
  3728 => x"050852bc",
  3729 => x"08880508",
  3730 => x"51f7a13f",
  3731 => x"b00870b0",
  3732 => x"0c54853d",
  3733 => x"0dbc0c04",
  3734 => x"803d0d86",
  3735 => x"5184963f",
  3736 => x"8151a1d3",
  3737 => x"3ffc3d0d",
  3738 => x"7670797b",
  3739 => x"55555555",
  3740 => x"8f72278c",
  3741 => x"38727507",
  3742 => x"83065170",
  3743 => x"802ea738",
  3744 => x"ff125271",
  3745 => x"ff2e9838",
  3746 => x"72708105",
  3747 => x"54337470",
  3748 => x"81055634",
  3749 => x"ff125271",
  3750 => x"ff2e0981",
  3751 => x"06ea3874",
  3752 => x"b00c863d",
  3753 => x"0d047451",
  3754 => x"72708405",
  3755 => x"54087170",
  3756 => x"8405530c",
  3757 => x"72708405",
  3758 => x"54087170",
  3759 => x"8405530c",
  3760 => x"72708405",
  3761 => x"54087170",
  3762 => x"8405530c",
  3763 => x"72708405",
  3764 => x"54087170",
  3765 => x"8405530c",
  3766 => x"f0125271",
  3767 => x"8f26c938",
  3768 => x"83722795",
  3769 => x"38727084",
  3770 => x"05540871",
  3771 => x"70840553",
  3772 => x"0cfc1252",
  3773 => x"718326ed",
  3774 => x"387054ff",
  3775 => x"8339fd3d",
  3776 => x"0d755384",
  3777 => x"d8130880",
  3778 => x"2e8a3880",
  3779 => x"5372b00c",
  3780 => x"853d0d04",
  3781 => x"81805272",
  3782 => x"518d9b3f",
  3783 => x"b00884d8",
  3784 => x"140cff53",
  3785 => x"b008802e",
  3786 => x"e438b008",
  3787 => x"549f5380",
  3788 => x"74708405",
  3789 => x"560cff13",
  3790 => x"53807324",
  3791 => x"ce388074",
  3792 => x"70840556",
  3793 => x"0cff1353",
  3794 => x"728025e3",
  3795 => x"38ffbc39",
  3796 => x"fd3d0d75",
  3797 => x"7755539f",
  3798 => x"74278d38",
  3799 => x"96730cff",
  3800 => x"5271b00c",
  3801 => x"853d0d04",
  3802 => x"84d81308",
  3803 => x"5271802e",
  3804 => x"93387310",
  3805 => x"10127008",
  3806 => x"79720c51",
  3807 => x"5271b00c",
  3808 => x"853d0d04",
  3809 => x"7251fef6",
  3810 => x"3fff52b0",
  3811 => x"08d33884",
  3812 => x"d8130874",
  3813 => x"10101170",
  3814 => x"087a720c",
  3815 => x"515152dd",
  3816 => x"39f93d0d",
  3817 => x"797b5856",
  3818 => x"769f2680",
  3819 => x"e83884d8",
  3820 => x"16085473",
  3821 => x"802eaa38",
  3822 => x"76101014",
  3823 => x"70085555",
  3824 => x"73802eba",
  3825 => x"38805873",
  3826 => x"812e8f38",
  3827 => x"73ff2ea3",
  3828 => x"3880750c",
  3829 => x"7651732d",
  3830 => x"805877b0",
  3831 => x"0c893d0d",
  3832 => x"047551fe",
  3833 => x"993fff58",
  3834 => x"b008ef38",
  3835 => x"84d81608",
  3836 => x"54c63996",
  3837 => x"760c810b",
  3838 => x"b00c893d",
  3839 => x"0d047551",
  3840 => x"81ed3f76",
  3841 => x"53b00852",
  3842 => x"755181ad",
  3843 => x"3fb008b0",
  3844 => x"0c893d0d",
  3845 => x"0496760c",
  3846 => x"ff0bb00c",
  3847 => x"893d0d04",
  3848 => x"fc3d0d76",
  3849 => x"785653ff",
  3850 => x"54749f26",
  3851 => x"b13884d8",
  3852 => x"13085271",
  3853 => x"802eae38",
  3854 => x"74101012",
  3855 => x"70085353",
  3856 => x"81547180",
  3857 => x"2e983882",
  3858 => x"5471ff2e",
  3859 => x"91388354",
  3860 => x"71812e8a",
  3861 => x"3880730c",
  3862 => x"7451712d",
  3863 => x"805473b0",
  3864 => x"0c863d0d",
  3865 => x"047251fd",
  3866 => x"953fb008",
  3867 => x"f13884d8",
  3868 => x"130852c4",
  3869 => x"39ff3d0d",
  3870 => x"735281bf",
  3871 => x"f80851fe",
  3872 => x"a03f833d",
  3873 => x"0d04fe3d",
  3874 => x"0d755374",
  3875 => x"5281bff8",
  3876 => x"0851fdbc",
  3877 => x"3f843d0d",
  3878 => x"04803d0d",
  3879 => x"81bff808",
  3880 => x"51fcdb3f",
  3881 => x"823d0d04",
  3882 => x"ff3d0d73",
  3883 => x"5281bff8",
  3884 => x"0851feec",
  3885 => x"3f833d0d",
  3886 => x"04fc3d0d",
  3887 => x"800b81e3",
  3888 => x"d40c7852",
  3889 => x"77519caa",
  3890 => x"3fb00854",
  3891 => x"b008ff2e",
  3892 => x"883873b0",
  3893 => x"0c863d0d",
  3894 => x"0481e3d4",
  3895 => x"08557480",
  3896 => x"2ef03876",
  3897 => x"75710c53",
  3898 => x"73b00c86",
  3899 => x"3d0d049b",
  3900 => x"fc3f04fc",
  3901 => x"3d0d7670",
  3902 => x"79707307",
  3903 => x"83065454",
  3904 => x"54557080",
  3905 => x"c3387170",
  3906 => x"08700970",
  3907 => x"f7fbfdff",
  3908 => x"130670f8",
  3909 => x"84828180",
  3910 => x"06515153",
  3911 => x"535470a6",
  3912 => x"38841472",
  3913 => x"74708405",
  3914 => x"560c7008",
  3915 => x"700970f7",
  3916 => x"fbfdff13",
  3917 => x"0670f884",
  3918 => x"82818006",
  3919 => x"51515353",
  3920 => x"5470802e",
  3921 => x"dc387352",
  3922 => x"71708105",
  3923 => x"53335170",
  3924 => x"73708105",
  3925 => x"553470f0",
  3926 => x"3874b00c",
  3927 => x"863d0d04",
  3928 => x"fd3d0d75",
  3929 => x"70718306",
  3930 => x"53555270",
  3931 => x"b8387170",
  3932 => x"087009f7",
  3933 => x"fbfdff12",
  3934 => x"0670f884",
  3935 => x"82818006",
  3936 => x"51515253",
  3937 => x"709d3884",
  3938 => x"13700870",
  3939 => x"09f7fbfd",
  3940 => x"ff120670",
  3941 => x"f8848281",
  3942 => x"80065151",
  3943 => x"52537080",
  3944 => x"2ee53872",
  3945 => x"52713351",
  3946 => x"70802e8a",
  3947 => x"38811270",
  3948 => x"33525270",
  3949 => x"f8387174",
  3950 => x"31b00c85",
  3951 => x"3d0d04fa",
  3952 => x"3d0d787a",
  3953 => x"7c705455",
  3954 => x"55527280",
  3955 => x"2e80d938",
  3956 => x"71740783",
  3957 => x"06517080",
  3958 => x"2e80d438",
  3959 => x"ff135372",
  3960 => x"ff2eb138",
  3961 => x"71337433",
  3962 => x"56517471",
  3963 => x"2e098106",
  3964 => x"a9387280",
  3965 => x"2e818738",
  3966 => x"7081ff06",
  3967 => x"5170802e",
  3968 => x"80fc3881",
  3969 => x"128115ff",
  3970 => x"15555552",
  3971 => x"72ff2e09",
  3972 => x"8106d138",
  3973 => x"71337433",
  3974 => x"56517081",
  3975 => x"ff067581",
  3976 => x"ff067171",
  3977 => x"31515252",
  3978 => x"70b00c88",
  3979 => x"3d0d0471",
  3980 => x"74575583",
  3981 => x"73278838",
  3982 => x"71087408",
  3983 => x"2e883874",
  3984 => x"765552ff",
  3985 => x"9739fc13",
  3986 => x"5372802e",
  3987 => x"b1387408",
  3988 => x"7009f7fb",
  3989 => x"fdff1206",
  3990 => x"70f88482",
  3991 => x"81800651",
  3992 => x"5151709a",
  3993 => x"38841584",
  3994 => x"17575583",
  3995 => x"7327d038",
  3996 => x"74087608",
  3997 => x"2ed03874",
  3998 => x"765552fe",
  3999 => x"df39800b",
  4000 => x"b00c883d",
  4001 => x"0d04f33d",
  4002 => x"0d606264",
  4003 => x"725a5a5e",
  4004 => x"5e805c76",
  4005 => x"70810558",
  4006 => x"3381bd99",
  4007 => x"11337083",
  4008 => x"2a708106",
  4009 => x"51555556",
  4010 => x"72e93875",
  4011 => x"ad2e8288",
  4012 => x"3875ab2e",
  4013 => x"82843877",
  4014 => x"30707907",
  4015 => x"80257990",
  4016 => x"32703070",
  4017 => x"72078025",
  4018 => x"73075357",
  4019 => x"57515372",
  4020 => x"802e8738",
  4021 => x"75b02e81",
  4022 => x"eb38778a",
  4023 => x"38885875",
  4024 => x"b02e8338",
  4025 => x"8a58810a",
  4026 => x"5a7b8438",
  4027 => x"fe0a5a77",
  4028 => x"527951f6",
  4029 => x"be3fb008",
  4030 => x"78537a52",
  4031 => x"5bf68f3f",
  4032 => x"b0085a80",
  4033 => x"7081bd99",
  4034 => x"18337082",
  4035 => x"2a708106",
  4036 => x"5156565a",
  4037 => x"5572802e",
  4038 => x"80c138d0",
  4039 => x"16567578",
  4040 => x"2580d738",
  4041 => x"80792475",
  4042 => x"7b260753",
  4043 => x"72933874",
  4044 => x"7a2e80eb",
  4045 => x"387a7625",
  4046 => x"80ed3872",
  4047 => x"802e80e7",
  4048 => x"38ff7770",
  4049 => x"81055933",
  4050 => x"575981bd",
  4051 => x"99163370",
  4052 => x"822a7081",
  4053 => x"06515454",
  4054 => x"72c13873",
  4055 => x"83065372",
  4056 => x"802e9738",
  4057 => x"738106c9",
  4058 => x"17555372",
  4059 => x"8538ffa9",
  4060 => x"16547356",
  4061 => x"777624ff",
  4062 => x"ab388079",
  4063 => x"2480f038",
  4064 => x"7b802e84",
  4065 => x"38743055",
  4066 => x"7c802e8c",
  4067 => x"38ff1753",
  4068 => x"7883387d",
  4069 => x"53727d0c",
  4070 => x"74b00c8f",
  4071 => x"3d0d0481",
  4072 => x"53757b24",
  4073 => x"ff953881",
  4074 => x"75792917",
  4075 => x"78708105",
  4076 => x"5a335856",
  4077 => x"59ff9339",
  4078 => x"815c7670",
  4079 => x"81055833",
  4080 => x"56fdf439",
  4081 => x"80773354",
  4082 => x"547280f8",
  4083 => x"2eb23872",
  4084 => x"80d83270",
  4085 => x"30708025",
  4086 => x"76075151",
  4087 => x"5372802e",
  4088 => x"fdf83881",
  4089 => x"17338218",
  4090 => x"58569058",
  4091 => x"fdf83981",
  4092 => x"0a557b84",
  4093 => x"38fe0a55",
  4094 => x"7f53a273",
  4095 => x"0cff8939",
  4096 => x"8154cc39",
  4097 => x"fd3d0d77",
  4098 => x"54765375",
  4099 => x"5281bff8",
  4100 => x"0851fcf2",
  4101 => x"3f853d0d",
  4102 => x"04f33d0d",
  4103 => x"60626472",
  4104 => x"5a5a5d5d",
  4105 => x"805e7670",
  4106 => x"81055833",
  4107 => x"81bd9911",
  4108 => x"3370832a",
  4109 => x"70810651",
  4110 => x"55555672",
  4111 => x"e93875ad",
  4112 => x"2e81ff38",
  4113 => x"75ab2e81",
  4114 => x"fb387730",
  4115 => x"70790780",
  4116 => x"25799032",
  4117 => x"70307072",
  4118 => x"07802573",
  4119 => x"07535757",
  4120 => x"51537280",
  4121 => x"2e873875",
  4122 => x"b02e81e2",
  4123 => x"38778a38",
  4124 => x"885875b0",
  4125 => x"2e83388a",
  4126 => x"587752ff",
  4127 => x"51f38f3f",
  4128 => x"b0087853",
  4129 => x"5aff51f3",
  4130 => x"aa3fb008",
  4131 => x"5b80705a",
  4132 => x"5581bd99",
  4133 => x"16337082",
  4134 => x"2a708106",
  4135 => x"51545472",
  4136 => x"802e80c1",
  4137 => x"38d01656",
  4138 => x"75782580",
  4139 => x"d7388079",
  4140 => x"24757b26",
  4141 => x"07537293",
  4142 => x"38747a2e",
  4143 => x"80eb387a",
  4144 => x"762580ed",
  4145 => x"3872802e",
  4146 => x"80e738ff",
  4147 => x"77708105",
  4148 => x"59335759",
  4149 => x"81bd9916",
  4150 => x"3370822a",
  4151 => x"70810651",
  4152 => x"545472c1",
  4153 => x"38738306",
  4154 => x"5372802e",
  4155 => x"97387381",
  4156 => x"06c91755",
  4157 => x"53728538",
  4158 => x"ffa91654",
  4159 => x"73567776",
  4160 => x"24ffab38",
  4161 => x"80792481",
  4162 => x"89387d80",
  4163 => x"2e843874",
  4164 => x"30557b80",
  4165 => x"2e8c38ff",
  4166 => x"17537883",
  4167 => x"387c5372",
  4168 => x"7c0c74b0",
  4169 => x"0c8f3d0d",
  4170 => x"04815375",
  4171 => x"7b24ff95",
  4172 => x"38817579",
  4173 => x"29177870",
  4174 => x"81055a33",
  4175 => x"585659ff",
  4176 => x"9339815e",
  4177 => x"76708105",
  4178 => x"583356fd",
  4179 => x"fd398077",
  4180 => x"33545472",
  4181 => x"80f82e80",
  4182 => x"c3387280",
  4183 => x"d8327030",
  4184 => x"70802576",
  4185 => x"07515153",
  4186 => x"72802efe",
  4187 => x"80388117",
  4188 => x"33821858",
  4189 => x"56907053",
  4190 => x"58ff51f1",
  4191 => x"913fb008",
  4192 => x"78535aff",
  4193 => x"51f1ac3f",
  4194 => x"b0085b80",
  4195 => x"705a55fe",
  4196 => x"8039ff60",
  4197 => x"5455a273",
  4198 => x"0cfef739",
  4199 => x"8154ffba",
  4200 => x"39fd3d0d",
  4201 => x"77547653",
  4202 => x"755281bf",
  4203 => x"f80851fc",
  4204 => x"e83f853d",
  4205 => x"0d04f33d",
  4206 => x"0d7f618b",
  4207 => x"1170f806",
  4208 => x"5c55555e",
  4209 => x"72962683",
  4210 => x"38905980",
  4211 => x"7924747a",
  4212 => x"26075380",
  4213 => x"5472742e",
  4214 => x"09810680",
  4215 => x"cb387d51",
  4216 => x"8bca3f78",
  4217 => x"83f72680",
  4218 => x"c6387883",
  4219 => x"2a701010",
  4220 => x"1081c7b4",
  4221 => x"058c1108",
  4222 => x"59595a76",
  4223 => x"782e83b0",
  4224 => x"38841708",
  4225 => x"fc06568c",
  4226 => x"17088818",
  4227 => x"08718c12",
  4228 => x"0c88120c",
  4229 => x"58751784",
  4230 => x"11088107",
  4231 => x"84120c53",
  4232 => x"7d518b89",
  4233 => x"3f881754",
  4234 => x"73b00c8f",
  4235 => x"3d0d0478",
  4236 => x"892a7983",
  4237 => x"2a5b5372",
  4238 => x"802ebf38",
  4239 => x"78862ab8",
  4240 => x"055a8473",
  4241 => x"27b43880",
  4242 => x"db135a94",
  4243 => x"7327ab38",
  4244 => x"788c2a80",
  4245 => x"ee055a80",
  4246 => x"d473279e",
  4247 => x"38788f2a",
  4248 => x"80f7055a",
  4249 => x"82d47327",
  4250 => x"91387892",
  4251 => x"2a80fc05",
  4252 => x"5a8ad473",
  4253 => x"27843880",
  4254 => x"fe5a7910",
  4255 => x"101081c7",
  4256 => x"b4058c11",
  4257 => x"08585576",
  4258 => x"752ea338",
  4259 => x"841708fc",
  4260 => x"06707a31",
  4261 => x"5556738f",
  4262 => x"2488d538",
  4263 => x"738025fe",
  4264 => x"e6388c17",
  4265 => x"08577675",
  4266 => x"2e098106",
  4267 => x"df38811a",
  4268 => x"5a81c7c4",
  4269 => x"08577681",
  4270 => x"c7bc2e82",
  4271 => x"c0388417",
  4272 => x"08fc0670",
  4273 => x"7a315556",
  4274 => x"738f2481",
  4275 => x"f93881c7",
  4276 => x"bc0b81c7",
  4277 => x"c80c81c7",
  4278 => x"bc0b81c7",
  4279 => x"c40c7380",
  4280 => x"25feb238",
  4281 => x"83ff7627",
  4282 => x"83df3875",
  4283 => x"892a7683",
  4284 => x"2a555372",
  4285 => x"802ebf38",
  4286 => x"75862ab8",
  4287 => x"05548473",
  4288 => x"27b43880",
  4289 => x"db135494",
  4290 => x"7327ab38",
  4291 => x"758c2a80",
  4292 => x"ee055480",
  4293 => x"d473279e",
  4294 => x"38758f2a",
  4295 => x"80f70554",
  4296 => x"82d47327",
  4297 => x"91387592",
  4298 => x"2a80fc05",
  4299 => x"548ad473",
  4300 => x"27843880",
  4301 => x"fe547310",
  4302 => x"101081c7",
  4303 => x"b4058811",
  4304 => x"08565874",
  4305 => x"782e86cf",
  4306 => x"38841508",
  4307 => x"fc065375",
  4308 => x"73278d38",
  4309 => x"88150855",
  4310 => x"74782e09",
  4311 => x"8106ea38",
  4312 => x"8c150881",
  4313 => x"c7b40b84",
  4314 => x"0508718c",
  4315 => x"1a0c7688",
  4316 => x"1a0c7888",
  4317 => x"130c788c",
  4318 => x"180c5d58",
  4319 => x"7953807a",
  4320 => x"2483e638",
  4321 => x"72822c81",
  4322 => x"712b5c53",
  4323 => x"7a7c2681",
  4324 => x"98387b7b",
  4325 => x"06537282",
  4326 => x"f13879fc",
  4327 => x"0684055a",
  4328 => x"7a10707d",
  4329 => x"06545b72",
  4330 => x"82e03884",
  4331 => x"1a5af139",
  4332 => x"88178c11",
  4333 => x"08585876",
  4334 => x"782e0981",
  4335 => x"06fcc238",
  4336 => x"821a5afd",
  4337 => x"ec397817",
  4338 => x"79810784",
  4339 => x"190c7081",
  4340 => x"c7c80c70",
  4341 => x"81c7c40c",
  4342 => x"81c7bc0b",
  4343 => x"8c120c8c",
  4344 => x"11088812",
  4345 => x"0c748107",
  4346 => x"84120c74",
  4347 => x"1175710c",
  4348 => x"51537d51",
  4349 => x"87b73f88",
  4350 => x"1754fcac",
  4351 => x"3981c7b4",
  4352 => x"0b840508",
  4353 => x"7a545c79",
  4354 => x"8025fef8",
  4355 => x"3882da39",
  4356 => x"7a097c06",
  4357 => x"7081c7b4",
  4358 => x"0b84050c",
  4359 => x"5c7a105b",
  4360 => x"7a7c2685",
  4361 => x"387a85b8",
  4362 => x"3881c7b4",
  4363 => x"0b880508",
  4364 => x"70841208",
  4365 => x"fc06707c",
  4366 => x"317c7226",
  4367 => x"8f722507",
  4368 => x"57575c5d",
  4369 => x"5572802e",
  4370 => x"80db3879",
  4371 => x"7a1681c7",
  4372 => x"ac081b90",
  4373 => x"115a5557",
  4374 => x"5b81c7a8",
  4375 => x"08ff2e88",
  4376 => x"38a08f13",
  4377 => x"e0800657",
  4378 => x"76527d51",
  4379 => x"86c03fb0",
  4380 => x"0854b008",
  4381 => x"ff2e9038",
  4382 => x"b0087627",
  4383 => x"82993874",
  4384 => x"81c7b42e",
  4385 => x"82913881",
  4386 => x"c7b40b88",
  4387 => x"05085584",
  4388 => x"1508fc06",
  4389 => x"707a317a",
  4390 => x"72268f72",
  4391 => x"25075255",
  4392 => x"537283e6",
  4393 => x"38747981",
  4394 => x"0784170c",
  4395 => x"79167081",
  4396 => x"c7b40b88",
  4397 => x"050c7581",
  4398 => x"0784120c",
  4399 => x"547e5257",
  4400 => x"85eb3f88",
  4401 => x"1754fae0",
  4402 => x"3975832a",
  4403 => x"70545480",
  4404 => x"7424819b",
  4405 => x"3872822c",
  4406 => x"81712b81",
  4407 => x"c7b80807",
  4408 => x"7081c7b4",
  4409 => x"0b84050c",
  4410 => x"75101010",
  4411 => x"81c7b405",
  4412 => x"88110858",
  4413 => x"5a5d5377",
  4414 => x"8c180c74",
  4415 => x"88180c76",
  4416 => x"88190c76",
  4417 => x"8c160cfc",
  4418 => x"f339797a",
  4419 => x"10101081",
  4420 => x"c7b40570",
  4421 => x"57595d8c",
  4422 => x"15085776",
  4423 => x"752ea338",
  4424 => x"841708fc",
  4425 => x"06707a31",
  4426 => x"5556738f",
  4427 => x"2483ca38",
  4428 => x"73802584",
  4429 => x"81388c17",
  4430 => x"08577675",
  4431 => x"2e098106",
  4432 => x"df388815",
  4433 => x"811b7083",
  4434 => x"06555b55",
  4435 => x"72c9387c",
  4436 => x"83065372",
  4437 => x"802efdb8",
  4438 => x"38ff1df8",
  4439 => x"19595d88",
  4440 => x"1808782e",
  4441 => x"ea38fdb5",
  4442 => x"39831a53",
  4443 => x"fc963983",
  4444 => x"1470822c",
  4445 => x"81712b81",
  4446 => x"c7b80807",
  4447 => x"7081c7b4",
  4448 => x"0b84050c",
  4449 => x"76101010",
  4450 => x"81c7b405",
  4451 => x"88110859",
  4452 => x"5b5e5153",
  4453 => x"fee13981",
  4454 => x"c6f80817",
  4455 => x"58b00876",
  4456 => x"2e818d38",
  4457 => x"81c7a808",
  4458 => x"ff2e83ec",
  4459 => x"38737631",
  4460 => x"1881c6f8",
  4461 => x"0c738706",
  4462 => x"70575372",
  4463 => x"802e8838",
  4464 => x"88733170",
  4465 => x"15555676",
  4466 => x"149fff06",
  4467 => x"a0807131",
  4468 => x"1770547f",
  4469 => x"53575383",
  4470 => x"d53fb008",
  4471 => x"53b008ff",
  4472 => x"2e81a038",
  4473 => x"81c6f808",
  4474 => x"167081c6",
  4475 => x"f80c7475",
  4476 => x"81c7b40b",
  4477 => x"88050c74",
  4478 => x"76311870",
  4479 => x"81075155",
  4480 => x"56587b81",
  4481 => x"c7b42e83",
  4482 => x"9c38798f",
  4483 => x"2682cb38",
  4484 => x"810b8415",
  4485 => x"0c841508",
  4486 => x"fc06707a",
  4487 => x"317a7226",
  4488 => x"8f722507",
  4489 => x"52555372",
  4490 => x"802efcf9",
  4491 => x"3880db39",
  4492 => x"b0089fff",
  4493 => x"065372fe",
  4494 => x"eb387781",
  4495 => x"c6f80c81",
  4496 => x"c7b40b88",
  4497 => x"05087b18",
  4498 => x"81078412",
  4499 => x"0c5581c7",
  4500 => x"a4087827",
  4501 => x"86387781",
  4502 => x"c7a40c81",
  4503 => x"c7a00878",
  4504 => x"27fcac38",
  4505 => x"7781c7a0",
  4506 => x"0c841508",
  4507 => x"fc06707a",
  4508 => x"317a7226",
  4509 => x"8f722507",
  4510 => x"52555372",
  4511 => x"802efca5",
  4512 => x"38883980",
  4513 => x"745456fe",
  4514 => x"db397d51",
  4515 => x"829f3f80",
  4516 => x"0bb00c8f",
  4517 => x"3d0d0473",
  4518 => x"53807424",
  4519 => x"a9387282",
  4520 => x"2c81712b",
  4521 => x"81c7b808",
  4522 => x"077081c7",
  4523 => x"b40b8405",
  4524 => x"0c5d5377",
  4525 => x"8c180c74",
  4526 => x"88180c76",
  4527 => x"88190c76",
  4528 => x"8c160cf9",
  4529 => x"b7398314",
  4530 => x"70822c81",
  4531 => x"712b81c7",
  4532 => x"b8080770",
  4533 => x"81c7b40b",
  4534 => x"84050c5e",
  4535 => x"5153d439",
  4536 => x"7b7b0653",
  4537 => x"72fca338",
  4538 => x"841a7b10",
  4539 => x"5c5af139",
  4540 => x"ff1a8111",
  4541 => x"515af7b9",
  4542 => x"39781779",
  4543 => x"81078419",
  4544 => x"0c8c1808",
  4545 => x"88190871",
  4546 => x"8c120c88",
  4547 => x"120c5970",
  4548 => x"81c7c80c",
  4549 => x"7081c7c4",
  4550 => x"0c81c7bc",
  4551 => x"0b8c120c",
  4552 => x"8c110888",
  4553 => x"120c7481",
  4554 => x"0784120c",
  4555 => x"74117571",
  4556 => x"0c5153f9",
  4557 => x"bd397517",
  4558 => x"84110881",
  4559 => x"0784120c",
  4560 => x"538c1708",
  4561 => x"88180871",
  4562 => x"8c120c88",
  4563 => x"120c587d",
  4564 => x"5180da3f",
  4565 => x"881754f5",
  4566 => x"cf397284",
  4567 => x"150cf41a",
  4568 => x"f8067084",
  4569 => x"1e088106",
  4570 => x"07841e0c",
  4571 => x"701d545b",
  4572 => x"850b8414",
  4573 => x"0c850b88",
  4574 => x"140c8f7b",
  4575 => x"27fdcf38",
  4576 => x"881c527d",
  4577 => x"5182903f",
  4578 => x"81c7b40b",
  4579 => x"88050881",
  4580 => x"c6f80859",
  4581 => x"55fdb739",
  4582 => x"7781c6f8",
  4583 => x"0c7381c7",
  4584 => x"a80cfc91",
  4585 => x"39728415",
  4586 => x"0cfda339",
  4587 => x"0404fd3d",
  4588 => x"0d800b81",
  4589 => x"e3d40c76",
  4590 => x"5186cb3f",
  4591 => x"b00853b0",
  4592 => x"08ff2e88",
  4593 => x"3872b00c",
  4594 => x"853d0d04",
  4595 => x"81e3d408",
  4596 => x"5473802e",
  4597 => x"f0387574",
  4598 => x"710c5272",
  4599 => x"b00c853d",
  4600 => x"0d04fb3d",
  4601 => x"0d777052",
  4602 => x"56c23f81",
  4603 => x"c7b40b88",
  4604 => x"05088411",
  4605 => x"08fc0670",
  4606 => x"7b319fef",
  4607 => x"05e08006",
  4608 => x"e0800556",
  4609 => x"5653a080",
  4610 => x"74249438",
  4611 => x"80527551",
  4612 => x"ff9c3f81",
  4613 => x"c7bc0815",
  4614 => x"5372b008",
  4615 => x"2e8f3875",
  4616 => x"51ff8a3f",
  4617 => x"805372b0",
  4618 => x"0c873d0d",
  4619 => x"04733052",
  4620 => x"7551fefa",
  4621 => x"3fb008ff",
  4622 => x"2ea83881",
  4623 => x"c7b40b88",
  4624 => x"05087575",
  4625 => x"31810784",
  4626 => x"120c5381",
  4627 => x"c6f80874",
  4628 => x"3181c6f8",
  4629 => x"0c7551fe",
  4630 => x"d43f810b",
  4631 => x"b00c873d",
  4632 => x"0d048052",
  4633 => x"7551fec6",
  4634 => x"3f81c7b4",
  4635 => x"0b880508",
  4636 => x"b0087131",
  4637 => x"56538f75",
  4638 => x"25ffa438",
  4639 => x"b00881c7",
  4640 => x"a8083181",
  4641 => x"c6f80c74",
  4642 => x"81078414",
  4643 => x"0c7551fe",
  4644 => x"9c3f8053",
  4645 => x"ff9039f6",
  4646 => x"3d0d7c7e",
  4647 => x"545b7280",
  4648 => x"2e828338",
  4649 => x"7a51fe84",
  4650 => x"3ff81384",
  4651 => x"110870fe",
  4652 => x"06701384",
  4653 => x"1108fc06",
  4654 => x"5d585954",
  4655 => x"5881c7bc",
  4656 => x"08752e82",
  4657 => x"de387884",
  4658 => x"160c8073",
  4659 => x"8106545a",
  4660 => x"727a2e81",
  4661 => x"d5387815",
  4662 => x"84110881",
  4663 => x"06515372",
  4664 => x"a0387817",
  4665 => x"577981e6",
  4666 => x"38881508",
  4667 => x"537281c7",
  4668 => x"bc2e82f9",
  4669 => x"388c1508",
  4670 => x"708c150c",
  4671 => x"7388120c",
  4672 => x"56768107",
  4673 => x"84190c76",
  4674 => x"1877710c",
  4675 => x"53798191",
  4676 => x"3883ff77",
  4677 => x"2781c838",
  4678 => x"76892a77",
  4679 => x"832a5653",
  4680 => x"72802ebf",
  4681 => x"3876862a",
  4682 => x"b8055584",
  4683 => x"7327b438",
  4684 => x"80db1355",
  4685 => x"947327ab",
  4686 => x"38768c2a",
  4687 => x"80ee0555",
  4688 => x"80d47327",
  4689 => x"9e38768f",
  4690 => x"2a80f705",
  4691 => x"5582d473",
  4692 => x"27913876",
  4693 => x"922a80fc",
  4694 => x"05558ad4",
  4695 => x"73278438",
  4696 => x"80fe5574",
  4697 => x"10101081",
  4698 => x"c7b40588",
  4699 => x"11085556",
  4700 => x"73762e82",
  4701 => x"b3388414",
  4702 => x"08fc0653",
  4703 => x"7673278d",
  4704 => x"38881408",
  4705 => x"5473762e",
  4706 => x"098106ea",
  4707 => x"388c1408",
  4708 => x"708c1a0c",
  4709 => x"74881a0c",
  4710 => x"7888120c",
  4711 => x"56778c15",
  4712 => x"0c7a51fc",
  4713 => x"883f8c3d",
  4714 => x"0d047708",
  4715 => x"78713159",
  4716 => x"77058819",
  4717 => x"08545772",
  4718 => x"81c7bc2e",
  4719 => x"80e0388c",
  4720 => x"1808708c",
  4721 => x"150c7388",
  4722 => x"120c56fe",
  4723 => x"89398815",
  4724 => x"088c1608",
  4725 => x"708c130c",
  4726 => x"5788170c",
  4727 => x"fea33976",
  4728 => x"832a7054",
  4729 => x"55807524",
  4730 => x"81983872",
  4731 => x"822c8171",
  4732 => x"2b81c7b8",
  4733 => x"080781c7",
  4734 => x"b40b8405",
  4735 => x"0c537410",
  4736 => x"101081c7",
  4737 => x"b4058811",
  4738 => x"08555675",
  4739 => x"8c190c73",
  4740 => x"88190c77",
  4741 => x"88170c77",
  4742 => x"8c150cff",
  4743 => x"8439815a",
  4744 => x"fdb43978",
  4745 => x"17738106",
  4746 => x"54577298",
  4747 => x"38770878",
  4748 => x"71315977",
  4749 => x"058c1908",
  4750 => x"881a0871",
  4751 => x"8c120c88",
  4752 => x"120c5757",
  4753 => x"76810784",
  4754 => x"190c7781",
  4755 => x"c7b40b88",
  4756 => x"050c81c7",
  4757 => x"b0087726",
  4758 => x"fec73881",
  4759 => x"c7ac0852",
  4760 => x"7a51fafe",
  4761 => x"3f7a51fa",
  4762 => x"c43ffeba",
  4763 => x"3981788c",
  4764 => x"150c7888",
  4765 => x"150c738c",
  4766 => x"1a0c7388",
  4767 => x"1a0c5afd",
  4768 => x"80398315",
  4769 => x"70822c81",
  4770 => x"712b81c7",
  4771 => x"b8080781",
  4772 => x"c7b40b84",
  4773 => x"050c5153",
  4774 => x"74101010",
  4775 => x"81c7b405",
  4776 => x"88110855",
  4777 => x"56fee439",
  4778 => x"74538075",
  4779 => x"24a73872",
  4780 => x"822c8171",
  4781 => x"2b81c7b8",
  4782 => x"080781c7",
  4783 => x"b40b8405",
  4784 => x"0c53758c",
  4785 => x"190c7388",
  4786 => x"190c7788",
  4787 => x"170c778c",
  4788 => x"150cfdcd",
  4789 => x"39831570",
  4790 => x"822c8171",
  4791 => x"2b81c7b8",
  4792 => x"080781c7",
  4793 => x"b40b8405",
  4794 => x"0c5153d6",
  4795 => x"39810bb0",
  4796 => x"0c04803d",
  4797 => x"0d72812e",
  4798 => x"8938800b",
  4799 => x"b00c823d",
  4800 => x"0d047351",
  4801 => x"b23ffe3d",
  4802 => x"0d81e3d0",
  4803 => x"0851708a",
  4804 => x"3881e3d8",
  4805 => x"7081e3d0",
  4806 => x"0c517075",
  4807 => x"125252ff",
  4808 => x"537087fb",
  4809 => x"80802688",
  4810 => x"387081e3",
  4811 => x"d00c7153",
  4812 => x"72b00c84",
  4813 => x"3d0d0400",
  4814 => x"ff390000",
  4815 => x"00000000",
  4816 => x"00000000",
  4817 => x"00000000",
  4818 => x"00000000",
  4819 => x"00cac5ca",
  4820 => x"c5c0c0c0",
  4821 => x"c0c0c0c0",
  4822 => x"c0c0c0cf",
  4823 => x"cfcfcf00",
  4824 => x"00000f0f",
  4825 => x"0f0f8f8f",
  4826 => x"cfcfcfcf",
  4827 => x"cfcf4f0f",
  4828 => x"0f0f0000",
  4829 => x"cfcfcfcf",
  4830 => x"0f0f0f0f",
  4831 => x"0f0f0f0f",
  4832 => x"0f0ffefe",
  4833 => x"fefc0000",
  4834 => x"cfcfcfcf",
  4835 => x"cfcfcfcf",
  4836 => x"cfcfcfcf",
  4837 => x"cfffff7e",
  4838 => x"7e000000",
  4839 => x"00000000",
  4840 => x"00000000",
  4841 => x"00000000",
  4842 => x"00003f3f",
  4843 => x"3f3f0101",
  4844 => x"01010101",
  4845 => x"01010101",
  4846 => x"3f3f3f3f",
  4847 => x"0000383c",
  4848 => x"3e3e3f3f",
  4849 => x"3f3b3b39",
  4850 => x"39383838",
  4851 => x"38383800",
  4852 => x"003f3f3f",
  4853 => x"3f383838",
  4854 => x"38383838",
  4855 => x"38383c3f",
  4856 => x"3f1f0f00",
  4857 => x"003f3f3f",
  4858 => x"3f030303",
  4859 => x"03030303",
  4860 => x"03033f3f",
  4861 => x"3f3e0000",
  4862 => x"00000000",
  4863 => x"00000000",
  4864 => x"00000000",
  4865 => x"00000000",
  4866 => x"00000000",
  4867 => x"00000000",
  4868 => x"00000000",
  4869 => x"00000000",
  4870 => x"00000000",
  4871 => x"00000000",
  4872 => x"00000000",
  4873 => x"00000000",
  4874 => x"00000000",
  4875 => x"00000000",
  4876 => x"00000000",
  4877 => x"00000000",
  4878 => x"00000000",
  4879 => x"00000000",
  4880 => x"00000000",
  4881 => x"00000000",
  4882 => x"00000000",
  4883 => x"00000000",
  4884 => x"00000000",
  4885 => x"00000000",
  4886 => x"8080c0c0",
  4887 => x"e0e06000",
  4888 => x"00000000",
  4889 => x"00000000",
  4890 => x"00000000",
  4891 => x"00000000",
  4892 => x"00000000",
  4893 => x"00000000",
  4894 => x"00000000",
  4895 => x"00000000",
  4896 => x"00000000",
  4897 => x"00000000",
  4898 => x"00000000",
  4899 => x"00000000",
  4900 => x"00000000",
  4901 => x"00000000",
  4902 => x"00000000",
  4903 => x"00000000",
  4904 => x"00000000",
  4905 => x"00000000",
  4906 => x"00000000",
  4907 => x"00000000",
  4908 => x"806098ee",
  4909 => x"77bbddec",
  4910 => x"ee6e0200",
  4911 => x"00000000",
  4912 => x"00e08080",
  4913 => x"e00000e0",
  4914 => x"a0a00000",
  4915 => x"e0000000",
  4916 => x"00e0c000",
  4917 => x"c0e00000",
  4918 => x"e08080e0",
  4919 => x"0000c020",
  4920 => x"20c00000",
  4921 => x"e0000000",
  4922 => x"20e02000",
  4923 => x"0020a060",
  4924 => x"20000000",
  4925 => x"00000000",
  4926 => x"00000000",
  4927 => x"00000000",
  4928 => x"00000000",
  4929 => x"00000000",
  4930 => x"00000000",
  4931 => x"00030007",
  4932 => x"00070701",
  4933 => x"00000000",
  4934 => x"00000000",
  4935 => x"00000300",
  4936 => x"c0030000",
  4937 => x"034242c0",
  4938 => x"00c34242",
  4939 => x"0000c380",
  4940 => x"01c00340",
  4941 => x"c04300c0",
  4942 => x"43408001",
  4943 => x"c20201c0",
  4944 => x"00c38202",
  4945 => x"80c00300",
  4946 => x"00c04342",
  4947 => x"8202c040",
  4948 => x"40800000",
  4949 => x"c0404000",
  4950 => x"80404000",
  4951 => x"00c04040",
  4952 => x"8000c040",
  4953 => x"4000c080",
  4954 => x"00c00000",
  4955 => x"00000000",
  4956 => x"00000000",
  4957 => x"00000000",
  4958 => x"00000000",
  4959 => x"00ff0000",
  4960 => x"0000c645",
  4961 => x"44800785",
  4962 => x"45408007",
  4963 => x"80424700",
  4964 => x"80474000",
  4965 => x"07c14344",
  4966 => x"00c38404",
  4967 => x"c30007c1",
  4968 => x"42418700",
  4969 => x"80404784",
  4970 => x"04c34047",
  4971 => x"8101c640",
  4972 => x"40070505",
  4973 => x"00040502",
  4974 => x"00000704",
  4975 => x"04030007",
  4976 => x"05050007",
  4977 => x"00020700",
  4978 => x"00000000",
  4979 => x"00000000",
  4980 => x"00000000",
  4981 => x"00000000",
  4982 => x"0000ff00",
  4983 => x"00000007",
  4984 => x"01030500",
  4985 => x"03040403",
  4986 => x"00040502",
  4987 => x"00040502",
  4988 => x"00000705",
  4989 => x"05000700",
  4990 => x"02070000",
  4991 => x"07040403",
  4992 => x"00030404",
  4993 => x"03000701",
  4994 => x"03050007",
  4995 => x"01010000",
  4996 => x"00000000",
  4997 => x"00000000",
  4998 => x"00000000",
  4999 => x"00000000",
  5000 => x"00000000",
  5001 => x"71756974",
  5002 => x"00000000",
  5003 => x"68656c70",
  5004 => x"00000000",
  5005 => x"30780000",
  5006 => x"0a307800",
  5007 => x"69326320",
  5008 => x"464d430a",
  5009 => x"00000000",
  5010 => x"61646472",
  5011 => x"6573733a",
  5012 => x"20307800",
  5013 => x"2020202d",
  5014 => x"2d3e2020",
  5015 => x"2041434b",
  5016 => x"0a000000",
  5017 => x"72656164",
  5018 => x"20646174",
  5019 => x"61202800",
  5020 => x"20627974",
  5021 => x"65732920",
  5022 => x"66726f6d",
  5023 => x"20493243",
  5024 => x"2d616464",
  5025 => x"72657373",
  5026 => x"20307800",
  5027 => x"0a0a0000",
  5028 => x"6e6f6163",
  5029 => x"6b200000",
  5030 => x"6368726f",
  5031 => x"6e74656c",
  5032 => x"20726567",
  5033 => x"20307800",
  5034 => x"3a203078",
  5035 => x"00000000",
  5036 => x"206e6163",
  5037 => x"6b000000",
  5038 => x"6572726f",
  5039 => x"7220286e",
  5040 => x"61636b29",
  5041 => x"0a000000",
  5042 => x"0a202063",
  5043 => x"68616e6e",
  5044 => x"656c2033",
  5045 => x"20696e70",
  5046 => x"7574206f",
  5047 => x"76657266",
  5048 => x"6c6f7700",
  5049 => x"0a202063",
  5050 => x"68616e6e",
  5051 => x"656c2032",
  5052 => x"20696e70",
  5053 => x"7574206f",
  5054 => x"76657266",
  5055 => x"6c6f7700",
  5056 => x"0a202063",
  5057 => x"68616e6e",
  5058 => x"656c2031",
  5059 => x"20696e70",
  5060 => x"7574206f",
  5061 => x"76657266",
  5062 => x"6c6f7700",
  5063 => x"0a202063",
  5064 => x"68616e6e",
  5065 => x"656c2030",
  5066 => x"20696e70",
  5067 => x"7574206f",
  5068 => x"76657266",
  5069 => x"6c6f7700",
  5070 => x"0a202063",
  5071 => x"68616e6e",
  5072 => x"656c2033",
  5073 => x"20717561",
  5074 => x"6473756d",
  5075 => x"206f7665",
  5076 => x"72666c6f",
  5077 => x"77000000",
  5078 => x"0a202063",
  5079 => x"68616e6e",
  5080 => x"656c2032",
  5081 => x"20717561",
  5082 => x"6473756d",
  5083 => x"206f7665",
  5084 => x"72666c6f",
  5085 => x"77000000",
  5086 => x"0a202063",
  5087 => x"68616e6e",
  5088 => x"656c2031",
  5089 => x"20717561",
  5090 => x"6473756d",
  5091 => x"206f7665",
  5092 => x"72666c6f",
  5093 => x"77000000",
  5094 => x"0a202063",
  5095 => x"68616e6e",
  5096 => x"656c2030",
  5097 => x"20717561",
  5098 => x"6473756d",
  5099 => x"206f7665",
  5100 => x"72666c6f",
  5101 => x"77000000",
  5102 => x"0a202073",
  5103 => x"756d2076",
  5104 => x"616c7565",
  5105 => x"20637574",
  5106 => x"74656400",
  5107 => x"0a202063",
  5108 => x"68616e6e",
  5109 => x"656c2033",
  5110 => x"20646976",
  5111 => x"6964656e",
  5112 => x"64206375",
  5113 => x"74746564",
  5114 => x"00000000",
  5115 => x"0a202063",
  5116 => x"68616e6e",
  5117 => x"656c2033",
  5118 => x"206e6f69",
  5119 => x"73652063",
  5120 => x"6f6d7065",
  5121 => x"6e736174",
  5122 => x"696f6e20",
  5123 => x"746f2062",
  5124 => x"69670000",
  5125 => x"0a202063",
  5126 => x"68616e6e",
  5127 => x"656c2033",
  5128 => x"206e6f69",
  5129 => x"73652076",
  5130 => x"616c7565",
  5131 => x"20637574",
  5132 => x"74656400",
  5133 => x"0a202063",
  5134 => x"68616e6e",
  5135 => x"656c2032",
  5136 => x"20646976",
  5137 => x"6964656e",
  5138 => x"64206375",
  5139 => x"74746564",
  5140 => x"00000000",
  5141 => x"0a202063",
  5142 => x"68616e6e",
  5143 => x"656c2032",
  5144 => x"206e6f69",
  5145 => x"73652063",
  5146 => x"6f6d7065",
  5147 => x"6e736174",
  5148 => x"696f6e20",
  5149 => x"746f2062",
  5150 => x"69670000",
  5151 => x"0a202063",
  5152 => x"68616e6e",
  5153 => x"656c2032",
  5154 => x"206e6f69",
  5155 => x"73652076",
  5156 => x"616c7565",
  5157 => x"20637574",
  5158 => x"74656400",
  5159 => x"0a202063",
  5160 => x"68616e6e",
  5161 => x"656c2031",
  5162 => x"20646976",
  5163 => x"6964656e",
  5164 => x"64206375",
  5165 => x"74746564",
  5166 => x"00000000",
  5167 => x"0a202063",
  5168 => x"68616e6e",
  5169 => x"656c2031",
  5170 => x"206e6f69",
  5171 => x"73652063",
  5172 => x"6f6d7065",
  5173 => x"6e736174",
  5174 => x"696f6e20",
  5175 => x"746f2062",
  5176 => x"69670000",
  5177 => x"0a202063",
  5178 => x"68616e6e",
  5179 => x"656c2031",
  5180 => x"206e6f69",
  5181 => x"73652076",
  5182 => x"616c7565",
  5183 => x"20637574",
  5184 => x"74656400",
  5185 => x"0a202063",
  5186 => x"68616e6e",
  5187 => x"656c2030",
  5188 => x"20646976",
  5189 => x"6964656e",
  5190 => x"64206375",
  5191 => x"74746564",
  5192 => x"00000000",
  5193 => x"0a202063",
  5194 => x"68616e6e",
  5195 => x"656c2030",
  5196 => x"206e6f69",
  5197 => x"73652063",
  5198 => x"6f6d7065",
  5199 => x"6e736174",
  5200 => x"696f6e20",
  5201 => x"746f2062",
  5202 => x"69670000",
  5203 => x"0a202063",
  5204 => x"68616e6e",
  5205 => x"656c2030",
  5206 => x"206e6f69",
  5207 => x"73652076",
  5208 => x"616c7565",
  5209 => x"20637574",
  5210 => x"74656400",
  5211 => x"0a202073",
  5212 => x"6f667477",
  5213 => x"61726520",
  5214 => x"6572726f",
  5215 => x"72000000",
  5216 => x"0a657874",
  5217 => x"65726e61",
  5218 => x"6c20636c",
  5219 => x"6f636b20",
  5220 => x"20202020",
  5221 => x"2020203a",
  5222 => x"20000000",
  5223 => x"61637469",
  5224 => x"76650000",
  5225 => x"0a6d6963",
  5226 => x"726f7075",
  5227 => x"6c736520",
  5228 => x"736f7572",
  5229 => x"63652020",
  5230 => x"2020203a",
  5231 => x"20000000",
  5232 => x"65787465",
  5233 => x"726e616c",
  5234 => x"00000000",
  5235 => x"0a6d6963",
  5236 => x"726f7075",
  5237 => x"6c736520",
  5238 => x"6576656e",
  5239 => x"74206c69",
  5240 => x"6d69743a",
  5241 => x"20000000",
  5242 => x"0a6d6561",
  5243 => x"73757265",
  5244 => x"6d656e74",
  5245 => x"206c656e",
  5246 => x"67746820",
  5247 => x"2020203a",
  5248 => x"20000000",
  5249 => x"0a626561",
  5250 => x"6d20706f",
  5251 => x"73697469",
  5252 => x"6f6e206d",
  5253 => x"6f6e6974",
  5254 => x"6f722072",
  5255 => x"65676973",
  5256 => x"74657273",
  5257 => x"00000000",
  5258 => x"0a202020",
  5259 => x"20202020",
  5260 => x"20202020",
  5261 => x"20202020",
  5262 => x"20202020",
  5263 => x"20202020",
  5264 => x"20636861",
  5265 => x"6e6e656c",
  5266 => x"20302020",
  5267 => x"20636861",
  5268 => x"6e6e656c",
  5269 => x"20312020",
  5270 => x"20636861",
  5271 => x"6e6e656c",
  5272 => x"20322020",
  5273 => x"20636861",
  5274 => x"6e6e656c",
  5275 => x"20330000",
  5276 => x"0a202020",
  5277 => x"20202020",
  5278 => x"20202020",
  5279 => x"20202020",
  5280 => x"20202020",
  5281 => x"20202020",
  5282 => x"202d2d2d",
  5283 => x"2d20686f",
  5284 => x"72697a6f",
  5285 => x"6e74616c",
  5286 => x"202d2d2d",
  5287 => x"2d2d2020",
  5288 => x"202d2d2d",
  5289 => x"2d2d2d20",
  5290 => x"76657274",
  5291 => x"6963616c",
  5292 => x"202d2d2d",
  5293 => x"2d2d0000",
  5294 => x"0a736361",
  5295 => x"6c657220",
  5296 => x"76616c75",
  5297 => x"65732020",
  5298 => x"20202020",
  5299 => x"20202020",
  5300 => x"20000000",
  5301 => x"0a6e6f69",
  5302 => x"73652063",
  5303 => x"6f6d7065",
  5304 => x"6e736174",
  5305 => x"696f6e20",
  5306 => x"20202020",
  5307 => x"20000000",
  5308 => x"0a6d6561",
  5309 => x"73757265",
  5310 => x"6d656e74",
  5311 => x"20202020",
  5312 => x"20202020",
  5313 => x"20202020",
  5314 => x"20000000",
  5315 => x"0a73616d",
  5316 => x"706c6573",
  5317 => x"20286469",
  5318 => x"7629203a",
  5319 => x"20000000",
  5320 => x"0a73756d",
  5321 => x"20636861",
  5322 => x"6e6e656c",
  5323 => x"2020203a",
  5324 => x"20000000",
  5325 => x"0a0a706f",
  5326 => x"73697469",
  5327 => x"6f6e2063",
  5328 => x"6f6d7075",
  5329 => x"74617469",
  5330 => x"6f6e0000",
  5331 => x"0a202073",
  5332 => x"63616c65",
  5333 => x"72207661",
  5334 => x"6c756573",
  5335 => x"20202020",
  5336 => x"20202020",
  5337 => x"20000000",
  5338 => x"0a20206f",
  5339 => x"66667365",
  5340 => x"74202020",
  5341 => x"20202020",
  5342 => x"20202020",
  5343 => x"20202020",
  5344 => x"20000000",
  5345 => x"0a6f7574",
  5346 => x"70757420",
  5347 => x"73656c65",
  5348 => x"6374203a",
  5349 => x"20000000",
  5350 => x"74657374",
  5351 => x"67656e00",
  5352 => x"4e4f5420",
  5353 => x"00000000",
  5354 => x"6368616e",
  5355 => x"6e656c20",
  5356 => x"30000000",
  5357 => x"0a63616c",
  5358 => x"63207374",
  5359 => x"61746520",
  5360 => x"2020203a",
  5361 => x"20307800",
  5362 => x"76657274",
  5363 => x"6963616c",
  5364 => x"00000000",
  5365 => x"686f7269",
  5366 => x"7a6f6e74",
  5367 => x"616c0000",
  5368 => x"73756d00",
  5369 => x"6368616e",
  5370 => x"6e656c20",
  5371 => x"33000000",
  5372 => x"6368616e",
  5373 => x"6e656c20",
  5374 => x"32000000",
  5375 => x"6368616e",
  5376 => x"6e656c20",
  5377 => x"31000000",
  5378 => x"786d6f64",
  5379 => x"656d2074",
  5380 => x"72616e73",
  5381 => x"6d69742e",
  5382 => x"2e2e0a00",
  5383 => x"20627974",
  5384 => x"65732074",
  5385 => x"72616e73",
  5386 => x"6d697474",
  5387 => x"65640a00",
  5388 => x"63616e63",
  5389 => x"656c0a00",
  5390 => x"72657472",
  5391 => x"79206f75",
  5392 => x"740a0000",
  5393 => x"786d6f64",
  5394 => x"656d2072",
  5395 => x"65636569",
  5396 => x"76652e2e",
  5397 => x"2e0a0000",
  5398 => x"20627974",
  5399 => x"65732072",
  5400 => x"65636569",
  5401 => x"7665640a",
  5402 => x"00000000",
  5403 => x"72782062",
  5404 => x"75666665",
  5405 => x"72206675",
  5406 => x"6c6c0a00",
  5407 => x"74696d65",
  5408 => x"206f7574",
  5409 => x"0a000000",
  5410 => x"64656275",
  5411 => x"67207265",
  5412 => x"67697374",
  5413 => x"65727300",
  5414 => x"0a6d6f64",
  5415 => x"65202020",
  5416 => x"20202020",
  5417 => x"203a2000",
  5418 => x"0a616464",
  5419 => x"72657373",
  5420 => x"20302020",
  5421 => x"203a2030",
  5422 => x"78000000",
  5423 => x"0a616464",
  5424 => x"72657373",
  5425 => x"20312020",
  5426 => x"203a2030",
  5427 => x"78000000",
  5428 => x"0a627566",
  5429 => x"66657220",
  5430 => x"73697a65",
  5431 => x"203a2000",
  5432 => x"6d61783a",
  5433 => x"20000000",
  5434 => x"6d696e3a",
  5435 => x"20000000",
  5436 => x"63683a20",
  5437 => x"00000000",
  5438 => x"73706c3a",
  5439 => x"20000000",
  5440 => x"73686f77",
  5441 => x"2042504d",
  5442 => x"20726567",
  5443 => x"69737465",
  5444 => x"72730000",
  5445 => x"62706d00",
  5446 => x"73656c65",
  5447 => x"6374206f",
  5448 => x"75747075",
  5449 => x"74206368",
  5450 => x"616e6e65",
  5451 => x"6c202830",
  5452 => x"2e2e3320",
  5453 => x"73756d20",
  5454 => x"68207629",
  5455 => x"00000000",
  5456 => x"73656c65",
  5457 => x"63740000",
  5458 => x"73797374",
  5459 => x"656d2072",
  5460 => x"65736574",
  5461 => x"00000000",
  5462 => x"72657365",
  5463 => x"74000000",
  5464 => x"73686f77",
  5465 => x"2f736574",
  5466 => x"20646562",
  5467 => x"75672072",
  5468 => x"65676973",
  5469 => x"74657273",
  5470 => x"203c7365",
  5471 => x"74206d6f",
  5472 => x"64653e00",
  5473 => x"64656275",
  5474 => x"67000000",
  5475 => x"636c6b20",
  5476 => x"736f7572",
  5477 => x"63653a20",
  5478 => x"2030203d",
  5479 => x"20696e74",
  5480 => x"2c203120",
  5481 => x"3d206578",
  5482 => x"74000000",
  5483 => x"636c6b00",
  5484 => x"6d696372",
  5485 => x"6f70756c",
  5486 => x"73652073",
  5487 => x"6f757263",
  5488 => x"653a2030",
  5489 => x"203d2069",
  5490 => x"6e742c20",
  5491 => x"31203d20",
  5492 => x"65787400",
  5493 => x"6d696372",
  5494 => x"6f000000",
  5495 => x"74657374",
  5496 => x"67656e65",
  5497 => x"7261746f",
  5498 => x"72203c73",
  5499 => x"63616c65",
  5500 => x"723e203c",
  5501 => x"72657374",
  5502 => x"6172743e",
  5503 => x"00000000",
  5504 => x"3c6d7574",
  5505 => x"655f6e3e",
  5506 => x"203c7273",
  5507 => x"745f6e3e",
  5508 => x"203c6270",
  5509 => x"625f6e3e",
  5510 => x"203c6f73",
  5511 => x"72313e20",
  5512 => x"3c6f7372",
  5513 => x"323e0000",
  5514 => x"64616363",
  5515 => x"6f6e6600",
  5516 => x"3c6d756c",
  5517 => x"7469706c",
  5518 => x"6965723e",
  5519 => x"20696e69",
  5520 => x"7469616c",
  5521 => x"697a6520",
  5522 => x"62756666",
  5523 => x"65720000",
  5524 => x"64616374",
  5525 => x"65737400",
  5526 => x"72657365",
  5527 => x"74206361",
  5528 => x"6c63756c",
  5529 => x"6174696f",
  5530 => x"6e206572",
  5531 => x"726f7273",
  5532 => x"00000000",
  5533 => x"63616c63",
  5534 => x"72657300",
  5535 => x"73686f77",
  5536 => x"20646562",
  5537 => x"75672062",
  5538 => x"75666665",
  5539 => x"72203c6c",
  5540 => x"656e6774",
  5541 => x"683e0000",
  5542 => x"636c6561",
  5543 => x"72206465",
  5544 => x"62756720",
  5545 => x"62756666",
  5546 => x"65720000",
  5547 => x"62636c65",
  5548 => x"61720000",
  5549 => x"62756666",
  5550 => x"6572206f",
  5551 => x"6e204c43",
  5552 => x"44203c63",
  5553 => x"683e203c",
  5554 => x"636f6d62",
  5555 => x"3e000000",
  5556 => x"73636f70",
  5557 => x"65000000",
  5558 => x"64656275",
  5559 => x"67207472",
  5560 => x"61636520",
  5561 => x"3c636c65",
  5562 => x"61723e00",
  5563 => x"74726163",
  5564 => x"65000000",
  5565 => x"73657475",
  5566 => x"70206368",
  5567 => x"616e6e65",
  5568 => x"6c207465",
  5569 => x"7374203c",
  5570 => x"63683e20",
  5571 => x"3c76616c",
  5572 => x"302e2e37",
  5573 => x"3e000000",
  5574 => x"63687465",
  5575 => x"73740000",
  5576 => x"72756e6e",
  5577 => x"696e6720",
  5578 => x"6c696768",
  5579 => x"74000000",
  5580 => x"72756e00",
  5581 => x"72756e20",
  5582 => x"64697370",
  5583 => x"6c617920",
  5584 => x"74657374",
  5585 => x"2066756e",
  5586 => x"6374696f",
  5587 => x"6e000000",
  5588 => x"64697370",
  5589 => x"6c617900",
  5590 => x"73657420",
  5591 => x"6261636b",
  5592 => x"6c696768",
  5593 => x"74203c30",
  5594 => x"2e2e3331",
  5595 => x"3e000000",
  5596 => x"6261636b",
  5597 => x"00000000",
  5598 => x"73686f77",
  5599 => x"206c6f67",
  5600 => x"6f206f6e",
  5601 => x"20676c63",
  5602 => x"64000000",
  5603 => x"6c6f676f",
  5604 => x"00000000",
  5605 => x"63686563",
  5606 => x"6b204932",
  5607 => x"43206164",
  5608 => x"64726573",
  5609 => x"73000000",
  5610 => x"69326300",
  5611 => x"72656164",
  5612 => x"20454550",
  5613 => x"524f4d20",
  5614 => x"3c627573",
  5615 => x"3e203c69",
  5616 => x"32635f61",
  5617 => x"6464723e",
  5618 => x"203c6c65",
  5619 => x"6e677468",
  5620 => x"3e000000",
  5621 => x"65657072",
  5622 => x"6f6d0000",
  5623 => x"41444320",
  5624 => x"72656769",
  5625 => x"73746572",
  5626 => x"20747261",
  5627 => x"6e736665",
  5628 => x"72203c76",
  5629 => x"616c7565",
  5630 => x"3e000000",
  5631 => x"61747261",
  5632 => x"6e730000",
  5633 => x"696e6974",
  5634 => x"20414443",
  5635 => x"20726567",
  5636 => x"69737465",
  5637 => x"72730000",
  5638 => x"61696e69",
  5639 => x"74000000",
  5640 => x"616c6961",
  5641 => x"7320666f",
  5642 => x"72207800",
  5643 => x"6d656d00",
  5644 => x"77726974",
  5645 => x"6520776f",
  5646 => x"7264203c",
  5647 => x"61646472",
  5648 => x"3e203c6c",
  5649 => x"656e6774",
  5650 => x"683e203c",
  5651 => x"76616c75",
  5652 => x"65287329",
  5653 => x"3e000000",
  5654 => x"776d656d",
  5655 => x"00000000",
  5656 => x"6558616d",
  5657 => x"696e6520",
  5658 => x"6d656d6f",
  5659 => x"7279203c",
  5660 => x"61646472",
  5661 => x"3e203c6c",
  5662 => x"656e6774",
  5663 => x"683e0000",
  5664 => x"636c6561",
  5665 => x"72207363",
  5666 => x"7265656e",
  5667 => x"00000000",
  5668 => x"636c6561",
  5669 => x"72000000",
  5670 => x"0a646562",
  5671 => x"75672074",
  5672 => x"72616365",
  5673 => x"206d656d",
  5674 => x"6f727900",
  5675 => x"0a74696d",
  5676 => x"65207374",
  5677 => x"616d7020",
  5678 => x"20202073",
  5679 => x"74617465",
  5680 => x"00000000",
  5681 => x"20203078",
  5682 => x"00000000",
  5683 => x"65787465",
  5684 => x"726e616c",
  5685 => x"20636c6f",
  5686 => x"636b2000",
  5687 => x"61637469",
  5688 => x"76650a00",
  5689 => x"73656c65",
  5690 => x"63746564",
  5691 => x"0a000000",
  5692 => x"6d696372",
  5693 => x"6f70756c",
  5694 => x"73652073",
  5695 => x"6f757263",
  5696 => x"653a2000",
  5697 => x"6265616d",
  5698 => x"20706f73",
  5699 => x"6974696f",
  5700 => x"6e206d6f",
  5701 => x"6e69746f",
  5702 => x"72000000",
  5703 => x"20286f6e",
  5704 => x"2073696d",
  5705 => x"290a0000",
  5706 => x"0a485720",
  5707 => x"73796e74",
  5708 => x"68657369",
  5709 => x"7a65643a",
  5710 => x"20000000",
  5711 => x"0a535720",
  5712 => x"636f6d70",
  5713 => x"696c6564",
  5714 => x"2020203a",
  5715 => x"20417567",
  5716 => x"20313620",
  5717 => x"32303131",
  5718 => x"20203134",
  5719 => x"3a30393a",
  5720 => x"30310000",
  5721 => x"0a737973",
  5722 => x"74656d20",
  5723 => x"636c6f63",
  5724 => x"6b20203a",
  5725 => x"20000000",
  5726 => x"204d487a",
  5727 => x"0a000000",
  5728 => x"44454255",
  5729 => x"47204d4f",
  5730 => x"44450000",
  5731 => x"204f4e0a",
  5732 => x"00000000",
  5733 => x"0000114f",
  5734 => x"000011b8",
  5735 => x"000011ad",
  5736 => x"000011a2",
  5737 => x"00001197",
  5738 => x"0000118d",
  5739 => x"00001183",
  5740 => x"000002c2",
  5741 => x"fc1902c4",
  5742 => x"fffefd3f",
  5743 => x"03e7fd3b",
  5744 => x"0000485d",
  5745 => x"999b4888",
  5746 => x"ffc4b7ce",
  5747 => x"6665b74e",
  5748 => x"3e200000",
  5749 => x"636f6d6d",
  5750 => x"616e6420",
  5751 => x"6e6f7420",
  5752 => x"666f756e",
  5753 => x"642e0a00",
  5754 => x"73757070",
  5755 => x"6f727465",
  5756 => x"6420636f",
  5757 => x"6d6d616e",
  5758 => x"64733a0a",
  5759 => x"0a000000",
  5760 => x"202d2000",
  5761 => x"04580808",
  5762 => x"20ff0000",
  5763 => x"00005a14",
  5764 => x"00005af4",
  5765 => x"02010305",
  5766 => x"05070501",
  5767 => x"03030505",
  5768 => x"02030104",
  5769 => x"05050505",
  5770 => x"05050505",
  5771 => x"05050101",
  5772 => x"04050404",
  5773 => x"07050505",
  5774 => x"05050505",
  5775 => x"05030405",
  5776 => x"05050505",
  5777 => x"05050505",
  5778 => x"05050505",
  5779 => x"05050503",
  5780 => x"04030505",
  5781 => x"02050504",
  5782 => x"05050405",
  5783 => x"04010204",
  5784 => x"02050404",
  5785 => x"05050404",
  5786 => x"04040507",
  5787 => x"05040404",
  5788 => x"02040500",
  5789 => x"04050200",
  5790 => x"04080303",
  5791 => x"04090003",
  5792 => x"06000000",
  5793 => x"00020204",
  5794 => x"04040400",
  5795 => x"04060003",
  5796 => x"05000000",
  5797 => x"00000404",
  5798 => x"05050204",
  5799 => x"05060305",
  5800 => x"04030705",
  5801 => x"04050303",
  5802 => x"02040502",
  5803 => x"03020405",
  5804 => x"06060604",
  5805 => x"05050505",
  5806 => x"05050504",
  5807 => x"04040404",
  5808 => x"03030303",
  5809 => x"05050505",
  5810 => x"05050505",
  5811 => x"05040404",
  5812 => x"04050404",
  5813 => x"04040404",
  5814 => x"04040503",
  5815 => x"04040404",
  5816 => x"02020303",
  5817 => x"04040404",
  5818 => x"04040405",
  5819 => x"04040404",
  5820 => x"04030303",
  5821 => x"00005f07",
  5822 => x"0007741c",
  5823 => x"771c172e",
  5824 => x"6a3e2b3a",
  5825 => x"06493608",
  5826 => x"36493036",
  5827 => x"49597648",
  5828 => x"073c4281",
  5829 => x"81423c0a",
  5830 => x"041f040a",
  5831 => x"08083e08",
  5832 => x"08806008",
  5833 => x"080840c0",
  5834 => x"300c033e",
  5835 => x"4141413e",
  5836 => x"44427f40",
  5837 => x"40466151",
  5838 => x"49462241",
  5839 => x"49493618",
  5840 => x"14127f10",
  5841 => x"27454545",
  5842 => x"393e4949",
  5843 => x"49300101",
  5844 => x"710d0336",
  5845 => x"49494936",
  5846 => x"06494929",
  5847 => x"1e36d008",
  5848 => x"14224114",
  5849 => x"14141414",
  5850 => x"41221408",
  5851 => x"02510906",
  5852 => x"3c4299a5",
  5853 => x"bd421c7c",
  5854 => x"1211127c",
  5855 => x"7f494949",
  5856 => x"363e4141",
  5857 => x"41227f41",
  5858 => x"41413e7f",
  5859 => x"49494941",
  5860 => x"7f090909",
  5861 => x"013e4149",
  5862 => x"497a7f08",
  5863 => x"08087f41",
  5864 => x"7f414041",
  5865 => x"413f7f08",
  5866 => x"1422417f",
  5867 => x"40404040",
  5868 => x"7f060c06",
  5869 => x"7f7f0608",
  5870 => x"307f3e41",
  5871 => x"41413e7f",
  5872 => x"09090906",
  5873 => x"3e4161c1",
  5874 => x"be7f0919",
  5875 => x"29462649",
  5876 => x"49493201",
  5877 => x"017f0101",
  5878 => x"3f404040",
  5879 => x"3f073840",
  5880 => x"38071f60",
  5881 => x"1f601f63",
  5882 => x"14081463",
  5883 => x"01067806",
  5884 => x"01615149",
  5885 => x"45437f41",
  5886 => x"41030c30",
  5887 => x"c041417f",
  5888 => x"04020102",
  5889 => x"04808080",
  5890 => x"80800102",
  5891 => x"20545454",
  5892 => x"787f4444",
  5893 => x"44383844",
  5894 => x"44443844",
  5895 => x"44447f38",
  5896 => x"54545458",
  5897 => x"087e0901",
  5898 => x"18a4a4a4",
  5899 => x"787f0404",
  5900 => x"787d807d",
  5901 => x"7f102844",
  5902 => x"3f407c04",
  5903 => x"7804787c",
  5904 => x"04047838",
  5905 => x"444438fc",
  5906 => x"24242418",
  5907 => x"18242424",
  5908 => x"fc7c0804",
  5909 => x"04485454",
  5910 => x"24043f44",
  5911 => x"403c4040",
  5912 => x"7c1c2040",
  5913 => x"201c1c60",
  5914 => x"601c6060",
  5915 => x"1c442810",
  5916 => x"28449ca0",
  5917 => x"601c6454",
  5918 => x"544c187e",
  5919 => x"8181ffff",
  5920 => x"81817e18",
  5921 => x"18040810",
  5922 => x"0c143e55",
  5923 => x"55ff8181",
  5924 => x"81ff8060",
  5925 => x"80608060",
  5926 => x"60600060",
  5927 => x"60006060",
  5928 => x"047f0414",
  5929 => x"7f140201",
  5930 => x"01024629",
  5931 => x"1608344a",
  5932 => x"31483000",
  5933 => x"18243e41",
  5934 => x"227f4941",
  5935 => x"03040403",
  5936 => x"03040304",
  5937 => x"04030403",
  5938 => x"183c3c18",
  5939 => x"08080808",
  5940 => x"03010203",
  5941 => x"020e020e",
  5942 => x"060e0048",
  5943 => x"30384438",
  5944 => x"54483844",
  5945 => x"fe44487e",
  5946 => x"49014438",
  5947 => x"28384403",
  5948 => x"147c1403",
  5949 => x"e7e74e55",
  5950 => x"55390101",
  5951 => x"0001011c",
  5952 => x"2a555522",
  5953 => x"1c1d151e",
  5954 => x"18240018",
  5955 => x"24080808",
  5956 => x"18080808",
  5957 => x"3c42bd95",
  5958 => x"a9423c01",
  5959 => x"01010101",
  5960 => x"06090906",
  5961 => x"44445f44",
  5962 => x"44191512",
  5963 => x"15150a02",
  5964 => x"01fc2020",
  5965 => x"1c0e7f01",
  5966 => x"7f011818",
  5967 => x"00804002",
  5968 => x"1f060909",
  5969 => x"06241800",
  5970 => x"2418824f",
  5971 => x"304c62f1",
  5972 => x"824f300c",
  5973 => x"d2b1955f",
  5974 => x"304c62f1",
  5975 => x"30484520",
  5976 => x"60392e38",
  5977 => x"6060382e",
  5978 => x"3960701d",
  5979 => x"131d7072",
  5980 => x"1d121e71",
  5981 => x"701d121d",
  5982 => x"70603b25",
  5983 => x"3b607e11",
  5984 => x"7f49411e",
  5985 => x"2161927c",
  5986 => x"5556447c",
  5987 => x"5655447c",
  5988 => x"5655467d",
  5989 => x"54544545",
  5990 => x"7e44447e",
  5991 => x"45467d46",
  5992 => x"457c4508",
  5993 => x"7f49413e",
  5994 => x"7e091222",
  5995 => x"7d384546",
  5996 => x"44383844",
  5997 => x"46453838",
  5998 => x"46454638",
  5999 => x"3a454546",
  6000 => x"39384544",
  6001 => x"45382214",
  6002 => x"081422bc",
  6003 => x"625a463d",
  6004 => x"3c41423c",
  6005 => x"3c42413c",
  6006 => x"3c42413e",
  6007 => x"3d40403d",
  6008 => x"0608f209",
  6009 => x"067f2222",
  6010 => x"1cfe0989",
  6011 => x"76205556",
  6012 => x"78205655",
  6013 => x"78225555",
  6014 => x"7a235556",
  6015 => x"7b205554",
  6016 => x"79275557",
  6017 => x"78205438",
  6018 => x"54483844",
  6019 => x"c4385556",
  6020 => x"58385655",
  6021 => x"583a5555",
  6022 => x"5a395454",
  6023 => x"59017a7a",
  6024 => x"01027902",
  6025 => x"02780260",
  6026 => x"91927c7b",
  6027 => x"090a7338",
  6028 => x"45463838",
  6029 => x"4645383a",
  6030 => x"45453a3b",
  6031 => x"45463b39",
  6032 => x"44443908",
  6033 => x"082a0808",
  6034 => x"b8644c3a",
  6035 => x"3c41427c",
  6036 => x"3c42417c",
  6037 => x"3a41417a",
  6038 => x"3d40407d",
  6039 => x"986219ff",
  6040 => x"423c9a60",
  6041 => x"1a000000",
  6042 => x"30622020",
  6043 => x"20202020",
  6044 => x"20202020",
  6045 => x"20202020",
  6046 => x"20202020",
  6047 => x"20202020",
  6048 => x"20202020",
  6049 => x"20202020",
  6050 => x"20200000",
  6051 => x"20202020",
  6052 => x"20202020",
  6053 => x"00000000",
  6054 => x"00202020",
  6055 => x"20202020",
  6056 => x"20202828",
  6057 => x"28282820",
  6058 => x"20202020",
  6059 => x"20202020",
  6060 => x"20202020",
  6061 => x"20202020",
  6062 => x"20881010",
  6063 => x"10101010",
  6064 => x"10101010",
  6065 => x"10101010",
  6066 => x"10040404",
  6067 => x"04040404",
  6068 => x"04040410",
  6069 => x"10101010",
  6070 => x"10104141",
  6071 => x"41414141",
  6072 => x"01010101",
  6073 => x"01010101",
  6074 => x"01010101",
  6075 => x"01010101",
  6076 => x"01010101",
  6077 => x"10101010",
  6078 => x"10104242",
  6079 => x"42424242",
  6080 => x"02020202",
  6081 => x"02020202",
  6082 => x"02020202",
  6083 => x"02020202",
  6084 => x"02020202",
  6085 => x"10101010",
  6086 => x"20000000",
  6087 => x"00000000",
  6088 => x"00000000",
  6089 => x"00000000",
  6090 => x"00000000",
  6091 => x"00000000",
  6092 => x"00000000",
  6093 => x"00000000",
  6094 => x"00000000",
  6095 => x"00000000",
  6096 => x"00000000",
  6097 => x"00000000",
  6098 => x"00000000",
  6099 => x"00000000",
  6100 => x"00000000",
  6101 => x"00000000",
  6102 => x"00000000",
  6103 => x"00000000",
  6104 => x"00000000",
  6105 => x"00000000",
  6106 => x"00000000",
  6107 => x"00000000",
  6108 => x"00000000",
  6109 => x"00000000",
  6110 => x"00000000",
  6111 => x"00000000",
  6112 => x"00000000",
  6113 => x"00000000",
  6114 => x"00000000",
  6115 => x"00000000",
  6116 => x"00000000",
  6117 => x"00000000",
  6118 => x"00000000",
  6119 => x"43000000",
  6120 => x"00000000",
  6121 => x"80000c00",
  6122 => x"80000b00",
  6123 => x"80000800",
  6124 => x"00000000",
  6125 => x"ff000000",
  6126 => x"00000000",
  6127 => x"00000000",
  6128 => x"00ffffff",
  6129 => x"ff00ffff",
  6130 => x"ffff00ff",
  6131 => x"ffffff00",
  6132 => x"00000000",
  6133 => x"00000000",
  6134 => x"80000a00",
  6135 => x"80000700",
  6136 => x"80000600",
  6137 => x"80000400",
  6138 => x"80000200",
  6139 => x"80000100",
  6140 => x"80000004",
  6141 => x"80000000",
  6142 => x"00005ffc",
  6143 => x"00000000",
  6144 => x"00006264",
  6145 => x"000062c0",
  6146 => x"0000631c",
  6147 => x"00000000",
  6148 => x"00000000",
  6149 => x"00000000",
  6150 => x"00000000",
  6151 => x"00000000",
  6152 => x"00000000",
  6153 => x"00000000",
  6154 => x"00000000",
  6155 => x"00000000",
  6156 => x"00005f9c",
  6157 => x"00000000",
  6158 => x"00000000",
  6159 => x"00000000",
  6160 => x"00000000",
  6161 => x"00000000",
  6162 => x"00000000",
  6163 => x"00000000",
  6164 => x"00000000",
  6165 => x"00000000",
  6166 => x"00000000",
  6167 => x"00000000",
  6168 => x"00000000",
  6169 => x"00000000",
  6170 => x"00000000",
  6171 => x"00000000",
  6172 => x"00000000",
  6173 => x"00000000",
  6174 => x"00000000",
  6175 => x"00000000",
  6176 => x"00000000",
  6177 => x"00000000",
  6178 => x"00000000",
  6179 => x"00000000",
  6180 => x"00000000",
  6181 => x"00000000",
  6182 => x"00000000",
  6183 => x"00000000",
  6184 => x"00000000",
  6185 => x"00000001",
  6186 => x"330eabcd",
  6187 => x"1234e66d",
  6188 => x"deec0005",
  6189 => x"000b0000",
  6190 => x"00000000",
  6191 => x"00000000",
  6192 => x"00000000",
  6193 => x"00000000",
  6194 => x"00000000",
  6195 => x"00000000",
  6196 => x"00000000",
  6197 => x"00000000",
  6198 => x"00000000",
  6199 => x"00000000",
  6200 => x"00000000",
  6201 => x"00000000",
  6202 => x"00000000",
  6203 => x"00000000",
  6204 => x"00000000",
  6205 => x"00000000",
  6206 => x"00000000",
  6207 => x"00000000",
  6208 => x"00000000",
  6209 => x"00000000",
  6210 => x"00000000",
  6211 => x"00000000",
  6212 => x"00000000",
  6213 => x"00000000",
  6214 => x"00000000",
  6215 => x"00000000",
  6216 => x"00000000",
  6217 => x"00000000",
  6218 => x"00000000",
  6219 => x"00000000",
  6220 => x"00000000",
  6221 => x"00000000",
  6222 => x"00000000",
  6223 => x"00000000",
  6224 => x"00000000",
  6225 => x"00000000",
  6226 => x"00000000",
  6227 => x"00000000",
  6228 => x"00000000",
  6229 => x"00000000",
  6230 => x"00000000",
  6231 => x"00000000",
  6232 => x"00000000",
  6233 => x"00000000",
  6234 => x"00000000",
  6235 => x"00000000",
  6236 => x"00000000",
  6237 => x"00000000",
  6238 => x"00000000",
  6239 => x"00000000",
  6240 => x"00000000",
  6241 => x"00000000",
  6242 => x"00000000",
  6243 => x"00000000",
  6244 => x"00000000",
  6245 => x"00000000",
  6246 => x"00000000",
  6247 => x"00000000",
  6248 => x"00000000",
  6249 => x"00000000",
  6250 => x"00000000",
  6251 => x"00000000",
  6252 => x"00000000",
  6253 => x"00000000",
  6254 => x"00000000",
  6255 => x"00000000",
  6256 => x"00000000",
  6257 => x"00000000",
  6258 => x"00000000",
  6259 => x"00000000",
  6260 => x"00000000",
  6261 => x"00000000",
  6262 => x"00000000",
  6263 => x"00000000",
  6264 => x"00000000",
  6265 => x"00000000",
  6266 => x"00000000",
  6267 => x"00000000",
  6268 => x"00000000",
  6269 => x"00000000",
  6270 => x"00000000",
  6271 => x"00000000",
  6272 => x"00000000",
  6273 => x"00000000",
  6274 => x"00000000",
  6275 => x"00000000",
  6276 => x"00000000",
  6277 => x"00000000",
  6278 => x"00000000",
  6279 => x"00000000",
  6280 => x"00000000",
  6281 => x"00000000",
  6282 => x"00000000",
  6283 => x"00000000",
  6284 => x"00000000",
  6285 => x"00000000",
  6286 => x"00000000",
  6287 => x"00000000",
  6288 => x"00000000",
  6289 => x"00000000",
  6290 => x"00000000",
  6291 => x"00000000",
  6292 => x"00000000",
  6293 => x"00000000",
  6294 => x"00000000",
  6295 => x"00000000",
  6296 => x"00000000",
  6297 => x"00000000",
  6298 => x"00000000",
  6299 => x"00000000",
  6300 => x"00000000",
  6301 => x"00000000",
  6302 => x"00000000",
  6303 => x"00000000",
  6304 => x"00000000",
  6305 => x"00000000",
  6306 => x"00000000",
  6307 => x"00000000",
  6308 => x"00000000",
  6309 => x"00000000",
  6310 => x"00000000",
  6311 => x"00000000",
  6312 => x"00000000",
  6313 => x"00000000",
  6314 => x"00000000",
  6315 => x"00000000",
  6316 => x"00000000",
  6317 => x"00000000",
  6318 => x"00000000",
  6319 => x"00000000",
  6320 => x"00000000",
  6321 => x"00000000",
  6322 => x"00000000",
  6323 => x"00000000",
  6324 => x"00000000",
  6325 => x"00000000",
  6326 => x"00000000",
  6327 => x"00000000",
  6328 => x"00000000",
  6329 => x"00000000",
  6330 => x"00000000",
  6331 => x"00000000",
  6332 => x"00000000",
  6333 => x"00000000",
  6334 => x"00000000",
  6335 => x"00000000",
  6336 => x"00000000",
  6337 => x"00000000",
  6338 => x"00000000",
  6339 => x"00000000",
  6340 => x"00000000",
  6341 => x"00000000",
  6342 => x"00000000",
  6343 => x"00000000",
  6344 => x"00000000",
  6345 => x"00000000",
  6346 => x"00000000",
  6347 => x"00000000",
  6348 => x"00000000",
  6349 => x"00000000",
  6350 => x"00000000",
  6351 => x"00000000",
  6352 => x"00000000",
  6353 => x"00000000",
  6354 => x"00000000",
  6355 => x"00000000",
  6356 => x"00000000",
  6357 => x"00000000",
  6358 => x"00000000",
  6359 => x"00000000",
  6360 => x"00000000",
  6361 => x"00000000",
  6362 => x"00000000",
  6363 => x"00000000",
  6364 => x"00000000",
  6365 => x"00000000",
  6366 => x"00000000",
  6367 => x"00000000",
  6368 => x"00000000",
  6369 => x"00000000",
  6370 => x"00000000",
  6371 => x"00000000",
  6372 => x"00000000",
  6373 => x"00000000",
  6374 => x"00000000",
  6375 => x"00000000",
  6376 => x"00000000",
  6377 => x"00000000",
  6378 => x"ffffffff",
  6379 => x"00000000",
  6380 => x"00020000",
  6381 => x"00000000",
  6382 => x"00000000",
  6383 => x"000063b4",
  6384 => x"000063b4",
  6385 => x"000063bc",
  6386 => x"000063bc",
  6387 => x"000063c4",
  6388 => x"000063c4",
  6389 => x"000063cc",
  6390 => x"000063cc",
  6391 => x"000063d4",
  6392 => x"000063d4",
  6393 => x"000063dc",
  6394 => x"000063dc",
  6395 => x"000063e4",
  6396 => x"000063e4",
  6397 => x"000063ec",
  6398 => x"000063ec",
  6399 => x"000063f4",
  6400 => x"000063f4",
  6401 => x"000063fc",
  6402 => x"000063fc",
  6403 => x"00006404",
  6404 => x"00006404",
  6405 => x"0000640c",
  6406 => x"0000640c",
  6407 => x"00006414",
  6408 => x"00006414",
  6409 => x"0000641c",
  6410 => x"0000641c",
  6411 => x"00006424",
  6412 => x"00006424",
  6413 => x"0000642c",
  6414 => x"0000642c",
  6415 => x"00006434",
  6416 => x"00006434",
  6417 => x"0000643c",
  6418 => x"0000643c",
  6419 => x"00006444",
  6420 => x"00006444",
  6421 => x"0000644c",
  6422 => x"0000644c",
  6423 => x"00006454",
  6424 => x"00006454",
  6425 => x"0000645c",
  6426 => x"0000645c",
  6427 => x"00006464",
  6428 => x"00006464",
  6429 => x"0000646c",
  6430 => x"0000646c",
  6431 => x"00006474",
  6432 => x"00006474",
  6433 => x"0000647c",
  6434 => x"0000647c",
  6435 => x"00006484",
  6436 => x"00006484",
  6437 => x"0000648c",
  6438 => x"0000648c",
  6439 => x"00006494",
  6440 => x"00006494",
  6441 => x"0000649c",
  6442 => x"0000649c",
  6443 => x"000064a4",
  6444 => x"000064a4",
  6445 => x"000064ac",
  6446 => x"000064ac",
  6447 => x"000064b4",
  6448 => x"000064b4",
  6449 => x"000064bc",
  6450 => x"000064bc",
  6451 => x"000064c4",
  6452 => x"000064c4",
  6453 => x"000064cc",
  6454 => x"000064cc",
  6455 => x"000064d4",
  6456 => x"000064d4",
  6457 => x"000064dc",
  6458 => x"000064dc",
  6459 => x"000064e4",
  6460 => x"000064e4",
  6461 => x"000064ec",
  6462 => x"000064ec",
  6463 => x"000064f4",
  6464 => x"000064f4",
  6465 => x"000064fc",
  6466 => x"000064fc",
  6467 => x"00006504",
  6468 => x"00006504",
  6469 => x"0000650c",
  6470 => x"0000650c",
  6471 => x"00006514",
  6472 => x"00006514",
  6473 => x"0000651c",
  6474 => x"0000651c",
  6475 => x"00006524",
  6476 => x"00006524",
  6477 => x"0000652c",
  6478 => x"0000652c",
  6479 => x"00006534",
  6480 => x"00006534",
  6481 => x"0000653c",
  6482 => x"0000653c",
  6483 => x"00006544",
  6484 => x"00006544",
  6485 => x"0000654c",
  6486 => x"0000654c",
  6487 => x"00006554",
  6488 => x"00006554",
  6489 => x"0000655c",
  6490 => x"0000655c",
  6491 => x"00006564",
  6492 => x"00006564",
  6493 => x"0000656c",
  6494 => x"0000656c",
  6495 => x"00006574",
  6496 => x"00006574",
  6497 => x"0000657c",
  6498 => x"0000657c",
  6499 => x"00006584",
  6500 => x"00006584",
  6501 => x"0000658c",
  6502 => x"0000658c",
  6503 => x"00006594",
  6504 => x"00006594",
  6505 => x"0000659c",
  6506 => x"0000659c",
  6507 => x"000065a4",
  6508 => x"000065a4",
  6509 => x"000065ac",
  6510 => x"000065ac",
  6511 => x"000065b4",
  6512 => x"000065b4",
  6513 => x"000065bc",
  6514 => x"000065bc",
  6515 => x"000065c4",
  6516 => x"000065c4",
  6517 => x"000065cc",
  6518 => x"000065cc",
  6519 => x"000065d4",
  6520 => x"000065d4",
  6521 => x"000065dc",
  6522 => x"000065dc",
  6523 => x"000065e4",
  6524 => x"000065e4",
  6525 => x"000065ec",
  6526 => x"000065ec",
  6527 => x"000065f4",
  6528 => x"000065f4",
  6529 => x"000065fc",
  6530 => x"000065fc",
  6531 => x"00006604",
  6532 => x"00006604",
  6533 => x"0000660c",
  6534 => x"0000660c",
  6535 => x"00006614",
  6536 => x"00006614",
  6537 => x"0000661c",
  6538 => x"0000661c",
  6539 => x"00006624",
  6540 => x"00006624",
  6541 => x"0000662c",
  6542 => x"0000662c",
  6543 => x"00006634",
  6544 => x"00006634",
  6545 => x"0000663c",
  6546 => x"0000663c",
  6547 => x"00006644",
  6548 => x"00006644",
  6549 => x"0000664c",
  6550 => x"0000664c",
  6551 => x"00006654",
  6552 => x"00006654",
  6553 => x"0000665c",
  6554 => x"0000665c",
  6555 => x"00006664",
  6556 => x"00006664",
  6557 => x"0000666c",
  6558 => x"0000666c",
  6559 => x"00006674",
  6560 => x"00006674",
  6561 => x"0000667c",
  6562 => x"0000667c",
  6563 => x"00006684",
  6564 => x"00006684",
  6565 => x"0000668c",
  6566 => x"0000668c",
  6567 => x"00006694",
  6568 => x"00006694",
  6569 => x"0000669c",
  6570 => x"0000669c",
  6571 => x"000066a4",
  6572 => x"000066a4",
  6573 => x"000066ac",
  6574 => x"000066ac",
  6575 => x"000066b4",
  6576 => x"000066b4",
  6577 => x"000066bc",
  6578 => x"000066bc",
  6579 => x"000066c4",
  6580 => x"000066c4",
  6581 => x"000066cc",
  6582 => x"000066cc",
  6583 => x"000066d4",
  6584 => x"000066d4",
  6585 => x"000066dc",
  6586 => x"000066dc",
  6587 => x"000066e4",
  6588 => x"000066e4",
  6589 => x"000066ec",
  6590 => x"000066ec",
  6591 => x"000066f4",
  6592 => x"000066f4",
  6593 => x"000066fc",
  6594 => x"000066fc",
  6595 => x"00006704",
  6596 => x"00006704",
  6597 => x"0000670c",
  6598 => x"0000670c",
  6599 => x"00006714",
  6600 => x"00006714",
  6601 => x"0000671c",
  6602 => x"0000671c",
  6603 => x"00006724",
  6604 => x"00006724",
  6605 => x"0000672c",
  6606 => x"0000672c",
  6607 => x"00006734",
  6608 => x"00006734",
  6609 => x"0000673c",
  6610 => x"0000673c",
  6611 => x"00006744",
  6612 => x"00006744",
  6613 => x"0000674c",
  6614 => x"0000674c",
  6615 => x"00006754",
  6616 => x"00006754",
  6617 => x"0000675c",
  6618 => x"0000675c",
  6619 => x"00006764",
  6620 => x"00006764",
  6621 => x"0000676c",
  6622 => x"0000676c",
  6623 => x"00006774",
  6624 => x"00006774",
  6625 => x"0000677c",
  6626 => x"0000677c",
  6627 => x"00006784",
  6628 => x"00006784",
  6629 => x"0000678c",
  6630 => x"0000678c",
  6631 => x"00006794",
  6632 => x"00006794",
  6633 => x"0000679c",
  6634 => x"0000679c",
  6635 => x"000067a4",
  6636 => x"000067a4",
  6637 => x"000067ac",
  6638 => x"000067ac",
	--others => x"aaaaaaaa" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
