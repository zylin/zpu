library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dram is
port (clk : in std_logic;
		mem_writeEnable : in std_logic;
		mem_readEnable : in std_logic;
		mem_addr : in std_logic_vector(maxAddrBit downto 0);
		mem_write : in std_logic_vector(wordSize-1 downto 0);
		mem_read : out std_logic_vector(wordSize-1 downto 0);
		mem_busy : out std_logic;
		mem_writeMask : in std_logic_vector(wordBytes-1 downto 0));
end dram;

architecture dram_arch of dram is


type ram_type is array(0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"0b0b0b0b",
1 => x"80700b0b",
2 => x"80d3900c",
3 => x"3a0b0b80",
4 => x"c8b20400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"80c8fb2d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80d2",
162 => x"fc738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0b8d",
171 => x"872d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0b8d",
179 => x"cb2d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80d38c0c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"83d93f80",
257 => x"ca953f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"ff3d0d0b",
281 => x"0b80e2f8",
282 => x"08528412",
283 => x"08708106",
284 => x"515170f6",
285 => x"38710881",
286 => x"ff06800c",
287 => x"833d0d04",
288 => x"ff3d0d0b",
289 => x"0b80e2f8",
290 => x"08528412",
291 => x"08700a10",
292 => x"0a708106",
293 => x"51515170",
294 => x"f1387372",
295 => x"0c833d0d",
296 => x"0480d38c",
297 => x"08802ea8",
298 => x"38838080",
299 => x"0b0b0b80",
300 => x"e2f80c82",
301 => x"a0800b0b",
302 => x"0b80e2fc",
303 => x"0c829080",
304 => x"0b80e38c",
305 => x"0c0b0b80",
306 => x"e3800b80",
307 => x"e3900c04",
308 => x"f8808080",
309 => x"a40b0b0b",
310 => x"80e2f80c",
311 => x"f8808082",
312 => x"800b0b0b",
313 => x"80e2fc0c",
314 => x"f8808084",
315 => x"800b80e3",
316 => x"8c0cf880",
317 => x"8080940b",
318 => x"80e3900c",
319 => x"f8808080",
320 => x"9c0b80e3",
321 => x"880cf880",
322 => x"8080a00b",
323 => x"80e3940c",
324 => x"04f23d0d",
325 => x"600b0b80",
326 => x"e2fc0856",
327 => x"5d82750c",
328 => x"8059805a",
329 => x"800b8f3d",
330 => x"71101017",
331 => x"70085957",
332 => x"5d5b8076",
333 => x"81ff067c",
334 => x"832b5658",
335 => x"5276537b",
336 => x"5181fa3f",
337 => x"7d7f7a72",
338 => x"077c7207",
339 => x"71716081",
340 => x"05415f5d",
341 => x"5b595755",
342 => x"7a8724bb",
343 => x"380b0b80",
344 => x"e2fc087b",
345 => x"10101170",
346 => x"08585155",
347 => x"807681ff",
348 => x"067c832b",
349 => x"56585276",
350 => x"537b5181",
351 => x"c03f7d7f",
352 => x"7a72077c",
353 => x"72077171",
354 => x"60810541",
355 => x"5f5d5b59",
356 => x"5755877b",
357 => x"25c73876",
358 => x"7d0c7784",
359 => x"1e0c7c80",
360 => x"0c903d0d",
361 => x"04ff3d0d",
362 => x"80e38433",
363 => x"5170a738",
364 => x"80d39808",
365 => x"70085252",
366 => x"70802e94",
367 => x"38841280",
368 => x"d3980c70",
369 => x"2d80d398",
370 => x"08700852",
371 => x"5270ee38",
372 => x"810b80e3",
373 => x"8434833d",
374 => x"0d040480",
375 => x"3d0d0b0b",
376 => x"80e2f408",
377 => x"802e8e38",
378 => x"0b0b0b0b",
379 => x"800b802e",
380 => x"09810685",
381 => x"38823d0d",
382 => x"040b0b80",
383 => x"e2f4510b",
384 => x"0b0bf3fc",
385 => x"3f823d0d",
386 => x"0404fe3d",
387 => x"0d89530b",
388 => x"0b80d2c8",
389 => x"51838d3f",
390 => x"0b0b80d2",
391 => x"d8518384",
392 => x"3f810a0b",
393 => x"80e3980c",
394 => x"ff0b80e3",
395 => x"9c0cff13",
396 => x"53728025",
397 => x"da387280",
398 => x"0c843d0d",
399 => x"04f93d0d",
400 => x"797b7d7f",
401 => x"56545254",
402 => x"72802ea0",
403 => x"38705771",
404 => x"58a07331",
405 => x"52807225",
406 => x"a1387770",
407 => x"742b5770",
408 => x"732a7875",
409 => x"2b075651",
410 => x"74765351",
411 => x"70740c71",
412 => x"84150c73",
413 => x"800c893d",
414 => x"0d048056",
415 => x"7772302b",
416 => x"55747653",
417 => x"51e639fb",
418 => x"3d0d7779",
419 => x"55558056",
420 => x"757524ab",
421 => x"38807424",
422 => x"9d388053",
423 => x"73527451",
424 => x"80e13f80",
425 => x"08547580",
426 => x"2e853880",
427 => x"08305473",
428 => x"800c873d",
429 => x"0d047330",
430 => x"76813257",
431 => x"54dc3974",
432 => x"30558156",
433 => x"738025d2",
434 => x"38ec39fa",
435 => x"3d0d787a",
436 => x"57558057",
437 => x"767524a4",
438 => x"38759f2c",
439 => x"54815375",
440 => x"74327431",
441 => x"5274519b",
442 => x"3f800854",
443 => x"76802e85",
444 => x"38800830",
445 => x"5473800c",
446 => x"883d0d04",
447 => x"74305581",
448 => x"57d739fc",
449 => x"3d0d7678",
450 => x"53548153",
451 => x"80747326",
452 => x"52557280",
453 => x"2e983870",
454 => x"802eab38",
455 => x"807224a6",
456 => x"38711073",
457 => x"10757226",
458 => x"53545272",
459 => x"ea387351",
460 => x"78833874",
461 => x"5170800c",
462 => x"863d0d04",
463 => x"720a100a",
464 => x"720a100a",
465 => x"53537280",
466 => x"2ee43871",
467 => x"7426ed38",
468 => x"73723175",
469 => x"7407740a",
470 => x"100a740a",
471 => x"100a5555",
472 => x"5654e339",
473 => x"f73d0d7c",
474 => x"70525380",
475 => x"f93f7254",
476 => x"80085580",
477 => x"d2e85681",
478 => x"57800881",
479 => x"055a8b3d",
480 => x"e4115953",
481 => x"8259f413",
482 => x"527b8811",
483 => x"08525381",
484 => x"b03f8008",
485 => x"30708008",
486 => x"079f2c8a",
487 => x"07800c53",
488 => x"8b3d0d04",
489 => x"f63d0d7c",
490 => x"80d39c08",
491 => x"71535553",
492 => x"b53f7255",
493 => x"80085680",
494 => x"d2e85781",
495 => x"58800881",
496 => x"055b8c3d",
497 => x"e4115a53",
498 => x"825af413",
499 => x"52881408",
500 => x"5180ee3f",
501 => x"80083070",
502 => x"8008079f",
503 => x"2c8a0780",
504 => x"0c548c3d",
505 => x"0d04fd3d",
506 => x"0d757071",
507 => x"83065355",
508 => x"5270b438",
509 => x"71700870",
510 => x"09f7fbfd",
511 => x"ff1206f8",
512 => x"84828180",
513 => x"06545253",
514 => x"719b3884",
515 => x"13700870",
516 => x"09f7fbfd",
517 => x"ff1206f8",
518 => x"84828180",
519 => x"06545253",
520 => x"71802ee7",
521 => x"38725271",
522 => x"33537280",
523 => x"2e8a3881",
524 => x"12703354",
525 => x"5272f838",
526 => x"71743180",
527 => x"0c853d0d",
528 => x"04f23d0d",
529 => x"60628811",
530 => x"08705856",
531 => x"5f5a7380",
532 => x"2e818c38",
533 => x"8c1a2270",
534 => x"832a8132",
535 => x"81065658",
536 => x"74863890",
537 => x"1a089138",
538 => x"795190b7",
539 => x"3fff5580",
540 => x"0880ec38",
541 => x"8c1a2258",
542 => x"7d085580",
543 => x"7883ffff",
544 => x"06700a10",
545 => x"0a810641",
546 => x"5c577e77",
547 => x"2e80d738",
548 => x"76903874",
549 => x"08841608",
550 => x"88175758",
551 => x"5676802e",
552 => x"f2387654",
553 => x"88807727",
554 => x"84388880",
555 => x"54735375",
556 => x"529c1a08",
557 => x"51a41a08",
558 => x"58772d80",
559 => x"0b800825",
560 => x"82e03880",
561 => x"08167780",
562 => x"08317f88",
563 => x"05088008",
564 => x"31706188",
565 => x"050c5b58",
566 => x"5678ffb4",
567 => x"38805574",
568 => x"800c903d",
569 => x"0d047a81",
570 => x"32810677",
571 => x"40567580",
572 => x"2e81bd38",
573 => x"76903874",
574 => x"08841608",
575 => x"88175758",
576 => x"5976802e",
577 => x"f238881a",
578 => x"087883ff",
579 => x"ff067089",
580 => x"2a810656",
581 => x"59567380",
582 => x"2e82f838",
583 => x"7577278b",
584 => x"3877872a",
585 => x"81065c7b",
586 => x"82b53876",
587 => x"76278338",
588 => x"76567553",
589 => x"78527908",
590 => x"5185833f",
591 => x"881a0876",
592 => x"31881b0c",
593 => x"7908167a",
594 => x"0c765675",
595 => x"19777731",
596 => x"7f880508",
597 => x"78317061",
598 => x"88050c41",
599 => x"58597e80",
600 => x"2efefa38",
601 => x"8c1a2258",
602 => x"ff8a3978",
603 => x"79547c53",
604 => x"7b525684",
605 => x"c93f881a",
606 => x"08793188",
607 => x"1b0c7908",
608 => x"197a0c7c",
609 => x"76315d7c",
610 => x"8e387951",
611 => x"8ff23f80",
612 => x"08818f38",
613 => x"80085f75",
614 => x"1c777731",
615 => x"7f880508",
616 => x"78317061",
617 => x"88050c5d",
618 => x"585c7a80",
619 => x"2efeae38",
620 => x"76818338",
621 => x"74088416",
622 => x"08881757",
623 => x"585c7680",
624 => x"2ef23876",
625 => x"538a527b",
626 => x"5182d33f",
627 => x"80087c31",
628 => x"81055d80",
629 => x"08843881",
630 => x"175d815f",
631 => x"7c59767d",
632 => x"27833876",
633 => x"59941a08",
634 => x"881b0811",
635 => x"5758807a",
636 => x"085c5490",
637 => x"1a087b27",
638 => x"83388154",
639 => x"75792584",
640 => x"3873ba38",
641 => x"777924fe",
642 => x"e2387753",
643 => x"7b529c1a",
644 => x"0851a41a",
645 => x"0859782d",
646 => x"80085680",
647 => x"088024fe",
648 => x"e2388c1a",
649 => x"2280c007",
650 => x"5e7d8c1b",
651 => x"23ff5574",
652 => x"800c903d",
653 => x"0d047eff",
654 => x"a338ff87",
655 => x"3975537b",
656 => x"527a5182",
657 => x"f93f7908",
658 => x"167a0c79",
659 => x"518eb13f",
660 => x"8008cf38",
661 => x"7c76315d",
662 => x"7cfebc38",
663 => x"feac3990",
664 => x"1a087a08",
665 => x"71317811",
666 => x"70565a57",
667 => x"5280d39c",
668 => x"08518494",
669 => x"3f800880",
670 => x"2effa738",
671 => x"8008901b",
672 => x"0c800816",
673 => x"7a0c7794",
674 => x"1b0c7688",
675 => x"1b0c7656",
676 => x"fd993979",
677 => x"0858901a",
678 => x"08782783",
679 => x"38815475",
680 => x"77278438",
681 => x"73b33894",
682 => x"1a085473",
683 => x"772680d3",
684 => x"38735378",
685 => x"529c1a08",
686 => x"51a41a08",
687 => x"58772d80",
688 => x"08568008",
689 => x"8024fd83",
690 => x"388c1a22",
691 => x"80c0075e",
692 => x"7d8c1b23",
693 => x"ff55fed7",
694 => x"39755378",
695 => x"52775181",
696 => x"dd3f7908",
697 => x"167a0c79",
698 => x"518d953f",
699 => x"8008802e",
700 => x"fcd9388c",
701 => x"1a2280c0",
702 => x"075e7d8c",
703 => x"1b23ff55",
704 => x"fead3976",
705 => x"77547953",
706 => x"78525681",
707 => x"b13f881a",
708 => x"08773188",
709 => x"1b0c7908",
710 => x"177a0cfc",
711 => x"ae39fa3d",
712 => x"0d7a7902",
713 => x"8805a705",
714 => x"33555354",
715 => x"83742780",
716 => x"df387183",
717 => x"06517080",
718 => x"d7387171",
719 => x"57558351",
720 => x"75828029",
721 => x"13ff1252",
722 => x"56708025",
723 => x"f3388374",
724 => x"27bc3874",
725 => x"08763270",
726 => x"09f7fbfd",
727 => x"ff1206f8",
728 => x"84828180",
729 => x"06515170",
730 => x"802e9838",
731 => x"74518052",
732 => x"70335772",
733 => x"772eb938",
734 => x"81118113",
735 => x"53518372",
736 => x"27ee38fc",
737 => x"14841656",
738 => x"54738326",
739 => x"c6387452",
740 => x"ff145170",
741 => x"ff2e9738",
742 => x"71335472",
743 => x"742e9838",
744 => x"8112ff12",
745 => x"525270ff",
746 => x"2e098106",
747 => x"eb388051",
748 => x"70800c88",
749 => x"3d0d0471",
750 => x"800c883d",
751 => x"0d04fa3d",
752 => x"0d787a7c",
753 => x"72727259",
754 => x"57555856",
755 => x"57747727",
756 => x"b2387515",
757 => x"51767127",
758 => x"aa387076",
759 => x"18ff1853",
760 => x"535370ff",
761 => x"2e9638ff",
762 => x"12ff1454",
763 => x"52723372",
764 => x"34ff1151",
765 => x"70ff2e09",
766 => x"8106ec38",
767 => x"76800c88",
768 => x"3d0d048f",
769 => x"762780e6",
770 => x"38747707",
771 => x"83065170",
772 => x"80dc3876",
773 => x"75525370",
774 => x"70840552",
775 => x"08737084",
776 => x"05550c72",
777 => x"71708405",
778 => x"53087170",
779 => x"8405530c",
780 => x"71708405",
781 => x"53087170",
782 => x"8405530c",
783 => x"71708405",
784 => x"53087170",
785 => x"8405530c",
786 => x"f0155553",
787 => x"738f26c7",
788 => x"38837427",
789 => x"95387070",
790 => x"84055208",
791 => x"73708405",
792 => x"550cfc14",
793 => x"54738326",
794 => x"ed387271",
795 => x"5452ff14",
796 => x"5170ff2e",
797 => x"ff863872",
798 => x"70810554",
799 => x"33727081",
800 => x"055434ff",
801 => x"1151ea39",
802 => x"ef3d0d63",
803 => x"6567405d",
804 => x"427b802e",
805 => x"85823861",
806 => x"51a9eb3f",
807 => x"f81c7084",
808 => x"120870fc",
809 => x"0670628b",
810 => x"0570f806",
811 => x"4159455c",
812 => x"5f415796",
813 => x"742782c5",
814 => x"38807b24",
815 => x"7e7c2607",
816 => x"58805477",
817 => x"742e0981",
818 => x"0682ab38",
819 => x"787b2581",
820 => x"fe387817",
821 => x"80dad80b",
822 => x"8805085b",
823 => x"5679762e",
824 => x"84c53884",
825 => x"160870fe",
826 => x"06178411",
827 => x"08810641",
828 => x"55557e82",
829 => x"8d3874fc",
830 => x"06587976",
831 => x"2e84e338",
832 => x"78185f7e",
833 => x"7b2581ff",
834 => x"387c8106",
835 => x"547382c1",
836 => x"38767708",
837 => x"31841108",
838 => x"fc065657",
839 => x"75802e91",
840 => x"3879762e",
841 => x"84f03874",
842 => x"18195877",
843 => x"7b258491",
844 => x"3876802e",
845 => x"829b3878",
846 => x"15567a76",
847 => x"24829238",
848 => x"8c170888",
849 => x"1808718c",
850 => x"120c8812",
851 => x"0c5e7559",
852 => x"881761fc",
853 => x"055b5679",
854 => x"a42685ff",
855 => x"387b7659",
856 => x"55937a27",
857 => x"80c9387b",
858 => x"7084055d",
859 => x"087c5676",
860 => x"0c747084",
861 => x"0556088c",
862 => x"180c9017",
863 => x"589b7a27",
864 => x"ae387470",
865 => x"84055608",
866 => x"780c7470",
867 => x"84055608",
868 => x"94180c98",
869 => x"1758a37a",
870 => x"27953874",
871 => x"70840556",
872 => x"08780c74",
873 => x"70840556",
874 => x"089c180c",
875 => x"a0175874",
876 => x"70840556",
877 => x"08755f78",
878 => x"7084055a",
879 => x"0c777e70",
880 => x"84054008",
881 => x"71708405",
882 => x"530c7e08",
883 => x"710c5d78",
884 => x"7b315675",
885 => x"8f2680c9",
886 => x"38841708",
887 => x"81067907",
888 => x"84180c78",
889 => x"17841108",
890 => x"81078412",
891 => x"0c5b6151",
892 => x"a7953f88",
893 => x"17547380",
894 => x"0c933d0d",
895 => x"04905bfd",
896 => x"b8397756",
897 => x"fe83398c",
898 => x"16088817",
899 => x"08718c12",
900 => x"0c88120c",
901 => x"587e707c",
902 => x"3157598f",
903 => x"7627ffb9",
904 => x"387a1784",
905 => x"18088106",
906 => x"7c078419",
907 => x"0c768107",
908 => x"84120c76",
909 => x"11841108",
910 => x"81078412",
911 => x"0c5b8805",
912 => x"5261518f",
913 => x"de3f6151",
914 => x"a6bd3f88",
915 => x"1754ffa6",
916 => x"397d5261",
917 => x"5197db3f",
918 => x"80085a80",
919 => x"08802e81",
920 => x"ab388008",
921 => x"f8056084",
922 => x"0508fe06",
923 => x"61055855",
924 => x"74772e83",
925 => x"f238fc19",
926 => x"5877a426",
927 => x"81b0387b",
928 => x"80085657",
929 => x"93782780",
930 => x"dc387b70",
931 => x"70840552",
932 => x"08800870",
933 => x"8405800c",
934 => x"0c800871",
935 => x"70840553",
936 => x"085d567b",
937 => x"76708405",
938 => x"580c579b",
939 => x"7827b638",
940 => x"76708405",
941 => x"58087570",
942 => x"8405570c",
943 => x"76708405",
944 => x"58087570",
945 => x"8405570c",
946 => x"a3782799",
947 => x"38767084",
948 => x"05580875",
949 => x"70840557",
950 => x"0c767084",
951 => x"05580875",
952 => x"70840557",
953 => x"0c767084",
954 => x"05580877",
955 => x"5e757084",
956 => x"05570c74",
957 => x"7d708405",
958 => x"5f087170",
959 => x"8405530c",
960 => x"7d08710c",
961 => x"5f7b5261",
962 => x"518e983f",
963 => x"6151a4f7",
964 => x"3f79800c",
965 => x"933d0d04",
966 => x"7d526151",
967 => x"96943f80",
968 => x"08800c93",
969 => x"3d0d0484",
970 => x"160855fb",
971 => x"c9397753",
972 => x"7b528008",
973 => x"51a2a93f",
974 => x"7b526151",
975 => x"8de53fcc",
976 => x"398c1608",
977 => x"88170871",
978 => x"8c120c88",
979 => x"120c5d8c",
980 => x"17088818",
981 => x"08718c12",
982 => x"0c88120c",
983 => x"597759fb",
984 => x"ef397818",
985 => x"901c4055",
986 => x"7e7524fb",
987 => x"9c387a17",
988 => x"7080dad8",
989 => x"0b88050c",
990 => x"757c3181",
991 => x"0784120c",
992 => x"56841708",
993 => x"81067b07",
994 => x"84180c61",
995 => x"51a3f83f",
996 => x"881754fc",
997 => x"e1397418",
998 => x"19901c5e",
999 => x"5a7c7a24",
1000 => x"fb8f388c",
1001 => x"17088818",
1002 => x"08718c12",
1003 => x"0c88120c",
1004 => x"5e881761",
1005 => x"fc055759",
1006 => x"75a42681",
1007 => x"b6387b79",
1008 => x"59559376",
1009 => x"2780c938",
1010 => x"7b708405",
1011 => x"5d087c56",
1012 => x"790c7470",
1013 => x"84055608",
1014 => x"8c180c90",
1015 => x"17589b76",
1016 => x"27ae3874",
1017 => x"70840556",
1018 => x"08780c74",
1019 => x"70840556",
1020 => x"0894180c",
1021 => x"981758a3",
1022 => x"76279538",
1023 => x"74708405",
1024 => x"5608780c",
1025 => x"74708405",
1026 => x"56089c18",
1027 => x"0ca01758",
1028 => x"74708405",
1029 => x"56087541",
1030 => x"78708405",
1031 => x"5a0c7760",
1032 => x"70840542",
1033 => x"08717084",
1034 => x"05530c60",
1035 => x"08710c5e",
1036 => x"7a177080",
1037 => x"dad80b88",
1038 => x"050c7a7c",
1039 => x"31810784",
1040 => x"120c5884",
1041 => x"17088106",
1042 => x"7b078418",
1043 => x"0c6151a2",
1044 => x"b63f7854",
1045 => x"73800c93",
1046 => x"3d0d0479",
1047 => x"537b5275",
1048 => x"519ffd3f",
1049 => x"fae93984",
1050 => x"1508fc06",
1051 => x"19605859",
1052 => x"fadd3975",
1053 => x"537b5278",
1054 => x"519fe53f",
1055 => x"7a177080",
1056 => x"dad80b88",
1057 => x"050c7a7c",
1058 => x"31810784",
1059 => x"120c5884",
1060 => x"17088106",
1061 => x"7b078418",
1062 => x"0c6151a1",
1063 => x"ea3f7854",
1064 => x"ffb239fa",
1065 => x"3d0d7880",
1066 => x"d39c0854",
1067 => x"55b81308",
1068 => x"802e81af",
1069 => x"388c1522",
1070 => x"7083ffff",
1071 => x"0670832a",
1072 => x"81328106",
1073 => x"55555672",
1074 => x"802e80da",
1075 => x"3873842a",
1076 => x"81328106",
1077 => x"57ff5376",
1078 => x"80f23873",
1079 => x"822a8106",
1080 => x"5473802e",
1081 => x"b938b015",
1082 => x"08547380",
1083 => x"2e9c3880",
1084 => x"c0155373",
1085 => x"732e8f38",
1086 => x"735280d3",
1087 => x"9c08518a",
1088 => x"a23f8c15",
1089 => x"225676b0",
1090 => x"160c75db",
1091 => x"0657768c",
1092 => x"1623800b",
1093 => x"84160c90",
1094 => x"1508750c",
1095 => x"76567588",
1096 => x"0754738c",
1097 => x"16239015",
1098 => x"08802ebf",
1099 => x"388c1522",
1100 => x"70810655",
1101 => x"53739c38",
1102 => x"720a100a",
1103 => x"81065675",
1104 => x"85389415",
1105 => x"08547388",
1106 => x"160c8053",
1107 => x"72800c88",
1108 => x"3d0d0480",
1109 => x"0b88160c",
1110 => x"94150830",
1111 => x"98160c80",
1112 => x"53ea3972",
1113 => x"5182a63f",
1114 => x"fecb3974",
1115 => x"518fc03f",
1116 => x"8c152270",
1117 => x"81065553",
1118 => x"73802eff",
1119 => x"bb38d439",
1120 => x"f83d0d7a",
1121 => x"5776802e",
1122 => x"81973880",
1123 => x"d39c0854",
1124 => x"b8140880",
1125 => x"2e80eb38",
1126 => x"8c172270",
1127 => x"902b7090",
1128 => x"2c70832a",
1129 => x"81328106",
1130 => x"5b5b5755",
1131 => x"7780cb38",
1132 => x"90170856",
1133 => x"75802e80",
1134 => x"c1387608",
1135 => x"76317678",
1136 => x"0c798306",
1137 => x"55557385",
1138 => x"38941708",
1139 => x"58778818",
1140 => x"0c807525",
1141 => x"a5387453",
1142 => x"75529c17",
1143 => x"0851a417",
1144 => x"0854732d",
1145 => x"800b8008",
1146 => x"2580c938",
1147 => x"80081675",
1148 => x"80083156",
1149 => x"56748024",
1150 => x"dd38800b",
1151 => x"800c8a3d",
1152 => x"0d047351",
1153 => x"81873f8c",
1154 => x"17227090",
1155 => x"2b70902c",
1156 => x"70832a81",
1157 => x"3281065b",
1158 => x"5b575577",
1159 => x"dd38ff90",
1160 => x"39a38052",
1161 => x"80d39c08",
1162 => x"518cd43f",
1163 => x"8008800c",
1164 => x"8a3d0d04",
1165 => x"8c172280",
1166 => x"c0075877",
1167 => x"8c1823ff",
1168 => x"0b800c8a",
1169 => x"3d0d04fa",
1170 => x"3d0d7970",
1171 => x"80dc298c",
1172 => x"11547a53",
1173 => x"56578fda",
1174 => x"3f800880",
1175 => x"08555680",
1176 => x"08802ea2",
1177 => x"3880088c",
1178 => x"0554800b",
1179 => x"80080c76",
1180 => x"80088405",
1181 => x"0c738008",
1182 => x"88050c74",
1183 => x"53805273",
1184 => x"519cf93f",
1185 => x"75547380",
1186 => x"0c883d0d",
1187 => x"04fe3d0d",
1188 => x"74aacc0b",
1189 => x"bc120c53",
1190 => x"810bb814",
1191 => x"0c800b84",
1192 => x"dc140c83",
1193 => x"0b84e014",
1194 => x"0c84e813",
1195 => x"84e4140c",
1196 => x"84130851",
1197 => x"8070720c",
1198 => x"7084130c",
1199 => x"7088130c",
1200 => x"52840b8c",
1201 => x"1223718e",
1202 => x"12237190",
1203 => x"120c7194",
1204 => x"120c7198",
1205 => x"120c709c",
1206 => x"120c80c3",
1207 => x"bc0ba012",
1208 => x"0c80c488",
1209 => x"0ba4120c",
1210 => x"80c5840b",
1211 => x"a8120c80",
1212 => x"c5d50bac",
1213 => x"120c8813",
1214 => x"0872710c",
1215 => x"7284120c",
1216 => x"7288120c",
1217 => x"51890b8c",
1218 => x"1223810b",
1219 => x"8e122371",
1220 => x"90120c71",
1221 => x"94120c71",
1222 => x"98120c70",
1223 => x"9c120c80",
1224 => x"c3bc0ba0",
1225 => x"120c80c4",
1226 => x"880ba412",
1227 => x"0c80c584",
1228 => x"0ba8120c",
1229 => x"80c5d50b",
1230 => x"ac120c8c",
1231 => x"13087271",
1232 => x"0c728412",
1233 => x"0c728812",
1234 => x"0c518a0b",
1235 => x"8c122382",
1236 => x"0b8e1223",
1237 => x"7190120c",
1238 => x"7194120c",
1239 => x"7198120c",
1240 => x"709c120c",
1241 => x"80c3bc0b",
1242 => x"a0120c80",
1243 => x"c4880ba4",
1244 => x"120c80c5",
1245 => x"840ba812",
1246 => x"0c80c5d5",
1247 => x"0bac120c",
1248 => x"843d0d04",
1249 => x"f83d0d7a",
1250 => x"80d39c08",
1251 => x"b8110857",
1252 => x"57587481",
1253 => x"ec38aacc",
1254 => x"0bbc170c",
1255 => x"810bb817",
1256 => x"0c7484dc",
1257 => x"170c830b",
1258 => x"84e0170c",
1259 => x"84e81684",
1260 => x"e4170c84",
1261 => x"16087571",
1262 => x"0c758412",
1263 => x"0c758812",
1264 => x"0c59840b",
1265 => x"8c1a2374",
1266 => x"8e1a2374",
1267 => x"901a0c74",
1268 => x"941a0c74",
1269 => x"981a0c78",
1270 => x"9c1a0c80",
1271 => x"c3bc0ba0",
1272 => x"1a0c80c4",
1273 => x"880ba41a",
1274 => x"0c80c584",
1275 => x"0ba81a0c",
1276 => x"80c5d50b",
1277 => x"ac1a0c88",
1278 => x"16087571",
1279 => x"0c758412",
1280 => x"0c758812",
1281 => x"0c57890b",
1282 => x"8c182381",
1283 => x"0b8e1823",
1284 => x"7490180c",
1285 => x"7494180c",
1286 => x"7498180c",
1287 => x"769c180c",
1288 => x"80c3bc0b",
1289 => x"a0180c80",
1290 => x"c4880ba4",
1291 => x"180c80c5",
1292 => x"840ba818",
1293 => x"0c80c5d5",
1294 => x"0bac180c",
1295 => x"8c160875",
1296 => x"710c7584",
1297 => x"120c7588",
1298 => x"120c548a",
1299 => x"0b8c1523",
1300 => x"820b8e15",
1301 => x"23749015",
1302 => x"0c749415",
1303 => x"0c749815",
1304 => x"0c739c15",
1305 => x"0c80c3bc",
1306 => x"0ba0150c",
1307 => x"80c4880b",
1308 => x"a4150c80",
1309 => x"c5840ba8",
1310 => x"150c80c5",
1311 => x"d50bac15",
1312 => x"0c84dc16",
1313 => x"88110884",
1314 => x"1208ff05",
1315 => x"57575780",
1316 => x"75249f38",
1317 => x"8c162270",
1318 => x"902b7090",
1319 => x"2c515559",
1320 => x"73802e80",
1321 => x"ed3880dc",
1322 => x"16ff1656",
1323 => x"56748025",
1324 => x"e3387608",
1325 => x"5574802e",
1326 => x"8f387488",
1327 => x"11088412",
1328 => x"08ff0557",
1329 => x"5757c839",
1330 => x"82fc5277",
1331 => x"518ae33f",
1332 => x"80088008",
1333 => x"55568008",
1334 => x"802ea338",
1335 => x"80088c05",
1336 => x"7580080c",
1337 => x"54840b80",
1338 => x"0884050c",
1339 => x"73800888",
1340 => x"050c82f0",
1341 => x"53745273",
1342 => x"5198813f",
1343 => x"75547374",
1344 => x"780c5573",
1345 => x"ffb4388c",
1346 => x"780c800b",
1347 => x"800c8a3d",
1348 => x"0d04810b",
1349 => x"8c172373",
1350 => x"760c7388",
1351 => x"170c7384",
1352 => x"170c7390",
1353 => x"170c7394",
1354 => x"170c7398",
1355 => x"170cff0b",
1356 => x"8e172373",
1357 => x"b0170c73",
1358 => x"b4170c73",
1359 => x"80c4170c",
1360 => x"7380c817",
1361 => x"0c75800c",
1362 => x"8a3d0d04",
1363 => x"ff3d0da3",
1364 => x"80527351",
1365 => x"86a93f83",
1366 => x"3d0d04ff",
1367 => x"3d0da380",
1368 => x"5280d39c",
1369 => x"08518697",
1370 => x"3f833d0d",
1371 => x"04fb3d0d",
1372 => x"77705256",
1373 => x"98903f80",
1374 => x"dad80b88",
1375 => x"05088411",
1376 => x"08fc0670",
1377 => x"7b319fef",
1378 => x"05e08006",
1379 => x"e0800552",
1380 => x"5555a080",
1381 => x"75249438",
1382 => x"80527551",
1383 => x"97ea3f80",
1384 => x"dae00814",
1385 => x"53728008",
1386 => x"2e8f3875",
1387 => x"5197d83f",
1388 => x"80537280",
1389 => x"0c873d0d",
1390 => x"04743052",
1391 => x"755197c8",
1392 => x"3f8008ff",
1393 => x"2ea83880",
1394 => x"dad80b88",
1395 => x"05087476",
1396 => x"31810784",
1397 => x"120c5380",
1398 => x"da9c0875",
1399 => x"3180da9c",
1400 => x"0c755197",
1401 => x"a23f810b",
1402 => x"800c873d",
1403 => x"0d048052",
1404 => x"75519794",
1405 => x"3f80dad8",
1406 => x"0b880508",
1407 => x"80087131",
1408 => x"54548f73",
1409 => x"25ffa438",
1410 => x"800880da",
1411 => x"cc083180",
1412 => x"da9c0c72",
1413 => x"81078415",
1414 => x"0c755196",
1415 => x"ea3f8053",
1416 => x"ff9039f7",
1417 => x"3d0d7b7d",
1418 => x"545a7280",
1419 => x"2e828338",
1420 => x"795196d2",
1421 => x"3ff81384",
1422 => x"110870fe",
1423 => x"06701384",
1424 => x"1108fc06",
1425 => x"5c575854",
1426 => x"5780dae0",
1427 => x"08742e82",
1428 => x"de387784",
1429 => x"150c8073",
1430 => x"81065659",
1431 => x"74792e81",
1432 => x"d5387714",
1433 => x"84110881",
1434 => x"06565374",
1435 => x"a0387716",
1436 => x"567881e6",
1437 => x"38881408",
1438 => x"557480da",
1439 => x"e02e82f9",
1440 => x"388c1408",
1441 => x"708c170c",
1442 => x"7588120c",
1443 => x"58758107",
1444 => x"84180c75",
1445 => x"1776710c",
1446 => x"54788191",
1447 => x"3883ff76",
1448 => x"2781c838",
1449 => x"75892a76",
1450 => x"832a5454",
1451 => x"73802ebf",
1452 => x"3875862a",
1453 => x"b8055384",
1454 => x"7427b438",
1455 => x"80db1453",
1456 => x"947427ab",
1457 => x"38758c2a",
1458 => x"80ee0553",
1459 => x"80d47427",
1460 => x"9e38758f",
1461 => x"2a80f705",
1462 => x"5382d474",
1463 => x"27913875",
1464 => x"922a80fc",
1465 => x"05538ad4",
1466 => x"74278438",
1467 => x"80fe5372",
1468 => x"10101080",
1469 => x"dad80588",
1470 => x"11085555",
1471 => x"73752e82",
1472 => x"bf388414",
1473 => x"08fc0659",
1474 => x"7579278d",
1475 => x"38881408",
1476 => x"5473752e",
1477 => x"098106ea",
1478 => x"388c1408",
1479 => x"708c190c",
1480 => x"7488190c",
1481 => x"7788120c",
1482 => x"55768c15",
1483 => x"0c795194",
1484 => x"d63f8b3d",
1485 => x"0d047608",
1486 => x"77713158",
1487 => x"76058818",
1488 => x"08565674",
1489 => x"80dae02e",
1490 => x"80e0388c",
1491 => x"1708708c",
1492 => x"170c7588",
1493 => x"120c53fe",
1494 => x"89398814",
1495 => x"088c1508",
1496 => x"708c130c",
1497 => x"5988190c",
1498 => x"fea33975",
1499 => x"832a7054",
1500 => x"54807424",
1501 => x"81983872",
1502 => x"822c8171",
1503 => x"2b80dadc",
1504 => x"080780da",
1505 => x"d80b8405",
1506 => x"0c741010",
1507 => x"1080dad8",
1508 => x"05881108",
1509 => x"718c1b0c",
1510 => x"70881b0c",
1511 => x"7988130c",
1512 => x"565a5576",
1513 => x"8c150cff",
1514 => x"84398159",
1515 => x"fdb43977",
1516 => x"16738106",
1517 => x"54557298",
1518 => x"38760877",
1519 => x"71315875",
1520 => x"058c1808",
1521 => x"88190871",
1522 => x"8c120c88",
1523 => x"120c5555",
1524 => x"74810784",
1525 => x"180c7680",
1526 => x"dad80b88",
1527 => x"050c80da",
1528 => x"d4087526",
1529 => x"fec73880",
1530 => x"dad00852",
1531 => x"7951fafd",
1532 => x"3f795193",
1533 => x"923ffeba",
1534 => x"3981778c",
1535 => x"170c7788",
1536 => x"170c758c",
1537 => x"190c7588",
1538 => x"190c59fd",
1539 => x"80398314",
1540 => x"70822c81",
1541 => x"712b80da",
1542 => x"dc080780",
1543 => x"dad80b84",
1544 => x"050c7510",
1545 => x"101080da",
1546 => x"d8058811",
1547 => x"08718c1c",
1548 => x"0c70881c",
1549 => x"0c7a8813",
1550 => x"0c575b56",
1551 => x"53fee439",
1552 => x"807324a3",
1553 => x"3872822c",
1554 => x"81712b80",
1555 => x"dadc0807",
1556 => x"80dad80b",
1557 => x"84050c58",
1558 => x"748c180c",
1559 => x"7388180c",
1560 => x"7688160c",
1561 => x"fdc33983",
1562 => x"1370822c",
1563 => x"81712b80",
1564 => x"dadc0807",
1565 => x"80dad80b",
1566 => x"84050c59",
1567 => x"53da39f9",
1568 => x"3d0d797b",
1569 => x"5853800b",
1570 => x"80d39c08",
1571 => x"53567272",
1572 => x"2ebc3884",
1573 => x"dc135574",
1574 => x"762eb338",
1575 => x"88150884",
1576 => x"1608ff05",
1577 => x"54548073",
1578 => x"2499388c",
1579 => x"14227090",
1580 => x"2b535871",
1581 => x"80d43880",
1582 => x"dc14ff14",
1583 => x"54547280",
1584 => x"25e93874",
1585 => x"085574d4",
1586 => x"3880d39c",
1587 => x"085284dc",
1588 => x"12557480",
1589 => x"2ead3888",
1590 => x"15088416",
1591 => x"08ff0554",
1592 => x"54807324",
1593 => x"98388c14",
1594 => x"2270902b",
1595 => x"535871ad",
1596 => x"3880dc14",
1597 => x"ff145454",
1598 => x"728025ea",
1599 => x"38740855",
1600 => x"74d53875",
1601 => x"800c893d",
1602 => x"0d047351",
1603 => x"762d7580",
1604 => x"080780dc",
1605 => x"15ff1555",
1606 => x"5556ffa2",
1607 => x"39735176",
1608 => x"2d758008",
1609 => x"0780dc15",
1610 => x"ff155555",
1611 => x"56ca39ea",
1612 => x"3d0d688c",
1613 => x"1122700a",
1614 => x"100a8106",
1615 => x"57585674",
1616 => x"80e4388e",
1617 => x"16227090",
1618 => x"2b70902c",
1619 => x"51555880",
1620 => x"7424b138",
1621 => x"983dc405",
1622 => x"53735280",
1623 => x"d39c0851",
1624 => x"93fb3f80",
1625 => x"0b800824",
1626 => x"97387983",
1627 => x"e0800654",
1628 => x"7380c080",
1629 => x"2e818f38",
1630 => x"73828080",
1631 => x"2e819138",
1632 => x"8c162257",
1633 => x"76908007",
1634 => x"54738c17",
1635 => x"23888052",
1636 => x"80d39c08",
1637 => x"51819b3f",
1638 => x"80089d38",
1639 => x"8c162282",
1640 => x"0755748c",
1641 => x"172380c3",
1642 => x"1670770c",
1643 => x"90170c81",
1644 => x"0b94170c",
1645 => x"983d0d04",
1646 => x"80d39c08",
1647 => x"aacc0bbc",
1648 => x"120c588c",
1649 => x"16228180",
1650 => x"0754738c",
1651 => x"17238008",
1652 => x"760c8008",
1653 => x"90170c88",
1654 => x"800b9417",
1655 => x"0c74802e",
1656 => x"d3388e16",
1657 => x"2270902b",
1658 => x"70902c53",
1659 => x"56549cd0",
1660 => x"3f800880",
1661 => x"2effbd38",
1662 => x"8c162281",
1663 => x"0757768c",
1664 => x"1723983d",
1665 => x"0d04810b",
1666 => x"8c172258",
1667 => x"55fef539",
1668 => x"a8160880",
1669 => x"c5842e09",
1670 => x"8106fee4",
1671 => x"388c1622",
1672 => x"88800754",
1673 => x"738c1723",
1674 => x"88800b80",
1675 => x"cc170cfe",
1676 => x"dc39f43d",
1677 => x"0d7e608b",
1678 => x"1170f806",
1679 => x"5b55555d",
1680 => x"72962683",
1681 => x"38905880",
1682 => x"78247479",
1683 => x"26075580",
1684 => x"5474742e",
1685 => x"09810680",
1686 => x"ca387c51",
1687 => x"8ea83f77",
1688 => x"83f72680",
1689 => x"c5387783",
1690 => x"2a701010",
1691 => x"1080dad8",
1692 => x"058c1108",
1693 => x"58585475",
1694 => x"772e81f0",
1695 => x"38841608",
1696 => x"fc068c17",
1697 => x"08881808",
1698 => x"718c120c",
1699 => x"88120c5b",
1700 => x"76058411",
1701 => x"08810784",
1702 => x"120c537c",
1703 => x"518de83f",
1704 => x"88165473",
1705 => x"800c8e3d",
1706 => x"0d047789",
1707 => x"2a78832a",
1708 => x"58547380",
1709 => x"2ebf3877",
1710 => x"862ab805",
1711 => x"57847427",
1712 => x"b43880db",
1713 => x"14579474",
1714 => x"27ab3877",
1715 => x"8c2a80ee",
1716 => x"055780d4",
1717 => x"74279e38",
1718 => x"778f2a80",
1719 => x"f7055782",
1720 => x"d4742791",
1721 => x"3877922a",
1722 => x"80fc0557",
1723 => x"8ad47427",
1724 => x"843880fe",
1725 => x"57761010",
1726 => x"1080dad8",
1727 => x"058c1108",
1728 => x"56537473",
1729 => x"2ea33884",
1730 => x"1508fc06",
1731 => x"70793155",
1732 => x"56738f24",
1733 => x"88e43873",
1734 => x"802588e6",
1735 => x"388c1508",
1736 => x"5574732e",
1737 => x"098106df",
1738 => x"38811759",
1739 => x"80dae808",
1740 => x"567580da",
1741 => x"e02e82cc",
1742 => x"38841608",
1743 => x"fc067079",
1744 => x"31555573",
1745 => x"8f24bb38",
1746 => x"80dae00b",
1747 => x"80daec0c",
1748 => x"80dae00b",
1749 => x"80dae80c",
1750 => x"80742480",
1751 => x"db387416",
1752 => x"84110881",
1753 => x"0784120c",
1754 => x"53feb039",
1755 => x"88168c11",
1756 => x"08575975",
1757 => x"792e0981",
1758 => x"06fe8238",
1759 => x"821459ff",
1760 => x"ab397716",
1761 => x"78810784",
1762 => x"180c7080",
1763 => x"daec0c70",
1764 => x"80dae80c",
1765 => x"80dae00b",
1766 => x"8c120c8c",
1767 => x"11088812",
1768 => x"0c748107",
1769 => x"84120c74",
1770 => x"0574710c",
1771 => x"5b7c518b",
1772 => x"d63f8816",
1773 => x"54fdec39",
1774 => x"83ff7527",
1775 => x"83913874",
1776 => x"892a7583",
1777 => x"2a545473",
1778 => x"802ebf38",
1779 => x"74862ab8",
1780 => x"05538474",
1781 => x"27b43880",
1782 => x"db145394",
1783 => x"7427ab38",
1784 => x"748c2a80",
1785 => x"ee055380",
1786 => x"d474279e",
1787 => x"38748f2a",
1788 => x"80f70553",
1789 => x"82d47427",
1790 => x"91387492",
1791 => x"2a80fc05",
1792 => x"538ad474",
1793 => x"27843880",
1794 => x"fe537210",
1795 => x"101080da",
1796 => x"d8058811",
1797 => x"08555773",
1798 => x"772e868b",
1799 => x"38841408",
1800 => x"fc065b74",
1801 => x"7b278d38",
1802 => x"88140854",
1803 => x"73772e09",
1804 => x"8106ea38",
1805 => x"8c140880",
1806 => x"dad80b84",
1807 => x"0508718c",
1808 => x"190c7588",
1809 => x"190c7788",
1810 => x"130c5c57",
1811 => x"758c150c",
1812 => x"78538079",
1813 => x"24839838",
1814 => x"72822c81",
1815 => x"712b5656",
1816 => x"747b2680",
1817 => x"ca387a75",
1818 => x"06577682",
1819 => x"a33878fc",
1820 => x"06840559",
1821 => x"7410707c",
1822 => x"06555573",
1823 => x"82923884",
1824 => x"1959f139",
1825 => x"80dad80b",
1826 => x"84050879",
1827 => x"545b7880",
1828 => x"25c63882",
1829 => x"da397409",
1830 => x"7b067080",
1831 => x"dad80b84",
1832 => x"050c5b74",
1833 => x"1055747b",
1834 => x"26853874",
1835 => x"85bc3880",
1836 => x"dad80b88",
1837 => x"05087084",
1838 => x"1208fc06",
1839 => x"707b317b",
1840 => x"72268f72",
1841 => x"25075d57",
1842 => x"5c5c5578",
1843 => x"802e80d9",
1844 => x"38791580",
1845 => x"dad00819",
1846 => x"90115954",
1847 => x"5680dacc",
1848 => x"08ff2e88",
1849 => x"38a08f13",
1850 => x"e0800657",
1851 => x"76527c51",
1852 => x"89963f80",
1853 => x"08548008",
1854 => x"ff2e9038",
1855 => x"80087627",
1856 => x"82a73874",
1857 => x"80dad82e",
1858 => x"829f3880",
1859 => x"dad80b88",
1860 => x"05085584",
1861 => x"1508fc06",
1862 => x"70793179",
1863 => x"72268f72",
1864 => x"25075d55",
1865 => x"5a7a83f2",
1866 => x"38778107",
1867 => x"84160c77",
1868 => x"157080da",
1869 => x"d80b8805",
1870 => x"0c748107",
1871 => x"84120c56",
1872 => x"7c5188c3",
1873 => x"3f881554",
1874 => x"73800c8e",
1875 => x"3d0d0474",
1876 => x"832a7054",
1877 => x"54807424",
1878 => x"819b3872",
1879 => x"822c8171",
1880 => x"2b80dadc",
1881 => x"08077080",
1882 => x"dad80b84",
1883 => x"050c7510",
1884 => x"101080da",
1885 => x"d8058811",
1886 => x"08718c1b",
1887 => x"0c70881b",
1888 => x"0c798813",
1889 => x"0c57555c",
1890 => x"55758c15",
1891 => x"0cfdc139",
1892 => x"78791010",
1893 => x"1080dad8",
1894 => x"0570565b",
1895 => x"5c8c1408",
1896 => x"5675742e",
1897 => x"a3388416",
1898 => x"08fc0670",
1899 => x"79315853",
1900 => x"768f2483",
1901 => x"f1387680",
1902 => x"2584af38",
1903 => x"8c160856",
1904 => x"75742e09",
1905 => x"8106df38",
1906 => x"8814811a",
1907 => x"70830655",
1908 => x"5a5472c9",
1909 => x"387b8306",
1910 => x"5675802e",
1911 => x"fdb838ff",
1912 => x"1cf81b5b",
1913 => x"5c881a08",
1914 => x"7a2eea38",
1915 => x"fdb53983",
1916 => x"1953fce4",
1917 => x"39831470",
1918 => x"822c8171",
1919 => x"2b80dadc",
1920 => x"08077080",
1921 => x"dad80b84",
1922 => x"050c7610",
1923 => x"101080da",
1924 => x"d8058811",
1925 => x"08718c1c",
1926 => x"0c70881c",
1927 => x"0c7a8813",
1928 => x"0c58535d",
1929 => x"5653fee1",
1930 => x"3980da9c",
1931 => x"08175980",
1932 => x"08762e81",
1933 => x"8b3880da",
1934 => x"cc08ff2e",
1935 => x"848e3873",
1936 => x"76311980",
1937 => x"da9c0c73",
1938 => x"87067056",
1939 => x"5372802e",
1940 => x"88388873",
1941 => x"31701555",
1942 => x"5576149f",
1943 => x"ff06a080",
1944 => x"71311670",
1945 => x"547e5351",
1946 => x"53869d3f",
1947 => x"80085680",
1948 => x"08ff2e81",
1949 => x"9e3880da",
1950 => x"9c081370",
1951 => x"80da9c0c",
1952 => x"747580da",
1953 => x"d80b8805",
1954 => x"0c777631",
1955 => x"15810755",
1956 => x"56597a80",
1957 => x"dad82e83",
1958 => x"c038798f",
1959 => x"2682ef38",
1960 => x"810b8415",
1961 => x"0c841508",
1962 => x"fc067079",
1963 => x"31797226",
1964 => x"8f722507",
1965 => x"5d555a7a",
1966 => x"802efced",
1967 => x"3880db39",
1968 => x"80089fff",
1969 => x"065574fe",
1970 => x"ed387880",
1971 => x"da9c0c80",
1972 => x"dad80b88",
1973 => x"05087a18",
1974 => x"81078412",
1975 => x"0c5580da",
1976 => x"c8087927",
1977 => x"86387880",
1978 => x"dac80c80",
1979 => x"dac40879",
1980 => x"27fca038",
1981 => x"7880dac4",
1982 => x"0c841508",
1983 => x"fc067079",
1984 => x"31797226",
1985 => x"8f722507",
1986 => x"5d555a7a",
1987 => x"802efc99",
1988 => x"38883980",
1989 => x"745753fe",
1990 => x"dd397c51",
1991 => x"84e93f80",
1992 => x"0b800c8e",
1993 => x"3d0d0480",
1994 => x"7324a538",
1995 => x"72822c81",
1996 => x"712b80da",
1997 => x"dc080770",
1998 => x"80dad80b",
1999 => x"84050c5c",
2000 => x"5a768c17",
2001 => x"0c738817",
2002 => x"0c758818",
2003 => x"0cf9fd39",
2004 => x"83137082",
2005 => x"2c81712b",
2006 => x"80dadc08",
2007 => x"077080da",
2008 => x"d80b8405",
2009 => x"0c5d5b53",
2010 => x"d8397a75",
2011 => x"065c7bfc",
2012 => x"9f388419",
2013 => x"75105659",
2014 => x"f139ff17",
2015 => x"810559f7",
2016 => x"ab398c15",
2017 => x"08881608",
2018 => x"718c120c",
2019 => x"88120c59",
2020 => x"75158411",
2021 => x"08810784",
2022 => x"120c587c",
2023 => x"5183e83f",
2024 => x"881554fb",
2025 => x"a3397716",
2026 => x"78810784",
2027 => x"180c8c17",
2028 => x"08881808",
2029 => x"718c120c",
2030 => x"88120c5c",
2031 => x"7080daec",
2032 => x"0c7080da",
2033 => x"e80c80da",
2034 => x"e00b8c12",
2035 => x"0c8c1108",
2036 => x"88120c77",
2037 => x"81078412",
2038 => x"0c770577",
2039 => x"710c557c",
2040 => x"5183a43f",
2041 => x"881654f5",
2042 => x"ba397216",
2043 => x"84110881",
2044 => x"0784120c",
2045 => x"588c1608",
2046 => x"88170871",
2047 => x"8c120c88",
2048 => x"120c577c",
2049 => x"5183803f",
2050 => x"881654f5",
2051 => x"96397284",
2052 => x"150cf41a",
2053 => x"f8067084",
2054 => x"1d088106",
2055 => x"07841d0c",
2056 => x"701c5556",
2057 => x"850b8415",
2058 => x"0c850b88",
2059 => x"150c8f76",
2060 => x"27fdab38",
2061 => x"881b527c",
2062 => x"51ebe83f",
2063 => x"80dad80b",
2064 => x"88050880",
2065 => x"da9c085a",
2066 => x"55fd9339",
2067 => x"7880da9c",
2068 => x"0c7380da",
2069 => x"cc0cfbef",
2070 => x"39728415",
2071 => x"0cfcff39",
2072 => x"fb3d0d77",
2073 => x"707a7c58",
2074 => x"5553568f",
2075 => x"752780e6",
2076 => x"38727607",
2077 => x"83065170",
2078 => x"80dc3875",
2079 => x"73525470",
2080 => x"70840552",
2081 => x"08747084",
2082 => x"05560c73",
2083 => x"71708405",
2084 => x"53087170",
2085 => x"8405530c",
2086 => x"71708405",
2087 => x"53087170",
2088 => x"8405530c",
2089 => x"71708405",
2090 => x"53087170",
2091 => x"8405530c",
2092 => x"f0165654",
2093 => x"748f26c7",
2094 => x"38837527",
2095 => x"95387070",
2096 => x"84055208",
2097 => x"74708405",
2098 => x"560cfc15",
2099 => x"55748326",
2100 => x"ed387371",
2101 => x"5452ff15",
2102 => x"5170ff2e",
2103 => x"98387270",
2104 => x"81055433",
2105 => x"72708105",
2106 => x"5434ff11",
2107 => x"5170ff2e",
2108 => x"098106ea",
2109 => x"3875800c",
2110 => x"873d0d04",
2111 => x"fb3d0d77",
2112 => x"7a71028c",
2113 => x"05a30533",
2114 => x"58545456",
2115 => x"83732780",
2116 => x"d4387583",
2117 => x"06517080",
2118 => x"cc387488",
2119 => x"2b750770",
2120 => x"71902b07",
2121 => x"55518f73",
2122 => x"27a73873",
2123 => x"72708405",
2124 => x"540c7174",
2125 => x"71708405",
2126 => x"530c7471",
2127 => x"70840553",
2128 => x"0c747170",
2129 => x"8405530c",
2130 => x"f0145452",
2131 => x"728f26db",
2132 => x"38837327",
2133 => x"90387372",
2134 => x"70840554",
2135 => x"0cfc1353",
2136 => x"728326f2",
2137 => x"38ff1351",
2138 => x"70ff2e93",
2139 => x"38747270",
2140 => x"81055434",
2141 => x"ff115170",
2142 => x"ff2e0981",
2143 => x"06ef3875",
2144 => x"800c873d",
2145 => x"0d040404",
2146 => x"fd3d0d80",
2147 => x"0b80e3a0",
2148 => x"0c765184",
2149 => x"ee3f8008",
2150 => x"538008ff",
2151 => x"2e883872",
2152 => x"800c853d",
2153 => x"0d0480e3",
2154 => x"a0085473",
2155 => x"802ef038",
2156 => x"7574710c",
2157 => x"5272800c",
2158 => x"853d0d04",
2159 => x"f93d0d79",
2160 => x"7c557b54",
2161 => x"8e112270",
2162 => x"902b7090",
2163 => x"2c555780",
2164 => x"d39c0853",
2165 => x"585683f3",
2166 => x"3f800857",
2167 => x"800b8008",
2168 => x"24933880",
2169 => x"d0160880",
2170 => x"080580d0",
2171 => x"170c7680",
2172 => x"0c893d0d",
2173 => x"048c1622",
2174 => x"83dfff06",
2175 => x"55748c17",
2176 => x"2376800c",
2177 => x"893d0d04",
2178 => x"fa3d0d78",
2179 => x"8c112270",
2180 => x"882a7081",
2181 => x"06515758",
2182 => x"5674a938",
2183 => x"8c162283",
2184 => x"dfff0655",
2185 => x"748c1723",
2186 => x"7a547953",
2187 => x"8e162270",
2188 => x"902b7090",
2189 => x"2c545680",
2190 => x"d39c0852",
2191 => x"5681b23f",
2192 => x"883d0d04",
2193 => x"82548053",
2194 => x"8e162270",
2195 => x"902b7090",
2196 => x"2c545680",
2197 => x"d39c0852",
2198 => x"5782b83f",
2199 => x"8c162283",
2200 => x"dfff0655",
2201 => x"748c1723",
2202 => x"7a547953",
2203 => x"8e162270",
2204 => x"902b7090",
2205 => x"2c545680",
2206 => x"d39c0852",
2207 => x"5680f23f",
2208 => x"883d0d04",
2209 => x"f93d0d79",
2210 => x"7c557b54",
2211 => x"8e112270",
2212 => x"902b7090",
2213 => x"2c555780",
2214 => x"d39c0853",
2215 => x"585681f3",
2216 => x"3f800857",
2217 => x"8008ff2e",
2218 => x"99388c16",
2219 => x"22a08007",
2220 => x"55748c17",
2221 => x"23800880",
2222 => x"d0170c76",
2223 => x"800c893d",
2224 => x"0d048c16",
2225 => x"2283dfff",
2226 => x"0655748c",
2227 => x"17237680",
2228 => x"0c893d0d",
2229 => x"04fe3d0d",
2230 => x"748e1122",
2231 => x"70902b70",
2232 => x"902c5551",
2233 => x"515380d3",
2234 => x"9c0851bd",
2235 => x"3f843d0d",
2236 => x"04fb3d0d",
2237 => x"800b80e3",
2238 => x"a00c7a53",
2239 => x"79527851",
2240 => x"82fc3f80",
2241 => x"08558008",
2242 => x"ff2e8838",
2243 => x"74800c87",
2244 => x"3d0d0480",
2245 => x"e3a00856",
2246 => x"75802ef0",
2247 => x"38777671",
2248 => x"0c547480",
2249 => x"0c873d0d",
2250 => x"04fd3d0d",
2251 => x"800b80e3",
2252 => x"a00c7651",
2253 => x"85853f80",
2254 => x"08538008",
2255 => x"ff2e8838",
2256 => x"72800c85",
2257 => x"3d0d0480",
2258 => x"e3a00854",
2259 => x"73802ef0",
2260 => x"38757471",
2261 => x"0c527280",
2262 => x"0c853d0d",
2263 => x"04fc3d0d",
2264 => x"800b80e3",
2265 => x"a00c7852",
2266 => x"775188b8",
2267 => x"3f800854",
2268 => x"8008ff2e",
2269 => x"88387380",
2270 => x"0c863d0d",
2271 => x"0480e3a0",
2272 => x"08557480",
2273 => x"2ef03876",
2274 => x"75710c53",
2275 => x"73800c86",
2276 => x"3d0d04fb",
2277 => x"3d0d800b",
2278 => x"80e3a00c",
2279 => x"7a537952",
2280 => x"78518593",
2281 => x"3f800855",
2282 => x"8008ff2e",
2283 => x"88387480",
2284 => x"0c873d0d",
2285 => x"0480e3a0",
2286 => x"08567580",
2287 => x"2ef03877",
2288 => x"76710c54",
2289 => x"74800c87",
2290 => x"3d0d04fb",
2291 => x"3d0d800b",
2292 => x"80e3a00c",
2293 => x"7a537952",
2294 => x"7851829a",
2295 => x"3f800855",
2296 => x"8008ff2e",
2297 => x"88387480",
2298 => x"0c873d0d",
2299 => x"0480e3a0",
2300 => x"08567580",
2301 => x"2ef03877",
2302 => x"76710c54",
2303 => x"74800c87",
2304 => x"3d0d04fe",
2305 => x"3d0d80e3",
2306 => x"a4085170",
2307 => x"8a3880e3",
2308 => x"ac7080e3",
2309 => x"a40c5174",
2310 => x"1152ff53",
2311 => x"7187fb80",
2312 => x"80268838",
2313 => x"7180e3a4",
2314 => x"0c705372",
2315 => x"800c843d",
2316 => x"0d04fd3d",
2317 => x"0d800b80",
2318 => x"d3900854",
2319 => x"5472812e",
2320 => x"9c387380",
2321 => x"e3a80cc0",
2322 => x"d83fffbf",
2323 => x"b33f80e2",
2324 => x"e0528151",
2325 => x"c3b43f80",
2326 => x"0851889b",
2327 => x"3f7280e3",
2328 => x"a80cc0bd",
2329 => x"3fffbf98",
2330 => x"3f80e2e0",
2331 => x"528151c3",
2332 => x"993f8008",
2333 => x"5188803f",
2334 => x"00ff3900",
2335 => x"ff39f53d",
2336 => x"0d7e6080",
2337 => x"e3a80870",
2338 => x"5b585b5b",
2339 => x"7580c538",
2340 => x"777a25a2",
2341 => x"38771b70",
2342 => x"337081ff",
2343 => x"06585859",
2344 => x"758a2e99",
2345 => x"387681ff",
2346 => x"0651ffbf",
2347 => x"d33f8118",
2348 => x"58797824",
2349 => x"e0387980",
2350 => x"0c8d3d0d",
2351 => x"048d51ff",
2352 => x"bfbe3f78",
2353 => x"337081ff",
2354 => x"065257ff",
2355 => x"bfb23f81",
2356 => x"1858de39",
2357 => x"79557a54",
2358 => x"7d538552",
2359 => x"8d3dfc05",
2360 => x"51ffbede",
2361 => x"3f800856",
2362 => x"87863f7b",
2363 => x"80080c75",
2364 => x"800c8d3d",
2365 => x"0d04f63d",
2366 => x"0d7d7f80",
2367 => x"e3a80870",
2368 => x"5a585a5a",
2369 => x"7580c438",
2370 => x"767925b2",
2371 => x"38761a58",
2372 => x"ffbecd3f",
2373 => x"80087834",
2374 => x"800b8008",
2375 => x"81ff0657",
2376 => x"58758a2e",
2377 => x"a238758d",
2378 => x"32703070",
2379 => x"80257a07",
2380 => x"51515675",
2381 => x"b8388117",
2382 => x"57787724",
2383 => x"d0387656",
2384 => x"75800c8c",
2385 => x"3d0d0481",
2386 => x"58dc3978",
2387 => x"5579547c",
2388 => x"5384528c",
2389 => x"3dfc0551",
2390 => x"ffbde73f",
2391 => x"80085686",
2392 => x"8f3f7a80",
2393 => x"080c7580",
2394 => x"0c8c3d0d",
2395 => x"04811756",
2396 => x"cf39f93d",
2397 => x"0d795780",
2398 => x"e3a80880",
2399 => x"2ead3876",
2400 => x"51c4e33f",
2401 => x"7b567a55",
2402 => x"80088105",
2403 => x"54765382",
2404 => x"52893dfc",
2405 => x"0551ffbd",
2406 => x"a93f8008",
2407 => x"5785d13f",
2408 => x"7780080c",
2409 => x"76800c89",
2410 => x"3d0d0485",
2411 => x"c33f850b",
2412 => x"80080cff",
2413 => x"0b800c89",
2414 => x"3d0d04fb",
2415 => x"3d0d80e3",
2416 => x"a8087056",
2417 => x"54738838",
2418 => x"74800c87",
2419 => x"3d0d0477",
2420 => x"53835287",
2421 => x"3dfc0551",
2422 => x"ffbce73f",
2423 => x"80085485",
2424 => x"8f3f7580",
2425 => x"080c7380",
2426 => x"0c873d0d",
2427 => x"04ff0b80",
2428 => x"0c04fb3d",
2429 => x"0d775580",
2430 => x"e3a80880",
2431 => x"2ea93874",
2432 => x"51c3e33f",
2433 => x"80088105",
2434 => x"54745387",
2435 => x"52873dfc",
2436 => x"0551ffbc",
2437 => x"ad3f8008",
2438 => x"5584d53f",
2439 => x"7580080c",
2440 => x"74800c87",
2441 => x"3d0d0484",
2442 => x"c73f850b",
2443 => x"80080cff",
2444 => x"0b800c87",
2445 => x"3d0d04fa",
2446 => x"3d0d80e3",
2447 => x"a808802e",
2448 => x"a3387a55",
2449 => x"79547853",
2450 => x"8652883d",
2451 => x"fc0551ff",
2452 => x"bbf03f80",
2453 => x"08568498",
2454 => x"3f768008",
2455 => x"0c75800c",
2456 => x"883d0d04",
2457 => x"848a3f9d",
2458 => x"0b80080c",
2459 => x"ff0b800c",
2460 => x"883d0d04",
2461 => x"f73d0d7b",
2462 => x"7d5b59bc",
2463 => x"53805279",
2464 => x"51f4f93f",
2465 => x"80705657",
2466 => x"98567419",
2467 => x"70337078",
2468 => x"2b790781",
2469 => x"18f81a5a",
2470 => x"58595558",
2471 => x"847524ea",
2472 => x"38767a23",
2473 => x"84195880",
2474 => x"70565798",
2475 => x"56741870",
2476 => x"3370782b",
2477 => x"79078118",
2478 => x"f81a5a58",
2479 => x"59515484",
2480 => x"7524ea38",
2481 => x"76821b23",
2482 => x"88195880",
2483 => x"70565798",
2484 => x"56741870",
2485 => x"3370782b",
2486 => x"79078118",
2487 => x"f81a5a58",
2488 => x"59515484",
2489 => x"7524ea38",
2490 => x"76841b0c",
2491 => x"8c195880",
2492 => x"70565798",
2493 => x"56741870",
2494 => x"3370782b",
2495 => x"79078118",
2496 => x"f81a5a58",
2497 => x"59515484",
2498 => x"7524ea38",
2499 => x"76881b23",
2500 => x"90195880",
2501 => x"70565798",
2502 => x"56741870",
2503 => x"3370782b",
2504 => x"79078118",
2505 => x"f81a5a58",
2506 => x"59515484",
2507 => x"7524ea38",
2508 => x"768a1b23",
2509 => x"94195880",
2510 => x"70565798",
2511 => x"56741870",
2512 => x"3370782b",
2513 => x"79078118",
2514 => x"f81a5a58",
2515 => x"59515484",
2516 => x"7524ea38",
2517 => x"768c1b23",
2518 => x"98195880",
2519 => x"70565798",
2520 => x"56741870",
2521 => x"3370782b",
2522 => x"79078118",
2523 => x"f81a5a58",
2524 => x"59515484",
2525 => x"7524ea38",
2526 => x"768e1b23",
2527 => x"9c195880",
2528 => x"705657b8",
2529 => x"56741870",
2530 => x"3370782b",
2531 => x"79078118",
2532 => x"f81a5a58",
2533 => x"595a5488",
2534 => x"7524ea38",
2535 => x"76901b0c",
2536 => x"8b3d0d04",
2537 => x"e93d0d6a",
2538 => x"80e3a808",
2539 => x"57577593",
2540 => x"3880c080",
2541 => x"0b84180c",
2542 => x"75ac180c",
2543 => x"75800c99",
2544 => x"3d0d0489",
2545 => x"3d70556a",
2546 => x"54558a52",
2547 => x"993dffbc",
2548 => x"0551ffb8",
2549 => x"ed3f8008",
2550 => x"77537552",
2551 => x"56fd953f",
2552 => x"818e3f77",
2553 => x"80080c75",
2554 => x"800c993d",
2555 => x"0d04e93d",
2556 => x"0d695780",
2557 => x"e3a80880",
2558 => x"2eb73876",
2559 => x"51ffbfe6",
2560 => x"3f893d70",
2561 => x"56800881",
2562 => x"05557754",
2563 => x"568f5299",
2564 => x"3dffbc05",
2565 => x"51ffb8aa",
2566 => x"3f80086b",
2567 => x"53765257",
2568 => x"fcd23f80",
2569 => x"cb3f7780",
2570 => x"080c7680",
2571 => x"0c993d0d",
2572 => x"04be3f85",
2573 => x"0b80080c",
2574 => x"ff0b800c",
2575 => x"993d0d04",
2576 => x"fc3d0d81",
2577 => x"5480e3a8",
2578 => x"08883873",
2579 => x"800c863d",
2580 => x"0d047653",
2581 => x"97b95286",
2582 => x"3dfc0551",
2583 => x"ffb7e33f",
2584 => x"8008548c",
2585 => x"3f748008",
2586 => x"0c73800c",
2587 => x"863d0d04",
2588 => x"80d39c08",
2589 => x"800c04f7",
2590 => x"3d0d7b80",
2591 => x"d39c0882",
2592 => x"c811085a",
2593 => x"545a7780",
2594 => x"2e80da38",
2595 => x"81881884",
2596 => x"1908ff05",
2597 => x"81712b59",
2598 => x"55598074",
2599 => x"2480ea38",
2600 => x"807424b5",
2601 => x"3873822b",
2602 => x"78118805",
2603 => x"56568180",
2604 => x"19087706",
2605 => x"5372802e",
2606 => x"b6387816",
2607 => x"70085353",
2608 => x"79517408",
2609 => x"53722dff",
2610 => x"14fc17fc",
2611 => x"1779812c",
2612 => x"5a575754",
2613 => x"738025d6",
2614 => x"38770858",
2615 => x"77ffad38",
2616 => x"80d39c08",
2617 => x"53bc1308",
2618 => x"a5387951",
2619 => x"f78a3f74",
2620 => x"0853722d",
2621 => x"ff14fc17",
2622 => x"fc177981",
2623 => x"2c5a5757",
2624 => x"54738025",
2625 => x"ffa838d1",
2626 => x"398057ff",
2627 => x"93397251",
2628 => x"bc130854",
2629 => x"732d7951",
2630 => x"f6de3fff",
2631 => x"3d0d80e2",
2632 => x"e80bfc05",
2633 => x"70085252",
2634 => x"70ff2e91",
2635 => x"38702dfc",
2636 => x"12700852",
2637 => x"5270ff2e",
2638 => x"098106f1",
2639 => x"38833d0d",
2640 => x"0404ffb8",
2641 => x"e03f0400",
2642 => x"48656c6c",
2643 => x"6f20776f",
2644 => x"726c6420",
2645 => x"310a0000",
2646 => x"48656c6c",
2647 => x"6f20776f",
2648 => x"726c6420",
2649 => x"320a0000",
2650 => x"0a000000",
2651 => x"43000000",
2652 => x"64756d6d",
2653 => x"792e6578",
2654 => x"65000000",
2655 => x"00ffffff",
2656 => x"ff00ffff",
2657 => x"ffff00ff",
2658 => x"ffffff00",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00003170",
2663 => x"000029a0",
2664 => x"00000000",
2665 => x"00002c08",
2666 => x"00002c64",
2667 => x"00002cc0",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"0000296c",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000001",
2707 => x"330eabcd",
2708 => x"1234e66d",
2709 => x"deec0005",
2710 => x"000b0000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"00000000",
2792 => x"00000000",
2793 => x"00000000",
2794 => x"00000000",
2795 => x"00000000",
2796 => x"00000000",
2797 => x"00000000",
2798 => x"00000000",
2799 => x"00000000",
2800 => x"00000000",
2801 => x"00000000",
2802 => x"00000000",
2803 => x"00000000",
2804 => x"00000000",
2805 => x"00000000",
2806 => x"00000000",
2807 => x"00000000",
2808 => x"00000000",
2809 => x"00000000",
2810 => x"00000000",
2811 => x"00000000",
2812 => x"00000000",
2813 => x"00000000",
2814 => x"00000000",
2815 => x"00000000",
2816 => x"00000000",
2817 => x"00000000",
2818 => x"00000000",
2819 => x"00000000",
2820 => x"00000000",
2821 => x"00000000",
2822 => x"00000000",
2823 => x"00000000",
2824 => x"00000000",
2825 => x"00000000",
2826 => x"00000000",
2827 => x"00000000",
2828 => x"00000000",
2829 => x"00000000",
2830 => x"00000000",
2831 => x"00000000",
2832 => x"00000000",
2833 => x"00000000",
2834 => x"00000000",
2835 => x"00000000",
2836 => x"00000000",
2837 => x"00000000",
2838 => x"00000000",
2839 => x"00000000",
2840 => x"00000000",
2841 => x"00000000",
2842 => x"00000000",
2843 => x"00000000",
2844 => x"00000000",
2845 => x"00000000",
2846 => x"00000000",
2847 => x"00000000",
2848 => x"00000000",
2849 => x"00000000",
2850 => x"00000000",
2851 => x"00000000",
2852 => x"00000000",
2853 => x"00000000",
2854 => x"00000000",
2855 => x"00000000",
2856 => x"00000000",
2857 => x"00000000",
2858 => x"00000000",
2859 => x"00000000",
2860 => x"00000000",
2861 => x"00000000",
2862 => x"00000000",
2863 => x"00000000",
2864 => x"00000000",
2865 => x"00000000",
2866 => x"00000000",
2867 => x"00000000",
2868 => x"00000000",
2869 => x"00000000",
2870 => x"00000000",
2871 => x"00000000",
2872 => x"00000000",
2873 => x"00000000",
2874 => x"00000000",
2875 => x"00000000",
2876 => x"00000000",
2877 => x"00000000",
2878 => x"00000000",
2879 => x"00000000",
2880 => x"00000000",
2881 => x"00000000",
2882 => x"00000000",
2883 => x"00000000",
2884 => x"00000000",
2885 => x"00000000",
2886 => x"00000000",
2887 => x"00000000",
2888 => x"00000000",
2889 => x"00000000",
2890 => x"00000000",
2891 => x"00000000",
2892 => x"00000000",
2893 => x"00000000",
2894 => x"00000000",
2895 => x"00000000",
2896 => x"00000000",
2897 => x"00000000",
2898 => x"00000000",
2899 => x"ffffffff",
2900 => x"00000000",
2901 => x"00020000",
2902 => x"00000000",
2903 => x"00000000",
2904 => x"00002d58",
2905 => x"00002d58",
2906 => x"00002d60",
2907 => x"00002d60",
2908 => x"00002d68",
2909 => x"00002d68",
2910 => x"00002d70",
2911 => x"00002d70",
2912 => x"00002d78",
2913 => x"00002d78",
2914 => x"00002d80",
2915 => x"00002d80",
2916 => x"00002d88",
2917 => x"00002d88",
2918 => x"00002d90",
2919 => x"00002d90",
2920 => x"00002d98",
2921 => x"00002d98",
2922 => x"00002da0",
2923 => x"00002da0",
2924 => x"00002da8",
2925 => x"00002da8",
2926 => x"00002db0",
2927 => x"00002db0",
2928 => x"00002db8",
2929 => x"00002db8",
2930 => x"00002dc0",
2931 => x"00002dc0",
2932 => x"00002dc8",
2933 => x"00002dc8",
2934 => x"00002dd0",
2935 => x"00002dd0",
2936 => x"00002dd8",
2937 => x"00002dd8",
2938 => x"00002de0",
2939 => x"00002de0",
2940 => x"00002de8",
2941 => x"00002de8",
2942 => x"00002df0",
2943 => x"00002df0",
2944 => x"00002df8",
2945 => x"00002df8",
2946 => x"00002e00",
2947 => x"00002e00",
2948 => x"00002e08",
2949 => x"00002e08",
2950 => x"00002e10",
2951 => x"00002e10",
2952 => x"00002e18",
2953 => x"00002e18",
2954 => x"00002e20",
2955 => x"00002e20",
2956 => x"00002e28",
2957 => x"00002e28",
2958 => x"00002e30",
2959 => x"00002e30",
2960 => x"00002e38",
2961 => x"00002e38",
2962 => x"00002e40",
2963 => x"00002e40",
2964 => x"00002e48",
2965 => x"00002e48",
2966 => x"00002e50",
2967 => x"00002e50",
2968 => x"00002e58",
2969 => x"00002e58",
2970 => x"00002e60",
2971 => x"00002e60",
2972 => x"00002e68",
2973 => x"00002e68",
2974 => x"00002e70",
2975 => x"00002e70",
2976 => x"00002e78",
2977 => x"00002e78",
2978 => x"00002e80",
2979 => x"00002e80",
2980 => x"00002e88",
2981 => x"00002e88",
2982 => x"00002e90",
2983 => x"00002e90",
2984 => x"00002e98",
2985 => x"00002e98",
2986 => x"00002ea0",
2987 => x"00002ea0",
2988 => x"00002ea8",
2989 => x"00002ea8",
2990 => x"00002eb0",
2991 => x"00002eb0",
2992 => x"00002eb8",
2993 => x"00002eb8",
2994 => x"00002ec0",
2995 => x"00002ec0",
2996 => x"00002ec8",
2997 => x"00002ec8",
2998 => x"00002ed0",
2999 => x"00002ed0",
3000 => x"00002ed8",
3001 => x"00002ed8",
3002 => x"00002ee0",
3003 => x"00002ee0",
3004 => x"00002ee8",
3005 => x"00002ee8",
3006 => x"00002ef0",
3007 => x"00002ef0",
3008 => x"00002ef8",
3009 => x"00002ef8",
3010 => x"00002f00",
3011 => x"00002f00",
3012 => x"00002f08",
3013 => x"00002f08",
3014 => x"00002f10",
3015 => x"00002f10",
3016 => x"00002f18",
3017 => x"00002f18",
3018 => x"00002f20",
3019 => x"00002f20",
3020 => x"00002f28",
3021 => x"00002f28",
3022 => x"00002f30",
3023 => x"00002f30",
3024 => x"00002f38",
3025 => x"00002f38",
3026 => x"00002f40",
3027 => x"00002f40",
3028 => x"00002f48",
3029 => x"00002f48",
3030 => x"00002f50",
3031 => x"00002f50",
3032 => x"00002f58",
3033 => x"00002f58",
3034 => x"00002f60",
3035 => x"00002f60",
3036 => x"00002f68",
3037 => x"00002f68",
3038 => x"00002f70",
3039 => x"00002f70",
3040 => x"00002f78",
3041 => x"00002f78",
3042 => x"00002f80",
3043 => x"00002f80",
3044 => x"00002f88",
3045 => x"00002f88",
3046 => x"00002f90",
3047 => x"00002f90",
3048 => x"00002f98",
3049 => x"00002f98",
3050 => x"00002fa0",
3051 => x"00002fa0",
3052 => x"00002fa8",
3053 => x"00002fa8",
3054 => x"00002fb0",
3055 => x"00002fb0",
3056 => x"00002fb8",
3057 => x"00002fb8",
3058 => x"00002fc0",
3059 => x"00002fc0",
3060 => x"00002fc8",
3061 => x"00002fc8",
3062 => x"00002fd0",
3063 => x"00002fd0",
3064 => x"00002fd8",
3065 => x"00002fd8",
3066 => x"00002fe0",
3067 => x"00002fe0",
3068 => x"00002fe8",
3069 => x"00002fe8",
3070 => x"00002ff0",
3071 => x"00002ff0",
3072 => x"00002ff8",
3073 => x"00002ff8",
3074 => x"00003000",
3075 => x"00003000",
3076 => x"00003008",
3077 => x"00003008",
3078 => x"00003010",
3079 => x"00003010",
3080 => x"00003018",
3081 => x"00003018",
3082 => x"00003020",
3083 => x"00003020",
3084 => x"00003028",
3085 => x"00003028",
3086 => x"00003030",
3087 => x"00003030",
3088 => x"00003038",
3089 => x"00003038",
3090 => x"00003040",
3091 => x"00003040",
3092 => x"00003048",
3093 => x"00003048",
3094 => x"00003050",
3095 => x"00003050",
3096 => x"00003058",
3097 => x"00003058",
3098 => x"00003060",
3099 => x"00003060",
3100 => x"00003068",
3101 => x"00003068",
3102 => x"00003070",
3103 => x"00003070",
3104 => x"00003078",
3105 => x"00003078",
3106 => x"00003080",
3107 => x"00003080",
3108 => x"00003088",
3109 => x"00003088",
3110 => x"00003090",
3111 => x"00003090",
3112 => x"00003098",
3113 => x"00003098",
3114 => x"000030a0",
3115 => x"000030a0",
3116 => x"000030a8",
3117 => x"000030a8",
3118 => x"000030b0",
3119 => x"000030b0",
3120 => x"000030b8",
3121 => x"000030b8",
3122 => x"000030c0",
3123 => x"000030c0",
3124 => x"000030c8",
3125 => x"000030c8",
3126 => x"000030d0",
3127 => x"000030d0",
3128 => x"000030d8",
3129 => x"000030d8",
3130 => x"000030e0",
3131 => x"000030e0",
3132 => x"000030e8",
3133 => x"000030e8",
3134 => x"000030f0",
3135 => x"000030f0",
3136 => x"000030f8",
3137 => x"000030f8",
3138 => x"00003100",
3139 => x"00003100",
3140 => x"00003108",
3141 => x"00003108",
3142 => x"00003110",
3143 => x"00003110",
3144 => x"00003118",
3145 => x"00003118",
3146 => x"00003120",
3147 => x"00003120",
3148 => x"00003128",
3149 => x"00003128",
3150 => x"00003130",
3151 => x"00003130",
3152 => x"00003138",
3153 => x"00003138",
3154 => x"00003140",
3155 => x"00003140",
3156 => x"00003148",
3157 => x"00003148",
3158 => x"00003150",
3159 => x"00003150",
3160 => x"00002970",
3161 => x"ffffffff",
3162 => x"00000000",
3163 => x"ffffffff",
3164 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		mem_busy<=mem_writeEnable or mem_readEnable;
		if (mem_writeEnable = '1') then
			ram(conv_integer(mem_addr(maxAddrBit downto minAddrBit))) := mem_write;
		end if;
		if (mem_readEnable = '1') then
			mem_read <= ram(conv_integer(mem_addr(maxAddrBit downto minAddrBit)));
		end if;
	end if;
end process;




end dram_arch;
