-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0ba7900c",
     3 => x"3a0b0b0b",
     4 => x"a4d80400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0ba5982d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba6",
   162 => x"fc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8a",
   171 => x"b12d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8b",
   179 => x"e32d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0ba78c0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f9e",
   257 => x"b83f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104a7",
   280 => x"8c08802e",
   281 => x"a138a790",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"b6f80c82",
   286 => x"a0800bb6",
   287 => x"fc0c8290",
   288 => x"800bb780",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0bb6",
   292 => x"f80cf880",
   293 => x"8082800b",
   294 => x"b6fc0cf8",
   295 => x"80808480",
   296 => x"0bb7800c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0bb6f8",
   300 => x"0c80c0a8",
   301 => x"80940bb6",
   302 => x"fc0c0b0b",
   303 => x"0ba6e80b",
   304 => x"b7800c04",
   305 => x"ff3d0db7",
   306 => x"84335170",
   307 => x"a338a798",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"a7980c70",
   312 => x"2da79808",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0bb78434",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0bb6",
   319 => x"f408802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0bb6f4",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"803d0df8",
   330 => x"80809080",
   331 => x"085183fd",
   332 => x"3f8c0802",
   333 => x"8c0cf93d",
   334 => x"0d800b8c",
   335 => x"08fc050c",
   336 => x"8c088805",
   337 => x"088025ab",
   338 => x"388c0888",
   339 => x"0508308c",
   340 => x"0888050c",
   341 => x"800b8c08",
   342 => x"f4050c8c",
   343 => x"08fc0508",
   344 => x"8838810b",
   345 => x"8c08f405",
   346 => x"0c8c08f4",
   347 => x"05088c08",
   348 => x"fc050c8c",
   349 => x"088c0508",
   350 => x"8025ab38",
   351 => x"8c088c05",
   352 => x"08308c08",
   353 => x"8c050c80",
   354 => x"0b8c08f0",
   355 => x"050c8c08",
   356 => x"fc050888",
   357 => x"38810b8c",
   358 => x"08f0050c",
   359 => x"8c08f005",
   360 => x"088c08fc",
   361 => x"050c8053",
   362 => x"8c088c05",
   363 => x"08528c08",
   364 => x"88050851",
   365 => x"81a73f80",
   366 => x"08708c08",
   367 => x"f8050c54",
   368 => x"8c08fc05",
   369 => x"08802e8c",
   370 => x"388c08f8",
   371 => x"0508308c",
   372 => x"08f8050c",
   373 => x"8c08f805",
   374 => x"0870800c",
   375 => x"54893d0d",
   376 => x"8c0c048c",
   377 => x"08028c0c",
   378 => x"fb3d0d80",
   379 => x"0b8c08fc",
   380 => x"050c8c08",
   381 => x"88050880",
   382 => x"2593388c",
   383 => x"08880508",
   384 => x"308c0888",
   385 => x"050c810b",
   386 => x"8c08fc05",
   387 => x"0c8c088c",
   388 => x"05088025",
   389 => x"8c388c08",
   390 => x"8c050830",
   391 => x"8c088c05",
   392 => x"0c81538c",
   393 => x"088c0508",
   394 => x"528c0888",
   395 => x"050851ad",
   396 => x"3f800870",
   397 => x"8c08f805",
   398 => x"0c548c08",
   399 => x"fc050880",
   400 => x"2e8c388c",
   401 => x"08f80508",
   402 => x"308c08f8",
   403 => x"050c8c08",
   404 => x"f8050870",
   405 => x"800c5487",
   406 => x"3d0d8c0c",
   407 => x"048c0802",
   408 => x"8c0cfd3d",
   409 => x"0d810b8c",
   410 => x"08fc050c",
   411 => x"800b8c08",
   412 => x"f8050c8c",
   413 => x"088c0508",
   414 => x"8c088805",
   415 => x"0827ac38",
   416 => x"8c08fc05",
   417 => x"08802ea3",
   418 => x"38800b8c",
   419 => x"088c0508",
   420 => x"2499388c",
   421 => x"088c0508",
   422 => x"108c088c",
   423 => x"050c8c08",
   424 => x"fc050810",
   425 => x"8c08fc05",
   426 => x"0cc9398c",
   427 => x"08fc0508",
   428 => x"802e80c9",
   429 => x"388c088c",
   430 => x"05088c08",
   431 => x"88050826",
   432 => x"a1388c08",
   433 => x"8805088c",
   434 => x"088c0508",
   435 => x"318c0888",
   436 => x"050c8c08",
   437 => x"f805088c",
   438 => x"08fc0508",
   439 => x"078c08f8",
   440 => x"050c8c08",
   441 => x"fc050881",
   442 => x"2a8c08fc",
   443 => x"050c8c08",
   444 => x"8c050881",
   445 => x"2a8c088c",
   446 => x"050cffaf",
   447 => x"398c0890",
   448 => x"0508802e",
   449 => x"8f388c08",
   450 => x"88050870",
   451 => x"8c08f405",
   452 => x"0c518d39",
   453 => x"8c08f805",
   454 => x"08708c08",
   455 => x"f4050c51",
   456 => x"8c08f405",
   457 => x"08800c85",
   458 => x"3d0d8c0c",
   459 => x"04803d0d",
   460 => x"865182fd",
   461 => x"3f815196",
   462 => x"dc3ffd3d",
   463 => x"0d755384",
   464 => x"d8130880",
   465 => x"2e8a3880",
   466 => x"5372800c",
   467 => x"853d0d04",
   468 => x"81805272",
   469 => x"5183d23f",
   470 => x"800884d8",
   471 => x"140cff53",
   472 => x"8008802e",
   473 => x"e4388008",
   474 => x"549f5380",
   475 => x"74708405",
   476 => x"560cff13",
   477 => x"53807324",
   478 => x"ce388074",
   479 => x"70840556",
   480 => x"0cff1353",
   481 => x"728025e3",
   482 => x"38ffbc39",
   483 => x"fd3d0d75",
   484 => x"7755539f",
   485 => x"74278d38",
   486 => x"96730cff",
   487 => x"5271800c",
   488 => x"853d0d04",
   489 => x"84d81308",
   490 => x"5271802e",
   491 => x"93387310",
   492 => x"10127008",
   493 => x"79720c51",
   494 => x"5271800c",
   495 => x"853d0d04",
   496 => x"7251fef6",
   497 => x"3fff5280",
   498 => x"08d33884",
   499 => x"d8130874",
   500 => x"10101170",
   501 => x"087a720c",
   502 => x"515152dd",
   503 => x"39f93d0d",
   504 => x"797b5856",
   505 => x"769f2680",
   506 => x"e83884d8",
   507 => x"16085473",
   508 => x"802eaa38",
   509 => x"76101014",
   510 => x"70085555",
   511 => x"73802eba",
   512 => x"38805873",
   513 => x"812e8f38",
   514 => x"73ff2ea3",
   515 => x"3880750c",
   516 => x"7651732d",
   517 => x"80587780",
   518 => x"0c893d0d",
   519 => x"047551fe",
   520 => x"993fff58",
   521 => x"8008ef38",
   522 => x"84d81608",
   523 => x"54c63996",
   524 => x"760c810b",
   525 => x"800c893d",
   526 => x"0d047551",
   527 => x"81e73f76",
   528 => x"53800852",
   529 => x"755181a9",
   530 => x"3f800880",
   531 => x"0c893d0d",
   532 => x"0496760c",
   533 => x"ff0b800c",
   534 => x"893d0d04",
   535 => x"fc3d0d76",
   536 => x"785653ff",
   537 => x"54749f26",
   538 => x"b13884d8",
   539 => x"13085271",
   540 => x"802eae38",
   541 => x"74101012",
   542 => x"70085353",
   543 => x"81547180",
   544 => x"2e983882",
   545 => x"5471ff2e",
   546 => x"91388354",
   547 => x"71812e8a",
   548 => x"3880730c",
   549 => x"7451712d",
   550 => x"80547380",
   551 => x"0c863d0d",
   552 => x"047251fd",
   553 => x"953f8008",
   554 => x"f13884d8",
   555 => x"130852c4",
   556 => x"39ff3d0d",
   557 => x"7352a79c",
   558 => x"0851fea1",
   559 => x"3f833d0d",
   560 => x"04fe3d0d",
   561 => x"75537452",
   562 => x"a79c0851",
   563 => x"fdbe3f84",
   564 => x"3d0d0480",
   565 => x"3d0da79c",
   566 => x"0851fcde",
   567 => x"3f823d0d",
   568 => x"04ff3d0d",
   569 => x"7352a79c",
   570 => x"0851fef0",
   571 => x"3f833d0d",
   572 => x"04fc3d0d",
   573 => x"800bb790",
   574 => x"0c785277",
   575 => x"5192973f",
   576 => x"80085480",
   577 => x"08ff2e88",
   578 => x"3873800c",
   579 => x"863d0d04",
   580 => x"b7900855",
   581 => x"74802ef1",
   582 => x"38767571",
   583 => x"0c537380",
   584 => x"0c863d0d",
   585 => x"0491ea3f",
   586 => x"04f33d0d",
   587 => x"7f618b11",
   588 => x"70f8065c",
   589 => x"55555e72",
   590 => x"96268338",
   591 => x"90598079",
   592 => x"24747a26",
   593 => x"07538054",
   594 => x"72742e09",
   595 => x"810680ca",
   596 => x"387d518b",
   597 => x"963f7883",
   598 => x"f72680c5",
   599 => x"3878832a",
   600 => x"70101010",
   601 => x"aed8058c",
   602 => x"11085959",
   603 => x"5a76782e",
   604 => x"83a73884",
   605 => x"1708fc06",
   606 => x"568c1708",
   607 => x"88180871",
   608 => x"8c120c88",
   609 => x"120c5875",
   610 => x"17841108",
   611 => x"81078412",
   612 => x"0c537d51",
   613 => x"8ad63f88",
   614 => x"17547380",
   615 => x"0c8f3d0d",
   616 => x"0478892a",
   617 => x"79832a5b",
   618 => x"5372802e",
   619 => x"bf387886",
   620 => x"2ab8055a",
   621 => x"847327b4",
   622 => x"3880db13",
   623 => x"5a947327",
   624 => x"ab38788c",
   625 => x"2a80ee05",
   626 => x"5a80d473",
   627 => x"279e3878",
   628 => x"8f2a80f7",
   629 => x"055a82d4",
   630 => x"73279138",
   631 => x"78922a80",
   632 => x"fc055a8a",
   633 => x"d4732784",
   634 => x"3880fe5a",
   635 => x"79101010",
   636 => x"aed8058c",
   637 => x"11085855",
   638 => x"76752ea3",
   639 => x"38841708",
   640 => x"fc06707a",
   641 => x"31555673",
   642 => x"8f2488aa",
   643 => x"38738025",
   644 => x"fee7388c",
   645 => x"17085776",
   646 => x"752e0981",
   647 => x"06df3881",
   648 => x"1a5aaee8",
   649 => x"085776ae",
   650 => x"e02e82b7",
   651 => x"38841708",
   652 => x"fc06707a",
   653 => x"31555673",
   654 => x"8f2481f3",
   655 => x"38aee00b",
   656 => x"aeec0cae",
   657 => x"e00baee8",
   658 => x"0c738025",
   659 => x"feb93883",
   660 => x"ff762783",
   661 => x"d2387589",
   662 => x"2a76832a",
   663 => x"55537280",
   664 => x"2ebf3875",
   665 => x"862ab805",
   666 => x"54847327",
   667 => x"b43880db",
   668 => x"13549473",
   669 => x"27ab3875",
   670 => x"8c2a80ee",
   671 => x"055480d4",
   672 => x"73279e38",
   673 => x"758f2a80",
   674 => x"f7055482",
   675 => x"d4732791",
   676 => x"3875922a",
   677 => x"80fc0554",
   678 => x"8ad47327",
   679 => x"843880fe",
   680 => x"54731010",
   681 => x"10aed805",
   682 => x"88110856",
   683 => x"5874782e",
   684 => x"86af3884",
   685 => x"1508fc06",
   686 => x"53757327",
   687 => x"8d388815",
   688 => x"08557478",
   689 => x"2e098106",
   690 => x"ea388c15",
   691 => x"08aed80b",
   692 => x"84050871",
   693 => x"8c1a0c76",
   694 => x"881a0c78",
   695 => x"88130c78",
   696 => x"8c180c5d",
   697 => x"58795380",
   698 => x"7a2483d7",
   699 => x"3872822c",
   700 => x"81712b5c",
   701 => x"537a7c26",
   702 => x"8193387b",
   703 => x"7b065372",
   704 => x"82e33879",
   705 => x"fc068405",
   706 => x"5a7a1070",
   707 => x"7d06545b",
   708 => x"7282d238",
   709 => x"841a5af1",
   710 => x"3988178c",
   711 => x"11085858",
   712 => x"76782e09",
   713 => x"8106fccb",
   714 => x"38821a5a",
   715 => x"fdf43978",
   716 => x"17798107",
   717 => x"84190c70",
   718 => x"aeec0c70",
   719 => x"aee80cae",
   720 => x"e00b8c12",
   721 => x"0c8c1108",
   722 => x"88120c74",
   723 => x"81078412",
   724 => x"0c741175",
   725 => x"710c5153",
   726 => x"7d518790",
   727 => x"3f881754",
   728 => x"fcb839ae",
   729 => x"d80b8405",
   730 => x"087a545c",
   731 => x"798025fe",
   732 => x"fc3882cf",
   733 => x"397a097c",
   734 => x"0670aed8",
   735 => x"0b84050c",
   736 => x"5c7a105b",
   737 => x"7a7c2685",
   738 => x"387a859a",
   739 => x"38aed80b",
   740 => x"88050870",
   741 => x"841208fc",
   742 => x"06707c31",
   743 => x"7c72268f",
   744 => x"72250757",
   745 => x"575c5d55",
   746 => x"72802e80",
   747 => x"d738797a",
   748 => x"16aed008",
   749 => x"1b90115a",
   750 => x"55575bae",
   751 => x"cc08ff2e",
   752 => x"8838a08f",
   753 => x"13e08006",
   754 => x"5776527d",
   755 => x"51869e3f",
   756 => x"80085480",
   757 => x"08ff2e8f",
   758 => x"38800876",
   759 => x"27828f38",
   760 => x"74aed82e",
   761 => x"828838ae",
   762 => x"d80b8805",
   763 => x"08558415",
   764 => x"08fc0670",
   765 => x"7a317a72",
   766 => x"268f7225",
   767 => x"07525553",
   768 => x"7283d138",
   769 => x"74798107",
   770 => x"84170c79",
   771 => x"1670aed8",
   772 => x"0b88050c",
   773 => x"75810784",
   774 => x"120c547e",
   775 => x"525785cc",
   776 => x"3f881754",
   777 => x"faf43975",
   778 => x"832a7054",
   779 => x"54807424",
   780 => x"81973872",
   781 => x"822c8171",
   782 => x"2baedc08",
   783 => x"0770aed8",
   784 => x"0b84050c",
   785 => x"75101010",
   786 => x"aed80588",
   787 => x"1108585a",
   788 => x"5d53778c",
   789 => x"180c7488",
   790 => x"180c7688",
   791 => x"190c768c",
   792 => x"160cfd81",
   793 => x"39797a10",
   794 => x"1010aed8",
   795 => x"05705759",
   796 => x"5d8c1508",
   797 => x"5776752e",
   798 => x"a3388417",
   799 => x"08fc0670",
   800 => x"7a315556",
   801 => x"738f2483",
   802 => x"b6387380",
   803 => x"2583ea38",
   804 => x"8c170857",
   805 => x"76752e09",
   806 => x"8106df38",
   807 => x"8815811b",
   808 => x"70830655",
   809 => x"5b5572c9",
   810 => x"387c8306",
   811 => x"5372802e",
   812 => x"fdc338ff",
   813 => x"1df81959",
   814 => x"5d881808",
   815 => x"782eea38",
   816 => x"fdbf3983",
   817 => x"1a53fca5",
   818 => x"39831470",
   819 => x"822c8171",
   820 => x"2baedc08",
   821 => x"0770aed8",
   822 => x"0b84050c",
   823 => x"76101010",
   824 => x"aed80588",
   825 => x"1108595b",
   826 => x"5e5153fe",
   827 => x"e539ae9c",
   828 => x"08175880",
   829 => x"08762e81",
   830 => x"8738aecc",
   831 => x"08ff2e83",
   832 => x"d8387376",
   833 => x"3118ae9c",
   834 => x"0c738706",
   835 => x"70575372",
   836 => x"802e8838",
   837 => x"88733170",
   838 => x"15555676",
   839 => x"149fff06",
   840 => x"a0807131",
   841 => x"1770547f",
   842 => x"53575383",
   843 => x"c03f8008",
   844 => x"538008ff",
   845 => x"2e819638",
   846 => x"ae9c0816",
   847 => x"70ae9c0c",
   848 => x"7475aed8",
   849 => x"0b88050c",
   850 => x"74763118",
   851 => x"70810751",
   852 => x"5556587b",
   853 => x"aed82e83",
   854 => x"8b38798f",
   855 => x"2682be38",
   856 => x"810b8415",
   857 => x"0c841508",
   858 => x"fc06707a",
   859 => x"317a7226",
   860 => x"8f722507",
   861 => x"52555372",
   862 => x"802efd88",
   863 => x"3880d539",
   864 => x"80089fff",
   865 => x"065372fe",
   866 => x"f13877ae",
   867 => x"9c0caed8",
   868 => x"0b880508",
   869 => x"7b188107",
   870 => x"84120c55",
   871 => x"aec80878",
   872 => x"27853877",
   873 => x"aec80cae",
   874 => x"c4087827",
   875 => x"fcc03877",
   876 => x"aec40c84",
   877 => x"1508fc06",
   878 => x"707a317a",
   879 => x"72268f72",
   880 => x"25075255",
   881 => x"5372802e",
   882 => x"fcba3888",
   883 => x"39807454",
   884 => x"56fee539",
   885 => x"7d518294",
   886 => x"3f800b80",
   887 => x"0c8f3d0d",
   888 => x"04735380",
   889 => x"7424a738",
   890 => x"72822c81",
   891 => x"712baedc",
   892 => x"080770ae",
   893 => x"d80b8405",
   894 => x"0c5d5377",
   895 => x"8c180c74",
   896 => x"88180c76",
   897 => x"88190c76",
   898 => x"8c160cf9",
   899 => x"d8398314",
   900 => x"70822c81",
   901 => x"712baedc",
   902 => x"080770ae",
   903 => x"d80b8405",
   904 => x"0c5e5153",
   905 => x"d6397b7b",
   906 => x"065372fc",
   907 => x"b838841a",
   908 => x"7b105c5a",
   909 => x"f139ff1a",
   910 => x"8111515a",
   911 => x"f7e43978",
   912 => x"17798107",
   913 => x"84190c8c",
   914 => x"18088819",
   915 => x"08718c12",
   916 => x"0c88120c",
   917 => x"5970aeec",
   918 => x"0c70aee8",
   919 => x"0caee00b",
   920 => x"8c120c8c",
   921 => x"11088812",
   922 => x"0c748107",
   923 => x"84120c74",
   924 => x"1175710c",
   925 => x"5153f9e0",
   926 => x"39751784",
   927 => x"11088107",
   928 => x"84120c53",
   929 => x"8c170888",
   930 => x"1808718c",
   931 => x"120c8812",
   932 => x"0c587d51",
   933 => x"80d63f88",
   934 => x"1754f5fe",
   935 => x"39728415",
   936 => x"0cf41af8",
   937 => x"0670841e",
   938 => x"08810607",
   939 => x"841e0c70",
   940 => x"1d545b85",
   941 => x"0b84140c",
   942 => x"850b8814",
   943 => x"0c8f7b27",
   944 => x"fdda3888",
   945 => x"1c527d51",
   946 => x"82823fae",
   947 => x"d80b8805",
   948 => x"08ae9c08",
   949 => x"5955fdc4",
   950 => x"3977ae9c",
   951 => x"0c73aecc",
   952 => x"0cfca639",
   953 => x"7284150c",
   954 => x"fdb23904",
   955 => x"04fd3d0d",
   956 => x"800bb790",
   957 => x"0c765186",
   958 => x"b23f8008",
   959 => x"538008ff",
   960 => x"2e883872",
   961 => x"800c853d",
   962 => x"0d04b790",
   963 => x"08547380",
   964 => x"2ef13875",
   965 => x"74710c52",
   966 => x"72800c85",
   967 => x"3d0d04fb",
   968 => x"3d0d7770",
   969 => x"5256c43f",
   970 => x"aed80b88",
   971 => x"05088411",
   972 => x"08fc0670",
   973 => x"7b319fef",
   974 => x"05e08006",
   975 => x"e0800556",
   976 => x"5653a080",
   977 => x"74249338",
   978 => x"80527551",
   979 => x"ff9f3fae",
   980 => x"e0081553",
   981 => x"7280082e",
   982 => x"8f387551",
   983 => x"ff8e3f80",
   984 => x"5372800c",
   985 => x"873d0d04",
   986 => x"73305275",
   987 => x"51fefe3f",
   988 => x"8008ff2e",
   989 => x"a538aed8",
   990 => x"0b880508",
   991 => x"75753181",
   992 => x"0784120c",
   993 => x"53ae9c08",
   994 => x"7431ae9c",
   995 => x"0c7551fe",
   996 => x"db3f810b",
   997 => x"800c873d",
   998 => x"0d048052",
   999 => x"7551fecd",
  1000 => x"3faed80b",
  1001 => x"88050880",
  1002 => x"08713156",
  1003 => x"538f7525",
  1004 => x"ffa83880",
  1005 => x"08aecc08",
  1006 => x"31ae9c0c",
  1007 => x"74810784",
  1008 => x"140c7551",
  1009 => x"fea63f80",
  1010 => x"53ff9639",
  1011 => x"f63d0d7c",
  1012 => x"7e545b72",
  1013 => x"802e8280",
  1014 => x"387a51fe",
  1015 => x"8e3ff813",
  1016 => x"84110870",
  1017 => x"fe067013",
  1018 => x"841108fc",
  1019 => x"065d5859",
  1020 => x"5458aee0",
  1021 => x"08752e82",
  1022 => x"d8387884",
  1023 => x"160c8073",
  1024 => x"8106545a",
  1025 => x"727a2e81",
  1026 => x"d3387815",
  1027 => x"84110881",
  1028 => x"06515372",
  1029 => x"9f387817",
  1030 => x"577981e3",
  1031 => x"38881508",
  1032 => x"5372aee0",
  1033 => x"2e82f138",
  1034 => x"8c150870",
  1035 => x"8c150c73",
  1036 => x"88120c56",
  1037 => x"76810784",
  1038 => x"190c7618",
  1039 => x"77710c53",
  1040 => x"79819038",
  1041 => x"83ff7727",
  1042 => x"81c63876",
  1043 => x"892a7783",
  1044 => x"2a565372",
  1045 => x"802ebf38",
  1046 => x"76862ab8",
  1047 => x"05558473",
  1048 => x"27b43880",
  1049 => x"db135594",
  1050 => x"7327ab38",
  1051 => x"768c2a80",
  1052 => x"ee055580",
  1053 => x"d473279e",
  1054 => x"38768f2a",
  1055 => x"80f70555",
  1056 => x"82d47327",
  1057 => x"91387692",
  1058 => x"2a80fc05",
  1059 => x"558ad473",
  1060 => x"27843880",
  1061 => x"fe557410",
  1062 => x"1010aed8",
  1063 => x"05881108",
  1064 => x"55567376",
  1065 => x"2e82a938",
  1066 => x"841408fc",
  1067 => x"06537673",
  1068 => x"278d3888",
  1069 => x"14085473",
  1070 => x"762e0981",
  1071 => x"06ea388c",
  1072 => x"1408708c",
  1073 => x"1a0c7488",
  1074 => x"1a0c7888",
  1075 => x"120c5677",
  1076 => x"8c150c7a",
  1077 => x"51fc953f",
  1078 => x"8c3d0d04",
  1079 => x"77087871",
  1080 => x"31597705",
  1081 => x"88190854",
  1082 => x"5772aee0",
  1083 => x"2e80dd38",
  1084 => x"8c180870",
  1085 => x"8c150c73",
  1086 => x"88120c56",
  1087 => x"fe8c3988",
  1088 => x"15088c16",
  1089 => x"08708c13",
  1090 => x"0c578817",
  1091 => x"0cfea539",
  1092 => x"76832a70",
  1093 => x"54558075",
  1094 => x"24819238",
  1095 => x"72822c81",
  1096 => x"712baedc",
  1097 => x"0807aed8",
  1098 => x"0b84050c",
  1099 => x"53741010",
  1100 => x"10aed805",
  1101 => x"88110855",
  1102 => x"56758c19",
  1103 => x"0c738819",
  1104 => x"0c778817",
  1105 => x"0c778c15",
  1106 => x"0cff8839",
  1107 => x"815afdba",
  1108 => x"39781773",
  1109 => x"81065457",
  1110 => x"72983877",
  1111 => x"08787131",
  1112 => x"5977058c",
  1113 => x"1908881a",
  1114 => x"08718c12",
  1115 => x"0c88120c",
  1116 => x"57577681",
  1117 => x"0784190c",
  1118 => x"77aed80b",
  1119 => x"88050cae",
  1120 => x"d4087726",
  1121 => x"fecd38ae",
  1122 => x"d008527a",
  1123 => x"51fb903f",
  1124 => x"7a51fad8",
  1125 => x"3ffec139",
  1126 => x"81788c15",
  1127 => x"0c788815",
  1128 => x"0c738c1a",
  1129 => x"0c73881a",
  1130 => x"0c5afd88",
  1131 => x"39831570",
  1132 => x"822c8171",
  1133 => x"2baedc08",
  1134 => x"07aed80b",
  1135 => x"84050c51",
  1136 => x"53741010",
  1137 => x"10aed805",
  1138 => x"88110855",
  1139 => x"56feea39",
  1140 => x"74538075",
  1141 => x"24a53872",
  1142 => x"822c8171",
  1143 => x"2baedc08",
  1144 => x"07aed80b",
  1145 => x"84050c53",
  1146 => x"758c190c",
  1147 => x"7388190c",
  1148 => x"7788170c",
  1149 => x"778c150c",
  1150 => x"fdd93983",
  1151 => x"1570822c",
  1152 => x"81712bae",
  1153 => x"dc0807ae",
  1154 => x"d80b8405",
  1155 => x"0c5153d8",
  1156 => x"39810b80",
  1157 => x"0c04803d",
  1158 => x"0d72812e",
  1159 => x"8938800b",
  1160 => x"800c823d",
  1161 => x"0d047351",
  1162 => x"80eb3ffe",
  1163 => x"3d0db788",
  1164 => x"08517088",
  1165 => x"38b79470",
  1166 => x"b7880c51",
  1167 => x"70751252",
  1168 => x"52ff5370",
  1169 => x"87fb8080",
  1170 => x"26873870",
  1171 => x"b7880c71",
  1172 => x"5372800c",
  1173 => x"843d0d04",
  1174 => x"fd3d0d80",
  1175 => x"0ba79008",
  1176 => x"54547281",
  1177 => x"2e983873",
  1178 => x"b78c0ce3",
  1179 => x"f23fe390",
  1180 => x"3fb6e052",
  1181 => x"8151e5ac",
  1182 => x"3f800851",
  1183 => x"9e3f72b7",
  1184 => x"8c0ce3db",
  1185 => x"3fe2f93f",
  1186 => x"b6e05281",
  1187 => x"51e5953f",
  1188 => x"80085187",
  1189 => x"3f00ff39",
  1190 => x"00ff39f7",
  1191 => x"3d0d7ba7",
  1192 => x"9c0882c8",
  1193 => x"11085a54",
  1194 => x"5a77802e",
  1195 => x"80d93881",
  1196 => x"88188419",
  1197 => x"08ff0581",
  1198 => x"712b5955",
  1199 => x"59807424",
  1200 => x"80e93880",
  1201 => x"7424b538",
  1202 => x"73822b78",
  1203 => x"11880556",
  1204 => x"56818019",
  1205 => x"08770653",
  1206 => x"72802eb5",
  1207 => x"38781670",
  1208 => x"08535379",
  1209 => x"51740853",
  1210 => x"722dff14",
  1211 => x"fc17fc17",
  1212 => x"79812c5a",
  1213 => x"57575473",
  1214 => x"8025d638",
  1215 => x"77085877",
  1216 => x"ffad38a7",
  1217 => x"9c0853bc",
  1218 => x"1308a538",
  1219 => x"7951ff85",
  1220 => x"3f740853",
  1221 => x"722dff14",
  1222 => x"fc17fc17",
  1223 => x"79812c5a",
  1224 => x"57575473",
  1225 => x"8025ffa9",
  1226 => x"38d23980",
  1227 => x"57ff9439",
  1228 => x"7251bc13",
  1229 => x"0853722d",
  1230 => x"7951fed9",
  1231 => x"3fff3d0d",
  1232 => x"b6e80bfc",
  1233 => x"05700852",
  1234 => x"5270ff2e",
  1235 => x"9138702d",
  1236 => x"fc127008",
  1237 => x"525270ff",
  1238 => x"2e098106",
  1239 => x"f138833d",
  1240 => x"0d0404e2",
  1241 => x"df3f0400",
  1242 => x"00000040",
  1243 => x"43000000",
  1244 => x"64756d6d",
  1245 => x"792e6578",
  1246 => x"65000000",
  1247 => x"00ffffff",
  1248 => x"ff00ffff",
  1249 => x"ffff00ff",
  1250 => x"ffffff00",
  1251 => x"00000000",
  1252 => x"00000000",
  1253 => x"00000000",
  1254 => x"00001b70",
  1255 => x"000013a0",
  1256 => x"00000000",
  1257 => x"00001608",
  1258 => x"00001664",
  1259 => x"000016c0",
  1260 => x"00000000",
  1261 => x"00000000",
  1262 => x"00000000",
  1263 => x"00000000",
  1264 => x"00000000",
  1265 => x"00000000",
  1266 => x"00000000",
  1267 => x"00000000",
  1268 => x"00000000",
  1269 => x"0000136c",
  1270 => x"00000000",
  1271 => x"00000000",
  1272 => x"00000000",
  1273 => x"00000000",
  1274 => x"00000000",
  1275 => x"00000000",
  1276 => x"00000000",
  1277 => x"00000000",
  1278 => x"00000000",
  1279 => x"00000000",
  1280 => x"00000000",
  1281 => x"00000000",
  1282 => x"00000000",
  1283 => x"00000000",
  1284 => x"00000000",
  1285 => x"00000000",
  1286 => x"00000000",
  1287 => x"00000000",
  1288 => x"00000000",
  1289 => x"00000000",
  1290 => x"00000000",
  1291 => x"00000000",
  1292 => x"00000000",
  1293 => x"00000000",
  1294 => x"00000000",
  1295 => x"00000000",
  1296 => x"00000000",
  1297 => x"00000000",
  1298 => x"00000001",
  1299 => x"330eabcd",
  1300 => x"1234e66d",
  1301 => x"deec0005",
  1302 => x"000b0000",
  1303 => x"00000000",
  1304 => x"00000000",
  1305 => x"00000000",
  1306 => x"00000000",
  1307 => x"00000000",
  1308 => x"00000000",
  1309 => x"00000000",
  1310 => x"00000000",
  1311 => x"00000000",
  1312 => x"00000000",
  1313 => x"00000000",
  1314 => x"00000000",
  1315 => x"00000000",
  1316 => x"00000000",
  1317 => x"00000000",
  1318 => x"00000000",
  1319 => x"00000000",
  1320 => x"00000000",
  1321 => x"00000000",
  1322 => x"00000000",
  1323 => x"00000000",
  1324 => x"00000000",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00000000",
  1329 => x"00000000",
  1330 => x"00000000",
  1331 => x"00000000",
  1332 => x"00000000",
  1333 => x"00000000",
  1334 => x"00000000",
  1335 => x"00000000",
  1336 => x"00000000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"00000000",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"00000000",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000000",
  1404 => x"00000000",
  1405 => x"00000000",
  1406 => x"00000000",
  1407 => x"00000000",
  1408 => x"00000000",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00000000",
  1414 => x"00000000",
  1415 => x"00000000",
  1416 => x"00000000",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"00000000",
  1420 => x"00000000",
  1421 => x"00000000",
  1422 => x"00000000",
  1423 => x"00000000",
  1424 => x"00000000",
  1425 => x"00000000",
  1426 => x"00000000",
  1427 => x"00000000",
  1428 => x"00000000",
  1429 => x"00000000",
  1430 => x"00000000",
  1431 => x"00000000",
  1432 => x"00000000",
  1433 => x"00000000",
  1434 => x"00000000",
  1435 => x"00000000",
  1436 => x"00000000",
  1437 => x"00000000",
  1438 => x"00000000",
  1439 => x"00000000",
  1440 => x"00000000",
  1441 => x"00000000",
  1442 => x"00000000",
  1443 => x"00000000",
  1444 => x"00000000",
  1445 => x"00000000",
  1446 => x"00000000",
  1447 => x"00000000",
  1448 => x"00000000",
  1449 => x"00000000",
  1450 => x"00000000",
  1451 => x"00000000",
  1452 => x"00000000",
  1453 => x"00000000",
  1454 => x"00000000",
  1455 => x"00000000",
  1456 => x"00000000",
  1457 => x"00000000",
  1458 => x"00000000",
  1459 => x"00000000",
  1460 => x"00000000",
  1461 => x"00000000",
  1462 => x"00000000",
  1463 => x"00000000",
  1464 => x"00000000",
  1465 => x"00000000",
  1466 => x"00000000",
  1467 => x"00000000",
  1468 => x"00000000",
  1469 => x"00000000",
  1470 => x"00000000",
  1471 => x"00000000",
  1472 => x"00000000",
  1473 => x"00000000",
  1474 => x"00000000",
  1475 => x"00000000",
  1476 => x"00000000",
  1477 => x"00000000",
  1478 => x"00000000",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000000",
  1483 => x"00000000",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"ffffffff",
  1492 => x"00000000",
  1493 => x"00020000",
  1494 => x"00000000",
  1495 => x"00000000",
  1496 => x"00001758",
  1497 => x"00001758",
  1498 => x"00001760",
  1499 => x"00001760",
  1500 => x"00001768",
  1501 => x"00001768",
  1502 => x"00001770",
  1503 => x"00001770",
  1504 => x"00001778",
  1505 => x"00001778",
  1506 => x"00001780",
  1507 => x"00001780",
  1508 => x"00001788",
  1509 => x"00001788",
  1510 => x"00001790",
  1511 => x"00001790",
  1512 => x"00001798",
  1513 => x"00001798",
  1514 => x"000017a0",
  1515 => x"000017a0",
  1516 => x"000017a8",
  1517 => x"000017a8",
  1518 => x"000017b0",
  1519 => x"000017b0",
  1520 => x"000017b8",
  1521 => x"000017b8",
  1522 => x"000017c0",
  1523 => x"000017c0",
  1524 => x"000017c8",
  1525 => x"000017c8",
  1526 => x"000017d0",
  1527 => x"000017d0",
  1528 => x"000017d8",
  1529 => x"000017d8",
  1530 => x"000017e0",
  1531 => x"000017e0",
  1532 => x"000017e8",
  1533 => x"000017e8",
  1534 => x"000017f0",
  1535 => x"000017f0",
  1536 => x"000017f8",
  1537 => x"000017f8",
  1538 => x"00001800",
  1539 => x"00001800",
  1540 => x"00001808",
  1541 => x"00001808",
  1542 => x"00001810",
  1543 => x"00001810",
  1544 => x"00001818",
  1545 => x"00001818",
  1546 => x"00001820",
  1547 => x"00001820",
  1548 => x"00001828",
  1549 => x"00001828",
  1550 => x"00001830",
  1551 => x"00001830",
  1552 => x"00001838",
  1553 => x"00001838",
  1554 => x"00001840",
  1555 => x"00001840",
  1556 => x"00001848",
  1557 => x"00001848",
  1558 => x"00001850",
  1559 => x"00001850",
  1560 => x"00001858",
  1561 => x"00001858",
  1562 => x"00001860",
  1563 => x"00001860",
  1564 => x"00001868",
  1565 => x"00001868",
  1566 => x"00001870",
  1567 => x"00001870",
  1568 => x"00001878",
  1569 => x"00001878",
  1570 => x"00001880",
  1571 => x"00001880",
  1572 => x"00001888",
  1573 => x"00001888",
  1574 => x"00001890",
  1575 => x"00001890",
  1576 => x"00001898",
  1577 => x"00001898",
  1578 => x"000018a0",
  1579 => x"000018a0",
  1580 => x"000018a8",
  1581 => x"000018a8",
  1582 => x"000018b0",
  1583 => x"000018b0",
  1584 => x"000018b8",
  1585 => x"000018b8",
  1586 => x"000018c0",
  1587 => x"000018c0",
  1588 => x"000018c8",
  1589 => x"000018c8",
  1590 => x"000018d0",
  1591 => x"000018d0",
  1592 => x"000018d8",
  1593 => x"000018d8",
  1594 => x"000018e0",
  1595 => x"000018e0",
  1596 => x"000018e8",
  1597 => x"000018e8",
  1598 => x"000018f0",
  1599 => x"000018f0",
  1600 => x"000018f8",
  1601 => x"000018f8",
  1602 => x"00001900",
  1603 => x"00001900",
  1604 => x"00001908",
  1605 => x"00001908",
  1606 => x"00001910",
  1607 => x"00001910",
  1608 => x"00001918",
  1609 => x"00001918",
  1610 => x"00001920",
  1611 => x"00001920",
  1612 => x"00001928",
  1613 => x"00001928",
  1614 => x"00001930",
  1615 => x"00001930",
  1616 => x"00001938",
  1617 => x"00001938",
  1618 => x"00001940",
  1619 => x"00001940",
  1620 => x"00001948",
  1621 => x"00001948",
  1622 => x"00001950",
  1623 => x"00001950",
  1624 => x"00001958",
  1625 => x"00001958",
  1626 => x"00001960",
  1627 => x"00001960",
  1628 => x"00001968",
  1629 => x"00001968",
  1630 => x"00001970",
  1631 => x"00001970",
  1632 => x"00001978",
  1633 => x"00001978",
  1634 => x"00001980",
  1635 => x"00001980",
  1636 => x"00001988",
  1637 => x"00001988",
  1638 => x"00001990",
  1639 => x"00001990",
  1640 => x"00001998",
  1641 => x"00001998",
  1642 => x"000019a0",
  1643 => x"000019a0",
  1644 => x"000019a8",
  1645 => x"000019a8",
  1646 => x"000019b0",
  1647 => x"000019b0",
  1648 => x"000019b8",
  1649 => x"000019b8",
  1650 => x"000019c0",
  1651 => x"000019c0",
  1652 => x"000019c8",
  1653 => x"000019c8",
  1654 => x"000019d0",
  1655 => x"000019d0",
  1656 => x"000019d8",
  1657 => x"000019d8",
  1658 => x"000019e0",
  1659 => x"000019e0",
  1660 => x"000019e8",
  1661 => x"000019e8",
  1662 => x"000019f0",
  1663 => x"000019f0",
  1664 => x"000019f8",
  1665 => x"000019f8",
  1666 => x"00001a00",
  1667 => x"00001a00",
  1668 => x"00001a08",
  1669 => x"00001a08",
  1670 => x"00001a10",
  1671 => x"00001a10",
  1672 => x"00001a18",
  1673 => x"00001a18",
  1674 => x"00001a20",
  1675 => x"00001a20",
  1676 => x"00001a28",
  1677 => x"00001a28",
  1678 => x"00001a30",
  1679 => x"00001a30",
  1680 => x"00001a38",
  1681 => x"00001a38",
  1682 => x"00001a40",
  1683 => x"00001a40",
  1684 => x"00001a48",
  1685 => x"00001a48",
  1686 => x"00001a50",
  1687 => x"00001a50",
  1688 => x"00001a58",
  1689 => x"00001a58",
  1690 => x"00001a60",
  1691 => x"00001a60",
  1692 => x"00001a68",
  1693 => x"00001a68",
  1694 => x"00001a70",
  1695 => x"00001a70",
  1696 => x"00001a78",
  1697 => x"00001a78",
  1698 => x"00001a80",
  1699 => x"00001a80",
  1700 => x"00001a88",
  1701 => x"00001a88",
  1702 => x"00001a90",
  1703 => x"00001a90",
  1704 => x"00001a98",
  1705 => x"00001a98",
  1706 => x"00001aa0",
  1707 => x"00001aa0",
  1708 => x"00001aa8",
  1709 => x"00001aa8",
  1710 => x"00001ab0",
  1711 => x"00001ab0",
  1712 => x"00001ab8",
  1713 => x"00001ab8",
  1714 => x"00001ac0",
  1715 => x"00001ac0",
  1716 => x"00001ac8",
  1717 => x"00001ac8",
  1718 => x"00001ad0",
  1719 => x"00001ad0",
  1720 => x"00001ad8",
  1721 => x"00001ad8",
  1722 => x"00001ae0",
  1723 => x"00001ae0",
  1724 => x"00001ae8",
  1725 => x"00001ae8",
  1726 => x"00001af0",
  1727 => x"00001af0",
  1728 => x"00001af8",
  1729 => x"00001af8",
  1730 => x"00001b00",
  1731 => x"00001b00",
  1732 => x"00001b08",
  1733 => x"00001b08",
  1734 => x"00001b10",
  1735 => x"00001b10",
  1736 => x"00001b18",
  1737 => x"00001b18",
  1738 => x"00001b20",
  1739 => x"00001b20",
  1740 => x"00001b28",
  1741 => x"00001b28",
  1742 => x"00001b30",
  1743 => x"00001b30",
  1744 => x"00001b38",
  1745 => x"00001b38",
  1746 => x"00001b40",
  1747 => x"00001b40",
  1748 => x"00001b48",
  1749 => x"00001b48",
  1750 => x"00001b50",
  1751 => x"00001b50",
  1752 => x"00001370",
  1753 => x"ffffffff",
  1754 => x"00000000",
  1755 => x"ffffffff",
  1756 => x"00000000",
  1757 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
