
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 14;
constant bytes : integer := 14184;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B0B0B";
    when 16#00001# => romdata <= X"82700B0B";
    when 16#00002# => romdata <= X"80DEE40C";
    when 16#00003# => romdata <= X"3A0B0B80";
    when 16#00004# => romdata <= X"CBDB0400";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"80088408";
    when 16#00009# => romdata <= X"88080B0B";
    when 16#0000A# => romdata <= X"0B91BF2D";
    when 16#0000B# => romdata <= X"880C840C";
    when 16#0000C# => romdata <= X"800C0400";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B0B88";
    when 16#00049# => romdata <= X"C4040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B0B88A7";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B80DE";
    when 16#000A2# => romdata <= X"D0738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B0B";
    when 16#000A5# => romdata <= X"88AA0400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"80088408";
    when 16#000A9# => romdata <= X"88087575";
    when 16#000AA# => romdata <= X"0B0B0BA9";
    when 16#000AB# => romdata <= X"922D5050";
    when 16#000AC# => romdata <= X"80085688";
    when 16#000AD# => romdata <= X"0C840C80";
    when 16#000AE# => romdata <= X"0C510400";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"80088408";
    when 16#000B1# => romdata <= X"88087575";
    when 16#000B2# => romdata <= X"0B0B0BAA";
    when 16#000B3# => romdata <= X"C42D5050";
    when 16#000B4# => romdata <= X"80085688";
    when 16#000B5# => romdata <= X"0C840C80";
    when 16#000B6# => romdata <= X"0C510400";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"80DEE00C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"82813F80";
    when 16#00101# => romdata <= X"C5C23F04";
    when 16#00102# => romdata <= X"10101010";
    when 16#00103# => romdata <= X"10101010";
    when 16#00104# => romdata <= X"10101010";
    when 16#00105# => romdata <= X"10101010";
    when 16#00106# => romdata <= X"10101010";
    when 16#00107# => romdata <= X"10101010";
    when 16#00108# => romdata <= X"10101010";
    when 16#00109# => romdata <= X"10101053";
    when 16#0010A# => romdata <= X"51047381";
    when 16#0010B# => romdata <= X"FF067383";
    when 16#0010C# => romdata <= X"06098105";
    when 16#0010D# => romdata <= X"83051010";
    when 16#0010E# => romdata <= X"102B0772";
    when 16#0010F# => romdata <= X"FC060C51";
    when 16#00110# => romdata <= X"51043C04";
    when 16#00111# => romdata <= X"72728072";
    when 16#00112# => romdata <= X"8106FF05";
    when 16#00113# => romdata <= X"09720605";
    when 16#00114# => romdata <= X"71105272";
    when 16#00115# => romdata <= X"0A100A53";
    when 16#00116# => romdata <= X"72ED3851";
    when 16#00117# => romdata <= X"51535104";
    when 16#00118# => romdata <= X"80DEE008";
    when 16#00119# => romdata <= X"802EA438";
    when 16#0011A# => romdata <= X"80DEE408";
    when 16#0011B# => romdata <= X"822EBD38";
    when 16#0011C# => romdata <= X"8380800B";
    when 16#0011D# => romdata <= X"0B0B80EE";
    when 16#0011E# => romdata <= X"E80C82A0";
    when 16#0011F# => romdata <= X"800B80EE";
    when 16#00120# => romdata <= X"EC0C8290";
    when 16#00121# => romdata <= X"800B80EE";
    when 16#00122# => romdata <= X"F00C04F8";
    when 16#00123# => romdata <= X"808080A4";
    when 16#00124# => romdata <= X"0B0B0B80";
    when 16#00125# => romdata <= X"EEE80CF8";
    when 16#00126# => romdata <= X"80808280";
    when 16#00127# => romdata <= X"0B80EEEC";
    when 16#00128# => romdata <= X"0CF88080";
    when 16#00129# => romdata <= X"84800B80";
    when 16#0012A# => romdata <= X"EEF00C04";
    when 16#0012B# => romdata <= X"80C0A880";
    when 16#0012C# => romdata <= X"8C0B0B0B";
    when 16#0012D# => romdata <= X"80EEE80C";
    when 16#0012E# => romdata <= X"80C0A880";
    when 16#0012F# => romdata <= X"940B80EE";
    when 16#00130# => romdata <= X"EC0C0B0B";
    when 16#00131# => romdata <= X"80CDF40B";
    when 16#00132# => romdata <= X"80EEF00C";
    when 16#00133# => romdata <= X"04FF3D0D";
    when 16#00134# => romdata <= X"80EEF433";
    when 16#00135# => romdata <= X"5170A738";
    when 16#00136# => romdata <= X"80DEEC08";
    when 16#00137# => romdata <= X"70085252";
    when 16#00138# => romdata <= X"70802E94";
    when 16#00139# => romdata <= X"38841280";
    when 16#0013A# => romdata <= X"DEEC0C70";
    when 16#0013B# => romdata <= X"2D80DEEC";
    when 16#0013C# => romdata <= X"08700852";
    when 16#0013D# => romdata <= X"5270EE38";
    when 16#0013E# => romdata <= X"810B80EE";
    when 16#0013F# => romdata <= X"F434833D";
    when 16#00140# => romdata <= X"0D040480";
    when 16#00141# => romdata <= X"3D0D0B0B";
    when 16#00142# => romdata <= X"80EEE408";
    when 16#00143# => romdata <= X"802E8E38";
    when 16#00144# => romdata <= X"0B0B0B0B";
    when 16#00145# => romdata <= X"800B802E";
    when 16#00146# => romdata <= X"09810685";
    when 16#00147# => romdata <= X"38823D0D";
    when 16#00148# => romdata <= X"040B0B80";
    when 16#00149# => romdata <= X"EEE4510B";
    when 16#0014A# => romdata <= X"0B0BF5D4";
    when 16#0014B# => romdata <= X"3F823D0D";
    when 16#0014C# => romdata <= X"0404FD3D";
    when 16#0014D# => romdata <= X"0D80DEF8";
    when 16#0014E# => romdata <= X"08881108";
    when 16#0014F# => romdata <= X"83DE8007";
    when 16#00150# => romdata <= X"88120C84";
    when 16#00151# => romdata <= X"1108FCA1";
    when 16#00152# => romdata <= X"FF068412";
    when 16#00153# => romdata <= X"0C538F51";
    when 16#00154# => romdata <= X"9AE03F80";
    when 16#00155# => romdata <= X"DEF80884";
    when 16#00156# => romdata <= X"1108E1FF";
    when 16#00157# => romdata <= X"0684120C";
    when 16#00158# => romdata <= X"84110886";
    when 16#00159# => romdata <= X"80078412";
    when 16#0015A# => romdata <= X"0C841108";
    when 16#0015B# => romdata <= X"80C08007";
    when 16#0015C# => romdata <= X"84120C53";
    when 16#0015D# => romdata <= X"81519A95";
    when 16#0015E# => romdata <= X"3F80DEF8";
    when 16#0015F# => romdata <= X"08841108";
    when 16#00160# => romdata <= X"FFBFFF06";
    when 16#00161# => romdata <= X"84120C53";
    when 16#00162# => romdata <= X"85519AA6";
    when 16#00163# => romdata <= X"3F80DEF8";
    when 16#00164# => romdata <= X"08841108";
    when 16#00165# => romdata <= X"80C08007";
    when 16#00166# => romdata <= X"84120C53";
    when 16#00167# => romdata <= X"815199ED";
    when 16#00168# => romdata <= X"3F80DEF8";
    when 16#00169# => romdata <= X"08841108";
    when 16#0016A# => romdata <= X"FFBFFF06";
    when 16#0016B# => romdata <= X"84120C53";
    when 16#0016C# => romdata <= X"815199FE";
    when 16#0016D# => romdata <= X"3F80DEF8";
    when 16#0016E# => romdata <= X"08841108";
    when 16#0016F# => romdata <= X"80C08007";
    when 16#00170# => romdata <= X"84120C53";
    when 16#00171# => romdata <= X"815199C5";
    when 16#00172# => romdata <= X"3F80DEF8";
    when 16#00173# => romdata <= X"08841108";
    when 16#00174# => romdata <= X"FFBFFF06";
    when 16#00175# => romdata <= X"84120C53";
    when 16#00176# => romdata <= X"815199D6";
    when 16#00177# => romdata <= X"3F80DEF8";
    when 16#00178# => romdata <= X"08841108";
    when 16#00179# => romdata <= X"E1FF0684";
    when 16#0017A# => romdata <= X"120C5384";
    when 16#0017B# => romdata <= X"800B8414";
    when 16#0017C# => romdata <= X"08707207";
    when 16#0017D# => romdata <= X"84160C53";
    when 16#0017E# => romdata <= X"84140870";
    when 16#0017F# => romdata <= X"80C08007";
    when 16#00180# => romdata <= X"84160C53";
    when 16#00181# => romdata <= X"54815199";
    when 16#00182# => romdata <= X"843F80DE";
    when 16#00183# => romdata <= X"F8088411";
    when 16#00184# => romdata <= X"0870FFBF";
    when 16#00185# => romdata <= X"FF068413";
    when 16#00186# => romdata <= X"0C535385";
    when 16#00187# => romdata <= X"5199933F";
    when 16#00188# => romdata <= X"80DEF808";
    when 16#00189# => romdata <= X"84110870";
    when 16#0018A# => romdata <= X"FEFFFF06";
    when 16#0018B# => romdata <= X"84130C53";
    when 16#0018C# => romdata <= X"84110870";
    when 16#0018D# => romdata <= X"E1FF0684";
    when 16#0018E# => romdata <= X"130C5384";
    when 16#0018F# => romdata <= X"11087076";
    when 16#00190# => romdata <= X"0784130C";
    when 16#00191# => romdata <= X"53841108";
    when 16#00192# => romdata <= X"80C08007";
    when 16#00193# => romdata <= X"84120C53";
    when 16#00194# => romdata <= X"815198B9";
    when 16#00195# => romdata <= X"3F80DEF8";
    when 16#00196# => romdata <= X"08841108";
    when 16#00197# => romdata <= X"FFBFFF06";
    when 16#00198# => romdata <= X"84120C84";
    when 16#00199# => romdata <= X"1108E1FF";
    when 16#0019A# => romdata <= X"0684120C";
    when 16#0019B# => romdata <= X"84110890";
    when 16#0019C# => romdata <= X"80078412";
    when 16#0019D# => romdata <= X"0C841108";
    when 16#0019E# => romdata <= X"80C08007";
    when 16#0019F# => romdata <= X"84120C54";
    when 16#001A0# => romdata <= X"81519889";
    when 16#001A1# => romdata <= X"3F80DEF8";
    when 16#001A2# => romdata <= X"08841108";
    when 16#001A3# => romdata <= X"FFBFFF06";
    when 16#001A4# => romdata <= X"84120C54";
    when 16#001A5# => romdata <= X"AA5197F5";
    when 16#001A6# => romdata <= X"3F80DEF8";
    when 16#001A7# => romdata <= X"08841108";
    when 16#001A8# => romdata <= X"FEFFFF06";
    when 16#001A9# => romdata <= X"84120C84";
    when 16#001AA# => romdata <= X"1108E1FF";
    when 16#001AB# => romdata <= X"0684120C";
    when 16#001AC# => romdata <= X"84110884";
    when 16#001AD# => romdata <= X"120C8411";
    when 16#001AE# => romdata <= X"0880C080";
    when 16#001AF# => romdata <= X"0784120C";
    when 16#001B0# => romdata <= X"54815197";
    when 16#001B1# => romdata <= X"C83F80DE";
    when 16#001B2# => romdata <= X"F8088411";
    when 16#001B3# => romdata <= X"08FFBFFF";
    when 16#001B4# => romdata <= X"0684120C";
    when 16#001B5# => romdata <= X"841108E1";
    when 16#001B6# => romdata <= X"FF068412";
    when 16#001B7# => romdata <= X"0C841108";
    when 16#001B8# => romdata <= X"98800784";
    when 16#001B9# => romdata <= X"120C8411";
    when 16#001BA# => romdata <= X"0880C080";
    when 16#001BB# => romdata <= X"0784120C";
    when 16#001BC# => romdata <= X"54815197";
    when 16#001BD# => romdata <= X"983F80DE";
    when 16#001BE# => romdata <= X"F8088411";
    when 16#001BF# => romdata <= X"08FFBFFF";
    when 16#001C0# => romdata <= X"0684120C";
    when 16#001C1# => romdata <= X"54AA5197";
    when 16#001C2# => romdata <= X"843F80DE";
    when 16#001C3# => romdata <= X"F8088411";
    when 16#001C4# => romdata <= X"08FEFFFF";
    when 16#001C5# => romdata <= X"0684120C";
    when 16#001C6# => romdata <= X"841108E1";
    when 16#001C7# => romdata <= X"FF068412";
    when 16#001C8# => romdata <= X"0C841108";
    when 16#001C9# => romdata <= X"84120C84";
    when 16#001CA# => romdata <= X"110880C0";
    when 16#001CB# => romdata <= X"80078412";
    when 16#001CC# => romdata <= X"0C548151";
    when 16#001CD# => romdata <= X"96D73F80";
    when 16#001CE# => romdata <= X"DEF80884";
    when 16#001CF# => romdata <= X"1108FFBF";
    when 16#001D0# => romdata <= X"FF068412";
    when 16#001D1# => romdata <= X"0C841108";
    when 16#001D2# => romdata <= X"E1FF0684";
    when 16#001D3# => romdata <= X"120C8411";
    when 16#001D4# => romdata <= X"088C8007";
    when 16#001D5# => romdata <= X"84120C84";
    when 16#001D6# => romdata <= X"110880C0";
    when 16#001D7# => romdata <= X"80078412";
    when 16#001D8# => romdata <= X"0C548151";
    when 16#001D9# => romdata <= X"96A73F80";
    when 16#001DA# => romdata <= X"DEF80884";
    when 16#001DB# => romdata <= X"1108FFBF";
    when 16#001DC# => romdata <= X"FF068412";
    when 16#001DD# => romdata <= X"0C54AA51";
    when 16#001DE# => romdata <= X"96933F81";
    when 16#001DF# => romdata <= X"0B80DEF8";
    when 16#001E0# => romdata <= X"08841108";
    when 16#001E1# => romdata <= X"70FEFFFF";
    when 16#001E2# => romdata <= X"0684130C";
    when 16#001E3# => romdata <= X"54841108";
    when 16#001E4# => romdata <= X"70E1FF06";
    when 16#001E5# => romdata <= X"84130C54";
    when 16#001E6# => romdata <= X"84110884";
    when 16#001E7# => romdata <= X"120C8411";
    when 16#001E8# => romdata <= X"087080C0";
    when 16#001E9# => romdata <= X"80078413";
    when 16#001EA# => romdata <= X"0C545470";
    when 16#001EB# => romdata <= X"525495DD";
    when 16#001EC# => romdata <= X"3F80DEF8";
    when 16#001ED# => romdata <= X"08841108";
    when 16#001EE# => romdata <= X"70FFBFFF";
    when 16#001EF# => romdata <= X"0684130C";
    when 16#001F0# => romdata <= X"53841108";
    when 16#001F1# => romdata <= X"70E1FF06";
    when 16#001F2# => romdata <= X"84130C53";
    when 16#001F3# => romdata <= X"84110870";
    when 16#001F4# => romdata <= X"82800784";
    when 16#001F5# => romdata <= X"130C5384";
    when 16#001F6# => romdata <= X"11087080";
    when 16#001F7# => romdata <= X"C0800784";
    when 16#001F8# => romdata <= X"130C5353";
    when 16#001F9# => romdata <= X"735195A5";
    when 16#001FA# => romdata <= X"3F80DEF8";
    when 16#001FB# => romdata <= X"08841108";
    when 16#001FC# => romdata <= X"FFBFFF06";
    when 16#001FD# => romdata <= X"84120C53";
    when 16#001FE# => romdata <= X"AA519591";
    when 16#001FF# => romdata <= X"3F825195";
    when 16#00200# => romdata <= X"B13F853D";
    when 16#00201# => romdata <= X"0D04FB3D";
    when 16#00202# => romdata <= X"0D777033";
    when 16#00203# => romdata <= X"53567180";
    when 16#00204# => romdata <= X"2E818F38";
    when 16#00205# => romdata <= X"71558116";
    when 16#00206# => romdata <= X"80DEF808";
    when 16#00207# => romdata <= X"84110881";
    when 16#00208# => romdata <= X"80800784";
    when 16#00209# => romdata <= X"120C8411";
    when 16#0020A# => romdata <= X"08E1FF06";
    when 16#0020B# => romdata <= X"84120C76";
    when 16#0020C# => romdata <= X"842B9E80";
    when 16#0020D# => romdata <= X"06841208";
    when 16#0020E# => romdata <= X"70720784";
    when 16#0020F# => romdata <= X"140C5584";
    when 16#00210# => romdata <= X"120880C0";
    when 16#00211# => romdata <= X"80078413";
    when 16#00212# => romdata <= X"0C565456";
    when 16#00213# => romdata <= X"815194BD";
    when 16#00214# => romdata <= X"3F80DEF8";
    when 16#00215# => romdata <= X"08841108";
    when 16#00216# => romdata <= X"FFBFFF06";
    when 16#00217# => romdata <= X"84120C84";
    when 16#00218# => romdata <= X"1108E1FF";
    when 16#00219# => romdata <= X"0684120C";
    when 16#0021A# => romdata <= X"75882B9E";
    when 16#0021B# => romdata <= X"80068412";
    when 16#0021C# => romdata <= X"08710784";
    when 16#0021D# => romdata <= X"130C8412";
    when 16#0021E# => romdata <= X"0880C080";
    when 16#0021F# => romdata <= X"0784130C";
    when 16#00220# => romdata <= X"55538151";
    when 16#00221# => romdata <= X"94873F80";
    when 16#00222# => romdata <= X"DEF80884";
    when 16#00223# => romdata <= X"1108FFBF";
    when 16#00224# => romdata <= X"FF068412";
    when 16#00225# => romdata <= X"0C53AE51";
    when 16#00226# => romdata <= X"93F33F75";
    when 16#00227# => romdata <= X"335574FE";
    when 16#00228# => romdata <= X"F538873D";
    when 16#00229# => romdata <= X"0D04FF3D";
    when 16#0022A# => romdata <= X"0D028F05";
    when 16#0022B# => romdata <= X"33705252";
    when 16#0022C# => romdata <= X"959F3F71";
    when 16#0022D# => romdata <= X"51968E3F";
    when 16#0022E# => romdata <= X"71800C83";
    when 16#0022F# => romdata <= X"3D0D04FF";
    when 16#00230# => romdata <= X"3D0D800B";
    when 16#00231# => romdata <= X"80EEFC08";
    when 16#00232# => romdata <= X"52527072";
    when 16#00233# => romdata <= X"2E098106";
    when 16#00234# => romdata <= X"83388152";
    when 16#00235# => romdata <= X"7180EEFC";
    when 16#00236# => romdata <= X"0C80DF80";
    when 16#00237# => romdata <= X"08528180";
    when 16#00238# => romdata <= X"0B8C130C";
    when 16#00239# => romdata <= X"833D0D04";
    when 16#0023A# => romdata <= X"FA3D0D02";
    when 16#0023B# => romdata <= X"A3053356";
    when 16#0023C# => romdata <= X"758D2E80";
    when 16#0023D# => romdata <= X"F3387588";
    when 16#0023E# => romdata <= X"32703077";
    when 16#0023F# => romdata <= X"80FF3270";
    when 16#00240# => romdata <= X"30728025";
    when 16#00241# => romdata <= X"71802507";
    when 16#00242# => romdata <= X"54515658";
    when 16#00243# => romdata <= X"55749438";
    when 16#00244# => romdata <= X"9F76278B";
    when 16#00245# => romdata <= X"3880F584";
    when 16#00246# => romdata <= X"33559E75";
    when 16#00247# => romdata <= X"27AE3888";
    when 16#00248# => romdata <= X"3D0D0480";
    when 16#00249# => romdata <= X"F5843356";
    when 16#0024A# => romdata <= X"75802EF3";
    when 16#0024B# => romdata <= X"38885190";
    when 16#0024C# => romdata <= X"FD3FA051";
    when 16#0024D# => romdata <= X"90F83F88";
    when 16#0024E# => romdata <= X"5190F33F";
    when 16#0024F# => romdata <= X"80F58433";
    when 16#00250# => romdata <= X"FF055776";
    when 16#00251# => romdata <= X"80F58434";
    when 16#00252# => romdata <= X"883D0D04";
    when 16#00253# => romdata <= X"755190DE";
    when 16#00254# => romdata <= X"3F80F584";
    when 16#00255# => romdata <= X"33811155";
    when 16#00256# => romdata <= X"577380F5";
    when 16#00257# => romdata <= X"84347580";
    when 16#00258# => romdata <= X"F4E01834";
    when 16#00259# => romdata <= X"883D0D04";
    when 16#0025A# => romdata <= X"8A5190C2";
    when 16#0025B# => romdata <= X"3F80F584";
    when 16#0025C# => romdata <= X"33811156";
    when 16#0025D# => romdata <= X"547480F5";
    when 16#0025E# => romdata <= X"8434800B";
    when 16#0025F# => romdata <= X"80F4E015";
    when 16#00260# => romdata <= X"34805680";
    when 16#00261# => romdata <= X"0B80F4E0";
    when 16#00262# => romdata <= X"17335654";
    when 16#00263# => romdata <= X"74A02E83";
    when 16#00264# => romdata <= X"38815474";
    when 16#00265# => romdata <= X"802E9038";
    when 16#00266# => romdata <= X"73802E8B";
    when 16#00267# => romdata <= X"38811670";
    when 16#00268# => romdata <= X"81FF0657";
    when 16#00269# => romdata <= X"57DD3975";
    when 16#0026A# => romdata <= X"802EBF38";
    when 16#0026B# => romdata <= X"800B80F5";
    when 16#0026C# => romdata <= X"80335555";
    when 16#0026D# => romdata <= X"747427AB";
    when 16#0026E# => romdata <= X"38735774";
    when 16#0026F# => romdata <= X"10101075";
    when 16#00270# => romdata <= X"10057654";
    when 16#00271# => romdata <= X"80F4E053";
    when 16#00272# => romdata <= X"80EF8005";
    when 16#00273# => romdata <= X"51A0A63F";
    when 16#00274# => romdata <= X"8008802E";
    when 16#00275# => romdata <= X"A6388115";
    when 16#00276# => romdata <= X"7081FF06";
    when 16#00277# => romdata <= X"56547675";
    when 16#00278# => romdata <= X"26D93880";
    when 16#00279# => romdata <= X"CE84518F";
    when 16#0027A# => romdata <= X"DF3F80CE";
    when 16#0027B# => romdata <= X"80518FD8";
    when 16#0027C# => romdata <= X"3F800B80";
    when 16#0027D# => romdata <= X"F5843488";
    when 16#0027E# => romdata <= X"3D0D0474";
    when 16#0027F# => romdata <= X"101080F4";
    when 16#00280# => romdata <= X"A0057008";
    when 16#00281# => romdata <= X"80F5880C";
    when 16#00282# => romdata <= X"56800B80";
    when 16#00283# => romdata <= X"F58434E7";
    when 16#00284# => romdata <= X"39FD3D0D";
    when 16#00285# => romdata <= X"8A518F96";
    when 16#00286# => romdata <= X"3F800B80";
    when 16#00287# => romdata <= X"F5843480";
    when 16#00288# => romdata <= X"0B80F580";
    when 16#00289# => romdata <= X"34800B80";
    when 16#0028A# => romdata <= X"F5880C80";
    when 16#0028B# => romdata <= X"CE985280";
    when 16#0028C# => romdata <= X"EF80519D";
    when 16#0028D# => romdata <= X"F43F80CE";
    when 16#0028E# => romdata <= X"9C5280F5";
    when 16#0028F# => romdata <= X"803370A0";
    when 16#00290# => romdata <= X"2980F0A0";
    when 16#00291# => romdata <= X"0552549D";
    when 16#00292# => romdata <= X"E03F80F5";
    when 16#00293# => romdata <= X"80337010";
    when 16#00294# => romdata <= X"1080F4A0";
    when 16#00295# => romdata <= X"0599C871";
    when 16#00296# => romdata <= X"0C548105";
    when 16#00297# => romdata <= X"537280F5";
    when 16#00298# => romdata <= X"803480CE";
    when 16#00299# => romdata <= X"A4527281";
    when 16#0029A# => romdata <= X"FF06708A";
    when 16#0029B# => romdata <= X"2980EF80";
    when 16#0029C# => romdata <= X"0552539D";
    when 16#0029D# => romdata <= X"B43F80CE";
    when 16#0029E# => romdata <= X"AC5280F5";
    when 16#0029F# => romdata <= X"803370A0";
    when 16#002A0# => romdata <= X"2980F0A0";
    when 16#002A1# => romdata <= X"0552549D";
    when 16#002A2# => romdata <= X"A03F80F5";
    when 16#002A3# => romdata <= X"80337010";
    when 16#002A4# => romdata <= X"1080F4A0";
    when 16#002A5# => romdata <= X"059D8A71";
    when 16#002A6# => romdata <= X"0C548105";
    when 16#002A7# => romdata <= X"537280F5";
    when 16#002A8# => romdata <= X"803480CF";
    when 16#002A9# => romdata <= X"D8527281";
    when 16#002AA# => romdata <= X"FF06708A";
    when 16#002AB# => romdata <= X"2980EF80";
    when 16#002AC# => romdata <= X"0552539C";
    when 16#002AD# => romdata <= X"F43F80CE";
    when 16#002AE# => romdata <= X"B85280F5";
    when 16#002AF# => romdata <= X"803370A0";
    when 16#002B0# => romdata <= X"2980F0A0";
    when 16#002B1# => romdata <= X"0552549C";
    when 16#002B2# => romdata <= X"E03F80F5";
    when 16#002B3# => romdata <= X"80337010";
    when 16#002B4# => romdata <= X"1080F4A0";
    when 16#002B5# => romdata <= X"0599C871";
    when 16#002B6# => romdata <= X"0C548105";
    when 16#002B7# => romdata <= X"537280F5";
    when 16#002B8# => romdata <= X"803480CE";
    when 16#002B9# => romdata <= X"C8527281";
    when 16#002BA# => romdata <= X"FF06708A";
    when 16#002BB# => romdata <= X"2980EF80";
    when 16#002BC# => romdata <= X"0552539C";
    when 16#002BD# => romdata <= X"B43F80CE";
    when 16#002BE# => romdata <= X"D05280F5";
    when 16#002BF# => romdata <= X"803370A0";
    when 16#002C0# => romdata <= X"2980F0A0";
    when 16#002C1# => romdata <= X"0552549C";
    when 16#002C2# => romdata <= X"A03F80F5";
    when 16#002C3# => romdata <= X"80337010";
    when 16#002C4# => romdata <= X"1080F4A0";
    when 16#002C5# => romdata <= X"059FDA71";
    when 16#002C6# => romdata <= X"0C548105";
    when 16#002C7# => romdata <= X"537280F5";
    when 16#002C8# => romdata <= X"803480CE";
    when 16#002C9# => romdata <= X"E0527281";
    when 16#002CA# => romdata <= X"FF06708A";
    when 16#002CB# => romdata <= X"2980EF80";
    when 16#002CC# => romdata <= X"0552539B";
    when 16#002CD# => romdata <= X"F43F80CE";
    when 16#002CE# => romdata <= X"E45280F5";
    when 16#002CF# => romdata <= X"803370A0";
    when 16#002D0# => romdata <= X"2980F0A0";
    when 16#002D1# => romdata <= X"0552549B";
    when 16#002D2# => romdata <= X"E03F80F5";
    when 16#002D3# => romdata <= X"80337010";
    when 16#002D4# => romdata <= X"1080F4A0";
    when 16#002D5# => romdata <= X"059FE671";
    when 16#002D6# => romdata <= X"0C548105";
    when 16#002D7# => romdata <= X"537280F5";
    when 16#002D8# => romdata <= X"803480CE";
    when 16#002D9# => romdata <= X"F4527281";
    when 16#002DA# => romdata <= X"FF06708A";
    when 16#002DB# => romdata <= X"2980EF80";
    when 16#002DC# => romdata <= X"0552539B";
    when 16#002DD# => romdata <= X"B43F80DC";
    when 16#002DE# => romdata <= X"885280F5";
    when 16#002DF# => romdata <= X"803370A0";
    when 16#002E0# => romdata <= X"2980F0A0";
    when 16#002E1# => romdata <= X"0552549B";
    when 16#002E2# => romdata <= X"A03F80F5";
    when 16#002E3# => romdata <= X"80337010";
    when 16#002E4# => romdata <= X"1080F4A0";
    when 16#002E5# => romdata <= X"0598B271";
    when 16#002E6# => romdata <= X"0C548105";
    when 16#002E7# => romdata <= X"537280F5";
    when 16#002E8# => romdata <= X"803480CD";
    when 16#002E9# => romdata <= X"F8527281";
    when 16#002EA# => romdata <= X"FF06708A";
    when 16#002EB# => romdata <= X"2980EF80";
    when 16#002EC# => romdata <= X"0552539A";
    when 16#002ED# => romdata <= X"F43F80DC";
    when 16#002EE# => romdata <= X"885280F5";
    when 16#002EF# => romdata <= X"803370A0";
    when 16#002F0# => romdata <= X"2980F0A0";
    when 16#002F1# => romdata <= X"0552549A";
    when 16#002F2# => romdata <= X"E03F80F5";
    when 16#002F3# => romdata <= X"80337010";
    when 16#002F4# => romdata <= X"1080F4A0";
    when 16#002F5# => romdata <= X"0598B971";
    when 16#002F6# => romdata <= X"0C548105";
    when 16#002F7# => romdata <= X"537280F5";
    when 16#002F8# => romdata <= X"803480CE";
    when 16#002F9# => romdata <= X"80518BE0";
    when 16#002FA# => romdata <= X"3F810B80";
    when 16#002FB# => romdata <= X"F58C348E";
    when 16#002FC# => romdata <= X"AB3F8008";
    when 16#002FD# => romdata <= X"AE3880F5";
    when 16#002FE# => romdata <= X"88085372";
    when 16#002FF# => romdata <= X"8D3880F5";
    when 16#00300# => romdata <= X"8C335372";
    when 16#00301# => romdata <= X"EA38853D";
    when 16#00302# => romdata <= X"0D04722D";
    when 16#00303# => romdata <= X"800B80F5";
    when 16#00304# => romdata <= X"880C80CE";
    when 16#00305# => romdata <= X"80518BB0";
    when 16#00306# => romdata <= X"3F80F58C";
    when 16#00307# => romdata <= X"335372CF";
    when 16#00308# => romdata <= X"38E4398E";
    when 16#00309# => romdata <= X"8A3F8008";
    when 16#0030A# => romdata <= X"81FF0651";
    when 16#0030B# => romdata <= X"F9BA3FFF";
    when 16#0030C# => romdata <= X"BE39800B";
    when 16#0030D# => romdata <= X"80F58C34";
    when 16#0030E# => romdata <= X"04FC3D0D";
    when 16#0030F# => romdata <= X"8A518AEE";
    when 16#00310# => romdata <= X"3F80CEFC";
    when 16#00311# => romdata <= X"518B813F";
    when 16#00312# => romdata <= X"800B80F5";
    when 16#00313# => romdata <= X"80335354";
    when 16#00314# => romdata <= X"73722780";
    when 16#00315# => romdata <= X"EA387310";
    when 16#00316# => romdata <= X"10107410";
    when 16#00317# => romdata <= X"0580EF80";
    when 16#00318# => romdata <= X"05705253";
    when 16#00319# => romdata <= X"8AE23F73";
    when 16#0031A# => romdata <= X"852B80F0";
    when 16#0031B# => romdata <= X"A0113353";
    when 16#0031C# => romdata <= X"5571802E";
    when 16#0031D# => romdata <= X"B2387251";
    when 16#0031E# => romdata <= X"9A9C3F80";
    when 16#0031F# => romdata <= X"0881FF06";
    when 16#00320# => romdata <= X"52718926";
    when 16#00321# => romdata <= X"9338A051";
    when 16#00322# => romdata <= X"8AA43F81";
    when 16#00323# => romdata <= X"127081FF";
    when 16#00324# => romdata <= X"06535389";
    when 16#00325# => romdata <= X"7227EF38";
    when 16#00326# => romdata <= X"80CF9451";
    when 16#00327# => romdata <= X"8AAA3F80";
    when 16#00328# => romdata <= X"F0A01551";
    when 16#00329# => romdata <= X"8AA23F8A";
    when 16#0032A# => romdata <= X"518A833F";
    when 16#0032B# => romdata <= X"81147081";
    when 16#0032C# => romdata <= X"FF0680F5";
    when 16#0032D# => romdata <= X"80335255";
    when 16#0032E# => romdata <= X"52717426";
    when 16#0032F# => romdata <= X"FF98388A";
    when 16#00330# => romdata <= X"5189EB3F";
    when 16#00331# => romdata <= X"863D0D04";
    when 16#00332# => romdata <= X"F63D0D80";
    when 16#00333# => romdata <= X"0B80F4E0";
    when 16#00334# => romdata <= X"3380F4E0";
    when 16#00335# => romdata <= X"59555673";
    when 16#00336# => romdata <= X"A02E0981";
    when 16#00337# => romdata <= X"06963881";
    when 16#00338# => romdata <= X"167081FF";
    when 16#00339# => romdata <= X"0680F4E0";
    when 16#0033A# => romdata <= X"11703353";
    when 16#0033B# => romdata <= X"59575473";
    when 16#0033C# => romdata <= X"A02EEC38";
    when 16#0033D# => romdata <= X"80588077";
    when 16#0033E# => romdata <= X"33565474";
    when 16#0033F# => romdata <= X"742E8338";
    when 16#00340# => romdata <= X"815474A0";
    when 16#00341# => romdata <= X"2E81CE38";
    when 16#00342# => romdata <= X"7381FB38";
    when 16#00343# => romdata <= X"74A02E81";
    when 16#00344# => romdata <= X"C4388118";
    when 16#00345# => romdata <= X"7081FF06";
    when 16#00346# => romdata <= X"59548178";
    when 16#00347# => romdata <= X"26D83890";
    when 16#00348# => romdata <= X"538C3DFC";
    when 16#00349# => romdata <= X"05527651";
    when 16#0034A# => romdata <= X"9E9A3F80";
    when 16#0034B# => romdata <= X"0859800B";
    when 16#0034C# => romdata <= X"80F4E033";
    when 16#0034D# => romdata <= X"80F4E059";
    when 16#0034E# => romdata <= X"555673A0";
    when 16#0034F# => romdata <= X"2E098106";
    when 16#00350# => romdata <= X"96388116";
    when 16#00351# => romdata <= X"7081FF06";
    when 16#00352# => romdata <= X"80F4E011";
    when 16#00353# => romdata <= X"70335759";
    when 16#00354# => romdata <= X"575873A0";
    when 16#00355# => romdata <= X"2EEC3880";
    when 16#00356# => romdata <= X"58807733";
    when 16#00357# => romdata <= X"56547474";
    when 16#00358# => romdata <= X"2E833881";
    when 16#00359# => romdata <= X"5474A02E";
    when 16#0035A# => romdata <= X"81AC3873";
    when 16#0035B# => romdata <= X"828C3874";
    when 16#0035C# => romdata <= X"A02E81A2";
    when 16#0035D# => romdata <= X"38811870";
    when 16#0035E# => romdata <= X"81FF0659";
    when 16#0035F# => romdata <= X"55827826";
    when 16#00360# => romdata <= X"D8389053";
    when 16#00361# => romdata <= X"8C3DF805";
    when 16#00362# => romdata <= X"5276519D";
    when 16#00363# => romdata <= X"B73F8008";
    when 16#00364# => romdata <= X"57800883";
    when 16#00365# => romdata <= X"38905778";
    when 16#00366# => romdata <= X"FC065580";
    when 16#00367# => romdata <= X"56757727";
    when 16#00368# => romdata <= X"AB387583";
    when 16#00369# => romdata <= X"06597880";
    when 16#0036A# => romdata <= X"2E819C38";
    when 16#0036B# => romdata <= X"80D1D851";
    when 16#0036C# => romdata <= X"88963F74";
    when 16#0036D# => romdata <= X"70840556";
    when 16#0036E# => romdata <= X"0852A051";
    when 16#0036F# => romdata <= X"88AD3FA0";
    when 16#00370# => romdata <= X"5187EB3F";
    when 16#00371# => romdata <= X"81165676";
    when 16#00372# => romdata <= X"7626D738";
    when 16#00373# => romdata <= X"8A5187DE";
    when 16#00374# => romdata <= X"3F8C3D0D";
    when 16#00375# => romdata <= X"04811670";
    when 16#00376# => romdata <= X"81FF0680";
    when 16#00377# => romdata <= X"F4E01170";
    when 16#00378# => romdata <= X"335C5257";
    when 16#00379# => romdata <= X"5778A02E";
    when 16#0037A# => romdata <= X"098106FE";
    when 16#0037B# => romdata <= X"A5388116";
    when 16#0037C# => romdata <= X"7081FF06";
    when 16#0037D# => romdata <= X"80F4E011";
    when 16#0037E# => romdata <= X"70335C52";
    when 16#0037F# => romdata <= X"575778A0";
    when 16#00380# => romdata <= X"2ED338FE";
    when 16#00381# => romdata <= X"8D398116";
    when 16#00382# => romdata <= X"7081FF06";
    when 16#00383# => romdata <= X"80F4E011";
    when 16#00384# => romdata <= X"595755FD";
    when 16#00385# => romdata <= X"E1398116";
    when 16#00386# => romdata <= X"7081FF06";
    when 16#00387# => romdata <= X"80F4E011";
    when 16#00388# => romdata <= X"70335752";
    when 16#00389# => romdata <= X"575773A0";
    when 16#0038A# => romdata <= X"2E098106";
    when 16#0038B# => romdata <= X"FEC73881";
    when 16#0038C# => romdata <= X"167081FF";
    when 16#0038D# => romdata <= X"0680F4E0";
    when 16#0038E# => romdata <= X"11703357";
    when 16#0038F# => romdata <= X"52575773";
    when 16#00390# => romdata <= X"A02ED338";
    when 16#00391# => romdata <= X"FEAF3980";
    when 16#00392# => romdata <= X"CF985186";
    when 16#00393# => romdata <= X"FB3F7452";
    when 16#00394# => romdata <= X"A0518797";
    when 16#00395# => romdata <= X"3F80CF9C";
    when 16#00396# => romdata <= X"5186ED3F";
    when 16#00397# => romdata <= X"80D1D851";
    when 16#00398# => romdata <= X"86E63F74";
    when 16#00399# => romdata <= X"70840556";
    when 16#0039A# => romdata <= X"0852A051";
    when 16#0039B# => romdata <= X"86FD3FA0";
    when 16#0039C# => romdata <= X"5186BB3F";
    when 16#0039D# => romdata <= X"811656FE";
    when 16#0039E# => romdata <= X"CE398116";
    when 16#0039F# => romdata <= X"7081FF06";
    when 16#003A0# => romdata <= X"80F4E011";
    when 16#003A1# => romdata <= X"595755FD";
    when 16#003A2# => romdata <= X"D039F63D";
    when 16#003A3# => romdata <= X"0D800B80";
    when 16#003A4# => romdata <= X"F4E03380";
    when 16#003A5# => romdata <= X"F4E05955";
    when 16#003A6# => romdata <= X"5673A02E";
    when 16#003A7# => romdata <= X"09810696";
    when 16#003A8# => romdata <= X"38811670";
    when 16#003A9# => romdata <= X"81FF0680";
    when 16#003AA# => romdata <= X"F4E01170";
    when 16#003AB# => romdata <= X"33535957";
    when 16#003AC# => romdata <= X"5473A02E";
    when 16#003AD# => romdata <= X"EC388058";
    when 16#003AE# => romdata <= X"80773356";
    when 16#003AF# => romdata <= X"5474742E";
    when 16#003B0# => romdata <= X"83388154";
    when 16#003B1# => romdata <= X"74A02E81";
    when 16#003B2# => romdata <= X"8F387381";
    when 16#003B3# => romdata <= X"BC3874A0";
    when 16#003B4# => romdata <= X"2E818538";
    when 16#003B5# => romdata <= X"81187081";
    when 16#003B6# => romdata <= X"FF065954";
    when 16#003B7# => romdata <= X"817826D8";
    when 16#003B8# => romdata <= X"3890538C";
    when 16#003B9# => romdata <= X"3DFC0552";
    when 16#003BA# => romdata <= X"76519AD8";
    when 16#003BB# => romdata <= X"3F800859";
    when 16#003BC# => romdata <= X"800B80F4";
    when 16#003BD# => romdata <= X"E03380F4";
    when 16#003BE# => romdata <= X"E0595556";
    when 16#003BF# => romdata <= X"73A02E09";
    when 16#003C0# => romdata <= X"81069638";
    when 16#003C1# => romdata <= X"81167081";
    when 16#003C2# => romdata <= X"FF0680F4";
    when 16#003C3# => romdata <= X"E0117033";
    when 16#003C4# => romdata <= X"57595758";
    when 16#003C5# => romdata <= X"73A02EEC";
    when 16#003C6# => romdata <= X"38805880";
    when 16#003C7# => romdata <= X"77335654";
    when 16#003C8# => romdata <= X"74742E83";
    when 16#003C9# => romdata <= X"38815474";
    when 16#003CA# => romdata <= X"A02E80ED";
    when 16#003CB# => romdata <= X"3873819A";
    when 16#003CC# => romdata <= X"3874A02E";
    when 16#003CD# => romdata <= X"80E33881";
    when 16#003CE# => romdata <= X"187081FF";
    when 16#003CF# => romdata <= X"06595582";
    when 16#003D0# => romdata <= X"7826D838";
    when 16#003D1# => romdata <= X"90538C3D";
    when 16#003D2# => romdata <= X"F8055276";
    when 16#003D3# => romdata <= X"5199F53F";
    when 16#003D4# => romdata <= X"8008790C";
    when 16#003D5# => romdata <= X"8C3D0D04";
    when 16#003D6# => romdata <= X"81167081";
    when 16#003D7# => romdata <= X"FF0680F4";
    when 16#003D8# => romdata <= X"E0117033";
    when 16#003D9# => romdata <= X"5C525757";
    when 16#003DA# => romdata <= X"78A02E09";
    when 16#003DB# => romdata <= X"8106FEE4";
    when 16#003DC# => romdata <= X"38811670";
    when 16#003DD# => romdata <= X"81FF0680";
    when 16#003DE# => romdata <= X"F4E01170";
    when 16#003DF# => romdata <= X"335C5257";
    when 16#003E0# => romdata <= X"5778A02E";
    when 16#003E1# => romdata <= X"D338FECC";
    when 16#003E2# => romdata <= X"39811670";
    when 16#003E3# => romdata <= X"81FF0680";
    when 16#003E4# => romdata <= X"F4E01159";
    when 16#003E5# => romdata <= X"5755FEA0";
    when 16#003E6# => romdata <= X"39811670";
    when 16#003E7# => romdata <= X"81FF0680";
    when 16#003E8# => romdata <= X"F4E01170";
    when 16#003E9# => romdata <= X"33575257";
    when 16#003EA# => romdata <= X"5773A02E";
    when 16#003EB# => romdata <= X"098106FF";
    when 16#003EC# => romdata <= X"86388116";
    when 16#003ED# => romdata <= X"7081FF06";
    when 16#003EE# => romdata <= X"80F4E011";
    when 16#003EF# => romdata <= X"70335752";
    when 16#003F0# => romdata <= X"575773A0";
    when 16#003F1# => romdata <= X"2ED338FE";
    when 16#003F2# => romdata <= X"EE398116";
    when 16#003F3# => romdata <= X"7081FF06";
    when 16#003F4# => romdata <= X"80F4E011";
    when 16#003F5# => romdata <= X"595755FE";
    when 16#003F6# => romdata <= X"C239803D";
    when 16#003F7# => romdata <= X"0D8C5183";
    when 16#003F8# => romdata <= X"CD3F823D";
    when 16#003F9# => romdata <= X"0D04FC3D";
    when 16#003FA# => romdata <= X"0DF881C0";
    when 16#003FB# => romdata <= X"8E80539F";
    when 16#003FC# => romdata <= X"0B80DEF8";
    when 16#003FD# => romdata <= X"087481FF";
    when 16#003FE# => romdata <= X"0684120C";
    when 16#003FF# => romdata <= X"80EEFC08";
    when 16#00400# => romdata <= X"54565471";
    when 16#00401# => romdata <= X"802E9F38";
    when 16#00402# => romdata <= X"729F2A73";
    when 16#00403# => romdata <= X"10075373";
    when 16#00404# => romdata <= X"802E9F38";
    when 16#00405# => romdata <= X"FF147381";
    when 16#00406# => romdata <= X"FF068417";
    when 16#00407# => romdata <= X"0C80EEFC";
    when 16#00408# => romdata <= X"08535471";
    when 16#00409# => romdata <= X"E338720A";
    when 16#0040A# => romdata <= X"100A739F";
    when 16#0040B# => romdata <= X"2B075373";
    when 16#0040C# => romdata <= X"E338863D";
    when 16#0040D# => romdata <= X"0D04F73D";
    when 16#0040E# => romdata <= X"0D80DEF8";
    when 16#0040F# => romdata <= X"08700881";
    when 16#00410# => romdata <= X"0A0680EE";
    when 16#00411# => romdata <= X"F80C5385";
    when 16#00412# => romdata <= X"8C3F85BA";
    when 16#00413# => romdata <= X"3FA39852";
    when 16#00414# => romdata <= X"80EEF808";
    when 16#00415# => romdata <= X"843891A6";
    when 16#00416# => romdata <= X"527180F5";
    when 16#00417# => romdata <= X"900CE9D2";
    when 16#00418# => romdata <= X"3F86BE3F";
    when 16#00419# => romdata <= X"80DEF008";
    when 16#0041A# => romdata <= X"53FAC98E";
    when 16#0041B# => romdata <= X"868C730C";
    when 16#0041C# => romdata <= X"72087084";
    when 16#0041D# => romdata <= X"2A810651";
    when 16#0041E# => romdata <= X"5473F538";
    when 16#0041F# => romdata <= X"80DEF808";
    when 16#00420# => romdata <= X"88110881";
    when 16#00421# => romdata <= X"FF078812";
    when 16#00422# => romdata <= X"0C7480EE";
    when 16#00423# => romdata <= X"FC0C9411";
    when 16#00424# => romdata <= X"08818007";
    when 16#00425# => romdata <= X"94120C8C";
    when 16#00426# => romdata <= X"11088180";
    when 16#00427# => romdata <= X"078C120C";
    when 16#00428# => romdata <= X"5380DF80";
    when 16#00429# => romdata <= X"08528180";
    when 16#0042A# => romdata <= X"0B80C013";
    when 16#0042B# => romdata <= X"0C80D294";
    when 16#0042C# => romdata <= X"5182953F";
    when 16#0042D# => romdata <= X"8C5181F6";
    when 16#0042E# => romdata <= X"3F80DBB8";
    when 16#0042F# => romdata <= X"5182893F";
    when 16#00430# => romdata <= X"80EEF808";
    when 16#00431# => romdata <= X"802E81A0";
    when 16#00432# => romdata <= X"3880DBC0";
    when 16#00433# => romdata <= X"5181F93F";
    when 16#00434# => romdata <= X"80DBCC51";
    when 16#00435# => romdata <= X"EEB03FF2";
    when 16#00436# => romdata <= X"B83FF881";
    when 16#00437# => romdata <= X"C08E8053";
    when 16#00438# => romdata <= X"9F0B80DE";
    when 16#00439# => romdata <= X"F8085555";
    when 16#0043A# => romdata <= X"80EEF808";
    when 16#0043B# => romdata <= X"802E80D3";
    when 16#0043C# => romdata <= X"387281FF";
    when 16#0043D# => romdata <= X"0684150C";
    when 16#0043E# => romdata <= X"80EEFC08";
    when 16#0043F# => romdata <= X"5271802E";
    when 16#00440# => romdata <= X"9F38729F";
    when 16#00441# => romdata <= X"2A731007";
    when 16#00442# => romdata <= X"5374802E";
    when 16#00443# => romdata <= X"9F38FF15";
    when 16#00444# => romdata <= X"7381FF06";
    when 16#00445# => romdata <= X"84160C80";
    when 16#00446# => romdata <= X"EEFC0853";
    when 16#00447# => romdata <= X"5571E338";
    when 16#00448# => romdata <= X"720A100A";
    when 16#00449# => romdata <= X"739F2B07";
    when 16#0044A# => romdata <= X"5374E338";
    when 16#0044B# => romdata <= X"8AE03F72";
    when 16#0044C# => romdata <= X"0A100A73";
    when 16#0044D# => romdata <= X"9F2B0753";
    when 16#0044E# => romdata <= X"80FD5182";
    when 16#0044F# => romdata <= X"F53F80DE";
    when 16#00450# => romdata <= X"F8085472";
    when 16#00451# => romdata <= X"81FF0684";
    when 16#00452# => romdata <= X"150C80EE";
    when 16#00453# => romdata <= X"FC085473";
    when 16#00454# => romdata <= X"802EDC38";
    when 16#00455# => romdata <= X"729F2A73";
    when 16#00456# => romdata <= X"10075380";
    when 16#00457# => romdata <= X"FD5182D2";
    when 16#00458# => romdata <= X"3F80DEF8";
    when 16#00459# => romdata <= X"0854DC39";
    when 16#0045A# => romdata <= X"80DBD851";
    when 16#0045B# => romdata <= X"80DA3F80";
    when 16#0045C# => romdata <= X"DBE85180";
    when 16#0045D# => romdata <= X"D33F80DB";
    when 16#0045E# => romdata <= X"CC51ED8A";
    when 16#0045F# => romdata <= X"3FF1923F";
    when 16#00460# => romdata <= X"F881C08E";
    when 16#00461# => romdata <= X"80539F0B";
    when 16#00462# => romdata <= X"80DEF808";
    when 16#00463# => romdata <= X"555580EE";
    when 16#00464# => romdata <= X"F808FEDD";
    when 16#00465# => romdata <= X"38FFAC39";
    when 16#00466# => romdata <= X"FF3D0D02";
    when 16#00467# => romdata <= X"8F053380";
    when 16#00468# => romdata <= X"DEF40852";
    when 16#00469# => romdata <= X"710C800B";
    when 16#0046A# => romdata <= X"800C833D";
    when 16#0046B# => romdata <= X"0D04FF3D";
    when 16#0046C# => romdata <= X"0D028F05";
    when 16#0046D# => romdata <= X"335180F5";
    when 16#0046E# => romdata <= X"90085271";
    when 16#0046F# => romdata <= X"2D800881";
    when 16#00470# => romdata <= X"FF06800C";
    when 16#00471# => romdata <= X"833D0D04";
    when 16#00472# => romdata <= X"FE3D0D74";
    when 16#00473# => romdata <= X"70335353";
    when 16#00474# => romdata <= X"71802E93";
    when 16#00475# => romdata <= X"38811372";
    when 16#00476# => romdata <= X"5280F590";
    when 16#00477# => romdata <= X"08535371";
    when 16#00478# => romdata <= X"2D723352";
    when 16#00479# => romdata <= X"71EF3884";
    when 16#0047A# => romdata <= X"3D0D04F4";
    when 16#0047B# => romdata <= X"3D0D7F02";
    when 16#0047C# => romdata <= X"8405BB05";
    when 16#0047D# => romdata <= X"33555788";
    when 16#0047E# => romdata <= X"0B8C3D5A";
    when 16#0047F# => romdata <= X"5A895380";
    when 16#00480# => romdata <= X"DCB05278";
    when 16#00481# => romdata <= X"5189943F";
    when 16#00482# => romdata <= X"737A2E80";
    when 16#00483# => romdata <= X"FA387956";
    when 16#00484# => romdata <= X"73902E80";
    when 16#00485# => romdata <= X"E73802A7";
    when 16#00486# => romdata <= X"0558768F";
    when 16#00487# => romdata <= X"06547389";
    when 16#00488# => romdata <= X"26BF3875";
    when 16#00489# => romdata <= X"18B01555";
    when 16#0048A# => romdata <= X"55737534";
    when 16#0048B# => romdata <= X"76842AFF";
    when 16#0048C# => romdata <= X"177081FF";
    when 16#0048D# => romdata <= X"06585557";
    when 16#0048E# => romdata <= X"75E03879";
    when 16#0048F# => romdata <= X"19557575";
    when 16#00490# => romdata <= X"34787033";
    when 16#00491# => romdata <= X"55557380";
    when 16#00492# => romdata <= X"2E933881";
    when 16#00493# => romdata <= X"15745280";
    when 16#00494# => romdata <= X"F5900857";
    when 16#00495# => romdata <= X"55752D74";
    when 16#00496# => romdata <= X"335473EF";
    when 16#00497# => romdata <= X"388E3D0D";
    when 16#00498# => romdata <= X"047518B7";
    when 16#00499# => romdata <= X"15555573";
    when 16#0049A# => romdata <= X"75347684";
    when 16#0049B# => romdata <= X"2AFF1770";
    when 16#0049C# => romdata <= X"81FF0658";
    when 16#0049D# => romdata <= X"555775FF";
    when 16#0049E# => romdata <= X"A138C039";
    when 16#0049F# => romdata <= X"8470575A";
    when 16#004A0# => romdata <= X"02A70558";
    when 16#004A1# => romdata <= X"FF943982";
    when 16#004A2# => romdata <= X"70575AF4";
    when 16#004A3# => romdata <= X"39FF3D0D";
    when 16#004A4# => romdata <= X"80DF8408";
    when 16#004A5# => romdata <= X"74101075";
    when 16#004A6# => romdata <= X"10059412";
    when 16#004A7# => romdata <= X"0C52850B";
    when 16#004A8# => romdata <= X"98130C98";
    when 16#004A9# => romdata <= X"12087081";
    when 16#004AA# => romdata <= X"06515170";
    when 16#004AB# => romdata <= X"F638833D";
    when 16#004AC# => romdata <= X"0D04FD3D";
    when 16#004AD# => romdata <= X"0D80DF84";
    when 16#004AE# => romdata <= X"0876B0EA";
    when 16#004AF# => romdata <= X"2994120C";
    when 16#004B0# => romdata <= X"54850B98";
    when 16#004B1# => romdata <= X"150C9814";
    when 16#004B2# => romdata <= X"08708106";
    when 16#004B3# => romdata <= X"515372F6";
    when 16#004B4# => romdata <= X"38853D0D";
    when 16#004B5# => romdata <= X"04803D0D";
    when 16#004B6# => romdata <= X"80DF8408";
    when 16#004B7# => romdata <= X"51870B84";
    when 16#004B8# => romdata <= X"120CFF0B";
    when 16#004B9# => romdata <= X"B4120CA7";
    when 16#004BA# => romdata <= X"0BB8120C";
    when 16#004BB# => romdata <= X"87E80BA4";
    when 16#004BC# => romdata <= X"120CA70B";
    when 16#004BD# => romdata <= X"A8120CB0";
    when 16#004BE# => romdata <= X"EA0B9412";
    when 16#004BF# => romdata <= X"0C870B98";
    when 16#004C0# => romdata <= X"120C823D";
    when 16#004C1# => romdata <= X"0D04803D";
    when 16#004C2# => romdata <= X"0D80DF88";
    when 16#004C3# => romdata <= X"0851B60B";
    when 16#004C4# => romdata <= X"8C120C83";
    when 16#004C5# => romdata <= X"0B88120C";
    when 16#004C6# => romdata <= X"823D0D04";
    when 16#004C7# => romdata <= X"803D0D80";
    when 16#004C8# => romdata <= X"DF880884";
    when 16#004C9# => romdata <= X"11088106";
    when 16#004CA# => romdata <= X"800C5182";
    when 16#004CB# => romdata <= X"3D0D04FF";
    when 16#004CC# => romdata <= X"3D0D80DF";
    when 16#004CD# => romdata <= X"88085284";
    when 16#004CE# => romdata <= X"12087081";
    when 16#004CF# => romdata <= X"06515170";
    when 16#004D0# => romdata <= X"802EF438";
    when 16#004D1# => romdata <= X"71087081";
    when 16#004D2# => romdata <= X"FF06800C";
    when 16#004D3# => romdata <= X"51833D0D";
    when 16#004D4# => romdata <= X"04FE3D0D";
    when 16#004D5# => romdata <= X"02930533";
    when 16#004D6# => romdata <= X"53728A2E";
    when 16#004D7# => romdata <= X"9C3880DF";
    when 16#004D8# => romdata <= X"88085284";
    when 16#004D9# => romdata <= X"12087089";
    when 16#004DA# => romdata <= X"2A708106";
    when 16#004DB# => romdata <= X"51515170";
    when 16#004DC# => romdata <= X"F2387272";
    when 16#004DD# => romdata <= X"0C843D0D";
    when 16#004DE# => romdata <= X"0480DF88";
    when 16#004DF# => romdata <= X"08528412";
    when 16#004E0# => romdata <= X"0870892A";
    when 16#004E1# => romdata <= X"70810651";
    when 16#004E2# => romdata <= X"515170F2";
    when 16#004E3# => romdata <= X"388D720C";
    when 16#004E4# => romdata <= X"84120870";
    when 16#004E5# => romdata <= X"892A7081";
    when 16#004E6# => romdata <= X"06515151";
    when 16#004E7# => romdata <= X"70C538D2";
    when 16#004E8# => romdata <= X"39803D0D";
    when 16#004E9# => romdata <= X"80DEFC08";
    when 16#004EA# => romdata <= X"51800B84";
    when 16#004EB# => romdata <= X"120C83FE";
    when 16#004EC# => romdata <= X"800B8812";
    when 16#004ED# => romdata <= X"0C800B80";
    when 16#004EE# => romdata <= X"F5943480";
    when 16#004EF# => romdata <= X"0B80F598";
    when 16#004F0# => romdata <= X"34823D0D";
    when 16#004F1# => romdata <= X"04FA3D0D";
    when 16#004F2# => romdata <= X"02A30533";
    when 16#004F3# => romdata <= X"80DEFC08";
    when 16#004F4# => romdata <= X"80F59433";
    when 16#004F5# => romdata <= X"7081FF06";
    when 16#004F6# => romdata <= X"70101011";
    when 16#004F7# => romdata <= X"80F59833";
    when 16#004F8# => romdata <= X"7081FF06";
    when 16#004F9# => romdata <= X"72902911";
    when 16#004FA# => romdata <= X"70882B78";
    when 16#004FB# => romdata <= X"07770C53";
    when 16#004FC# => romdata <= X"5B5B5555";
    when 16#004FD# => romdata <= X"59545473";
    when 16#004FE# => romdata <= X"8A2E9838";
    when 16#004FF# => romdata <= X"7480CF2E";
    when 16#00500# => romdata <= X"9238738C";
    when 16#00501# => romdata <= X"2EA43881";
    when 16#00502# => romdata <= X"16537280";
    when 16#00503# => romdata <= X"F5983488";
    when 16#00504# => romdata <= X"3D0D0471";
    when 16#00505# => romdata <= X"A326A338";
    when 16#00506# => romdata <= X"81175271";
    when 16#00507# => romdata <= X"80F59434";
    when 16#00508# => romdata <= X"800B80F5";
    when 16#00509# => romdata <= X"9834883D";
    when 16#0050A# => romdata <= X"0D048052";
    when 16#0050B# => romdata <= X"71882B73";
    when 16#0050C# => romdata <= X"0C811252";
    when 16#0050D# => romdata <= X"97907226";
    when 16#0050E# => romdata <= X"F338800B";
    when 16#0050F# => romdata <= X"80F59434";
    when 16#00510# => romdata <= X"800B80F5";
    when 16#00511# => romdata <= X"9834DF39";
    when 16#00512# => romdata <= X"8C08028C";
    when 16#00513# => romdata <= X"0CFD3D0D";
    when 16#00514# => romdata <= X"80538C08";
    when 16#00515# => romdata <= X"8C050852";
    when 16#00516# => romdata <= X"8C088805";
    when 16#00517# => romdata <= X"085182DE";
    when 16#00518# => romdata <= X"3F800870";
    when 16#00519# => romdata <= X"800C5485";
    when 16#0051A# => romdata <= X"3D0D8C0C";
    when 16#0051B# => romdata <= X"048C0802";
    when 16#0051C# => romdata <= X"8C0CFD3D";
    when 16#0051D# => romdata <= X"0D81538C";
    when 16#0051E# => romdata <= X"088C0508";
    when 16#0051F# => romdata <= X"528C0888";
    when 16#00520# => romdata <= X"05085182";
    when 16#00521# => romdata <= X"B93F8008";
    when 16#00522# => romdata <= X"70800C54";
    when 16#00523# => romdata <= X"853D0D8C";
    when 16#00524# => romdata <= X"0C048C08";
    when 16#00525# => romdata <= X"028C0CF9";
    when 16#00526# => romdata <= X"3D0D800B";
    when 16#00527# => romdata <= X"8C08FC05";
    when 16#00528# => romdata <= X"0C8C0888";
    when 16#00529# => romdata <= X"05088025";
    when 16#0052A# => romdata <= X"AB388C08";
    when 16#0052B# => romdata <= X"88050830";
    when 16#0052C# => romdata <= X"8C088805";
    when 16#0052D# => romdata <= X"0C800B8C";
    when 16#0052E# => romdata <= X"08F4050C";
    when 16#0052F# => romdata <= X"8C08FC05";
    when 16#00530# => romdata <= X"08883881";
    when 16#00531# => romdata <= X"0B8C08F4";
    when 16#00532# => romdata <= X"050C8C08";
    when 16#00533# => romdata <= X"F405088C";
    when 16#00534# => romdata <= X"08FC050C";
    when 16#00535# => romdata <= X"8C088C05";
    when 16#00536# => romdata <= X"088025AB";
    when 16#00537# => romdata <= X"388C088C";
    when 16#00538# => romdata <= X"0508308C";
    when 16#00539# => romdata <= X"088C050C";
    when 16#0053A# => romdata <= X"800B8C08";
    when 16#0053B# => romdata <= X"F0050C8C";
    when 16#0053C# => romdata <= X"08FC0508";
    when 16#0053D# => romdata <= X"8838810B";
    when 16#0053E# => romdata <= X"8C08F005";
    when 16#0053F# => romdata <= X"0C8C08F0";
    when 16#00540# => romdata <= X"05088C08";
    when 16#00541# => romdata <= X"FC050C80";
    when 16#00542# => romdata <= X"538C088C";
    when 16#00543# => romdata <= X"0508528C";
    when 16#00544# => romdata <= X"08880508";
    when 16#00545# => romdata <= X"5181A73F";
    when 16#00546# => romdata <= X"8008708C";
    when 16#00547# => romdata <= X"08F8050C";
    when 16#00548# => romdata <= X"548C08FC";
    when 16#00549# => romdata <= X"0508802E";
    when 16#0054A# => romdata <= X"8C388C08";
    when 16#0054B# => romdata <= X"F8050830";
    when 16#0054C# => romdata <= X"8C08F805";
    when 16#0054D# => romdata <= X"0C8C08F8";
    when 16#0054E# => romdata <= X"05087080";
    when 16#0054F# => romdata <= X"0C54893D";
    when 16#00550# => romdata <= X"0D8C0C04";
    when 16#00551# => romdata <= X"8C08028C";
    when 16#00552# => romdata <= X"0CFB3D0D";
    when 16#00553# => romdata <= X"800B8C08";
    when 16#00554# => romdata <= X"FC050C8C";
    when 16#00555# => romdata <= X"08880508";
    when 16#00556# => romdata <= X"80259338";
    when 16#00557# => romdata <= X"8C088805";
    when 16#00558# => romdata <= X"08308C08";
    when 16#00559# => romdata <= X"88050C81";
    when 16#0055A# => romdata <= X"0B8C08FC";
    when 16#0055B# => romdata <= X"050C8C08";
    when 16#0055C# => romdata <= X"8C050880";
    when 16#0055D# => romdata <= X"258C388C";
    when 16#0055E# => romdata <= X"088C0508";
    when 16#0055F# => romdata <= X"308C088C";
    when 16#00560# => romdata <= X"050C8153";
    when 16#00561# => romdata <= X"8C088C05";
    when 16#00562# => romdata <= X"08528C08";
    when 16#00563# => romdata <= X"88050851";
    when 16#00564# => romdata <= X"AD3F8008";
    when 16#00565# => romdata <= X"708C08F8";
    when 16#00566# => romdata <= X"050C548C";
    when 16#00567# => romdata <= X"08FC0508";
    when 16#00568# => romdata <= X"802E8C38";
    when 16#00569# => romdata <= X"8C08F805";
    when 16#0056A# => romdata <= X"08308C08";
    when 16#0056B# => romdata <= X"F8050C8C";
    when 16#0056C# => romdata <= X"08F80508";
    when 16#0056D# => romdata <= X"70800C54";
    when 16#0056E# => romdata <= X"873D0D8C";
    when 16#0056F# => romdata <= X"0C048C08";
    when 16#00570# => romdata <= X"028C0CFD";
    when 16#00571# => romdata <= X"3D0D810B";
    when 16#00572# => romdata <= X"8C08FC05";
    when 16#00573# => romdata <= X"0C800B8C";
    when 16#00574# => romdata <= X"08F8050C";
    when 16#00575# => romdata <= X"8C088C05";
    when 16#00576# => romdata <= X"088C0888";
    when 16#00577# => romdata <= X"050827AC";
    when 16#00578# => romdata <= X"388C08FC";
    when 16#00579# => romdata <= X"0508802E";
    when 16#0057A# => romdata <= X"A338800B";
    when 16#0057B# => romdata <= X"8C088C05";
    when 16#0057C# => romdata <= X"08249938";
    when 16#0057D# => romdata <= X"8C088C05";
    when 16#0057E# => romdata <= X"08108C08";
    when 16#0057F# => romdata <= X"8C050C8C";
    when 16#00580# => romdata <= X"08FC0508";
    when 16#00581# => romdata <= X"108C08FC";
    when 16#00582# => romdata <= X"050CC939";
    when 16#00583# => romdata <= X"8C08FC05";
    when 16#00584# => romdata <= X"08802E80";
    when 16#00585# => romdata <= X"C9388C08";
    when 16#00586# => romdata <= X"8C05088C";
    when 16#00587# => romdata <= X"08880508";
    when 16#00588# => romdata <= X"26A1388C";
    when 16#00589# => romdata <= X"08880508";
    when 16#0058A# => romdata <= X"8C088C05";
    when 16#0058B# => romdata <= X"08318C08";
    when 16#0058C# => romdata <= X"88050C8C";
    when 16#0058D# => romdata <= X"08F80508";
    when 16#0058E# => romdata <= X"8C08FC05";
    when 16#0058F# => romdata <= X"08078C08";
    when 16#00590# => romdata <= X"F8050C8C";
    when 16#00591# => romdata <= X"08FC0508";
    when 16#00592# => romdata <= X"812A8C08";
    when 16#00593# => romdata <= X"FC050C8C";
    when 16#00594# => romdata <= X"088C0508";
    when 16#00595# => romdata <= X"812A8C08";
    when 16#00596# => romdata <= X"8C050CFF";
    when 16#00597# => romdata <= X"AF398C08";
    when 16#00598# => romdata <= X"90050880";
    when 16#00599# => romdata <= X"2E8F388C";
    when 16#0059A# => romdata <= X"08880508";
    when 16#0059B# => romdata <= X"708C08F4";
    when 16#0059C# => romdata <= X"050C518D";
    when 16#0059D# => romdata <= X"398C08F8";
    when 16#0059E# => romdata <= X"0508708C";
    when 16#0059F# => romdata <= X"08F4050C";
    when 16#005A0# => romdata <= X"518C08F4";
    when 16#005A1# => romdata <= X"0508800C";
    when 16#005A2# => romdata <= X"853D0D8C";
    when 16#005A3# => romdata <= X"0C04803D";
    when 16#005A4# => romdata <= X"0D865184";
    when 16#005A5# => romdata <= X"963F8151";
    when 16#005A6# => romdata <= X"9F873FFC";
    when 16#005A7# => romdata <= X"3D0D7670";
    when 16#005A8# => romdata <= X"797B5555";
    when 16#005A9# => romdata <= X"55558F72";
    when 16#005AA# => romdata <= X"278C3872";
    when 16#005AB# => romdata <= X"75078306";
    when 16#005AC# => romdata <= X"5170802E";
    when 16#005AD# => romdata <= X"A738FF12";
    when 16#005AE# => romdata <= X"5271FF2E";
    when 16#005AF# => romdata <= X"98387270";
    when 16#005B0# => romdata <= X"81055433";
    when 16#005B1# => romdata <= X"74708105";
    when 16#005B2# => romdata <= X"5634FF12";
    when 16#005B3# => romdata <= X"5271FF2E";
    when 16#005B4# => romdata <= X"098106EA";
    when 16#005B5# => romdata <= X"3874800C";
    when 16#005B6# => romdata <= X"863D0D04";
    when 16#005B7# => romdata <= X"74517270";
    when 16#005B8# => romdata <= X"84055408";
    when 16#005B9# => romdata <= X"71708405";
    when 16#005BA# => romdata <= X"530C7270";
    when 16#005BB# => romdata <= X"84055408";
    when 16#005BC# => romdata <= X"71708405";
    when 16#005BD# => romdata <= X"530C7270";
    when 16#005BE# => romdata <= X"84055408";
    when 16#005BF# => romdata <= X"71708405";
    when 16#005C0# => romdata <= X"530C7270";
    when 16#005C1# => romdata <= X"84055408";
    when 16#005C2# => romdata <= X"71708405";
    when 16#005C3# => romdata <= X"530CF012";
    when 16#005C4# => romdata <= X"52718F26";
    when 16#005C5# => romdata <= X"C9388372";
    when 16#005C6# => romdata <= X"27953872";
    when 16#005C7# => romdata <= X"70840554";
    when 16#005C8# => romdata <= X"08717084";
    when 16#005C9# => romdata <= X"05530CFC";
    when 16#005CA# => romdata <= X"12527183";
    when 16#005CB# => romdata <= X"26ED3870";
    when 16#005CC# => romdata <= X"54FF8339";
    when 16#005CD# => romdata <= X"FD3D0D75";
    when 16#005CE# => romdata <= X"5384D813";
    when 16#005CF# => romdata <= X"08802E8A";
    when 16#005D0# => romdata <= X"38805372";
    when 16#005D1# => romdata <= X"800C853D";
    when 16#005D2# => romdata <= X"0D048180";
    when 16#005D3# => romdata <= X"5272518A";
    when 16#005D4# => romdata <= X"883F8008";
    when 16#005D5# => romdata <= X"84D8140C";
    when 16#005D6# => romdata <= X"FF538008";
    when 16#005D7# => romdata <= X"802EE438";
    when 16#005D8# => romdata <= X"8008549F";
    when 16#005D9# => romdata <= X"53807470";
    when 16#005DA# => romdata <= X"8405560C";
    when 16#005DB# => romdata <= X"FF135380";
    when 16#005DC# => romdata <= X"7324CE38";
    when 16#005DD# => romdata <= X"80747084";
    when 16#005DE# => romdata <= X"05560CFF";
    when 16#005DF# => romdata <= X"13537280";
    when 16#005E0# => romdata <= X"25E338FF";
    when 16#005E1# => romdata <= X"BC39FD3D";
    when 16#005E2# => romdata <= X"0D757755";
    when 16#005E3# => romdata <= X"539F7427";
    when 16#005E4# => romdata <= X"8D389673";
    when 16#005E5# => romdata <= X"0CFF5271";
    when 16#005E6# => romdata <= X"800C853D";
    when 16#005E7# => romdata <= X"0D0484D8";
    when 16#005E8# => romdata <= X"13085271";
    when 16#005E9# => romdata <= X"802E9338";
    when 16#005EA# => romdata <= X"73101012";
    when 16#005EB# => romdata <= X"70087972";
    when 16#005EC# => romdata <= X"0C515271";
    when 16#005ED# => romdata <= X"800C853D";
    when 16#005EE# => romdata <= X"0D047251";
    when 16#005EF# => romdata <= X"FEF63FFF";
    when 16#005F0# => romdata <= X"528008D3";
    when 16#005F1# => romdata <= X"3884D813";
    when 16#005F2# => romdata <= X"08741010";
    when 16#005F3# => romdata <= X"1170087A";
    when 16#005F4# => romdata <= X"720C5151";
    when 16#005F5# => romdata <= X"52DD39F9";
    when 16#005F6# => romdata <= X"3D0D797B";
    when 16#005F7# => romdata <= X"5856769F";
    when 16#005F8# => romdata <= X"2680E838";
    when 16#005F9# => romdata <= X"84D81608";
    when 16#005FA# => romdata <= X"5473802E";
    when 16#005FB# => romdata <= X"AA387610";
    when 16#005FC# => romdata <= X"10147008";
    when 16#005FD# => romdata <= X"55557380";
    when 16#005FE# => romdata <= X"2EBA3880";
    when 16#005FF# => romdata <= X"5873812E";
    when 16#00600# => romdata <= X"8F3873FF";
    when 16#00601# => romdata <= X"2EA33880";
    when 16#00602# => romdata <= X"750C7651";
    when 16#00603# => romdata <= X"732D8058";
    when 16#00604# => romdata <= X"77800C89";
    when 16#00605# => romdata <= X"3D0D0475";
    when 16#00606# => romdata <= X"51FE993F";
    when 16#00607# => romdata <= X"FF588008";
    when 16#00608# => romdata <= X"EF3884D8";
    when 16#00609# => romdata <= X"160854C6";
    when 16#0060A# => romdata <= X"3996760C";
    when 16#0060B# => romdata <= X"810B800C";
    when 16#0060C# => romdata <= X"893D0D04";
    when 16#0060D# => romdata <= X"755181ED";
    when 16#0060E# => romdata <= X"3F765380";
    when 16#0060F# => romdata <= X"08527551";
    when 16#00610# => romdata <= X"81AD3F80";
    when 16#00611# => romdata <= X"08800C89";
    when 16#00612# => romdata <= X"3D0D0496";
    when 16#00613# => romdata <= X"760CFF0B";
    when 16#00614# => romdata <= X"800C893D";
    when 16#00615# => romdata <= X"0D04FC3D";
    when 16#00616# => romdata <= X"0D767856";
    when 16#00617# => romdata <= X"53FF5474";
    when 16#00618# => romdata <= X"9F26B138";
    when 16#00619# => romdata <= X"84D81308";
    when 16#0061A# => romdata <= X"5271802E";
    when 16#0061B# => romdata <= X"AE387410";
    when 16#0061C# => romdata <= X"10127008";
    when 16#0061D# => romdata <= X"53538154";
    when 16#0061E# => romdata <= X"71802E98";
    when 16#0061F# => romdata <= X"38825471";
    when 16#00620# => romdata <= X"FF2E9138";
    when 16#00621# => romdata <= X"83547181";
    when 16#00622# => romdata <= X"2E8A3880";
    when 16#00623# => romdata <= X"730C7451";
    when 16#00624# => romdata <= X"712D8054";
    when 16#00625# => romdata <= X"73800C86";
    when 16#00626# => romdata <= X"3D0D0472";
    when 16#00627# => romdata <= X"51FD953F";
    when 16#00628# => romdata <= X"8008F138";
    when 16#00629# => romdata <= X"84D81308";
    when 16#0062A# => romdata <= X"52C439FF";
    when 16#0062B# => romdata <= X"3D0D7352";
    when 16#0062C# => romdata <= X"80DF8C08";
    when 16#0062D# => romdata <= X"51FEA03F";
    when 16#0062E# => romdata <= X"833D0D04";
    when 16#0062F# => romdata <= X"FE3D0D75";
    when 16#00630# => romdata <= X"53745280";
    when 16#00631# => romdata <= X"DF8C0851";
    when 16#00632# => romdata <= X"FDBC3F84";
    when 16#00633# => romdata <= X"3D0D0480";
    when 16#00634# => romdata <= X"3D0D80DF";
    when 16#00635# => romdata <= X"8C0851FC";
    when 16#00636# => romdata <= X"DB3F823D";
    when 16#00637# => romdata <= X"0D04FF3D";
    when 16#00638# => romdata <= X"0D735280";
    when 16#00639# => romdata <= X"DF8C0851";
    when 16#0063A# => romdata <= X"FEEC3F83";
    when 16#0063B# => romdata <= X"3D0D04FC";
    when 16#0063C# => romdata <= X"3D0D800B";
    when 16#0063D# => romdata <= X"80F5A40C";
    when 16#0063E# => romdata <= X"78527751";
    when 16#0063F# => romdata <= X"99973F80";
    when 16#00640# => romdata <= X"08548008";
    when 16#00641# => romdata <= X"FF2E8838";
    when 16#00642# => romdata <= X"73800C86";
    when 16#00643# => romdata <= X"3D0D0480";
    when 16#00644# => romdata <= X"F5A40855";
    when 16#00645# => romdata <= X"74802EF0";
    when 16#00646# => romdata <= X"38767571";
    when 16#00647# => romdata <= X"0C537380";
    when 16#00648# => romdata <= X"0C863D0D";
    when 16#00649# => romdata <= X"0498E93F";
    when 16#0064A# => romdata <= X"04FC3D0D";
    when 16#0064B# => romdata <= X"76707970";
    when 16#0064C# => romdata <= X"73078306";
    when 16#0064D# => romdata <= X"54545455";
    when 16#0064E# => romdata <= X"7080C338";
    when 16#0064F# => romdata <= X"71700870";
    when 16#00650# => romdata <= X"0970F7FB";
    when 16#00651# => romdata <= X"FDFF1306";
    when 16#00652# => romdata <= X"70F88482";
    when 16#00653# => romdata <= X"81800651";
    when 16#00654# => romdata <= X"51535354";
    when 16#00655# => romdata <= X"70A63884";
    when 16#00656# => romdata <= X"14727470";
    when 16#00657# => romdata <= X"8405560C";
    when 16#00658# => romdata <= X"70087009";
    when 16#00659# => romdata <= X"70F7FBFD";
    when 16#0065A# => romdata <= X"FF130670";
    when 16#0065B# => romdata <= X"F8848281";
    when 16#0065C# => romdata <= X"80065151";
    when 16#0065D# => romdata <= X"53535470";
    when 16#0065E# => romdata <= X"802EDC38";
    when 16#0065F# => romdata <= X"73527170";
    when 16#00660# => romdata <= X"81055333";
    when 16#00661# => romdata <= X"51707370";
    when 16#00662# => romdata <= X"81055534";
    when 16#00663# => romdata <= X"70F03874";
    when 16#00664# => romdata <= X"800C863D";
    when 16#00665# => romdata <= X"0D04FD3D";
    when 16#00666# => romdata <= X"0D757071";
    when 16#00667# => romdata <= X"83065355";
    when 16#00668# => romdata <= X"5270B838";
    when 16#00669# => romdata <= X"71700870";
    when 16#0066A# => romdata <= X"09F7FBFD";
    when 16#0066B# => romdata <= X"FF120670";
    when 16#0066C# => romdata <= X"F8848281";
    when 16#0066D# => romdata <= X"80065151";
    when 16#0066E# => romdata <= X"5253709D";
    when 16#0066F# => romdata <= X"38841370";
    when 16#00670# => romdata <= X"087009F7";
    when 16#00671# => romdata <= X"FBFDFF12";
    when 16#00672# => romdata <= X"0670F884";
    when 16#00673# => romdata <= X"82818006";
    when 16#00674# => romdata <= X"51515253";
    when 16#00675# => romdata <= X"70802EE5";
    when 16#00676# => romdata <= X"38725271";
    when 16#00677# => romdata <= X"33517080";
    when 16#00678# => romdata <= X"2E8A3881";
    when 16#00679# => romdata <= X"12703352";
    when 16#0067A# => romdata <= X"5270F838";
    when 16#0067B# => romdata <= X"71743180";
    when 16#0067C# => romdata <= X"0C853D0D";
    when 16#0067D# => romdata <= X"04FA3D0D";
    when 16#0067E# => romdata <= X"787A7C70";
    when 16#0067F# => romdata <= X"54555552";
    when 16#00680# => romdata <= X"72802E80";
    when 16#00681# => romdata <= X"D9387174";
    when 16#00682# => romdata <= X"07830651";
    when 16#00683# => romdata <= X"70802E80";
    when 16#00684# => romdata <= X"D438FF13";
    when 16#00685# => romdata <= X"5372FF2E";
    when 16#00686# => romdata <= X"B1387133";
    when 16#00687# => romdata <= X"74335651";
    when 16#00688# => romdata <= X"74712E09";
    when 16#00689# => romdata <= X"8106A938";
    when 16#0068A# => romdata <= X"72802E81";
    when 16#0068B# => romdata <= X"87387081";
    when 16#0068C# => romdata <= X"FF065170";
    when 16#0068D# => romdata <= X"802E80FC";
    when 16#0068E# => romdata <= X"38811281";
    when 16#0068F# => romdata <= X"15FF1555";
    when 16#00690# => romdata <= X"555272FF";
    when 16#00691# => romdata <= X"2E098106";
    when 16#00692# => romdata <= X"D1387133";
    when 16#00693# => romdata <= X"74335651";
    when 16#00694# => romdata <= X"7081FF06";
    when 16#00695# => romdata <= X"7581FF06";
    when 16#00696# => romdata <= X"71713151";
    when 16#00697# => romdata <= X"52527080";
    when 16#00698# => romdata <= X"0C883D0D";
    when 16#00699# => romdata <= X"04717457";
    when 16#0069A# => romdata <= X"55837327";
    when 16#0069B# => romdata <= X"88387108";
    when 16#0069C# => romdata <= X"74082E88";
    when 16#0069D# => romdata <= X"38747655";
    when 16#0069E# => romdata <= X"52FF9739";
    when 16#0069F# => romdata <= X"FC135372";
    when 16#006A0# => romdata <= X"802EB138";
    when 16#006A1# => romdata <= X"74087009";
    when 16#006A2# => romdata <= X"F7FBFDFF";
    when 16#006A3# => romdata <= X"120670F8";
    when 16#006A4# => romdata <= X"84828180";
    when 16#006A5# => romdata <= X"06515151";
    when 16#006A6# => romdata <= X"709A3884";
    when 16#006A7# => romdata <= X"15841757";
    when 16#006A8# => romdata <= X"55837327";
    when 16#006A9# => romdata <= X"D0387408";
    when 16#006AA# => romdata <= X"76082ED0";
    when 16#006AB# => romdata <= X"38747655";
    when 16#006AC# => romdata <= X"52FEDF39";
    when 16#006AD# => romdata <= X"800B800C";
    when 16#006AE# => romdata <= X"883D0D04";
    when 16#006AF# => romdata <= X"F33D0D60";
    when 16#006B0# => romdata <= X"6264725A";
    when 16#006B1# => romdata <= X"5A5D5D80";
    when 16#006B2# => romdata <= X"5E767081";
    when 16#006B3# => romdata <= X"05583380";
    when 16#006B4# => romdata <= X"DCBD1133";
    when 16#006B5# => romdata <= X"70832A70";
    when 16#006B6# => romdata <= X"81065155";
    when 16#006B7# => romdata <= X"555672E9";
    when 16#006B8# => romdata <= X"3875AD2E";
    when 16#006B9# => romdata <= X"81FF3875";
    when 16#006BA# => romdata <= X"AB2E81FB";
    when 16#006BB# => romdata <= X"38773070";
    when 16#006BC# => romdata <= X"79078025";
    when 16#006BD# => romdata <= X"79903270";
    when 16#006BE# => romdata <= X"30707207";
    when 16#006BF# => romdata <= X"80257307";
    when 16#006C0# => romdata <= X"53575751";
    when 16#006C1# => romdata <= X"5372802E";
    when 16#006C2# => romdata <= X"873875B0";
    when 16#006C3# => romdata <= X"2E81E238";
    when 16#006C4# => romdata <= X"778A3888";
    when 16#006C5# => romdata <= X"5875B02E";
    when 16#006C6# => romdata <= X"83388A58";
    when 16#006C7# => romdata <= X"7752FF51";
    when 16#006C8# => romdata <= X"F2A63F80";
    when 16#006C9# => romdata <= X"0878535A";
    when 16#006CA# => romdata <= X"FF51F2C1";
    when 16#006CB# => romdata <= X"3F80085B";
    when 16#006CC# => romdata <= X"80705A55";
    when 16#006CD# => romdata <= X"80DCBD16";
    when 16#006CE# => romdata <= X"3370822A";
    when 16#006CF# => romdata <= X"70810651";
    when 16#006D0# => romdata <= X"54547280";
    when 16#006D1# => romdata <= X"2E80C138";
    when 16#006D2# => romdata <= X"D0165675";
    when 16#006D3# => romdata <= X"782580D7";
    when 16#006D4# => romdata <= X"38807924";
    when 16#006D5# => romdata <= X"757B2607";
    when 16#006D6# => romdata <= X"53729338";
    when 16#006D7# => romdata <= X"747A2E80";
    when 16#006D8# => romdata <= X"EB387A76";
    when 16#006D9# => romdata <= X"2580ED38";
    when 16#006DA# => romdata <= X"72802E80";
    when 16#006DB# => romdata <= X"E738FF77";
    when 16#006DC# => romdata <= X"70810559";
    when 16#006DD# => romdata <= X"33575980";
    when 16#006DE# => romdata <= X"DCBD1633";
    when 16#006DF# => romdata <= X"70822A70";
    when 16#006E0# => romdata <= X"81065154";
    when 16#006E1# => romdata <= X"5472C138";
    when 16#006E2# => romdata <= X"73830653";
    when 16#006E3# => romdata <= X"72802E97";
    when 16#006E4# => romdata <= X"38738106";
    when 16#006E5# => romdata <= X"C9175553";
    when 16#006E6# => romdata <= X"728538FF";
    when 16#006E7# => romdata <= X"A9165473";
    when 16#006E8# => romdata <= X"56777624";
    when 16#006E9# => romdata <= X"FFAB3880";
    when 16#006EA# => romdata <= X"79248189";
    when 16#006EB# => romdata <= X"387D802E";
    when 16#006EC# => romdata <= X"84387430";
    when 16#006ED# => romdata <= X"557B802E";
    when 16#006EE# => romdata <= X"8C38FF17";
    when 16#006EF# => romdata <= X"53788338";
    when 16#006F0# => romdata <= X"7C53727C";
    when 16#006F1# => romdata <= X"0C74800C";
    when 16#006F2# => romdata <= X"8F3D0D04";
    when 16#006F3# => romdata <= X"8153757B";
    when 16#006F4# => romdata <= X"24FF9538";
    when 16#006F5# => romdata <= X"81757929";
    when 16#006F6# => romdata <= X"17787081";
    when 16#006F7# => romdata <= X"055A3358";
    when 16#006F8# => romdata <= X"5659FF93";
    when 16#006F9# => romdata <= X"39815E76";
    when 16#006FA# => romdata <= X"70810558";
    when 16#006FB# => romdata <= X"3356FDFD";
    when 16#006FC# => romdata <= X"39807733";
    when 16#006FD# => romdata <= X"54547280";
    when 16#006FE# => romdata <= X"F82E80C3";
    when 16#006FF# => romdata <= X"387280D8";
    when 16#00700# => romdata <= X"32703070";
    when 16#00701# => romdata <= X"80257607";
    when 16#00702# => romdata <= X"51515372";
    when 16#00703# => romdata <= X"802EFE80";
    when 16#00704# => romdata <= X"38811733";
    when 16#00705# => romdata <= X"82185856";
    when 16#00706# => romdata <= X"90705358";
    when 16#00707# => romdata <= X"FF51F0A8";
    when 16#00708# => romdata <= X"3F800878";
    when 16#00709# => romdata <= X"535AFF51";
    when 16#0070A# => romdata <= X"F0C33F80";
    when 16#0070B# => romdata <= X"085B8070";
    when 16#0070C# => romdata <= X"5A55FE80";
    when 16#0070D# => romdata <= X"39FF6054";
    when 16#0070E# => romdata <= X"55A2730C";
    when 16#0070F# => romdata <= X"FEF73981";
    when 16#00710# => romdata <= X"54FFBA39";
    when 16#00711# => romdata <= X"FD3D0D77";
    when 16#00712# => romdata <= X"54765375";
    when 16#00713# => romdata <= X"5280DF8C";
    when 16#00714# => romdata <= X"0851FCE8";
    when 16#00715# => romdata <= X"3F853D0D";
    when 16#00716# => romdata <= X"04F33D0D";
    when 16#00717# => romdata <= X"7F618B11";
    when 16#00718# => romdata <= X"70F8065C";
    when 16#00719# => romdata <= X"55555E72";
    when 16#0071A# => romdata <= X"96268338";
    when 16#0071B# => romdata <= X"90598079";
    when 16#0071C# => romdata <= X"24747A26";
    when 16#0071D# => romdata <= X"07538054";
    when 16#0071E# => romdata <= X"72742E09";
    when 16#0071F# => romdata <= X"810680CB";
    when 16#00720# => romdata <= X"387D518B";
    when 16#00721# => romdata <= X"CA3F7883";
    when 16#00722# => romdata <= X"F72680C6";
    when 16#00723# => romdata <= X"3878832A";
    when 16#00724# => romdata <= X"70101010";
    when 16#00725# => romdata <= X"80E6C805";
    when 16#00726# => romdata <= X"8C110859";
    when 16#00727# => romdata <= X"595A7678";
    when 16#00728# => romdata <= X"2E83B038";
    when 16#00729# => romdata <= X"841708FC";
    when 16#0072A# => romdata <= X"06568C17";
    when 16#0072B# => romdata <= X"08881808";
    when 16#0072C# => romdata <= X"718C120C";
    when 16#0072D# => romdata <= X"88120C58";
    when 16#0072E# => romdata <= X"75178411";
    when 16#0072F# => romdata <= X"08810784";
    when 16#00730# => romdata <= X"120C537D";
    when 16#00731# => romdata <= X"518B893F";
    when 16#00732# => romdata <= X"88175473";
    when 16#00733# => romdata <= X"800C8F3D";
    when 16#00734# => romdata <= X"0D047889";
    when 16#00735# => romdata <= X"2A79832A";
    when 16#00736# => romdata <= X"5B537280";
    when 16#00737# => romdata <= X"2EBF3878";
    when 16#00738# => romdata <= X"862AB805";
    when 16#00739# => romdata <= X"5A847327";
    when 16#0073A# => romdata <= X"B43880DB";
    when 16#0073B# => romdata <= X"135A9473";
    when 16#0073C# => romdata <= X"27AB3878";
    when 16#0073D# => romdata <= X"8C2A80EE";
    when 16#0073E# => romdata <= X"055A80D4";
    when 16#0073F# => romdata <= X"73279E38";
    when 16#00740# => romdata <= X"788F2A80";
    when 16#00741# => romdata <= X"F7055A82";
    when 16#00742# => romdata <= X"D4732791";
    when 16#00743# => romdata <= X"3878922A";
    when 16#00744# => romdata <= X"80FC055A";
    when 16#00745# => romdata <= X"8AD47327";
    when 16#00746# => romdata <= X"843880FE";
    when 16#00747# => romdata <= X"5A791010";
    when 16#00748# => romdata <= X"1080E6C8";
    when 16#00749# => romdata <= X"058C1108";
    when 16#0074A# => romdata <= X"58557675";
    when 16#0074B# => romdata <= X"2EA33884";
    when 16#0074C# => romdata <= X"1708FC06";
    when 16#0074D# => romdata <= X"707A3155";
    when 16#0074E# => romdata <= X"56738F24";
    when 16#0074F# => romdata <= X"88D53873";
    when 16#00750# => romdata <= X"8025FEE6";
    when 16#00751# => romdata <= X"388C1708";
    when 16#00752# => romdata <= X"5776752E";
    when 16#00753# => romdata <= X"098106DF";
    when 16#00754# => romdata <= X"38811A5A";
    when 16#00755# => romdata <= X"80E6D808";
    when 16#00756# => romdata <= X"577680E6";
    when 16#00757# => romdata <= X"D02E82C0";
    when 16#00758# => romdata <= X"38841708";
    when 16#00759# => romdata <= X"FC06707A";
    when 16#0075A# => romdata <= X"31555673";
    when 16#0075B# => romdata <= X"8F2481F9";
    when 16#0075C# => romdata <= X"3880E6D0";
    when 16#0075D# => romdata <= X"0B80E6DC";
    when 16#0075E# => romdata <= X"0C80E6D0";
    when 16#0075F# => romdata <= X"0B80E6D8";
    when 16#00760# => romdata <= X"0C738025";
    when 16#00761# => romdata <= X"FEB23883";
    when 16#00762# => romdata <= X"FF762783";
    when 16#00763# => romdata <= X"DF387589";
    when 16#00764# => romdata <= X"2A76832A";
    when 16#00765# => romdata <= X"55537280";
    when 16#00766# => romdata <= X"2EBF3875";
    when 16#00767# => romdata <= X"862AB805";
    when 16#00768# => romdata <= X"54847327";
    when 16#00769# => romdata <= X"B43880DB";
    when 16#0076A# => romdata <= X"13549473";
    when 16#0076B# => romdata <= X"27AB3875";
    when 16#0076C# => romdata <= X"8C2A80EE";
    when 16#0076D# => romdata <= X"055480D4";
    when 16#0076E# => romdata <= X"73279E38";
    when 16#0076F# => romdata <= X"758F2A80";
    when 16#00770# => romdata <= X"F7055482";
    when 16#00771# => romdata <= X"D4732791";
    when 16#00772# => romdata <= X"3875922A";
    when 16#00773# => romdata <= X"80FC0554";
    when 16#00774# => romdata <= X"8AD47327";
    when 16#00775# => romdata <= X"843880FE";
    when 16#00776# => romdata <= X"54731010";
    when 16#00777# => romdata <= X"1080E6C8";
    when 16#00778# => romdata <= X"05881108";
    when 16#00779# => romdata <= X"56587478";
    when 16#0077A# => romdata <= X"2E86CF38";
    when 16#0077B# => romdata <= X"841508FC";
    when 16#0077C# => romdata <= X"06537573";
    when 16#0077D# => romdata <= X"278D3888";
    when 16#0077E# => romdata <= X"15085574";
    when 16#0077F# => romdata <= X"782E0981";
    when 16#00780# => romdata <= X"06EA388C";
    when 16#00781# => romdata <= X"150880E6";
    when 16#00782# => romdata <= X"C80B8405";
    when 16#00783# => romdata <= X"08718C1A";
    when 16#00784# => romdata <= X"0C76881A";
    when 16#00785# => romdata <= X"0C788813";
    when 16#00786# => romdata <= X"0C788C18";
    when 16#00787# => romdata <= X"0C5D5879";
    when 16#00788# => romdata <= X"53807A24";
    when 16#00789# => romdata <= X"83E63872";
    when 16#0078A# => romdata <= X"822C8171";
    when 16#0078B# => romdata <= X"2B5C537A";
    when 16#0078C# => romdata <= X"7C268198";
    when 16#0078D# => romdata <= X"387B7B06";
    when 16#0078E# => romdata <= X"537282F1";
    when 16#0078F# => romdata <= X"3879FC06";
    when 16#00790# => romdata <= X"84055A7A";
    when 16#00791# => romdata <= X"10707D06";
    when 16#00792# => romdata <= X"545B7282";
    when 16#00793# => romdata <= X"E038841A";
    when 16#00794# => romdata <= X"5AF13988";
    when 16#00795# => romdata <= X"178C1108";
    when 16#00796# => romdata <= X"58587678";
    when 16#00797# => romdata <= X"2E098106";
    when 16#00798# => romdata <= X"FCC23882";
    when 16#00799# => romdata <= X"1A5AFDEC";
    when 16#0079A# => romdata <= X"39781779";
    when 16#0079B# => romdata <= X"81078419";
    when 16#0079C# => romdata <= X"0C7080E6";
    when 16#0079D# => romdata <= X"DC0C7080";
    when 16#0079E# => romdata <= X"E6D80C80";
    when 16#0079F# => romdata <= X"E6D00B8C";
    when 16#007A0# => romdata <= X"120C8C11";
    when 16#007A1# => romdata <= X"0888120C";
    when 16#007A2# => romdata <= X"74810784";
    when 16#007A3# => romdata <= X"120C7411";
    when 16#007A4# => romdata <= X"75710C51";
    when 16#007A5# => romdata <= X"537D5187";
    when 16#007A6# => romdata <= X"B73F8817";
    when 16#007A7# => romdata <= X"54FCAC39";
    when 16#007A8# => romdata <= X"80E6C80B";
    when 16#007A9# => romdata <= X"8405087A";
    when 16#007AA# => romdata <= X"545C7980";
    when 16#007AB# => romdata <= X"25FEF838";
    when 16#007AC# => romdata <= X"82DA397A";
    when 16#007AD# => romdata <= X"097C0670";
    when 16#007AE# => romdata <= X"80E6C80B";
    when 16#007AF# => romdata <= X"84050C5C";
    when 16#007B0# => romdata <= X"7A105B7A";
    when 16#007B1# => romdata <= X"7C268538";
    when 16#007B2# => romdata <= X"7A85B838";
    when 16#007B3# => romdata <= X"80E6C80B";
    when 16#007B4# => romdata <= X"88050870";
    when 16#007B5# => romdata <= X"841208FC";
    when 16#007B6# => romdata <= X"06707C31";
    when 16#007B7# => romdata <= X"7C72268F";
    when 16#007B8# => romdata <= X"72250757";
    when 16#007B9# => romdata <= X"575C5D55";
    when 16#007BA# => romdata <= X"72802E80";
    when 16#007BB# => romdata <= X"DB38797A";
    when 16#007BC# => romdata <= X"1680E6C0";
    when 16#007BD# => romdata <= X"081B9011";
    when 16#007BE# => romdata <= X"5A55575B";
    when 16#007BF# => romdata <= X"80E6BC08";
    when 16#007C0# => romdata <= X"FF2E8838";
    when 16#007C1# => romdata <= X"A08F13E0";
    when 16#007C2# => romdata <= X"80065776";
    when 16#007C3# => romdata <= X"527D5186";
    when 16#007C4# => romdata <= X"C03F8008";
    when 16#007C5# => romdata <= X"548008FF";
    when 16#007C6# => romdata <= X"2E903880";
    when 16#007C7# => romdata <= X"08762782";
    when 16#007C8# => romdata <= X"99387480";
    when 16#007C9# => romdata <= X"E6C82E82";
    when 16#007CA# => romdata <= X"913880E6";
    when 16#007CB# => romdata <= X"C80B8805";
    when 16#007CC# => romdata <= X"08558415";
    when 16#007CD# => romdata <= X"08FC0670";
    when 16#007CE# => romdata <= X"7A317A72";
    when 16#007CF# => romdata <= X"268F7225";
    when 16#007D0# => romdata <= X"07525553";
    when 16#007D1# => romdata <= X"7283E638";
    when 16#007D2# => romdata <= X"74798107";
    when 16#007D3# => romdata <= X"84170C79";
    when 16#007D4# => romdata <= X"167080E6";
    when 16#007D5# => romdata <= X"C80B8805";
    when 16#007D6# => romdata <= X"0C758107";
    when 16#007D7# => romdata <= X"84120C54";
    when 16#007D8# => romdata <= X"7E525785";
    when 16#007D9# => romdata <= X"EB3F8817";
    when 16#007DA# => romdata <= X"54FAE039";
    when 16#007DB# => romdata <= X"75832A70";
    when 16#007DC# => romdata <= X"54548074";
    when 16#007DD# => romdata <= X"24819B38";
    when 16#007DE# => romdata <= X"72822C81";
    when 16#007DF# => romdata <= X"712B80E6";
    when 16#007E0# => romdata <= X"CC080770";
    when 16#007E1# => romdata <= X"80E6C80B";
    when 16#007E2# => romdata <= X"84050C75";
    when 16#007E3# => romdata <= X"10101080";
    when 16#007E4# => romdata <= X"E6C80588";
    when 16#007E5# => romdata <= X"1108585A";
    when 16#007E6# => romdata <= X"5D53778C";
    when 16#007E7# => romdata <= X"180C7488";
    when 16#007E8# => romdata <= X"180C7688";
    when 16#007E9# => romdata <= X"190C768C";
    when 16#007EA# => romdata <= X"160CFCF3";
    when 16#007EB# => romdata <= X"39797A10";
    when 16#007EC# => romdata <= X"101080E6";
    when 16#007ED# => romdata <= X"C8057057";
    when 16#007EE# => romdata <= X"595D8C15";
    when 16#007EF# => romdata <= X"08577675";
    when 16#007F0# => romdata <= X"2EA33884";
    when 16#007F1# => romdata <= X"1708FC06";
    when 16#007F2# => romdata <= X"707A3155";
    when 16#007F3# => romdata <= X"56738F24";
    when 16#007F4# => romdata <= X"83CA3873";
    when 16#007F5# => romdata <= X"80258481";
    when 16#007F6# => romdata <= X"388C1708";
    when 16#007F7# => romdata <= X"5776752E";
    when 16#007F8# => romdata <= X"098106DF";
    when 16#007F9# => romdata <= X"38881581";
    when 16#007FA# => romdata <= X"1B708306";
    when 16#007FB# => romdata <= X"555B5572";
    when 16#007FC# => romdata <= X"C9387C83";
    when 16#007FD# => romdata <= X"06537280";
    when 16#007FE# => romdata <= X"2EFDB838";
    when 16#007FF# => romdata <= X"FF1DF819";
    when 16#00800# => romdata <= X"595D8818";
    when 16#00801# => romdata <= X"08782EEA";
    when 16#00802# => romdata <= X"38FDB539";
    when 16#00803# => romdata <= X"831A53FC";
    when 16#00804# => romdata <= X"96398314";
    when 16#00805# => romdata <= X"70822C81";
    when 16#00806# => romdata <= X"712B80E6";
    when 16#00807# => romdata <= X"CC080770";
    when 16#00808# => romdata <= X"80E6C80B";
    when 16#00809# => romdata <= X"84050C76";
    when 16#0080A# => romdata <= X"10101080";
    when 16#0080B# => romdata <= X"E6C80588";
    when 16#0080C# => romdata <= X"1108595B";
    when 16#0080D# => romdata <= X"5E5153FE";
    when 16#0080E# => romdata <= X"E13980E6";
    when 16#0080F# => romdata <= X"8C081758";
    when 16#00810# => romdata <= X"8008762E";
    when 16#00811# => romdata <= X"818D3880";
    when 16#00812# => romdata <= X"E6BC08FF";
    when 16#00813# => romdata <= X"2E83EC38";
    when 16#00814# => romdata <= X"73763118";
    when 16#00815# => romdata <= X"80E68C0C";
    when 16#00816# => romdata <= X"73870670";
    when 16#00817# => romdata <= X"57537280";
    when 16#00818# => romdata <= X"2E883888";
    when 16#00819# => romdata <= X"73317015";
    when 16#0081A# => romdata <= X"55567614";
    when 16#0081B# => romdata <= X"9FFF06A0";
    when 16#0081C# => romdata <= X"80713117";
    when 16#0081D# => romdata <= X"70547F53";
    when 16#0081E# => romdata <= X"575383D5";
    when 16#0081F# => romdata <= X"3F800853";
    when 16#00820# => romdata <= X"8008FF2E";
    when 16#00821# => romdata <= X"81A03880";
    when 16#00822# => romdata <= X"E68C0816";
    when 16#00823# => romdata <= X"7080E68C";
    when 16#00824# => romdata <= X"0C747580";
    when 16#00825# => romdata <= X"E6C80B88";
    when 16#00826# => romdata <= X"050C7476";
    when 16#00827# => romdata <= X"31187081";
    when 16#00828# => romdata <= X"07515556";
    when 16#00829# => romdata <= X"587B80E6";
    when 16#0082A# => romdata <= X"C82E839C";
    when 16#0082B# => romdata <= X"38798F26";
    when 16#0082C# => romdata <= X"82CB3881";
    when 16#0082D# => romdata <= X"0B84150C";
    when 16#0082E# => romdata <= X"841508FC";
    when 16#0082F# => romdata <= X"06707A31";
    when 16#00830# => romdata <= X"7A72268F";
    when 16#00831# => romdata <= X"72250752";
    when 16#00832# => romdata <= X"55537280";
    when 16#00833# => romdata <= X"2EFCF938";
    when 16#00834# => romdata <= X"80DB3980";
    when 16#00835# => romdata <= X"089FFF06";
    when 16#00836# => romdata <= X"5372FEEB";
    when 16#00837# => romdata <= X"387780E6";
    when 16#00838# => romdata <= X"8C0C80E6";
    when 16#00839# => romdata <= X"C80B8805";
    when 16#0083A# => romdata <= X"087B1881";
    when 16#0083B# => romdata <= X"0784120C";
    when 16#0083C# => romdata <= X"5580E6B8";
    when 16#0083D# => romdata <= X"08782786";
    when 16#0083E# => romdata <= X"387780E6";
    when 16#0083F# => romdata <= X"B80C80E6";
    when 16#00840# => romdata <= X"B4087827";
    when 16#00841# => romdata <= X"FCAC3877";
    when 16#00842# => romdata <= X"80E6B40C";
    when 16#00843# => romdata <= X"841508FC";
    when 16#00844# => romdata <= X"06707A31";
    when 16#00845# => romdata <= X"7A72268F";
    when 16#00846# => romdata <= X"72250752";
    when 16#00847# => romdata <= X"55537280";
    when 16#00848# => romdata <= X"2EFCA538";
    when 16#00849# => romdata <= X"88398074";
    when 16#0084A# => romdata <= X"5456FEDB";
    when 16#0084B# => romdata <= X"397D5182";
    when 16#0084C# => romdata <= X"9F3F800B";
    when 16#0084D# => romdata <= X"800C8F3D";
    when 16#0084E# => romdata <= X"0D047353";
    when 16#0084F# => romdata <= X"807424A9";
    when 16#00850# => romdata <= X"3872822C";
    when 16#00851# => romdata <= X"81712B80";
    when 16#00852# => romdata <= X"E6CC0807";
    when 16#00853# => romdata <= X"7080E6C8";
    when 16#00854# => romdata <= X"0B84050C";
    when 16#00855# => romdata <= X"5D53778C";
    when 16#00856# => romdata <= X"180C7488";
    when 16#00857# => romdata <= X"180C7688";
    when 16#00858# => romdata <= X"190C768C";
    when 16#00859# => romdata <= X"160CF9B7";
    when 16#0085A# => romdata <= X"39831470";
    when 16#0085B# => romdata <= X"822C8171";
    when 16#0085C# => romdata <= X"2B80E6CC";
    when 16#0085D# => romdata <= X"08077080";
    when 16#0085E# => romdata <= X"E6C80B84";
    when 16#0085F# => romdata <= X"050C5E51";
    when 16#00860# => romdata <= X"53D4397B";
    when 16#00861# => romdata <= X"7B065372";
    when 16#00862# => romdata <= X"FCA33884";
    when 16#00863# => romdata <= X"1A7B105C";
    when 16#00864# => romdata <= X"5AF139FF";
    when 16#00865# => romdata <= X"1A811151";
    when 16#00866# => romdata <= X"5AF7B939";
    when 16#00867# => romdata <= X"78177981";
    when 16#00868# => romdata <= X"0784190C";
    when 16#00869# => romdata <= X"8C180888";
    when 16#0086A# => romdata <= X"1908718C";
    when 16#0086B# => romdata <= X"120C8812";
    when 16#0086C# => romdata <= X"0C597080";
    when 16#0086D# => romdata <= X"E6DC0C70";
    when 16#0086E# => romdata <= X"80E6D80C";
    when 16#0086F# => romdata <= X"80E6D00B";
    when 16#00870# => romdata <= X"8C120C8C";
    when 16#00871# => romdata <= X"11088812";
    when 16#00872# => romdata <= X"0C748107";
    when 16#00873# => romdata <= X"84120C74";
    when 16#00874# => romdata <= X"1175710C";
    when 16#00875# => romdata <= X"5153F9BD";
    when 16#00876# => romdata <= X"39751784";
    when 16#00877# => romdata <= X"11088107";
    when 16#00878# => romdata <= X"84120C53";
    when 16#00879# => romdata <= X"8C170888";
    when 16#0087A# => romdata <= X"1808718C";
    when 16#0087B# => romdata <= X"120C8812";
    when 16#0087C# => romdata <= X"0C587D51";
    when 16#0087D# => romdata <= X"80DA3F88";
    when 16#0087E# => romdata <= X"1754F5CF";
    when 16#0087F# => romdata <= X"39728415";
    when 16#00880# => romdata <= X"0CF41AF8";
    when 16#00881# => romdata <= X"0670841E";
    when 16#00882# => romdata <= X"08810607";
    when 16#00883# => romdata <= X"841E0C70";
    when 16#00884# => romdata <= X"1D545B85";
    when 16#00885# => romdata <= X"0B84140C";
    when 16#00886# => romdata <= X"850B8814";
    when 16#00887# => romdata <= X"0C8F7B27";
    when 16#00888# => romdata <= X"FDCF3888";
    when 16#00889# => romdata <= X"1C527D51";
    when 16#0088A# => romdata <= X"82903F80";
    when 16#0088B# => romdata <= X"E6C80B88";
    when 16#0088C# => romdata <= X"050880E6";
    when 16#0088D# => romdata <= X"8C085955";
    when 16#0088E# => romdata <= X"FDB73977";
    when 16#0088F# => romdata <= X"80E68C0C";
    when 16#00890# => romdata <= X"7380E6BC";
    when 16#00891# => romdata <= X"0CFC9139";
    when 16#00892# => romdata <= X"7284150C";
    when 16#00893# => romdata <= X"FDA33904";
    when 16#00894# => romdata <= X"04FD3D0D";
    when 16#00895# => romdata <= X"800B80F5";
    when 16#00896# => romdata <= X"A40C7651";
    when 16#00897# => romdata <= X"86CC3F80";
    when 16#00898# => romdata <= X"08538008";
    when 16#00899# => romdata <= X"FF2E8838";
    when 16#0089A# => romdata <= X"72800C85";
    when 16#0089B# => romdata <= X"3D0D0480";
    when 16#0089C# => romdata <= X"F5A40854";
    when 16#0089D# => romdata <= X"73802EF0";
    when 16#0089E# => romdata <= X"38757471";
    when 16#0089F# => romdata <= X"0C527280";
    when 16#008A0# => romdata <= X"0C853D0D";
    when 16#008A1# => romdata <= X"04FB3D0D";
    when 16#008A2# => romdata <= X"77705256";
    when 16#008A3# => romdata <= X"C23F80E6";
    when 16#008A4# => romdata <= X"C80B8805";
    when 16#008A5# => romdata <= X"08841108";
    when 16#008A6# => romdata <= X"FC06707B";
    when 16#008A7# => romdata <= X"319FEF05";
    when 16#008A8# => romdata <= X"E08006E0";
    when 16#008A9# => romdata <= X"80055656";
    when 16#008AA# => romdata <= X"53A08074";
    when 16#008AB# => romdata <= X"24943880";
    when 16#008AC# => romdata <= X"527551FF";
    when 16#008AD# => romdata <= X"9C3F80E6";
    when 16#008AE# => romdata <= X"D0081553";
    when 16#008AF# => romdata <= X"7280082E";
    when 16#008B0# => romdata <= X"8F387551";
    when 16#008B1# => romdata <= X"FF8A3F80";
    when 16#008B2# => romdata <= X"5372800C";
    when 16#008B3# => romdata <= X"873D0D04";
    when 16#008B4# => romdata <= X"73305275";
    when 16#008B5# => romdata <= X"51FEFA3F";
    when 16#008B6# => romdata <= X"8008FF2E";
    when 16#008B7# => romdata <= X"A83880E6";
    when 16#008B8# => romdata <= X"C80B8805";
    when 16#008B9# => romdata <= X"08757531";
    when 16#008BA# => romdata <= X"81078412";
    when 16#008BB# => romdata <= X"0C5380E6";
    when 16#008BC# => romdata <= X"8C087431";
    when 16#008BD# => romdata <= X"80E68C0C";
    when 16#008BE# => romdata <= X"7551FED4";
    when 16#008BF# => romdata <= X"3F810B80";
    when 16#008C0# => romdata <= X"0C873D0D";
    when 16#008C1# => romdata <= X"04805275";
    when 16#008C2# => romdata <= X"51FEC63F";
    when 16#008C3# => romdata <= X"80E6C80B";
    when 16#008C4# => romdata <= X"88050880";
    when 16#008C5# => romdata <= X"08713156";
    when 16#008C6# => romdata <= X"538F7525";
    when 16#008C7# => romdata <= X"FFA43880";
    when 16#008C8# => romdata <= X"0880E6BC";
    when 16#008C9# => romdata <= X"083180E6";
    when 16#008CA# => romdata <= X"8C0C7481";
    when 16#008CB# => romdata <= X"0784140C";
    when 16#008CC# => romdata <= X"7551FE9C";
    when 16#008CD# => romdata <= X"3F8053FF";
    when 16#008CE# => romdata <= X"9039F63D";
    when 16#008CF# => romdata <= X"0D7C7E54";
    when 16#008D0# => romdata <= X"5B72802E";
    when 16#008D1# => romdata <= X"8283387A";
    when 16#008D2# => romdata <= X"51FE843F";
    when 16#008D3# => romdata <= X"F8138411";
    when 16#008D4# => romdata <= X"0870FE06";
    when 16#008D5# => romdata <= X"70138411";
    when 16#008D6# => romdata <= X"08FC065D";
    when 16#008D7# => romdata <= X"58595458";
    when 16#008D8# => romdata <= X"80E6D008";
    when 16#008D9# => romdata <= X"752E82DE";
    when 16#008DA# => romdata <= X"38788416";
    when 16#008DB# => romdata <= X"0C807381";
    when 16#008DC# => romdata <= X"06545A72";
    when 16#008DD# => romdata <= X"7A2E81D5";
    when 16#008DE# => romdata <= X"38781584";
    when 16#008DF# => romdata <= X"11088106";
    when 16#008E0# => romdata <= X"515372A0";
    when 16#008E1# => romdata <= X"38781757";
    when 16#008E2# => romdata <= X"7981E638";
    when 16#008E3# => romdata <= X"88150853";
    when 16#008E4# => romdata <= X"7280E6D0";
    when 16#008E5# => romdata <= X"2E82F938";
    when 16#008E6# => romdata <= X"8C150870";
    when 16#008E7# => romdata <= X"8C150C73";
    when 16#008E8# => romdata <= X"88120C56";
    when 16#008E9# => romdata <= X"76810784";
    when 16#008EA# => romdata <= X"190C7618";
    when 16#008EB# => romdata <= X"77710C53";
    when 16#008EC# => romdata <= X"79819138";
    when 16#008ED# => romdata <= X"83FF7727";
    when 16#008EE# => romdata <= X"81C83876";
    when 16#008EF# => romdata <= X"892A7783";
    when 16#008F0# => romdata <= X"2A565372";
    when 16#008F1# => romdata <= X"802EBF38";
    when 16#008F2# => romdata <= X"76862AB8";
    when 16#008F3# => romdata <= X"05558473";
    when 16#008F4# => romdata <= X"27B43880";
    when 16#008F5# => romdata <= X"DB135594";
    when 16#008F6# => romdata <= X"7327AB38";
    when 16#008F7# => romdata <= X"768C2A80";
    when 16#008F8# => romdata <= X"EE055580";
    when 16#008F9# => romdata <= X"D473279E";
    when 16#008FA# => romdata <= X"38768F2A";
    when 16#008FB# => romdata <= X"80F70555";
    when 16#008FC# => romdata <= X"82D47327";
    when 16#008FD# => romdata <= X"91387692";
    when 16#008FE# => romdata <= X"2A80FC05";
    when 16#008FF# => romdata <= X"558AD473";
    when 16#00900# => romdata <= X"27843880";
    when 16#00901# => romdata <= X"FE557410";
    when 16#00902# => romdata <= X"101080E6";
    when 16#00903# => romdata <= X"C8058811";
    when 16#00904# => romdata <= X"08555673";
    when 16#00905# => romdata <= X"762E82B3";
    when 16#00906# => romdata <= X"38841408";
    when 16#00907# => romdata <= X"FC065376";
    when 16#00908# => romdata <= X"73278D38";
    when 16#00909# => romdata <= X"88140854";
    when 16#0090A# => romdata <= X"73762E09";
    when 16#0090B# => romdata <= X"8106EA38";
    when 16#0090C# => romdata <= X"8C140870";
    when 16#0090D# => romdata <= X"8C1A0C74";
    when 16#0090E# => romdata <= X"881A0C78";
    when 16#0090F# => romdata <= X"88120C56";
    when 16#00910# => romdata <= X"778C150C";
    when 16#00911# => romdata <= X"7A51FC88";
    when 16#00912# => romdata <= X"3F8C3D0D";
    when 16#00913# => romdata <= X"04770878";
    when 16#00914# => romdata <= X"71315977";
    when 16#00915# => romdata <= X"05881908";
    when 16#00916# => romdata <= X"54577280";
    when 16#00917# => romdata <= X"E6D02E80";
    when 16#00918# => romdata <= X"E0388C18";
    when 16#00919# => romdata <= X"08708C15";
    when 16#0091A# => romdata <= X"0C738812";
    when 16#0091B# => romdata <= X"0C56FE89";
    when 16#0091C# => romdata <= X"39881508";
    when 16#0091D# => romdata <= X"8C160870";
    when 16#0091E# => romdata <= X"8C130C57";
    when 16#0091F# => romdata <= X"88170CFE";
    when 16#00920# => romdata <= X"A3397683";
    when 16#00921# => romdata <= X"2A705455";
    when 16#00922# => romdata <= X"80752481";
    when 16#00923# => romdata <= X"98387282";
    when 16#00924# => romdata <= X"2C81712B";
    when 16#00925# => romdata <= X"80E6CC08";
    when 16#00926# => romdata <= X"0780E6C8";
    when 16#00927# => romdata <= X"0B84050C";
    when 16#00928# => romdata <= X"53741010";
    when 16#00929# => romdata <= X"1080E6C8";
    when 16#0092A# => romdata <= X"05881108";
    when 16#0092B# => romdata <= X"5556758C";
    when 16#0092C# => romdata <= X"190C7388";
    when 16#0092D# => romdata <= X"190C7788";
    when 16#0092E# => romdata <= X"170C778C";
    when 16#0092F# => romdata <= X"150CFF84";
    when 16#00930# => romdata <= X"39815AFD";
    when 16#00931# => romdata <= X"B4397817";
    when 16#00932# => romdata <= X"73810654";
    when 16#00933# => romdata <= X"57729838";
    when 16#00934# => romdata <= X"77087871";
    when 16#00935# => romdata <= X"31597705";
    when 16#00936# => romdata <= X"8C190888";
    when 16#00937# => romdata <= X"1A08718C";
    when 16#00938# => romdata <= X"120C8812";
    when 16#00939# => romdata <= X"0C575776";
    when 16#0093A# => romdata <= X"81078419";
    when 16#0093B# => romdata <= X"0C7780E6";
    when 16#0093C# => romdata <= X"C80B8805";
    when 16#0093D# => romdata <= X"0C80E6C4";
    when 16#0093E# => romdata <= X"087726FE";
    when 16#0093F# => romdata <= X"C73880E6";
    when 16#00940# => romdata <= X"C008527A";
    when 16#00941# => romdata <= X"51FAFE3F";
    when 16#00942# => romdata <= X"7A51FAC4";
    when 16#00943# => romdata <= X"3FFEBA39";
    when 16#00944# => romdata <= X"81788C15";
    when 16#00945# => romdata <= X"0C788815";
    when 16#00946# => romdata <= X"0C738C1A";
    when 16#00947# => romdata <= X"0C73881A";
    when 16#00948# => romdata <= X"0C5AFD80";
    when 16#00949# => romdata <= X"39831570";
    when 16#0094A# => romdata <= X"822C8171";
    when 16#0094B# => romdata <= X"2B80E6CC";
    when 16#0094C# => romdata <= X"080780E6";
    when 16#0094D# => romdata <= X"C80B8405";
    when 16#0094E# => romdata <= X"0C515374";
    when 16#0094F# => romdata <= X"10101080";
    when 16#00950# => romdata <= X"E6C80588";
    when 16#00951# => romdata <= X"11085556";
    when 16#00952# => romdata <= X"FEE43974";
    when 16#00953# => romdata <= X"53807524";
    when 16#00954# => romdata <= X"A7387282";
    when 16#00955# => romdata <= X"2C81712B";
    when 16#00956# => romdata <= X"80E6CC08";
    when 16#00957# => romdata <= X"0780E6C8";
    when 16#00958# => romdata <= X"0B84050C";
    when 16#00959# => romdata <= X"53758C19";
    when 16#0095A# => romdata <= X"0C738819";
    when 16#0095B# => romdata <= X"0C778817";
    when 16#0095C# => romdata <= X"0C778C15";
    when 16#0095D# => romdata <= X"0CFDCD39";
    when 16#0095E# => romdata <= X"83157082";
    when 16#0095F# => romdata <= X"2C81712B";
    when 16#00960# => romdata <= X"80E6CC08";
    when 16#00961# => romdata <= X"0780E6C8";
    when 16#00962# => romdata <= X"0B84050C";
    when 16#00963# => romdata <= X"5153D639";
    when 16#00964# => romdata <= X"810B800C";
    when 16#00965# => romdata <= X"04803D0D";
    when 16#00966# => romdata <= X"72812E89";
    when 16#00967# => romdata <= X"38800B80";
    when 16#00968# => romdata <= X"0C823D0D";
    when 16#00969# => romdata <= X"04735180";
    when 16#0096A# => romdata <= X"F83FFE3D";
    when 16#0096B# => romdata <= X"0D80F59C";
    when 16#0096C# => romdata <= X"0851708A";
    when 16#0096D# => romdata <= X"3880F5A8";
    when 16#0096E# => romdata <= X"7080F59C";
    when 16#0096F# => romdata <= X"0C517075";
    when 16#00970# => romdata <= X"125252FF";
    when 16#00971# => romdata <= X"537087FB";
    when 16#00972# => romdata <= X"80802688";
    when 16#00973# => romdata <= X"387080F5";
    when 16#00974# => romdata <= X"9C0C7153";
    when 16#00975# => romdata <= X"72800C84";
    when 16#00976# => romdata <= X"3D0D04FD";
    when 16#00977# => romdata <= X"3D0D800B";
    when 16#00978# => romdata <= X"80DEE408";
    when 16#00979# => romdata <= X"54547281";
    when 16#0097A# => romdata <= X"2E9C3873";
    when 16#0097B# => romdata <= X"80F5A00C";
    when 16#0097C# => romdata <= X"FFBCED3F";
    when 16#0097D# => romdata <= X"FFBC893F";
    when 16#0097E# => romdata <= X"80EED052";
    when 16#0097F# => romdata <= X"8151D4B6";
    when 16#00980# => romdata <= X"3F800851";
    when 16#00981# => romdata <= X"9F3F7280";
    when 16#00982# => romdata <= X"F5A00CFF";
    when 16#00983# => romdata <= X"BCD23FFF";
    when 16#00984# => romdata <= X"BBEE3F80";
    when 16#00985# => romdata <= X"EED05281";
    when 16#00986# => romdata <= X"51D49B3F";
    when 16#00987# => romdata <= X"80085184";
    when 16#00988# => romdata <= X"3F00FF39";
    when 16#00989# => romdata <= X"F73D0D7B";
    when 16#0098A# => romdata <= X"80DF8C08";
    when 16#0098B# => romdata <= X"82C81108";
    when 16#0098C# => romdata <= X"5A545A77";
    when 16#0098D# => romdata <= X"802E80DA";
    when 16#0098E# => romdata <= X"38818818";
    when 16#0098F# => romdata <= X"841908FF";
    when 16#00990# => romdata <= X"0581712B";
    when 16#00991# => romdata <= X"59555980";
    when 16#00992# => romdata <= X"742480EA";
    when 16#00993# => romdata <= X"38807424";
    when 16#00994# => romdata <= X"B5387382";
    when 16#00995# => romdata <= X"2B781188";
    when 16#00996# => romdata <= X"05565681";
    when 16#00997# => romdata <= X"80190877";
    when 16#00998# => romdata <= X"06537280";
    when 16#00999# => romdata <= X"2EB63878";
    when 16#0099A# => romdata <= X"16700853";
    when 16#0099B# => romdata <= X"53795174";
    when 16#0099C# => romdata <= X"0853722D";
    when 16#0099D# => romdata <= X"FF14FC17";
    when 16#0099E# => romdata <= X"FC177981";
    when 16#0099F# => romdata <= X"2C5A5757";
    when 16#009A0# => romdata <= X"54738025";
    when 16#009A1# => romdata <= X"D6387708";
    when 16#009A2# => romdata <= X"5877FFAD";
    when 16#009A3# => romdata <= X"3880DF8C";
    when 16#009A4# => romdata <= X"0853BC13";
    when 16#009A5# => romdata <= X"08A53879";
    when 16#009A6# => romdata <= X"51FF863F";
    when 16#009A7# => romdata <= X"74085372";
    when 16#009A8# => romdata <= X"2DFF14FC";
    when 16#009A9# => romdata <= X"17FC1779";
    when 16#009AA# => romdata <= X"812C5A57";
    when 16#009AB# => romdata <= X"57547380";
    when 16#009AC# => romdata <= X"25FFA838";
    when 16#009AD# => romdata <= X"D1398057";
    when 16#009AE# => romdata <= X"FF933972";
    when 16#009AF# => romdata <= X"51BC1308";
    when 16#009B0# => romdata <= X"53722D79";
    when 16#009B1# => romdata <= X"51FEDA3F";
    when 16#009B2# => romdata <= X"FF3D0D80";
    when 16#009B3# => romdata <= X"EED80BFC";
    when 16#009B4# => romdata <= X"05700852";
    when 16#009B5# => romdata <= X"5270FF2E";
    when 16#009B6# => romdata <= X"9138702D";
    when 16#009B7# => romdata <= X"FC127008";
    when 16#009B8# => romdata <= X"525270FF";
    when 16#009B9# => romdata <= X"2E098106";
    when 16#009BA# => romdata <= X"F138833D";
    when 16#009BB# => romdata <= X"0D0404FF";
    when 16#009BC# => romdata <= X"BBDB3F04";
    when 16#009BD# => romdata <= X"00000040";
    when 16#009BE# => romdata <= X"68656C70";
    when 16#009BF# => romdata <= X"00000000";
    when 16#009C0# => romdata <= X"3E200000";
    when 16#009C1# => romdata <= X"636F6D6D";
    when 16#009C2# => romdata <= X"616E6420";
    when 16#009C3# => romdata <= X"6E6F7420";
    when 16#009C4# => romdata <= X"666F756E";
    when 16#009C5# => romdata <= X"642E0A00";
    when 16#009C6# => romdata <= X"6D656D00";
    when 16#009C7# => romdata <= X"6C696B65";
    when 16#009C8# => romdata <= X"20780000";
    when 16#009C9# => romdata <= X"776D656D";
    when 16#009CA# => romdata <= X"00000000";
    when 16#009CB# => romdata <= X"77726974";
    when 16#009CC# => romdata <= X"6520776F";
    when 16#009CD# => romdata <= X"72640000";
    when 16#009CE# => romdata <= X"6558616D";
    when 16#009CF# => romdata <= X"696E6520";
    when 16#009D0# => romdata <= X"6D656D6F";
    when 16#009D1# => romdata <= X"72790000";
    when 16#009D2# => romdata <= X"636C6561";
    when 16#009D3# => romdata <= X"72000000";
    when 16#009D4# => romdata <= X"636C6561";
    when 16#009D5# => romdata <= X"72207363";
    when 16#009D6# => romdata <= X"7265656E";
    when 16#009D7# => romdata <= X"00000000";
    when 16#009D8# => romdata <= X"6C656400";
    when 16#009D9# => romdata <= X"73746172";
    when 16#009DA# => romdata <= X"74204C45";
    when 16#009DB# => romdata <= X"44207465";
    when 16#009DC# => romdata <= X"73740000";
    when 16#009DD# => romdata <= X"71756974";
    when 16#009DE# => romdata <= X"00000000";
    when 16#009DF# => romdata <= X"73757070";
    when 16#009E0# => romdata <= X"6F727465";
    when 16#009E1# => romdata <= X"6420636F";
    when 16#009E2# => romdata <= X"6D6D616E";
    when 16#009E3# => romdata <= X"64733A0A";
    when 16#009E4# => romdata <= X"0A000000";
    when 16#009E5# => romdata <= X"202D2000";
    when 16#009E6# => romdata <= X"0A307800";
    when 16#009E7# => romdata <= X"203A2000";
    when 16#009E8# => romdata <= X"0A677265";
    when 16#009E9# => romdata <= X"74682072";
    when 16#009EA# => romdata <= X"65676973";
    when 16#009EB# => romdata <= X"74657273";
    when 16#009EC# => romdata <= X"3A000000";
    when 16#009ED# => romdata <= X"0A636F6E";
    when 16#009EE# => romdata <= X"74726F6C";
    when 16#009EF# => romdata <= X"3A202020";
    when 16#009F0# => romdata <= X"20202030";
    when 16#009F1# => romdata <= X"78000000";
    when 16#009F2# => romdata <= X"0A737461";
    when 16#009F3# => romdata <= X"7475733A";
    when 16#009F4# => romdata <= X"20202020";
    when 16#009F5# => romdata <= X"20202030";
    when 16#009F6# => romdata <= X"78000000";
    when 16#009F7# => romdata <= X"0A6D6163";
    when 16#009F8# => romdata <= X"5F6D7362";
    when 16#009F9# => romdata <= X"3A202020";
    when 16#009FA# => romdata <= X"20202030";
    when 16#009FB# => romdata <= X"78000000";
    when 16#009FC# => romdata <= X"0A6D6163";
    when 16#009FD# => romdata <= X"5F6C7362";
    when 16#009FE# => romdata <= X"3A202020";
    when 16#009FF# => romdata <= X"20202030";
    when 16#00A00# => romdata <= X"78000000";
    when 16#00A01# => romdata <= X"0A6D6469";
    when 16#00A02# => romdata <= X"6F5F636F";
    when 16#00A03# => romdata <= X"6E74726F";
    when 16#00A04# => romdata <= X"6C3A2030";
    when 16#00A05# => romdata <= X"78000000";
    when 16#00A06# => romdata <= X"0A74785F";
    when 16#00A07# => romdata <= X"706F696E";
    when 16#00A08# => romdata <= X"7465723A";
    when 16#00A09# => romdata <= X"20202030";
    when 16#00A0A# => romdata <= X"78000000";
    when 16#00A0B# => romdata <= X"0A72785F";
    when 16#00A0C# => romdata <= X"706F696E";
    when 16#00A0D# => romdata <= X"7465723A";
    when 16#00A0E# => romdata <= X"20202030";
    when 16#00A0F# => romdata <= X"78000000";
    when 16#00A10# => romdata <= X"0A656463";
    when 16#00A11# => romdata <= X"6C5F6970";
    when 16#00A12# => romdata <= X"3A202020";
    when 16#00A13# => romdata <= X"20202030";
    when 16#00A14# => romdata <= X"78000000";
    when 16#00A15# => romdata <= X"0A686173";
    when 16#00A16# => romdata <= X"685F6D73";
    when 16#00A17# => romdata <= X"623A2020";
    when 16#00A18# => romdata <= X"20202030";
    when 16#00A19# => romdata <= X"78000000";
    when 16#00A1A# => romdata <= X"0A686173";
    when 16#00A1B# => romdata <= X"685F6C73";
    when 16#00A1C# => romdata <= X"623A2020";
    when 16#00A1D# => romdata <= X"20202030";
    when 16#00A1E# => romdata <= X"78000000";
    when 16#00A1F# => romdata <= X"0A6D6469";
    when 16#00A20# => romdata <= X"6F207068";
    when 16#00A21# => romdata <= X"79207265";
    when 16#00A22# => romdata <= X"67697374";
    when 16#00A23# => romdata <= X"65727300";
    when 16#00A24# => romdata <= X"0A206D64";
    when 16#00A25# => romdata <= X"696F2070";
    when 16#00A26# => romdata <= X"68793A20";
    when 16#00A27# => romdata <= X"30780000";
    when 16#00A28# => romdata <= X"0A202072";
    when 16#00A29# => romdata <= X"65673A20";
    when 16#00A2A# => romdata <= X"00000000";
    when 16#00A2B# => romdata <= X"2D3E2030";
    when 16#00A2C# => romdata <= X"78000000";
    when 16#00A2D# => romdata <= X"67726574";
    when 16#00A2E# => romdata <= X"682D3E63";
    when 16#00A2F# => romdata <= X"6F6E7472";
    when 16#00A30# => romdata <= X"6F6C3A20";
    when 16#00A31# => romdata <= X"30780000";
    when 16#00A32# => romdata <= X"67726574";
    when 16#00A33# => romdata <= X"682D3E73";
    when 16#00A34# => romdata <= X"74617475";
    when 16#00A35# => romdata <= X"73203A20";
    when 16#00A36# => romdata <= X"30780000";
    when 16#00A37# => romdata <= X"64657363";
    when 16#00A38# => romdata <= X"722D3E63";
    when 16#00A39# => romdata <= X"6F6E7472";
    when 16#00A3A# => romdata <= X"6F6C3A20";
    when 16#00A3B# => romdata <= X"30780000";
    when 16#00A3C# => romdata <= X"77726974";
    when 16#00A3D# => romdata <= X"65206164";
    when 16#00A3E# => romdata <= X"64726573";
    when 16#00A3F# => romdata <= X"733A2030";
    when 16#00A40# => romdata <= X"78000000";
    when 16#00A41# => romdata <= X"20206C65";
    when 16#00A42# => romdata <= X"6E677468";
    when 16#00A43# => romdata <= X"3A203078";
    when 16#00A44# => romdata <= X"00000000";
    when 16#00A45# => romdata <= X"0A0A0000";
    when 16#00A46# => romdata <= X"72656164";
    when 16#00A47# => romdata <= X"20206164";
    when 16#00A48# => romdata <= X"64726573";
    when 16#00A49# => romdata <= X"733A2030";
    when 16#00A4A# => romdata <= X"78000000";
    when 16#00A4B# => romdata <= X"20206578";
    when 16#00A4C# => romdata <= X"70656374";
    when 16#00A4D# => romdata <= X"3A203078";
    when 16#00A4E# => romdata <= X"00000000";
    when 16#00A4F# => romdata <= X"2020676F";
    when 16#00A50# => romdata <= X"743A2030";
    when 16#00A51# => romdata <= X"78000000";
    when 16#00A52# => romdata <= X"20657272";
    when 16#00A53# => romdata <= X"6F720000";
    when 16#00A54# => romdata <= X"206F6B00";
    when 16#00A55# => romdata <= X"6D656D6F";
    when 16#00A56# => romdata <= X"72792074";
    when 16#00A57# => romdata <= X"65737420";
    when 16#00A58# => romdata <= X"696E6974";
    when 16#00A59# => romdata <= X"00000000";
    when 16#00A5A# => romdata <= X"70686173";
    when 16#00A5B# => romdata <= X"65207368";
    when 16#00A5C# => romdata <= X"69667420";
    when 16#00A5D# => romdata <= X"202D2020";
    when 16#00A5E# => romdata <= X"76616C75";
    when 16#00A5F# => romdata <= X"653A2000";
    when 16#00A60# => romdata <= X"20207374";
    when 16#00A61# => romdata <= X"61747573";
    when 16#00A62# => romdata <= X"3A203078";
    when 16#00A63# => romdata <= X"00000000";
    when 16#00A64# => romdata <= X"20202020";
    when 16#00A65# => romdata <= X"20000000";
    when 16#00A66# => romdata <= X"6F6B2020";
    when 16#00A67# => romdata <= X"00000000";
    when 16#00A68# => romdata <= X"4641494C";
    when 16#00A69# => romdata <= X"00000000";
    when 16#00A6A# => romdata <= X"44445220";
    when 16#00A6B# => romdata <= X"6D656D6F";
    when 16#00A6C# => romdata <= X"72792069";
    when 16#00A6D# => romdata <= X"6E666F00";
    when 16#00A6E# => romdata <= X"0A0A6175";
    when 16#00A6F# => romdata <= X"746F2074";
    when 16#00A70# => romdata <= X"5F524552";
    when 16#00A71# => romdata <= X"45534820";
    when 16#00A72# => romdata <= X"3A000000";
    when 16#00A73# => romdata <= X"0A636C6F";
    when 16#00A74# => romdata <= X"636B2065";
    when 16#00A75# => romdata <= X"6E61626C";
    when 16#00A76# => romdata <= X"6520203A";
    when 16#00A77# => romdata <= X"30780000";
    when 16#00A78# => romdata <= X"0A696E69";
    when 16#00A79# => romdata <= X"74616C69";
    when 16#00A7A# => romdata <= X"7A652020";
    when 16#00A7B# => romdata <= X"2020203A";
    when 16#00A7C# => romdata <= X"30780000";
    when 16#00A7D# => romdata <= X"0A636F6C";
    when 16#00A7E# => romdata <= X"756D6E20";
    when 16#00A7F# => romdata <= X"73697A65";
    when 16#00A80# => romdata <= X"2020203A";
    when 16#00A81# => romdata <= X"00000000";
    when 16#00A82# => romdata <= X"0A62616E";
    when 16#00A83# => romdata <= X"6B73697A";
    when 16#00A84# => romdata <= X"65202020";
    when 16#00A85# => romdata <= X"2020203A";
    when 16#00A86# => romdata <= X"00000000";
    when 16#00A87# => romdata <= X"4D627974";
    when 16#00A88# => romdata <= X"65000000";
    when 16#00A89# => romdata <= X"0A745F52";
    when 16#00A8A# => romdata <= X"43442020";
    when 16#00A8B# => romdata <= X"20202020";
    when 16#00A8C# => romdata <= X"2020203A";
    when 16#00A8D# => romdata <= X"00000000";
    when 16#00A8E# => romdata <= X"0A745F52";
    when 16#00A8F# => romdata <= X"46432020";
    when 16#00A90# => romdata <= X"20202020";
    when 16#00A91# => romdata <= X"2020203A";
    when 16#00A92# => romdata <= X"00000000";
    when 16#00A93# => romdata <= X"0A745F52";
    when 16#00A94# => romdata <= X"50202020";
    when 16#00A95# => romdata <= X"20202020";
    when 16#00A96# => romdata <= X"2020203A";
    when 16#00A97# => romdata <= X"00000000";
    when 16#00A98# => romdata <= X"0A726566";
    when 16#00A99# => romdata <= X"72657368";
    when 16#00A9A# => romdata <= X"20656E2E";
    when 16#00A9B# => romdata <= X"2020203A";
    when 16#00A9C# => romdata <= X"30780000";
    when 16#00A9D# => romdata <= X"0A0A4444";
    when 16#00A9E# => romdata <= X"52206672";
    when 16#00A9F# => romdata <= X"65717565";
    when 16#00AA0# => romdata <= X"6E637920";
    when 16#00AA1# => romdata <= X"3A000000";
    when 16#00AA2# => romdata <= X"0A444452";
    when 16#00AA3# => romdata <= X"20646174";
    when 16#00AA4# => romdata <= X"61207769";
    when 16#00AA5# => romdata <= X"6474683A";
    when 16#00AA6# => romdata <= X"00000000";
    when 16#00AA7# => romdata <= X"0A6D6F62";
    when 16#00AA8# => romdata <= X"696C6520";
    when 16#00AA9# => romdata <= X"73757070";
    when 16#00AAA# => romdata <= X"6F72743A";
    when 16#00AAB# => romdata <= X"30780000";
    when 16#00AAC# => romdata <= X"0A0A7374";
    when 16#00AAD# => romdata <= X"61747573";
    when 16#00AAE# => romdata <= X"20726561";
    when 16#00AAF# => romdata <= X"64202020";
    when 16#00AB0# => romdata <= X"3A307800";
    when 16#00AB1# => romdata <= X"0A0A7365";
    when 16#00AB2# => romdata <= X"6C662072";
    when 16#00AB3# => romdata <= X"65667265";
    when 16#00AB4# => romdata <= X"73682020";
    when 16#00AB5# => romdata <= X"3A000000";
    when 16#00AB6# => romdata <= X"20353132";
    when 16#00AB7# => romdata <= X"00000000";
    when 16#00AB8# => romdata <= X"34303639";
    when 16#00AB9# => romdata <= X"00000000";
    when 16#00ABA# => romdata <= X"312F3800";
    when 16#00ABB# => romdata <= X"20617272";
    when 16#00ABC# => romdata <= X"61790000";
    when 16#00ABD# => romdata <= X"0A74656D";
    when 16#00ABE# => romdata <= X"702D636F";
    when 16#00ABF# => romdata <= X"6D702072";
    when 16#00AC0# => romdata <= X"6566723A";
    when 16#00AC1# => romdata <= X"00000000";
    when 16#00AC2# => romdata <= X"C2B04300";
    when 16#00AC3# => romdata <= X"0A647269";
    when 16#00AC4# => romdata <= X"76652073";
    when 16#00AC5# => romdata <= X"7472656E";
    when 16#00AC6# => romdata <= X"6774683A";
    when 16#00AC7# => romdata <= X"00000000";
    when 16#00AC8# => romdata <= X"0A706F77";
    when 16#00AC9# => romdata <= X"65722073";
    when 16#00ACA# => romdata <= X"6176696E";
    when 16#00ACB# => romdata <= X"6720203A";
    when 16#00ACC# => romdata <= X"00000000";
    when 16#00ACD# => romdata <= X"756E6B6E";
    when 16#00ACE# => romdata <= X"6F776E00";
    when 16#00ACF# => romdata <= X"0A745F58";
    when 16#00AD0# => romdata <= X"50202020";
    when 16#00AD1# => romdata <= X"20202020";
    when 16#00AD2# => romdata <= X"2020203A";
    when 16#00AD3# => romdata <= X"00000000";
    when 16#00AD4# => romdata <= X"0A745F58";
    when 16#00AD5# => romdata <= X"53522020";
    when 16#00AD6# => romdata <= X"20202020";
    when 16#00AD7# => romdata <= X"2020203A";
    when 16#00AD8# => romdata <= X"00000000";
    when 16#00AD9# => romdata <= X"0A745F43";
    when 16#00ADA# => romdata <= X"4B452020";
    when 16#00ADB# => romdata <= X"20202020";
    when 16#00ADC# => romdata <= X"2020203A";
    when 16#00ADD# => romdata <= X"00000000";
    when 16#00ADE# => romdata <= X"0A434153";
    when 16#00ADF# => romdata <= X"206C6174";
    when 16#00AE0# => romdata <= X"656E6379";
    when 16#00AE1# => romdata <= X"2020203A";
    when 16#00AE2# => romdata <= X"00000000";
    when 16#00AE3# => romdata <= X"0A6D6F62";
    when 16#00AE4# => romdata <= X"696C6520";
    when 16#00AE5# => romdata <= X"656E6162";
    when 16#00AE6# => romdata <= X"6C65643A";
    when 16#00AE7# => romdata <= X"30780000";
    when 16#00AE8# => romdata <= X"0A0A7068";
    when 16#00AE9# => romdata <= X"7920636F";
    when 16#00AEA# => romdata <= X"6E666967";
    when 16#00AEB# => romdata <= X"20302020";
    when 16#00AEC# => romdata <= X"3A307800";
    when 16#00AED# => romdata <= X"0A0A7068";
    when 16#00AEE# => romdata <= X"7920636F";
    when 16#00AEF# => romdata <= X"6E666967";
    when 16#00AF0# => romdata <= X"20312020";
    when 16#00AF1# => romdata <= X"3A307800";
    when 16#00AF2# => romdata <= X"31303234";
    when 16#00AF3# => romdata <= X"00000000";
    when 16#00AF4# => romdata <= X"32303438";
    when 16#00AF5# => romdata <= X"00000000";
    when 16#00AF6# => romdata <= X"66756C6C";
    when 16#00AF7# => romdata <= X"00000000";
    when 16#00AF8# => romdata <= X"37300000";
    when 16#00AF9# => romdata <= X"64656570";
    when 16#00AFA# => romdata <= X"20706F77";
    when 16#00AFB# => romdata <= X"65722064";
    when 16#00AFC# => romdata <= X"6F776E00";
    when 16#00AFD# => romdata <= X"636C6F63";
    when 16#00AFE# => romdata <= X"6B207374";
    when 16#00AFF# => romdata <= X"6F700000";
    when 16#00B00# => romdata <= X"73656C66";
    when 16#00B01# => romdata <= X"20726566";
    when 16#00B02# => romdata <= X"72657368";
    when 16#00B03# => romdata <= X"00000000";
    when 16#00B04# => romdata <= X"706F7765";
    when 16#00B05# => romdata <= X"7220646F";
    when 16#00B06# => romdata <= X"776E0000";
    when 16#00B07# => romdata <= X"6E6F6E65";
    when 16#00B08# => romdata <= X"00000000";
    when 16#00B09# => romdata <= X"312F3200";
    when 16#00B0A# => romdata <= X"312F3400";
    when 16#00B0B# => romdata <= X"312F3100";
    when 16#00B0C# => romdata <= X"332F3400";
    when 16#00B0D# => romdata <= X"38350000";
    when 16#00B0E# => romdata <= X"34350000";
    when 16#00B0F# => romdata <= X"68616C66";
    when 16#00B10# => romdata <= X"00000000";
    when 16#00B11# => romdata <= X"31350000";
    when 16#00B12# => romdata <= X"61646472";
    when 16#00B13# => romdata <= X"6573733A";
    when 16#00B14# => romdata <= X"20307800";
    when 16#00B15# => romdata <= X"20646174";
    when 16#00B16# => romdata <= X"613A2030";
    when 16#00B17# => romdata <= X"78000000";
    when 16#00B18# => romdata <= X"0A0A4443";
    when 16#00B19# => romdata <= X"4D207068";
    when 16#00B1A# => romdata <= X"61736520";
    when 16#00B1B# => romdata <= X"73686966";
    when 16#00B1C# => romdata <= X"74207465";
    when 16#00B1D# => romdata <= X"7374696E";
    when 16#00B1E# => romdata <= X"67000000";
    when 16#00B1F# => romdata <= X"0A696E69";
    when 16#00B20# => romdata <= X"7469616C";
    when 16#00B21# => romdata <= X"3A200000";
    when 16#00B22# => romdata <= X"676F2064";
    when 16#00B23# => romdata <= X"6F776E00";
    when 16#00B24# => romdata <= X"7363616E";
    when 16#00B25# => romdata <= X"2072616E";
    when 16#00B26# => romdata <= X"67650000";
    when 16#00B27# => romdata <= X"09000000";
    when 16#00B28# => romdata <= X"676F2074";
    when 16#00B29# => romdata <= X"6F206579";
    when 16#00B2A# => romdata <= X"65000000";
    when 16#00B2B# => romdata <= X"6C6F7720";
    when 16#00B2C# => romdata <= X"666F756E";
    when 16#00B2D# => romdata <= X"64000000";
    when 16#00B2E# => romdata <= X"68696768";
    when 16#00B2F# => romdata <= X"20666F75";
    when 16#00B30# => romdata <= X"6E640000";
    when 16#00B31# => romdata <= X"0A6C6F77";
    when 16#00B32# => romdata <= X"3A202020";
    when 16#00B33# => romdata <= X"20202020";
    when 16#00B34# => romdata <= X"20200000";
    when 16#00B35# => romdata <= X"0A686967";
    when 16#00B36# => romdata <= X"683A2020";
    when 16#00B37# => romdata <= X"20202020";
    when 16#00B38# => romdata <= X"20200000";
    when 16#00B39# => romdata <= X"0A646966";
    when 16#00B3A# => romdata <= X"663A2020";
    when 16#00B3B# => romdata <= X"20202020";
    when 16#00B3C# => romdata <= X"20200000";
    when 16#00B3D# => romdata <= X"0A6D696E";
    when 16#00B3E# => romdata <= X"5F657272";
    when 16#00B3F# => romdata <= X"3A202020";
    when 16#00B40# => romdata <= X"20200000";
    when 16#00B41# => romdata <= X"0A6D696E";
    when 16#00B42# => romdata <= X"5F657272";
    when 16#00B43# => romdata <= X"5F706F73";
    when 16#00B44# => romdata <= X"3A200000";
    when 16#00B45# => romdata <= X"676F206D";
    when 16#00B46# => romdata <= X"696E5F65";
    when 16#00B47# => romdata <= X"72726F72";
    when 16#00B48# => romdata <= X"00000000";
    when 16#00B49# => romdata <= X"0A66696E";
    when 16#00B4A# => romdata <= X"616C3A20";
    when 16#00B4B# => romdata <= X"20202020";
    when 16#00B4C# => romdata <= X"20200000";
    when 16#00B4D# => romdata <= X"64636D5F";
    when 16#00B4E# => romdata <= X"74657374";
    when 16#00B4F# => romdata <= X"5F707320";
    when 16#00B50# => romdata <= X"646F6E65";
    when 16#00B51# => romdata <= X"00000000";
    when 16#00B52# => romdata <= X"6C6F7720";
    when 16#00B53# => romdata <= X"4E4F5420";
    when 16#00B54# => romdata <= X"666F756E";
    when 16#00B55# => romdata <= X"64000000";
    when 16#00B56# => romdata <= X"68696768";
    when 16#00B57# => romdata <= X"204E4F54";
    when 16#00B58# => romdata <= X"20666F75";
    when 16#00B59# => romdata <= X"6E640000";
    when 16#00B5A# => romdata <= X"676F207A";
    when 16#00B5B# => romdata <= X"65726F00";
    when 16#00B5C# => romdata <= X"64617461";
    when 16#00B5D# => romdata <= X"2076616C";
    when 16#00B5E# => romdata <= X"69640000";
    when 16#00B5F# => romdata <= X"6C6F7720";
    when 16#00B60# => romdata <= X"20666F75";
    when 16#00B61# => romdata <= X"6E640000";
    when 16#00B62# => romdata <= X"0A646966";
    when 16#00B63# => romdata <= X"662F323A";
    when 16#00B64# => romdata <= X"20202020";
    when 16#00B65# => romdata <= X"20200000";
    when 16#00B66# => romdata <= X"6C6F7720";
    when 16#00B67# => romdata <= X"204E4F54";
    when 16#00B68# => romdata <= X"20666F75";
    when 16#00B69# => romdata <= X"6E640000";
    when 16#00B6A# => romdata <= X"64617461";
    when 16#00B6B# => romdata <= X"204E4F54";
    when 16#00B6C# => romdata <= X"2076616C";
    when 16#00B6D# => romdata <= X"69640000";
    when 16#00B6E# => romdata <= X"74657374";
    when 16#00B6F# => romdata <= X"2E632000";
    when 16#00B70# => romdata <= X"286F6E20";
    when 16#00B71# => romdata <= X"73696D29";
    when 16#00B72# => romdata <= X"0A000000";
    when 16#00B73# => romdata <= X"696E6974";
    when 16#00B74# => romdata <= X"20646F6E";
    when 16#00B75# => romdata <= X"652E0000";
    when 16#00B76# => romdata <= X"286F6E20";
    when 16#00B77# => romdata <= X"68617264";
    when 16#00B78# => romdata <= X"77617265";
    when 16#00B79# => romdata <= X"290A0000";
    when 16#00B7A# => romdata <= X"636F6D70";
    when 16#00B7B# => romdata <= X"696C6564";
    when 16#00B7C# => romdata <= X"3A204A61";
    when 16#00B7D# => romdata <= X"6E203234";
    when 16#00B7E# => romdata <= X"20323031";
    when 16#00B7F# => romdata <= X"31202031";
    when 16#00B80# => romdata <= X"333A3535";
    when 16#00B81# => romdata <= X"3A33330A";
    when 16#00B82# => romdata <= X"00000000";
    when 16#00B83# => romdata <= X"30622020";
    when 16#00B84# => romdata <= X"20202020";
    when 16#00B85# => romdata <= X"20202020";
    when 16#00B86# => romdata <= X"20202020";
    when 16#00B87# => romdata <= X"20202020";
    when 16#00B88# => romdata <= X"20202020";
    when 16#00B89# => romdata <= X"20202020";
    when 16#00B8A# => romdata <= X"20202020";
    when 16#00B8B# => romdata <= X"20200000";
    when 16#00B8C# => romdata <= X"20202020";
    when 16#00B8D# => romdata <= X"20202020";
    when 16#00B8E# => romdata <= X"00000000";
    when 16#00B8F# => romdata <= X"00202020";
    when 16#00B90# => romdata <= X"20202020";
    when 16#00B91# => romdata <= X"20202828";
    when 16#00B92# => romdata <= X"28282820";
    when 16#00B93# => romdata <= X"20202020";
    when 16#00B94# => romdata <= X"20202020";
    when 16#00B95# => romdata <= X"20202020";
    when 16#00B96# => romdata <= X"20202020";
    when 16#00B97# => romdata <= X"20881010";
    when 16#00B98# => romdata <= X"10101010";
    when 16#00B99# => romdata <= X"10101010";
    when 16#00B9A# => romdata <= X"10101010";
    when 16#00B9B# => romdata <= X"10040404";
    when 16#00B9C# => romdata <= X"04040404";
    when 16#00B9D# => romdata <= X"04040410";
    when 16#00B9E# => romdata <= X"10101010";
    when 16#00B9F# => romdata <= X"10104141";
    when 16#00BA0# => romdata <= X"41414141";
    when 16#00BA1# => romdata <= X"01010101";
    when 16#00BA2# => romdata <= X"01010101";
    when 16#00BA3# => romdata <= X"01010101";
    when 16#00BA4# => romdata <= X"01010101";
    when 16#00BA5# => romdata <= X"01010101";
    when 16#00BA6# => romdata <= X"10101010";
    when 16#00BA7# => romdata <= X"10104242";
    when 16#00BA8# => romdata <= X"42424242";
    when 16#00BA9# => romdata <= X"02020202";
    when 16#00BAA# => romdata <= X"02020202";
    when 16#00BAB# => romdata <= X"02020202";
    when 16#00BAC# => romdata <= X"02020202";
    when 16#00BAD# => romdata <= X"02020202";
    when 16#00BAE# => romdata <= X"10101010";
    when 16#00BAF# => romdata <= X"20000000";
    when 16#00BB0# => romdata <= X"00000000";
    when 16#00BB1# => romdata <= X"00000000";
    when 16#00BB2# => romdata <= X"00000000";
    when 16#00BB3# => romdata <= X"00000000";
    when 16#00BB4# => romdata <= X"00000000";
    when 16#00BB5# => romdata <= X"00000000";
    when 16#00BB6# => romdata <= X"00000000";
    when 16#00BB7# => romdata <= X"00000000";
    when 16#00BB8# => romdata <= X"00000000";
    when 16#00BB9# => romdata <= X"00000000";
    when 16#00BBA# => romdata <= X"00000000";
    when 16#00BBB# => romdata <= X"00000000";
    when 16#00BBC# => romdata <= X"00000000";
    when 16#00BBD# => romdata <= X"00000000";
    when 16#00BBE# => romdata <= X"00000000";
    when 16#00BBF# => romdata <= X"00000000";
    when 16#00BC0# => romdata <= X"00000000";
    when 16#00BC1# => romdata <= X"00000000";
    when 16#00BC2# => romdata <= X"00000000";
    when 16#00BC3# => romdata <= X"00000000";
    when 16#00BC4# => romdata <= X"00000000";
    when 16#00BC5# => romdata <= X"00000000";
    when 16#00BC6# => romdata <= X"00000000";
    when 16#00BC7# => romdata <= X"00000000";
    when 16#00BC8# => romdata <= X"00000000";
    when 16#00BC9# => romdata <= X"00000000";
    when 16#00BCA# => romdata <= X"00000000";
    when 16#00BCB# => romdata <= X"00000000";
    when 16#00BCC# => romdata <= X"00000000";
    when 16#00BCD# => romdata <= X"00000000";
    when 16#00BCE# => romdata <= X"00000000";
    when 16#00BCF# => romdata <= X"00000000";
    when 16#00BD0# => romdata <= X"43000000";
    when 16#00BD1# => romdata <= X"64756D6D";
    when 16#00BD2# => romdata <= X"792E6578";
    when 16#00BD3# => romdata <= X"65000000";
    when 16#00BD4# => romdata <= X"00FFFFFF";
    when 16#00BD5# => romdata <= X"FF00FFFF";
    when 16#00BD6# => romdata <= X"FFFF00FF";
    when 16#00BD7# => romdata <= X"FFFFFF00";
    when 16#00BD8# => romdata <= X"00000000";
    when 16#00BD9# => romdata <= X"00000000";
    when 16#00BDA# => romdata <= X"00000000";
    when 16#00BDB# => romdata <= X"00003760";
    when 16#00BDC# => romdata <= X"FFF00000";
    when 16#00BDD# => romdata <= X"80000D00";
    when 16#00BDE# => romdata <= X"80000800";
    when 16#00BDF# => romdata <= X"80000600";
    when 16#00BE0# => romdata <= X"80000300";
    when 16#00BE1# => romdata <= X"80000200";
    when 16#00BE2# => romdata <= X"80000100";
    when 16#00BE3# => romdata <= X"00002F90";
    when 16#00BE4# => romdata <= X"00000000";
    when 16#00BE5# => romdata <= X"000031F8";
    when 16#00BE6# => romdata <= X"00003254";
    when 16#00BE7# => romdata <= X"000032B0";
    when 16#00BE8# => romdata <= X"00000000";
    when 16#00BE9# => romdata <= X"00000000";
    when 16#00BEA# => romdata <= X"00000000";
    when 16#00BEB# => romdata <= X"00000000";
    when 16#00BEC# => romdata <= X"00000000";
    when 16#00BED# => romdata <= X"00000000";
    when 16#00BEE# => romdata <= X"00000000";
    when 16#00BEF# => romdata <= X"00000000";
    when 16#00BF0# => romdata <= X"00000000";
    when 16#00BF1# => romdata <= X"00002F40";
    when 16#00BF2# => romdata <= X"00000000";
    when 16#00BF3# => romdata <= X"00000000";
    when 16#00BF4# => romdata <= X"00000000";
    when 16#00BF5# => romdata <= X"00000000";
    when 16#00BF6# => romdata <= X"00000000";
    when 16#00BF7# => romdata <= X"00000000";
    when 16#00BF8# => romdata <= X"00000000";
    when 16#00BF9# => romdata <= X"00000000";
    when 16#00BFA# => romdata <= X"00000000";
    when 16#00BFB# => romdata <= X"00000000";
    when 16#00BFC# => romdata <= X"00000000";
    when 16#00BFD# => romdata <= X"00000000";
    when 16#00BFE# => romdata <= X"00000000";
    when 16#00BFF# => romdata <= X"00000000";
    when 16#00C00# => romdata <= X"00000000";
    when 16#00C01# => romdata <= X"00000000";
    when 16#00C02# => romdata <= X"00000000";
    when 16#00C03# => romdata <= X"00000000";
    when 16#00C04# => romdata <= X"00000000";
    when 16#00C05# => romdata <= X"00000000";
    when 16#00C06# => romdata <= X"00000000";
    when 16#00C07# => romdata <= X"00000000";
    when 16#00C08# => romdata <= X"00000000";
    when 16#00C09# => romdata <= X"00000000";
    when 16#00C0A# => romdata <= X"00000000";
    when 16#00C0B# => romdata <= X"00000000";
    when 16#00C0C# => romdata <= X"00000000";
    when 16#00C0D# => romdata <= X"00000000";
    when 16#00C0E# => romdata <= X"00000001";
    when 16#00C0F# => romdata <= X"330EABCD";
    when 16#00C10# => romdata <= X"1234E66D";
    when 16#00C11# => romdata <= X"DEEC0005";
    when 16#00C12# => romdata <= X"000B0000";
    when 16#00C13# => romdata <= X"00000000";
    when 16#00C14# => romdata <= X"00000000";
    when 16#00C15# => romdata <= X"00000000";
    when 16#00C16# => romdata <= X"00000000";
    when 16#00C17# => romdata <= X"00000000";
    when 16#00C18# => romdata <= X"00000000";
    when 16#00C19# => romdata <= X"00000000";
    when 16#00C1A# => romdata <= X"00000000";
    when 16#00C1B# => romdata <= X"00000000";
    when 16#00C1C# => romdata <= X"00000000";
    when 16#00C1D# => romdata <= X"00000000";
    when 16#00C1E# => romdata <= X"00000000";
    when 16#00C1F# => romdata <= X"00000000";
    when 16#00C20# => romdata <= X"00000000";
    when 16#00C21# => romdata <= X"00000000";
    when 16#00C22# => romdata <= X"00000000";
    when 16#00C23# => romdata <= X"00000000";
    when 16#00C24# => romdata <= X"00000000";
    when 16#00C25# => romdata <= X"00000000";
    when 16#00C26# => romdata <= X"00000000";
    when 16#00C27# => romdata <= X"00000000";
    when 16#00C28# => romdata <= X"00000000";
    when 16#00C29# => romdata <= X"00000000";
    when 16#00C2A# => romdata <= X"00000000";
    when 16#00C2B# => romdata <= X"00000000";
    when 16#00C2C# => romdata <= X"00000000";
    when 16#00C2D# => romdata <= X"00000000";
    when 16#00C2E# => romdata <= X"00000000";
    when 16#00C2F# => romdata <= X"00000000";
    when 16#00C30# => romdata <= X"00000000";
    when 16#00C31# => romdata <= X"00000000";
    when 16#00C32# => romdata <= X"00000000";
    when 16#00C33# => romdata <= X"00000000";
    when 16#00C34# => romdata <= X"00000000";
    when 16#00C35# => romdata <= X"00000000";
    when 16#00C36# => romdata <= X"00000000";
    when 16#00C37# => romdata <= X"00000000";
    when 16#00C38# => romdata <= X"00000000";
    when 16#00C39# => romdata <= X"00000000";
    when 16#00C3A# => romdata <= X"00000000";
    when 16#00C3B# => romdata <= X"00000000";
    when 16#00C3C# => romdata <= X"00000000";
    when 16#00C3D# => romdata <= X"00000000";
    when 16#00C3E# => romdata <= X"00000000";
    when 16#00C3F# => romdata <= X"00000000";
    when 16#00C40# => romdata <= X"00000000";
    when 16#00C41# => romdata <= X"00000000";
    when 16#00C42# => romdata <= X"00000000";
    when 16#00C43# => romdata <= X"00000000";
    when 16#00C44# => romdata <= X"00000000";
    when 16#00C45# => romdata <= X"00000000";
    when 16#00C46# => romdata <= X"00000000";
    when 16#00C47# => romdata <= X"00000000";
    when 16#00C48# => romdata <= X"00000000";
    when 16#00C49# => romdata <= X"00000000";
    when 16#00C4A# => romdata <= X"00000000";
    when 16#00C4B# => romdata <= X"00000000";
    when 16#00C4C# => romdata <= X"00000000";
    when 16#00C4D# => romdata <= X"00000000";
    when 16#00C4E# => romdata <= X"00000000";
    when 16#00C4F# => romdata <= X"00000000";
    when 16#00C50# => romdata <= X"00000000";
    when 16#00C51# => romdata <= X"00000000";
    when 16#00C52# => romdata <= X"00000000";
    when 16#00C53# => romdata <= X"00000000";
    when 16#00C54# => romdata <= X"00000000";
    when 16#00C55# => romdata <= X"00000000";
    when 16#00C56# => romdata <= X"00000000";
    when 16#00C57# => romdata <= X"00000000";
    when 16#00C58# => romdata <= X"00000000";
    when 16#00C59# => romdata <= X"00000000";
    when 16#00C5A# => romdata <= X"00000000";
    when 16#00C5B# => romdata <= X"00000000";
    when 16#00C5C# => romdata <= X"00000000";
    when 16#00C5D# => romdata <= X"00000000";
    when 16#00C5E# => romdata <= X"00000000";
    when 16#00C5F# => romdata <= X"00000000";
    when 16#00C60# => romdata <= X"00000000";
    when 16#00C61# => romdata <= X"00000000";
    when 16#00C62# => romdata <= X"00000000";
    when 16#00C63# => romdata <= X"00000000";
    when 16#00C64# => romdata <= X"00000000";
    when 16#00C65# => romdata <= X"00000000";
    when 16#00C66# => romdata <= X"00000000";
    when 16#00C67# => romdata <= X"00000000";
    when 16#00C68# => romdata <= X"00000000";
    when 16#00C69# => romdata <= X"00000000";
    when 16#00C6A# => romdata <= X"00000000";
    when 16#00C6B# => romdata <= X"00000000";
    when 16#00C6C# => romdata <= X"00000000";
    when 16#00C6D# => romdata <= X"00000000";
    when 16#00C6E# => romdata <= X"00000000";
    when 16#00C6F# => romdata <= X"00000000";
    when 16#00C70# => romdata <= X"00000000";
    when 16#00C71# => romdata <= X"00000000";
    when 16#00C72# => romdata <= X"00000000";
    when 16#00C73# => romdata <= X"00000000";
    when 16#00C74# => romdata <= X"00000000";
    when 16#00C75# => romdata <= X"00000000";
    when 16#00C76# => romdata <= X"00000000";
    when 16#00C77# => romdata <= X"00000000";
    when 16#00C78# => romdata <= X"00000000";
    when 16#00C79# => romdata <= X"00000000";
    when 16#00C7A# => romdata <= X"00000000";
    when 16#00C7B# => romdata <= X"00000000";
    when 16#00C7C# => romdata <= X"00000000";
    when 16#00C7D# => romdata <= X"00000000";
    when 16#00C7E# => romdata <= X"00000000";
    when 16#00C7F# => romdata <= X"00000000";
    when 16#00C80# => romdata <= X"00000000";
    when 16#00C81# => romdata <= X"00000000";
    when 16#00C82# => romdata <= X"00000000";
    when 16#00C83# => romdata <= X"00000000";
    when 16#00C84# => romdata <= X"00000000";
    when 16#00C85# => romdata <= X"00000000";
    when 16#00C86# => romdata <= X"00000000";
    when 16#00C87# => romdata <= X"00000000";
    when 16#00C88# => romdata <= X"00000000";
    when 16#00C89# => romdata <= X"00000000";
    when 16#00C8A# => romdata <= X"00000000";
    when 16#00C8B# => romdata <= X"00000000";
    when 16#00C8C# => romdata <= X"00000000";
    when 16#00C8D# => romdata <= X"00000000";
    when 16#00C8E# => romdata <= X"00000000";
    when 16#00C8F# => romdata <= X"00000000";
    when 16#00C90# => romdata <= X"00000000";
    when 16#00C91# => romdata <= X"00000000";
    when 16#00C92# => romdata <= X"00000000";
    when 16#00C93# => romdata <= X"00000000";
    when 16#00C94# => romdata <= X"00000000";
    when 16#00C95# => romdata <= X"00000000";
    when 16#00C96# => romdata <= X"00000000";
    when 16#00C97# => romdata <= X"00000000";
    when 16#00C98# => romdata <= X"00000000";
    when 16#00C99# => romdata <= X"00000000";
    when 16#00C9A# => romdata <= X"00000000";
    when 16#00C9B# => romdata <= X"00000000";
    when 16#00C9C# => romdata <= X"00000000";
    when 16#00C9D# => romdata <= X"00000000";
    when 16#00C9E# => romdata <= X"00000000";
    when 16#00C9F# => romdata <= X"00000000";
    when 16#00CA0# => romdata <= X"00000000";
    when 16#00CA1# => romdata <= X"00000000";
    when 16#00CA2# => romdata <= X"00000000";
    when 16#00CA3# => romdata <= X"00000000";
    when 16#00CA4# => romdata <= X"00000000";
    when 16#00CA5# => romdata <= X"00000000";
    when 16#00CA6# => romdata <= X"00000000";
    when 16#00CA7# => romdata <= X"00000000";
    when 16#00CA8# => romdata <= X"00000000";
    when 16#00CA9# => romdata <= X"00000000";
    when 16#00CAA# => romdata <= X"00000000";
    when 16#00CAB# => romdata <= X"00000000";
    when 16#00CAC# => romdata <= X"00000000";
    when 16#00CAD# => romdata <= X"00000000";
    when 16#00CAE# => romdata <= X"00000000";
    when 16#00CAF# => romdata <= X"00000000";
    when 16#00CB0# => romdata <= X"00000000";
    when 16#00CB1# => romdata <= X"00000000";
    when 16#00CB2# => romdata <= X"00000000";
    when 16#00CB3# => romdata <= X"00000000";
    when 16#00CB4# => romdata <= X"00000000";
    when 16#00CB5# => romdata <= X"00000000";
    when 16#00CB6# => romdata <= X"00000000";
    when 16#00CB7# => romdata <= X"00000000";
    when 16#00CB8# => romdata <= X"00000000";
    when 16#00CB9# => romdata <= X"00000000";
    when 16#00CBA# => romdata <= X"00000000";
    when 16#00CBB# => romdata <= X"00000000";
    when 16#00CBC# => romdata <= X"00000000";
    when 16#00CBD# => romdata <= X"00000000";
    when 16#00CBE# => romdata <= X"00000000";
    when 16#00CBF# => romdata <= X"00000000";
    when 16#00CC0# => romdata <= X"00000000";
    when 16#00CC1# => romdata <= X"00000000";
    when 16#00CC2# => romdata <= X"00000000";
    when 16#00CC3# => romdata <= X"00000000";
    when 16#00CC4# => romdata <= X"00000000";
    when 16#00CC5# => romdata <= X"00000000";
    when 16#00CC6# => romdata <= X"00000000";
    when 16#00CC7# => romdata <= X"00000000";
    when 16#00CC8# => romdata <= X"00000000";
    when 16#00CC9# => romdata <= X"00000000";
    when 16#00CCA# => romdata <= X"00000000";
    when 16#00CCB# => romdata <= X"00000000";
    when 16#00CCC# => romdata <= X"00000000";
    when 16#00CCD# => romdata <= X"00000000";
    when 16#00CCE# => romdata <= X"00000000";
    when 16#00CCF# => romdata <= X"FFFFFFFF";
    when 16#00CD0# => romdata <= X"00000000";
    when 16#00CD1# => romdata <= X"00020000";
    when 16#00CD2# => romdata <= X"00000000";
    when 16#00CD3# => romdata <= X"00000000";
    when 16#00CD4# => romdata <= X"00003348";
    when 16#00CD5# => romdata <= X"00003348";
    when 16#00CD6# => romdata <= X"00003350";
    when 16#00CD7# => romdata <= X"00003350";
    when 16#00CD8# => romdata <= X"00003358";
    when 16#00CD9# => romdata <= X"00003358";
    when 16#00CDA# => romdata <= X"00003360";
    when 16#00CDB# => romdata <= X"00003360";
    when 16#00CDC# => romdata <= X"00003368";
    when 16#00CDD# => romdata <= X"00003368";
    when 16#00CDE# => romdata <= X"00003370";
    when 16#00CDF# => romdata <= X"00003370";
    when 16#00CE0# => romdata <= X"00003378";
    when 16#00CE1# => romdata <= X"00003378";
    when 16#00CE2# => romdata <= X"00003380";
    when 16#00CE3# => romdata <= X"00003380";
    when 16#00CE4# => romdata <= X"00003388";
    when 16#00CE5# => romdata <= X"00003388";
    when 16#00CE6# => romdata <= X"00003390";
    when 16#00CE7# => romdata <= X"00003390";
    when 16#00CE8# => romdata <= X"00003398";
    when 16#00CE9# => romdata <= X"00003398";
    when 16#00CEA# => romdata <= X"000033A0";
    when 16#00CEB# => romdata <= X"000033A0";
    when 16#00CEC# => romdata <= X"000033A8";
    when 16#00CED# => romdata <= X"000033A8";
    when 16#00CEE# => romdata <= X"000033B0";
    when 16#00CEF# => romdata <= X"000033B0";
    when 16#00CF0# => romdata <= X"000033B8";
    when 16#00CF1# => romdata <= X"000033B8";
    when 16#00CF2# => romdata <= X"000033C0";
    when 16#00CF3# => romdata <= X"000033C0";
    when 16#00CF4# => romdata <= X"000033C8";
    when 16#00CF5# => romdata <= X"000033C8";
    when 16#00CF6# => romdata <= X"000033D0";
    when 16#00CF7# => romdata <= X"000033D0";
    when 16#00CF8# => romdata <= X"000033D8";
    when 16#00CF9# => romdata <= X"000033D8";
    when 16#00CFA# => romdata <= X"000033E0";
    when 16#00CFB# => romdata <= X"000033E0";
    when 16#00CFC# => romdata <= X"000033E8";
    when 16#00CFD# => romdata <= X"000033E8";
    when 16#00CFE# => romdata <= X"000033F0";
    when 16#00CFF# => romdata <= X"000033F0";
    when 16#00D00# => romdata <= X"000033F8";
    when 16#00D01# => romdata <= X"000033F8";
    when 16#00D02# => romdata <= X"00003400";
    when 16#00D03# => romdata <= X"00003400";
    when 16#00D04# => romdata <= X"00003408";
    when 16#00D05# => romdata <= X"00003408";
    when 16#00D06# => romdata <= X"00003410";
    when 16#00D07# => romdata <= X"00003410";
    when 16#00D08# => romdata <= X"00003418";
    when 16#00D09# => romdata <= X"00003418";
    when 16#00D0A# => romdata <= X"00003420";
    when 16#00D0B# => romdata <= X"00003420";
    when 16#00D0C# => romdata <= X"00003428";
    when 16#00D0D# => romdata <= X"00003428";
    when 16#00D0E# => romdata <= X"00003430";
    when 16#00D0F# => romdata <= X"00003430";
    when 16#00D10# => romdata <= X"00003438";
    when 16#00D11# => romdata <= X"00003438";
    when 16#00D12# => romdata <= X"00003440";
    when 16#00D13# => romdata <= X"00003440";
    when 16#00D14# => romdata <= X"00003448";
    when 16#00D15# => romdata <= X"00003448";
    when 16#00D16# => romdata <= X"00003450";
    when 16#00D17# => romdata <= X"00003450";
    when 16#00D18# => romdata <= X"00003458";
    when 16#00D19# => romdata <= X"00003458";
    when 16#00D1A# => romdata <= X"00003460";
    when 16#00D1B# => romdata <= X"00003460";
    when 16#00D1C# => romdata <= X"00003468";
    when 16#00D1D# => romdata <= X"00003468";
    when 16#00D1E# => romdata <= X"00003470";
    when 16#00D1F# => romdata <= X"00003470";
    when 16#00D20# => romdata <= X"00003478";
    when 16#00D21# => romdata <= X"00003478";
    when 16#00D22# => romdata <= X"00003480";
    when 16#00D23# => romdata <= X"00003480";
    when 16#00D24# => romdata <= X"00003488";
    when 16#00D25# => romdata <= X"00003488";
    when 16#00D26# => romdata <= X"00003490";
    when 16#00D27# => romdata <= X"00003490";
    when 16#00D28# => romdata <= X"00003498";
    when 16#00D29# => romdata <= X"00003498";
    when 16#00D2A# => romdata <= X"000034A0";
    when 16#00D2B# => romdata <= X"000034A0";
    when 16#00D2C# => romdata <= X"000034A8";
    when 16#00D2D# => romdata <= X"000034A8";
    when 16#00D2E# => romdata <= X"000034B0";
    when 16#00D2F# => romdata <= X"000034B0";
    when 16#00D30# => romdata <= X"000034B8";
    when 16#00D31# => romdata <= X"000034B8";
    when 16#00D32# => romdata <= X"000034C0";
    when 16#00D33# => romdata <= X"000034C0";
    when 16#00D34# => romdata <= X"000034C8";
    when 16#00D35# => romdata <= X"000034C8";
    when 16#00D36# => romdata <= X"000034D0";
    when 16#00D37# => romdata <= X"000034D0";
    when 16#00D38# => romdata <= X"000034D8";
    when 16#00D39# => romdata <= X"000034D8";
    when 16#00D3A# => romdata <= X"000034E0";
    when 16#00D3B# => romdata <= X"000034E0";
    when 16#00D3C# => romdata <= X"000034E8";
    when 16#00D3D# => romdata <= X"000034E8";
    when 16#00D3E# => romdata <= X"000034F0";
    when 16#00D3F# => romdata <= X"000034F0";
    when 16#00D40# => romdata <= X"000034F8";
    when 16#00D41# => romdata <= X"000034F8";
    when 16#00D42# => romdata <= X"00003500";
    when 16#00D43# => romdata <= X"00003500";
    when 16#00D44# => romdata <= X"00003508";
    when 16#00D45# => romdata <= X"00003508";
    when 16#00D46# => romdata <= X"00003510";
    when 16#00D47# => romdata <= X"00003510";
    when 16#00D48# => romdata <= X"00003518";
    when 16#00D49# => romdata <= X"00003518";
    when 16#00D4A# => romdata <= X"00003520";
    when 16#00D4B# => romdata <= X"00003520";
    when 16#00D4C# => romdata <= X"00003528";
    when 16#00D4D# => romdata <= X"00003528";
    when 16#00D4E# => romdata <= X"00003530";
    when 16#00D4F# => romdata <= X"00003530";
    when 16#00D50# => romdata <= X"00003538";
    when 16#00D51# => romdata <= X"00003538";
    when 16#00D52# => romdata <= X"00003540";
    when 16#00D53# => romdata <= X"00003540";
    when 16#00D54# => romdata <= X"00003548";
    when 16#00D55# => romdata <= X"00003548";
    when 16#00D56# => romdata <= X"00003550";
    when 16#00D57# => romdata <= X"00003550";
    when 16#00D58# => romdata <= X"00003558";
    when 16#00D59# => romdata <= X"00003558";
    when 16#00D5A# => romdata <= X"00003560";
    when 16#00D5B# => romdata <= X"00003560";
    when 16#00D5C# => romdata <= X"00003568";
    when 16#00D5D# => romdata <= X"00003568";
    when 16#00D5E# => romdata <= X"00003570";
    when 16#00D5F# => romdata <= X"00003570";
    when 16#00D60# => romdata <= X"00003578";
    when 16#00D61# => romdata <= X"00003578";
    when 16#00D62# => romdata <= X"00003580";
    when 16#00D63# => romdata <= X"00003580";
    when 16#00D64# => romdata <= X"00003588";
    when 16#00D65# => romdata <= X"00003588";
    when 16#00D66# => romdata <= X"00003590";
    when 16#00D67# => romdata <= X"00003590";
    when 16#00D68# => romdata <= X"00003598";
    when 16#00D69# => romdata <= X"00003598";
    when 16#00D6A# => romdata <= X"000035A0";
    when 16#00D6B# => romdata <= X"000035A0";
    when 16#00D6C# => romdata <= X"000035A8";
    when 16#00D6D# => romdata <= X"000035A8";
    when 16#00D6E# => romdata <= X"000035B0";
    when 16#00D6F# => romdata <= X"000035B0";
    when 16#00D70# => romdata <= X"000035B8";
    when 16#00D71# => romdata <= X"000035B8";
    when 16#00D72# => romdata <= X"000035C0";
    when 16#00D73# => romdata <= X"000035C0";
    when 16#00D74# => romdata <= X"000035C8";
    when 16#00D75# => romdata <= X"000035C8";
    when 16#00D76# => romdata <= X"000035D0";
    when 16#00D77# => romdata <= X"000035D0";
    when 16#00D78# => romdata <= X"000035D8";
    when 16#00D79# => romdata <= X"000035D8";
    when 16#00D7A# => romdata <= X"000035E0";
    when 16#00D7B# => romdata <= X"000035E0";
    when 16#00D7C# => romdata <= X"000035E8";
    when 16#00D7D# => romdata <= X"000035E8";
    when 16#00D7E# => romdata <= X"000035F0";
    when 16#00D7F# => romdata <= X"000035F0";
    when 16#00D80# => romdata <= X"000035F8";
    when 16#00D81# => romdata <= X"000035F8";
    when 16#00D82# => romdata <= X"00003600";
    when 16#00D83# => romdata <= X"00003600";
    when 16#00D84# => romdata <= X"00003608";
    when 16#00D85# => romdata <= X"00003608";
    when 16#00D86# => romdata <= X"00003610";
    when 16#00D87# => romdata <= X"00003610";
    when 16#00D88# => romdata <= X"00003618";
    when 16#00D89# => romdata <= X"00003618";
    when 16#00D8A# => romdata <= X"00003620";
    when 16#00D8B# => romdata <= X"00003620";
    when 16#00D8C# => romdata <= X"00003628";
    when 16#00D8D# => romdata <= X"00003628";
    when 16#00D8E# => romdata <= X"00003630";
    when 16#00D8F# => romdata <= X"00003630";
    when 16#00D90# => romdata <= X"00003638";
    when 16#00D91# => romdata <= X"00003638";
    when 16#00D92# => romdata <= X"00003640";
    when 16#00D93# => romdata <= X"00003640";
    when 16#00D94# => romdata <= X"00003648";
    when 16#00D95# => romdata <= X"00003648";
    when 16#00D96# => romdata <= X"00003650";
    when 16#00D97# => romdata <= X"00003650";
    when 16#00D98# => romdata <= X"00003658";
    when 16#00D99# => romdata <= X"00003658";
    when 16#00D9A# => romdata <= X"00003660";
    when 16#00D9B# => romdata <= X"00003660";
    when 16#00D9C# => romdata <= X"00003668";
    when 16#00D9D# => romdata <= X"00003668";
    when 16#00D9E# => romdata <= X"00003670";
    when 16#00D9F# => romdata <= X"00003670";
    when 16#00DA0# => romdata <= X"00003678";
    when 16#00DA1# => romdata <= X"00003678";
    when 16#00DA2# => romdata <= X"00003680";
    when 16#00DA3# => romdata <= X"00003680";
    when 16#00DA4# => romdata <= X"00003688";
    when 16#00DA5# => romdata <= X"00003688";
    when 16#00DA6# => romdata <= X"00003690";
    when 16#00DA7# => romdata <= X"00003690";
    when 16#00DA8# => romdata <= X"00003698";
    when 16#00DA9# => romdata <= X"00003698";
    when 16#00DAA# => romdata <= X"000036A0";
    when 16#00DAB# => romdata <= X"000036A0";
    when 16#00DAC# => romdata <= X"000036A8";
    when 16#00DAD# => romdata <= X"000036A8";
    when 16#00DAE# => romdata <= X"000036B0";
    when 16#00DAF# => romdata <= X"000036B0";
    when 16#00DB0# => romdata <= X"000036B8";
    when 16#00DB1# => romdata <= X"000036B8";
    when 16#00DB2# => romdata <= X"000036C0";
    when 16#00DB3# => romdata <= X"000036C0";
    when 16#00DB4# => romdata <= X"000036C8";
    when 16#00DB5# => romdata <= X"000036C8";
    when 16#00DB6# => romdata <= X"000036D0";
    when 16#00DB7# => romdata <= X"000036D0";
    when 16#00DB8# => romdata <= X"000036D8";
    when 16#00DB9# => romdata <= X"000036D8";
    when 16#00DBA# => romdata <= X"000036E0";
    when 16#00DBB# => romdata <= X"000036E0";
    when 16#00DBC# => romdata <= X"000036E8";
    when 16#00DBD# => romdata <= X"000036E8";
    when 16#00DBE# => romdata <= X"000036F0";
    when 16#00DBF# => romdata <= X"000036F0";
    when 16#00DC0# => romdata <= X"000036F8";
    when 16#00DC1# => romdata <= X"000036F8";
    when 16#00DC2# => romdata <= X"00003700";
    when 16#00DC3# => romdata <= X"00003700";
    when 16#00DC4# => romdata <= X"00003708";
    when 16#00DC5# => romdata <= X"00003708";
    when 16#00DC6# => romdata <= X"00003710";
    when 16#00DC7# => romdata <= X"00003710";
    when 16#00DC8# => romdata <= X"00003718";
    when 16#00DC9# => romdata <= X"00003718";
    when 16#00DCA# => romdata <= X"00003720";
    when 16#00DCB# => romdata <= X"00003720";
    when 16#00DCC# => romdata <= X"00003728";
    when 16#00DCD# => romdata <= X"00003728";
    when 16#00DCE# => romdata <= X"00003730";
    when 16#00DCF# => romdata <= X"00003730";
    when 16#00DD0# => romdata <= X"00003738";
    when 16#00DD1# => romdata <= X"00003738";
    when 16#00DD2# => romdata <= X"00003740";
    when 16#00DD3# => romdata <= X"00003740";
    when 16#00DD4# => romdata <= X"00002F44";
    when 16#00DD5# => romdata <= X"FFFFFFFF";
    when 16#00DD6# => romdata <= X"00000000";
    when 16#00DD7# => romdata <= X"FFFFFFFF";
    when 16#00DD8# => romdata <= X"00000000";
    when 16#00DD9# => romdata <= X"00000000";
    when 16#00DDA# => romdata <= X"00000000";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
