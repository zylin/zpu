package version is

    constant version_time_c : string( 1 to 21) := "Nov 07 2011  11:21:56";

end package version;
