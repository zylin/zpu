library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

library zylin;
use zylin.zpu_config.all;
use zylin.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"800b0b0b",
1 => x"0b0b8070",
2 => x"0b0b80d6",
3 => x"f00c3a0b",
4 => x"0b80cd92",
5 => x"04000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"80cde02d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b0b2a",
20 => x"83ffff06",
21 => x"52040000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b0b2b09",
29 => x"067383ff",
30 => x"ff0b0b0b",
31 => x"0b83a504",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"72728072",
73 => x"8106ff05",
74 => x"09720605",
75 => x"71105272",
76 => x"0a100a53",
77 => x"72ed3851",
78 => x"51535104",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"04067383",
106 => x"06098105",
107 => x"8205832b",
108 => x"0b2b0772",
109 => x"fc060c51",
110 => x"51040000",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04098105",
139 => x"83051010",
140 => x"102b0772",
141 => x"fc060c51",
142 => x"51040000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80d6",
162 => x"dc738306",
163 => x"10100508",
164 => x"067381ff",
165 => x"06738306",
166 => x"0b0b0b84",
167 => x"a9040000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0b8e",
171 => x"fd2d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0b90",
179 => x"af2d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07535050",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075350",
199 => x"50040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80d6ec0c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"04000000",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"839f3f80",
257 => x"cdf83f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51043c04",
267 => x"70700b0b",
268 => x"80e6d808",
269 => x"52841208",
270 => x"70810651",
271 => x"5170f638",
272 => x"710881ff",
273 => x"06800c50",
274 => x"50047070",
275 => x"0b0b80e6",
276 => x"d8085284",
277 => x"1208700a",
278 => x"100a7081",
279 => x"06515151",
280 => x"70f13873",
281 => x"720c5050",
282 => x"0480d6ec",
283 => x"08802ea8",
284 => x"38838080",
285 => x"0b0b0b80",
286 => x"e6d80c82",
287 => x"a0800b0b",
288 => x"0b80e6dc",
289 => x"0c829080",
290 => x"0b80e6ec",
291 => x"0c0b0b80",
292 => x"e6e00b80",
293 => x"e6f00c04",
294 => x"f8808080",
295 => x"a40b0b0b",
296 => x"80e6d80c",
297 => x"f8808082",
298 => x"800b0b0b",
299 => x"80e6dc0c",
300 => x"f8808084",
301 => x"800b80e6",
302 => x"ec0cf880",
303 => x"8080940b",
304 => x"80e6f00c",
305 => x"f8808080",
306 => x"9c0b80e6",
307 => x"e80cf880",
308 => x"8080a00b",
309 => x"80e6f40c",
310 => x"04f23d0d",
311 => x"600b0b80",
312 => x"e6dc0856",
313 => x"5d82750c",
314 => x"8059805a",
315 => x"800b8f3d",
316 => x"71101017",
317 => x"70085a57",
318 => x"5d5b8077",
319 => x"81ff067c",
320 => x"832b5658",
321 => x"5276537b",
322 => x"5182fc3f",
323 => x"7d7f7a72",
324 => x"077c7207",
325 => x"71716081",
326 => x"05415f5d",
327 => x"5b595755",
328 => x"7a8724bb",
329 => x"380b0b80",
330 => x"e6dc087b",
331 => x"10101170",
332 => x"08595155",
333 => x"807781ff",
334 => x"067c832b",
335 => x"56585276",
336 => x"537b5182",
337 => x"c23f7d7f",
338 => x"7a72077c",
339 => x"72077171",
340 => x"60810541",
341 => x"5f5d5b59",
342 => x"5755877b",
343 => x"25c73876",
344 => x"7d0c7784",
345 => x"1e0c7c80",
346 => x"0c903d0d",
347 => x"04707080",
348 => x"e6e43351",
349 => x"70a73880",
350 => x"d6f80870",
351 => x"08525270",
352 => x"802e9438",
353 => x"841280d6",
354 => x"f80c702d",
355 => x"80d6f808",
356 => x"70085252",
357 => x"70ee3881",
358 => x"0b80e6e4",
359 => x"34505004",
360 => x"04700b0b",
361 => x"80e6d408",
362 => x"802e8e38",
363 => x"0b0b0b0b",
364 => x"800b802e",
365 => x"09810683",
366 => x"3850040b",
367 => x"0b80e6d4",
368 => x"510b0b0b",
369 => x"f4ba3f50",
370 => x"04048c08",
371 => x"028c0c70",
372 => x"70707080",
373 => x"0b8c08fc",
374 => x"050c8c08",
375 => x"fc050889",
376 => x"24818e38",
377 => x"0b0b80d6",
378 => x"a85188f3",
379 => x"3f0b0b80",
380 => x"d6b85188",
381 => x"ea3ffc0b",
382 => x"80e6f80c",
383 => x"80e6f808",
384 => x"812c5372",
385 => x"fe2e8438",
386 => x"86f13f8a",
387 => x"0b80e6fc",
388 => x"0c80e6fc",
389 => x"0880e6f8",
390 => x"08295372",
391 => x"d82e8438",
392 => x"86d93f8a",
393 => x"0b80e6f8",
394 => x"0c84e2ad",
395 => x"800b80e6",
396 => x"fc0c80e6",
397 => x"fc0880e6",
398 => x"f8082953",
399 => x"72afd7c2",
400 => x"802e8438",
401 => x"86b53f81",
402 => x"0a0b80e6",
403 => x"f80cff0b",
404 => x"80e6fc0c",
405 => x"80e6fc08",
406 => x"80e6f808",
407 => x"25843886",
408 => x"9a3f8c08",
409 => x"fc050881",
410 => x"058c08fc",
411 => x"050cfeea",
412 => x"398c08fc",
413 => x"05088a2e",
414 => x"843885ff",
415 => x"3f72800c",
416 => x"50505050",
417 => x"8c0c048c",
418 => x"08028c0c",
419 => x"f53d0d8c",
420 => x"08940508",
421 => x"9d388c08",
422 => x"8c05088c",
423 => x"08900508",
424 => x"8c088805",
425 => x"08585654",
426 => x"73760c74",
427 => x"84170c81",
428 => x"bf39800b",
429 => x"8c08f005",
430 => x"0c800b8c",
431 => x"08f4050c",
432 => x"8c088c05",
433 => x"088c0890",
434 => x"05085654",
435 => x"738c08f0",
436 => x"050c748c",
437 => x"08f4050c",
438 => x"8c08f805",
439 => x"8c08f005",
440 => x"56568870",
441 => x"54755376",
442 => x"5254859a",
443 => x"3fa00b8c",
444 => x"08940508",
445 => x"318c08ec",
446 => x"050c8c08",
447 => x"ec050880",
448 => x"249d3880",
449 => x"0b8c08f4",
450 => x"050c8c08",
451 => x"ec050830",
452 => x"8c08fc05",
453 => x"08712b8c",
454 => x"08f0050c",
455 => x"54b9398c",
456 => x"08fc0508",
457 => x"8c08ec05",
458 => x"082a8c08",
459 => x"e8050c8c",
460 => x"08fc0508",
461 => x"8c089405",
462 => x"082b8c08",
463 => x"f4050c8c",
464 => x"08f80508",
465 => x"8c089405",
466 => x"082b708c",
467 => x"08e80508",
468 => x"078c08f0",
469 => x"050c548c",
470 => x"08f00508",
471 => x"8c08f405",
472 => x"088c0888",
473 => x"05085856",
474 => x"5473760c",
475 => x"7484170c",
476 => x"8c088805",
477 => x"08800c8d",
478 => x"3d0d8c0c",
479 => x"048c0802",
480 => x"8c0cf93d",
481 => x"0d800b8c",
482 => x"08fc050c",
483 => x"8c088805",
484 => x"088025ab",
485 => x"388c0888",
486 => x"0508308c",
487 => x"0888050c",
488 => x"800b8c08",
489 => x"f4050c8c",
490 => x"08fc0508",
491 => x"8838810b",
492 => x"8c08f405",
493 => x"0c8c08f4",
494 => x"05088c08",
495 => x"fc050c8c",
496 => x"088c0508",
497 => x"8025ab38",
498 => x"8c088c05",
499 => x"08308c08",
500 => x"8c050c80",
501 => x"0b8c08f0",
502 => x"050c8c08",
503 => x"fc050888",
504 => x"38810b8c",
505 => x"08f0050c",
506 => x"8c08f005",
507 => x"088c08fc",
508 => x"050c8053",
509 => x"8c088c05",
510 => x"08528c08",
511 => x"88050851",
512 => x"81a73f80",
513 => x"08708c08",
514 => x"f8050c54",
515 => x"8c08fc05",
516 => x"08802e8c",
517 => x"388c08f8",
518 => x"0508308c",
519 => x"08f8050c",
520 => x"8c08f805",
521 => x"0870800c",
522 => x"54893d0d",
523 => x"8c0c048c",
524 => x"08028c0c",
525 => x"fb3d0d80",
526 => x"0b8c08fc",
527 => x"050c8c08",
528 => x"88050880",
529 => x"2593388c",
530 => x"08880508",
531 => x"308c0888",
532 => x"050c810b",
533 => x"8c08fc05",
534 => x"0c8c088c",
535 => x"05088025",
536 => x"8c388c08",
537 => x"8c050830",
538 => x"8c088c05",
539 => x"0c81538c",
540 => x"088c0508",
541 => x"528c0888",
542 => x"050851ad",
543 => x"3f800870",
544 => x"8c08f805",
545 => x"0c548c08",
546 => x"fc050880",
547 => x"2e8c388c",
548 => x"08f80508",
549 => x"308c08f8",
550 => x"050c8c08",
551 => x"f8050870",
552 => x"800c5487",
553 => x"3d0d8c0c",
554 => x"048c0802",
555 => x"8c0c7070",
556 => x"7070810b",
557 => x"8c08fc05",
558 => x"0c800b8c",
559 => x"08f8050c",
560 => x"8c088c05",
561 => x"088c0888",
562 => x"050827ac",
563 => x"388c08fc",
564 => x"0508802e",
565 => x"a338800b",
566 => x"8c088c05",
567 => x"08249938",
568 => x"8c088c05",
569 => x"08108c08",
570 => x"8c050c8c",
571 => x"08fc0508",
572 => x"108c08fc",
573 => x"050cc939",
574 => x"8c08fc05",
575 => x"08802e80",
576 => x"c9388c08",
577 => x"8c05088c",
578 => x"08880508",
579 => x"26a1388c",
580 => x"08880508",
581 => x"8c088c05",
582 => x"08318c08",
583 => x"88050c8c",
584 => x"08f80508",
585 => x"8c08fc05",
586 => x"08078c08",
587 => x"f8050c8c",
588 => x"08fc0508",
589 => x"812a8c08",
590 => x"fc050c8c",
591 => x"088c0508",
592 => x"812a8c08",
593 => x"8c050cff",
594 => x"af398c08",
595 => x"90050880",
596 => x"2e8f388c",
597 => x"08880508",
598 => x"708c08f4",
599 => x"050c518d",
600 => x"398c08f8",
601 => x"0508708c",
602 => x"08f4050c",
603 => x"518c08f4",
604 => x"0508800c",
605 => x"50505050",
606 => x"8c0c0470",
607 => x"865184ea",
608 => x"3f8151ba",
609 => x"d83ffc3d",
610 => x"0d767079",
611 => x"7b555555",
612 => x"558f7227",
613 => x"8c387275",
614 => x"07830651",
615 => x"70802ea7",
616 => x"38ff1252",
617 => x"71ff2e98",
618 => x"38727081",
619 => x"05543374",
620 => x"70810556",
621 => x"34ff1252",
622 => x"71ff2e09",
623 => x"8106ea38",
624 => x"74800c86",
625 => x"3d0d0474",
626 => x"51727084",
627 => x"05540871",
628 => x"70840553",
629 => x"0c727084",
630 => x"05540871",
631 => x"70840553",
632 => x"0c727084",
633 => x"05540871",
634 => x"70840553",
635 => x"0c727084",
636 => x"05540871",
637 => x"70840553",
638 => x"0cf01252",
639 => x"718f26c9",
640 => x"38837227",
641 => x"95387270",
642 => x"84055408",
643 => x"71708405",
644 => x"530cfc12",
645 => x"52718326",
646 => x"ed387054",
647 => x"ff8339f7",
648 => x"3d0d7c70",
649 => x"525384b8",
650 => x"3f725480",
651 => x"085580d6",
652 => x"c8568157",
653 => x"80088105",
654 => x"5a8b3de4",
655 => x"11595382",
656 => x"59f41352",
657 => x"7b881108",
658 => x"525384f5",
659 => x"3f800830",
660 => x"70800807",
661 => x"9f2c8a07",
662 => x"800c538b",
663 => x"3d0d0470",
664 => x"70735280",
665 => x"d6fc0851",
666 => x"ffb53f50",
667 => x"50047070",
668 => x"70707553",
669 => x"84d81308",
670 => x"802e8b38",
671 => x"80537280",
672 => x"0c505050",
673 => x"50048180",
674 => x"5272518a",
675 => x"9b3f8008",
676 => x"84d8140c",
677 => x"ff538008",
678 => x"802ee338",
679 => x"8008549f",
680 => x"53807470",
681 => x"8405560c",
682 => x"ff135380",
683 => x"7324cd38",
684 => x"80747084",
685 => x"05560cff",
686 => x"13537280",
687 => x"25e338ff",
688 => x"bb397070",
689 => x"70707577",
690 => x"55539f74",
691 => x"278e3896",
692 => x"730cff52",
693 => x"71800c50",
694 => x"50505004",
695 => x"84d81308",
696 => x"5271802e",
697 => x"94387310",
698 => x"10127008",
699 => x"79720c51",
700 => x"5271800c",
701 => x"50505050",
702 => x"047251fe",
703 => x"f13fff52",
704 => x"8008d138",
705 => x"84d81308",
706 => x"74101011",
707 => x"70087a72",
708 => x"0c515152",
709 => x"dc39f93d",
710 => x"0d797b58",
711 => x"56769f26",
712 => x"80e83884",
713 => x"d8160854",
714 => x"73802eaa",
715 => x"38761010",
716 => x"14700855",
717 => x"5573802e",
718 => x"ba388058",
719 => x"73812e8f",
720 => x"3873ff2e",
721 => x"a3388075",
722 => x"0c765173",
723 => x"2d805877",
724 => x"800c893d",
725 => x"0d047551",
726 => x"fe943fff",
727 => x"588008ef",
728 => x"3884d816",
729 => x"0854c639",
730 => x"96760c81",
731 => x"0b800c89",
732 => x"3d0d0475",
733 => x"5181e53f",
734 => x"76538008",
735 => x"52755181",
736 => x"a53f8008",
737 => x"800c893d",
738 => x"0d049676",
739 => x"0cff0b80",
740 => x"0c893d0d",
741 => x"04fc3d0d",
742 => x"76785653",
743 => x"ff54749f",
744 => x"26b13884",
745 => x"d8130852",
746 => x"71802eae",
747 => x"38741010",
748 => x"12700853",
749 => x"53815471",
750 => x"802e9838",
751 => x"825471ff",
752 => x"2e913883",
753 => x"5471812e",
754 => x"8a388073",
755 => x"0c745171",
756 => x"2d805473",
757 => x"800c863d",
758 => x"0d047251",
759 => x"fd903f80",
760 => x"08f13884",
761 => x"d8130852",
762 => x"c4397070",
763 => x"735280d6",
764 => x"fc0851fe",
765 => x"a13f5050",
766 => x"04707070",
767 => x"75537452",
768 => x"80d6fc08",
769 => x"51fdbb3f",
770 => x"50505004",
771 => x"7080d6fc",
772 => x"0851fcda",
773 => x"3f500470",
774 => x"70735280",
775 => x"d6fc0851",
776 => x"fef33f50",
777 => x"5004fc3d",
778 => x"0d800b80",
779 => x"e7800c78",
780 => x"527751b4",
781 => x"9b3f8008",
782 => x"548008ff",
783 => x"2e883873",
784 => x"800c863d",
785 => x"0d0480e7",
786 => x"80085574",
787 => x"802ef038",
788 => x"7675710c",
789 => x"5373800c",
790 => x"863d0d04",
791 => x"b3ed3f04",
792 => x"70707070",
793 => x"75707183",
794 => x"06535552",
795 => x"70b83871",
796 => x"70087009",
797 => x"f7fbfdff",
798 => x"120670f8",
799 => x"84828180",
800 => x"06515152",
801 => x"53709d38",
802 => x"84137008",
803 => x"7009f7fb",
804 => x"fdff1206",
805 => x"70f88482",
806 => x"81800651",
807 => x"51525370",
808 => x"802ee538",
809 => x"72527133",
810 => x"5170802e",
811 => x"8a388112",
812 => x"70335252",
813 => x"70f83871",
814 => x"7431800c",
815 => x"50505050",
816 => x"04f23d0d",
817 => x"60628811",
818 => x"08705757",
819 => x"5f5a7480",
820 => x"2e819038",
821 => x"8c1a2270",
822 => x"832a8132",
823 => x"70810651",
824 => x"55587386",
825 => x"38901a08",
826 => x"91387951",
827 => x"9cd03fff",
828 => x"54800880",
829 => x"ee388c1a",
830 => x"22587d08",
831 => x"57807883",
832 => x"ffff0670",
833 => x"0a100a70",
834 => x"81065156",
835 => x"57557375",
836 => x"2e80d738",
837 => x"74903876",
838 => x"08841808",
839 => x"88195956",
840 => x"5974802e",
841 => x"f2387454",
842 => x"88807527",
843 => x"84388880",
844 => x"54735378",
845 => x"529c1a08",
846 => x"51a41a08",
847 => x"54732d80",
848 => x"0b800825",
849 => x"82e63880",
850 => x"08197580",
851 => x"08317f88",
852 => x"05088008",
853 => x"31706188",
854 => x"050c5656",
855 => x"5973ffb4",
856 => x"38805473",
857 => x"800c903d",
858 => x"0d047581",
859 => x"32708106",
860 => x"76415154",
861 => x"73802e81",
862 => x"c1387490",
863 => x"38760884",
864 => x"18088819",
865 => x"59565974",
866 => x"802ef238",
867 => x"881a0878",
868 => x"83ffff06",
869 => x"70892a70",
870 => x"81065156",
871 => x"59567380",
872 => x"2e82fa38",
873 => x"7575278d",
874 => x"3877872a",
875 => x"70810651",
876 => x"547382b5",
877 => x"38747627",
878 => x"83387456",
879 => x"75537852",
880 => x"79085190",
881 => x"f83f881a",
882 => x"08763188",
883 => x"1b0c7908",
884 => x"167a0c74",
885 => x"56751975",
886 => x"77317f88",
887 => x"05087831",
888 => x"70618805",
889 => x"0c565659",
890 => x"73802efe",
891 => x"f4388c1a",
892 => x"2258ff86",
893 => x"39777854",
894 => x"79537b52",
895 => x"5690be3f",
896 => x"881a0878",
897 => x"31881b0c",
898 => x"7908187a",
899 => x"0c7c7631",
900 => x"5d7c8e38",
901 => x"79519c8a",
902 => x"3f800881",
903 => x"8f388008",
904 => x"5f751975",
905 => x"77317f88",
906 => x"05087831",
907 => x"70618805",
908 => x"0c565659",
909 => x"73802efe",
910 => x"a8387481",
911 => x"83387608",
912 => x"84180888",
913 => x"19595659",
914 => x"74802ef2",
915 => x"3874538a",
916 => x"5278518e",
917 => x"c93f8008",
918 => x"79318105",
919 => x"5d800884",
920 => x"3881155d",
921 => x"815f7c58",
922 => x"747d2783",
923 => x"38745894",
924 => x"1a08881b",
925 => x"0811575c",
926 => x"807a085c",
927 => x"54901a08",
928 => x"7b278338",
929 => x"81547578",
930 => x"25843873",
931 => x"ba387b78",
932 => x"24fee238",
933 => x"7b537852",
934 => x"9c1a0851",
935 => x"a41a0854",
936 => x"732d8008",
937 => x"56800880",
938 => x"24fee238",
939 => x"8c1a2280",
940 => x"c0075473",
941 => x"8c1b23ff",
942 => x"5473800c",
943 => x"903d0d04",
944 => x"7effa338",
945 => x"ff873975",
946 => x"5378527a",
947 => x"518eee3f",
948 => x"7908167a",
949 => x"0c79519a",
950 => x"c93f8008",
951 => x"cf387c76",
952 => x"315d7cfe",
953 => x"bc38feac",
954 => x"39901a08",
955 => x"7a087131",
956 => x"76117056",
957 => x"5a575280",
958 => x"d6fc0851",
959 => x"90843f80",
960 => x"08802eff",
961 => x"a7388008",
962 => x"901b0c80",
963 => x"08167a0c",
964 => x"77941b0c",
965 => x"74881b0c",
966 => x"7456fd99",
967 => x"39790858",
968 => x"901a0878",
969 => x"27833881",
970 => x"54757527",
971 => x"843873b3",
972 => x"38941a08",
973 => x"56757526",
974 => x"80d33875",
975 => x"5378529c",
976 => x"1a0851a4",
977 => x"1a085473",
978 => x"2d800856",
979 => x"80088024",
980 => x"fd83388c",
981 => x"1a2280c0",
982 => x"0754738c",
983 => x"1b23ff54",
984 => x"fed73975",
985 => x"53785277",
986 => x"518dd23f",
987 => x"7908167a",
988 => x"0c795199",
989 => x"ad3f8008",
990 => x"802efcd9",
991 => x"388c1a22",
992 => x"80c00754",
993 => x"738c1b23",
994 => x"ff54fead",
995 => x"39747554",
996 => x"79537852",
997 => x"568da63f",
998 => x"881a0875",
999 => x"31881b0c",
1000 => x"7908157a",
1001 => x"0cfcae39",
1002 => x"f33d0d7f",
1003 => x"618b1170",
1004 => x"f8065c55",
1005 => x"555e7296",
1006 => x"26833890",
1007 => x"59807924",
1008 => x"747a2607",
1009 => x"53805472",
1010 => x"742e0981",
1011 => x"0680cb38",
1012 => x"7d518eac",
1013 => x"3f7883f7",
1014 => x"2680c638",
1015 => x"78832a70",
1016 => x"10101080",
1017 => x"deb8058c",
1018 => x"11085959",
1019 => x"5a76782e",
1020 => x"83b03884",
1021 => x"1708fc06",
1022 => x"568c1708",
1023 => x"88180871",
1024 => x"8c120c88",
1025 => x"120c5875",
1026 => x"17841108",
1027 => x"81078412",
1028 => x"0c537d51",
1029 => x"8deb3f88",
1030 => x"17547380",
1031 => x"0c8f3d0d",
1032 => x"0478892a",
1033 => x"79832a5b",
1034 => x"5372802e",
1035 => x"bf387886",
1036 => x"2ab8055a",
1037 => x"847327b4",
1038 => x"3880db13",
1039 => x"5a947327",
1040 => x"ab38788c",
1041 => x"2a80ee05",
1042 => x"5a80d473",
1043 => x"279e3878",
1044 => x"8f2a80f7",
1045 => x"055a82d4",
1046 => x"73279138",
1047 => x"78922a80",
1048 => x"fc055a8a",
1049 => x"d4732784",
1050 => x"3880fe5a",
1051 => x"79101010",
1052 => x"80deb805",
1053 => x"8c110858",
1054 => x"5576752e",
1055 => x"a3388417",
1056 => x"08fc0670",
1057 => x"7a315556",
1058 => x"738f2488",
1059 => x"d5387380",
1060 => x"25fee638",
1061 => x"8c170857",
1062 => x"76752e09",
1063 => x"8106df38",
1064 => x"811a5a80",
1065 => x"dec80857",
1066 => x"7680dec0",
1067 => x"2e82c038",
1068 => x"841708fc",
1069 => x"06707a31",
1070 => x"5556738f",
1071 => x"2481f938",
1072 => x"80dec00b",
1073 => x"80decc0c",
1074 => x"80dec00b",
1075 => x"80dec80c",
1076 => x"738025fe",
1077 => x"b23883ff",
1078 => x"762783df",
1079 => x"3875892a",
1080 => x"76832a55",
1081 => x"5372802e",
1082 => x"bf387586",
1083 => x"2ab80554",
1084 => x"847327b4",
1085 => x"3880db13",
1086 => x"54947327",
1087 => x"ab38758c",
1088 => x"2a80ee05",
1089 => x"5480d473",
1090 => x"279e3875",
1091 => x"8f2a80f7",
1092 => x"055482d4",
1093 => x"73279138",
1094 => x"75922a80",
1095 => x"fc05548a",
1096 => x"d4732784",
1097 => x"3880fe54",
1098 => x"73101010",
1099 => x"80deb805",
1100 => x"88110856",
1101 => x"5874782e",
1102 => x"86cf3884",
1103 => x"1508fc06",
1104 => x"53757327",
1105 => x"8d388815",
1106 => x"08557478",
1107 => x"2e098106",
1108 => x"ea388c15",
1109 => x"0880deb8",
1110 => x"0b840508",
1111 => x"718c1a0c",
1112 => x"76881a0c",
1113 => x"7888130c",
1114 => x"788c180c",
1115 => x"5d587953",
1116 => x"807a2483",
1117 => x"e6387282",
1118 => x"2c81712b",
1119 => x"5c537a7c",
1120 => x"26819838",
1121 => x"7b7b0653",
1122 => x"7282f138",
1123 => x"79fc0684",
1124 => x"055a7a10",
1125 => x"707d0654",
1126 => x"5b7282e0",
1127 => x"38841a5a",
1128 => x"f1398817",
1129 => x"8c110858",
1130 => x"5876782e",
1131 => x"098106fc",
1132 => x"c238821a",
1133 => x"5afdec39",
1134 => x"78177981",
1135 => x"0784190c",
1136 => x"7080decc",
1137 => x"0c7080de",
1138 => x"c80c80de",
1139 => x"c00b8c12",
1140 => x"0c8c1108",
1141 => x"88120c74",
1142 => x"81078412",
1143 => x"0c741175",
1144 => x"710c5153",
1145 => x"7d518a99",
1146 => x"3f881754",
1147 => x"fcac3980",
1148 => x"deb80b84",
1149 => x"05087a54",
1150 => x"5c798025",
1151 => x"fef83882",
1152 => x"da397a09",
1153 => x"7c067080",
1154 => x"deb80b84",
1155 => x"050c5c7a",
1156 => x"105b7a7c",
1157 => x"2685387a",
1158 => x"85b83880",
1159 => x"deb80b88",
1160 => x"05087084",
1161 => x"1208fc06",
1162 => x"707c317c",
1163 => x"72268f72",
1164 => x"25075757",
1165 => x"5c5d5572",
1166 => x"802e80db",
1167 => x"38797a16",
1168 => x"80deb008",
1169 => x"1b90115a",
1170 => x"55575b80",
1171 => x"deac08ff",
1172 => x"2e8838a0",
1173 => x"8f13e080",
1174 => x"06577652",
1175 => x"7d5191a7",
1176 => x"3f800854",
1177 => x"8008ff2e",
1178 => x"90388008",
1179 => x"76278299",
1180 => x"387480de",
1181 => x"b82e8291",
1182 => x"3880deb8",
1183 => x"0b880508",
1184 => x"55841508",
1185 => x"fc06707a",
1186 => x"317a7226",
1187 => x"8f722507",
1188 => x"52555372",
1189 => x"83e63874",
1190 => x"79810784",
1191 => x"170c7916",
1192 => x"7080deb8",
1193 => x"0b88050c",
1194 => x"75810784",
1195 => x"120c547e",
1196 => x"525788cd",
1197 => x"3f881754",
1198 => x"fae03975",
1199 => x"832a7054",
1200 => x"54807424",
1201 => x"819b3872",
1202 => x"822c8171",
1203 => x"2b80debc",
1204 => x"08077080",
1205 => x"deb80b84",
1206 => x"050c7510",
1207 => x"101080de",
1208 => x"b8058811",
1209 => x"08585a5d",
1210 => x"53778c18",
1211 => x"0c748818",
1212 => x"0c768819",
1213 => x"0c768c16",
1214 => x"0cfcf339",
1215 => x"797a1010",
1216 => x"1080deb8",
1217 => x"05705759",
1218 => x"5d8c1508",
1219 => x"5776752e",
1220 => x"a3388417",
1221 => x"08fc0670",
1222 => x"7a315556",
1223 => x"738f2483",
1224 => x"ca387380",
1225 => x"25848138",
1226 => x"8c170857",
1227 => x"76752e09",
1228 => x"8106df38",
1229 => x"8815811b",
1230 => x"70830655",
1231 => x"5b5572c9",
1232 => x"387c8306",
1233 => x"5372802e",
1234 => x"fdb838ff",
1235 => x"1df81959",
1236 => x"5d881808",
1237 => x"782eea38",
1238 => x"fdb53983",
1239 => x"1a53fc96",
1240 => x"39831470",
1241 => x"822c8171",
1242 => x"2b80debc",
1243 => x"08077080",
1244 => x"deb80b84",
1245 => x"050c7610",
1246 => x"101080de",
1247 => x"b8058811",
1248 => x"08595b5e",
1249 => x"5153fee1",
1250 => x"3980ddfc",
1251 => x"08175880",
1252 => x"08762e81",
1253 => x"8d3880de",
1254 => x"ac08ff2e",
1255 => x"83ec3873",
1256 => x"76311880",
1257 => x"ddfc0c73",
1258 => x"87067057",
1259 => x"5372802e",
1260 => x"88388873",
1261 => x"31701555",
1262 => x"5676149f",
1263 => x"ff06a080",
1264 => x"71311770",
1265 => x"547f5357",
1266 => x"538ebc3f",
1267 => x"80085380",
1268 => x"08ff2e81",
1269 => x"a03880dd",
1270 => x"fc081670",
1271 => x"80ddfc0c",
1272 => x"747580de",
1273 => x"b80b8805",
1274 => x"0c747631",
1275 => x"18708107",
1276 => x"51555658",
1277 => x"7b80deb8",
1278 => x"2e839c38",
1279 => x"798f2682",
1280 => x"cb38810b",
1281 => x"84150c84",
1282 => x"1508fc06",
1283 => x"707a317a",
1284 => x"72268f72",
1285 => x"25075255",
1286 => x"5372802e",
1287 => x"fcf93880",
1288 => x"db398008",
1289 => x"9fff0653",
1290 => x"72feeb38",
1291 => x"7780ddfc",
1292 => x"0c80deb8",
1293 => x"0b880508",
1294 => x"7b188107",
1295 => x"84120c55",
1296 => x"80dea808",
1297 => x"78278638",
1298 => x"7780dea8",
1299 => x"0c80dea4",
1300 => x"087827fc",
1301 => x"ac387780",
1302 => x"dea40c84",
1303 => x"1508fc06",
1304 => x"707a317a",
1305 => x"72268f72",
1306 => x"25075255",
1307 => x"5372802e",
1308 => x"fca53888",
1309 => x"39807454",
1310 => x"56fedb39",
1311 => x"7d518581",
1312 => x"3f800b80",
1313 => x"0c8f3d0d",
1314 => x"04735380",
1315 => x"7424a938",
1316 => x"72822c81",
1317 => x"712b80de",
1318 => x"bc080770",
1319 => x"80deb80b",
1320 => x"84050c5d",
1321 => x"53778c18",
1322 => x"0c748818",
1323 => x"0c768819",
1324 => x"0c768c16",
1325 => x"0cf9b739",
1326 => x"83147082",
1327 => x"2c81712b",
1328 => x"80debc08",
1329 => x"077080de",
1330 => x"b80b8405",
1331 => x"0c5e5153",
1332 => x"d4397b7b",
1333 => x"065372fc",
1334 => x"a338841a",
1335 => x"7b105c5a",
1336 => x"f139ff1a",
1337 => x"8111515a",
1338 => x"f7b93978",
1339 => x"17798107",
1340 => x"84190c8c",
1341 => x"18088819",
1342 => x"08718c12",
1343 => x"0c88120c",
1344 => x"597080de",
1345 => x"cc0c7080",
1346 => x"dec80c80",
1347 => x"dec00b8c",
1348 => x"120c8c11",
1349 => x"0888120c",
1350 => x"74810784",
1351 => x"120c7411",
1352 => x"75710c51",
1353 => x"53f9bd39",
1354 => x"75178411",
1355 => x"08810784",
1356 => x"120c538c",
1357 => x"17088818",
1358 => x"08718c12",
1359 => x"0c88120c",
1360 => x"587d5183",
1361 => x"bc3f8817",
1362 => x"54f5cf39",
1363 => x"7284150c",
1364 => x"f41af806",
1365 => x"70841e08",
1366 => x"81060784",
1367 => x"1e0c701d",
1368 => x"545b850b",
1369 => x"84140c85",
1370 => x"0b88140c",
1371 => x"8f7b27fd",
1372 => x"cf38881c",
1373 => x"527d5193",
1374 => x"e73f80de",
1375 => x"b80b8805",
1376 => x"0880ddfc",
1377 => x"085955fd",
1378 => x"b7397780",
1379 => x"ddfc0c73",
1380 => x"80deac0c",
1381 => x"fc913972",
1382 => x"84150cfd",
1383 => x"a339fa3d",
1384 => x"0d7a7902",
1385 => x"8805a705",
1386 => x"33565253",
1387 => x"8373278a",
1388 => x"38708306",
1389 => x"5271802e",
1390 => x"a838ff13",
1391 => x"5372ff2e",
1392 => x"97387033",
1393 => x"5273722e",
1394 => x"91388111",
1395 => x"ff145451",
1396 => x"72ff2e09",
1397 => x"8106eb38",
1398 => x"80517080",
1399 => x"0c883d0d",
1400 => x"04707257",
1401 => x"55835175",
1402 => x"82802914",
1403 => x"ff125256",
1404 => x"708025f3",
1405 => x"38837327",
1406 => x"bf387408",
1407 => x"76327009",
1408 => x"f7fbfdff",
1409 => x"120670f8",
1410 => x"84828180",
1411 => x"06515151",
1412 => x"70802e99",
1413 => x"38745180",
1414 => x"52703357",
1415 => x"73772eff",
1416 => x"b9388111",
1417 => x"81135351",
1418 => x"837227ed",
1419 => x"38fc1384",
1420 => x"16565372",
1421 => x"8326c338",
1422 => x"7451fefe",
1423 => x"39fa3d0d",
1424 => x"787a7c72",
1425 => x"72725757",
1426 => x"57595656",
1427 => x"747627b2",
1428 => x"38761551",
1429 => x"757127aa",
1430 => x"38707717",
1431 => x"ff145455",
1432 => x"5371ff2e",
1433 => x"9638ff14",
1434 => x"ff145454",
1435 => x"72337434",
1436 => x"ff125271",
1437 => x"ff2e0981",
1438 => x"06ec3875",
1439 => x"800c883d",
1440 => x"0d04768f",
1441 => x"269738ff",
1442 => x"125271ff",
1443 => x"2eed3872",
1444 => x"70810554",
1445 => x"33747081",
1446 => x"055634eb",
1447 => x"39747607",
1448 => x"83065170",
1449 => x"e2387575",
1450 => x"54517270",
1451 => x"84055408",
1452 => x"71708405",
1453 => x"530c7270",
1454 => x"84055408",
1455 => x"71708405",
1456 => x"530c7270",
1457 => x"84055408",
1458 => x"71708405",
1459 => x"530c7270",
1460 => x"84055408",
1461 => x"71708405",
1462 => x"530cf012",
1463 => x"52718f26",
1464 => x"c9388372",
1465 => x"27953872",
1466 => x"70840554",
1467 => x"08717084",
1468 => x"05530cfc",
1469 => x"12527183",
1470 => x"26ed3870",
1471 => x"54ff8839",
1472 => x"0404ef3d",
1473 => x"0d636567",
1474 => x"405d427b",
1475 => x"802e84f9",
1476 => x"386151ec",
1477 => x"3ff81c70",
1478 => x"84120870",
1479 => x"fc067062",
1480 => x"8b0570f8",
1481 => x"06415945",
1482 => x"5b5c4157",
1483 => x"96742782",
1484 => x"c338807b",
1485 => x"247e7c26",
1486 => x"07598054",
1487 => x"78742e09",
1488 => x"810682a9",
1489 => x"38777b25",
1490 => x"81fc3877",
1491 => x"1780deb8",
1492 => x"0b880508",
1493 => x"5e567c76",
1494 => x"2e84bd38",
1495 => x"84160870",
1496 => x"fe061784",
1497 => x"11088106",
1498 => x"51555573",
1499 => x"828b3874",
1500 => x"fc06597c",
1501 => x"762e84dd",
1502 => x"3877195f",
1503 => x"7e7b2581",
1504 => x"fd387981",
1505 => x"06547382",
1506 => x"bf387677",
1507 => x"08318411",
1508 => x"08fc0656",
1509 => x"5a75802e",
1510 => x"91387c76",
1511 => x"2e84ea38",
1512 => x"74191859",
1513 => x"787b2584",
1514 => x"89387980",
1515 => x"2e829938",
1516 => x"7715567a",
1517 => x"76248290",
1518 => x"388c1a08",
1519 => x"881b0871",
1520 => x"8c120c88",
1521 => x"120c5579",
1522 => x"76595788",
1523 => x"1761fc05",
1524 => x"575975a4",
1525 => x"2685ef38",
1526 => x"7b795555",
1527 => x"93762780",
1528 => x"c9387b70",
1529 => x"84055d08",
1530 => x"7c56790c",
1531 => x"74708405",
1532 => x"56088c18",
1533 => x"0c901754",
1534 => x"9b7627ae",
1535 => x"38747084",
1536 => x"05560874",
1537 => x"0c747084",
1538 => x"05560894",
1539 => x"180c9817",
1540 => x"54a37627",
1541 => x"95387470",
1542 => x"84055608",
1543 => x"740c7470",
1544 => x"84055608",
1545 => x"9c180ca0",
1546 => x"17547470",
1547 => x"84055608",
1548 => x"74708405",
1549 => x"560c7470",
1550 => x"84055608",
1551 => x"74708405",
1552 => x"560c7408",
1553 => x"740c777b",
1554 => x"3156758f",
1555 => x"2680c938",
1556 => x"84170881",
1557 => x"06780784",
1558 => x"180c7717",
1559 => x"84110881",
1560 => x"0784120c",
1561 => x"546151fd",
1562 => x"983f8817",
1563 => x"5473800c",
1564 => x"933d0d04",
1565 => x"905bfdba",
1566 => x"397856fe",
1567 => x"85398c16",
1568 => x"08881708",
1569 => x"718c120c",
1570 => x"88120c55",
1571 => x"7e707c31",
1572 => x"57588f76",
1573 => x"27ffb938",
1574 => x"7a178418",
1575 => x"0881067c",
1576 => x"0784190c",
1577 => x"76810784",
1578 => x"120c7611",
1579 => x"84110881",
1580 => x"0784120c",
1581 => x"55880552",
1582 => x"61518da4",
1583 => x"3f6151fc",
1584 => x"c03f8817",
1585 => x"54ffa639",
1586 => x"7d526151",
1587 => x"edda3f80",
1588 => x"08598008",
1589 => x"802e81a3",
1590 => x"388008f8",
1591 => x"05608405",
1592 => x"08fe0661",
1593 => x"05555776",
1594 => x"742e83e6",
1595 => x"38fc1856",
1596 => x"75a42681",
1597 => x"aa387b80",
1598 => x"08555593",
1599 => x"762780d8",
1600 => x"38747084",
1601 => x"05560880",
1602 => x"08708405",
1603 => x"800c0c80",
1604 => x"08757084",
1605 => x"05570871",
1606 => x"70840553",
1607 => x"0c549b76",
1608 => x"27b63874",
1609 => x"70840556",
1610 => x"08747084",
1611 => x"05560c74",
1612 => x"70840556",
1613 => x"08747084",
1614 => x"05560ca3",
1615 => x"76279938",
1616 => x"74708405",
1617 => x"56087470",
1618 => x"8405560c",
1619 => x"74708405",
1620 => x"56087470",
1621 => x"8405560c",
1622 => x"74708405",
1623 => x"56087470",
1624 => x"8405560c",
1625 => x"74708405",
1626 => x"56087470",
1627 => x"8405560c",
1628 => x"7408740c",
1629 => x"7b526151",
1630 => x"8be63f61",
1631 => x"51fb823f",
1632 => x"78547380",
1633 => x"0c933d0d",
1634 => x"047d5261",
1635 => x"51ec993f",
1636 => x"8008800c",
1637 => x"933d0d04",
1638 => x"84160855",
1639 => x"fbd13975",
1640 => x"537b5280",
1641 => x"0851dfde",
1642 => x"3f7b5261",
1643 => x"518bb13f",
1644 => x"ca398c16",
1645 => x"08881708",
1646 => x"718c120c",
1647 => x"88120c55",
1648 => x"8c1a0888",
1649 => x"1b08718c",
1650 => x"120c8812",
1651 => x"0c557979",
1652 => x"5957fbf7",
1653 => x"39771990",
1654 => x"1c555573",
1655 => x"7524fba2",
1656 => x"387a1770",
1657 => x"80deb80b",
1658 => x"88050c75",
1659 => x"7c318107",
1660 => x"84120c5d",
1661 => x"84170881",
1662 => x"067b0784",
1663 => x"180c6151",
1664 => x"f9ff3f88",
1665 => x"1754fce5",
1666 => x"39741918",
1667 => x"901c555d",
1668 => x"737d24fb",
1669 => x"95388c1a",
1670 => x"08881b08",
1671 => x"718c120c",
1672 => x"88120c55",
1673 => x"881a61fc",
1674 => x"05575975",
1675 => x"a42681ae",
1676 => x"387b7955",
1677 => x"55937627",
1678 => x"80c9387b",
1679 => x"7084055d",
1680 => x"087c5679",
1681 => x"0c747084",
1682 => x"0556088c",
1683 => x"1b0c901a",
1684 => x"549b7627",
1685 => x"ae387470",
1686 => x"84055608",
1687 => x"740c7470",
1688 => x"84055608",
1689 => x"941b0c98",
1690 => x"1a54a376",
1691 => x"27953874",
1692 => x"70840556",
1693 => x"08740c74",
1694 => x"70840556",
1695 => x"089c1b0c",
1696 => x"a01a5474",
1697 => x"70840556",
1698 => x"08747084",
1699 => x"05560c74",
1700 => x"70840556",
1701 => x"08747084",
1702 => x"05560c74",
1703 => x"08740c7a",
1704 => x"1a7080de",
1705 => x"b80b8805",
1706 => x"0c7d7c31",
1707 => x"81078412",
1708 => x"0c54841a",
1709 => x"0881067b",
1710 => x"07841b0c",
1711 => x"6151f8c1",
1712 => x"3f7854fd",
1713 => x"bd397553",
1714 => x"7b527851",
1715 => x"ddb83ffa",
1716 => x"f5398417",
1717 => x"08fc0618",
1718 => x"605858fa",
1719 => x"e9397553",
1720 => x"7b527851",
1721 => x"dda03f7a",
1722 => x"1a7080de",
1723 => x"b80b8805",
1724 => x"0c7d7c31",
1725 => x"81078412",
1726 => x"0c54841a",
1727 => x"0881067b",
1728 => x"07841b0c",
1729 => x"ffb63970",
1730 => x"70707080",
1731 => x"0b80e780",
1732 => x"0c765196",
1733 => x"cc3f8008",
1734 => x"538008ff",
1735 => x"2e893872",
1736 => x"800c5050",
1737 => x"50500480",
1738 => x"e7800854",
1739 => x"73802eef",
1740 => x"38757471",
1741 => x"0c527280",
1742 => x"0c505050",
1743 => x"5004fa3d",
1744 => x"0d7880d6",
1745 => x"fc085455",
1746 => x"b8130880",
1747 => x"2e81b638",
1748 => x"8c152270",
1749 => x"83ffff06",
1750 => x"70832a81",
1751 => x"32708106",
1752 => x"51555556",
1753 => x"72802e80",
1754 => x"dc387384",
1755 => x"2a813281",
1756 => x"0657ff53",
1757 => x"7680f738",
1758 => x"73822a70",
1759 => x"81065153",
1760 => x"72802eb9",
1761 => x"38b01508",
1762 => x"5473802e",
1763 => x"9c3880c0",
1764 => x"15537373",
1765 => x"2e8f3873",
1766 => x"5280d6fc",
1767 => x"085187c0",
1768 => x"3f8c1522",
1769 => x"5676b016",
1770 => x"0c75db06",
1771 => x"53728c16",
1772 => x"23800b84",
1773 => x"160c9015",
1774 => x"08750c72",
1775 => x"56758807",
1776 => x"53728c16",
1777 => x"23901508",
1778 => x"802e80c1",
1779 => x"388c1522",
1780 => x"70810655",
1781 => x"53739e38",
1782 => x"720a100a",
1783 => x"70810651",
1784 => x"53728538",
1785 => x"94150854",
1786 => x"7388160c",
1787 => x"80537280",
1788 => x"0c883d0d",
1789 => x"04800b88",
1790 => x"160c9415",
1791 => x"08309816",
1792 => x"0c8053ea",
1793 => x"39725182",
1794 => x"f73ffec4",
1795 => x"3974518c",
1796 => x"de3f8c15",
1797 => x"22708106",
1798 => x"55537380",
1799 => x"2effb938",
1800 => x"d439f83d",
1801 => x"0d7a5877",
1802 => x"802e8199",
1803 => x"3880d6fc",
1804 => x"0854b814",
1805 => x"08802e80",
1806 => x"ed388c18",
1807 => x"2270902b",
1808 => x"70902c70",
1809 => x"832a8132",
1810 => x"81065c51",
1811 => x"57547880",
1812 => x"cd389018",
1813 => x"08577680",
1814 => x"2e80c338",
1815 => x"77087731",
1816 => x"77790c76",
1817 => x"83067a58",
1818 => x"55557385",
1819 => x"38941808",
1820 => x"56758819",
1821 => x"0c807525",
1822 => x"a5387453",
1823 => x"76529c18",
1824 => x"0851a418",
1825 => x"0854732d",
1826 => x"800b8008",
1827 => x"2580c938",
1828 => x"80081775",
1829 => x"80083156",
1830 => x"57748024",
1831 => x"dd38800b",
1832 => x"800c8a3d",
1833 => x"0d047351",
1834 => x"81d63f8c",
1835 => x"18227090",
1836 => x"2b70902c",
1837 => x"70832a81",
1838 => x"3281065c",
1839 => x"51575478",
1840 => x"dd38ff8e",
1841 => x"39b8a252",
1842 => x"80d6fc08",
1843 => x"5189e73f",
1844 => x"8008800c",
1845 => x"8a3d0d04",
1846 => x"8c182280",
1847 => x"c0075473",
1848 => x"8c1923ff",
1849 => x"0b800c8a",
1850 => x"3d0d0470",
1851 => x"72518071",
1852 => x"0c800b84",
1853 => x"120c800b",
1854 => x"88120c02",
1855 => x"8e05228c",
1856 => x"12230292",
1857 => x"05228e12",
1858 => x"23800b90",
1859 => x"120c800b",
1860 => x"94120c80",
1861 => x"0b98120c",
1862 => x"709c120c",
1863 => x"80c8810b",
1864 => x"a0120c80",
1865 => x"c8cd0ba4",
1866 => x"120c80c9",
1867 => x"c90ba812",
1868 => x"0c80ca9a",
1869 => x"0bac120c",
1870 => x"5004fa3d",
1871 => x"0d797080",
1872 => x"dc298c11",
1873 => x"547a5356",
1874 => x"57e4dd3f",
1875 => x"80088008",
1876 => x"55568008",
1877 => x"802ea238",
1878 => x"80088c05",
1879 => x"54800b80",
1880 => x"080c7680",
1881 => x"0884050c",
1882 => x"73800888",
1883 => x"050c7453",
1884 => x"80527351",
1885 => x"8bfc3f75",
1886 => x"5473800c",
1887 => x"883d0d04",
1888 => x"fc3d0d76",
1889 => x"bd930bbc",
1890 => x"120c5581",
1891 => x"0bb8160c",
1892 => x"800b84dc",
1893 => x"160c830b",
1894 => x"84e0160c",
1895 => x"84e81584",
1896 => x"e4160c74",
1897 => x"54805384",
1898 => x"52841508",
1899 => x"51febc3f",
1900 => x"74548153",
1901 => x"89528815",
1902 => x"0851feaf",
1903 => x"3f745482",
1904 => x"538a528c",
1905 => x"150851fe",
1906 => x"a23f863d",
1907 => x"0d04f93d",
1908 => x"0d7980d6",
1909 => x"fc085457",
1910 => x"b8130880",
1911 => x"2e80c838",
1912 => x"84dc1356",
1913 => x"88160884",
1914 => x"1708ff05",
1915 => x"55558074",
1916 => x"249f388c",
1917 => x"15227090",
1918 => x"2b70902c",
1919 => x"51545872",
1920 => x"802e80ca",
1921 => x"3880dc15",
1922 => x"ff155555",
1923 => x"738025e3",
1924 => x"38750853",
1925 => x"72802e9f",
1926 => x"38725688",
1927 => x"16088417",
1928 => x"08ff0555",
1929 => x"55c83972",
1930 => x"51fed53f",
1931 => x"80d6fc08",
1932 => x"84dc0556",
1933 => x"ffae3984",
1934 => x"527651fd",
1935 => x"fd3f8008",
1936 => x"760c8008",
1937 => x"802e80c0",
1938 => x"38800856",
1939 => x"ce39810b",
1940 => x"8c162372",
1941 => x"750c7288",
1942 => x"160c7284",
1943 => x"160c7290",
1944 => x"160c7294",
1945 => x"160c7298",
1946 => x"160cff0b",
1947 => x"8e162372",
1948 => x"b0160c72",
1949 => x"b4160c72",
1950 => x"80c4160c",
1951 => x"7280c816",
1952 => x"0c74800c",
1953 => x"893d0d04",
1954 => x"8c770c80",
1955 => x"0b800c89",
1956 => x"3d0d0470",
1957 => x"70b8a252",
1958 => x"7351869a",
1959 => x"3f505004",
1960 => x"7080d6fc",
1961 => x"0851ec3f",
1962 => x"5004fb3d",
1963 => x"0d777052",
1964 => x"56f0cd3f",
1965 => x"80deb80b",
1966 => x"88050884",
1967 => x"1108fc06",
1968 => x"707b319f",
1969 => x"ef05e080",
1970 => x"06e08005",
1971 => x"565653a0",
1972 => x"80742494",
1973 => x"38805275",
1974 => x"51f8ac3f",
1975 => x"80dec008",
1976 => x"15537280",
1977 => x"082e8f38",
1978 => x"7551f095",
1979 => x"3f805372",
1980 => x"800c873d",
1981 => x"0d047330",
1982 => x"527551f8",
1983 => x"8a3f8008",
1984 => x"ff2ea838",
1985 => x"80deb80b",
1986 => x"88050875",
1987 => x"75318107",
1988 => x"84120c53",
1989 => x"80ddfc08",
1990 => x"743180dd",
1991 => x"fc0c7551",
1992 => x"efdf3f81",
1993 => x"0b800c87",
1994 => x"3d0d0480",
1995 => x"527551f7",
1996 => x"d63f80de",
1997 => x"b80b8805",
1998 => x"08800871",
1999 => x"3156538f",
2000 => x"7525ffa4",
2001 => x"38800880",
2002 => x"deac0831",
2003 => x"80ddfc0c",
2004 => x"74810784",
2005 => x"140c7551",
2006 => x"efa73f80",
2007 => x"53ff9039",
2008 => x"f63d0d7c",
2009 => x"7e545b72",
2010 => x"802e8283",
2011 => x"387a51ef",
2012 => x"8f3ff813",
2013 => x"84110870",
2014 => x"fe067013",
2015 => x"841108fc",
2016 => x"065d5859",
2017 => x"545880de",
2018 => x"c008752e",
2019 => x"82de3878",
2020 => x"84160c80",
2021 => x"73810654",
2022 => x"5a727a2e",
2023 => x"81d53878",
2024 => x"15841108",
2025 => x"81065153",
2026 => x"72a03878",
2027 => x"17577981",
2028 => x"e6388815",
2029 => x"08537280",
2030 => x"dec02e82",
2031 => x"f9388c15",
2032 => x"08708c15",
2033 => x"0c738812",
2034 => x"0c567681",
2035 => x"0784190c",
2036 => x"76187771",
2037 => x"0c537981",
2038 => x"913883ff",
2039 => x"772781c8",
2040 => x"3876892a",
2041 => x"77832a56",
2042 => x"5372802e",
2043 => x"bf387686",
2044 => x"2ab80555",
2045 => x"847327b4",
2046 => x"3880db13",
2047 => x"55947327",
2048 => x"ab38768c",
2049 => x"2a80ee05",
2050 => x"5580d473",
2051 => x"279e3876",
2052 => x"8f2a80f7",
2053 => x"055582d4",
2054 => x"73279138",
2055 => x"76922a80",
2056 => x"fc05558a",
2057 => x"d4732784",
2058 => x"3880fe55",
2059 => x"74101010",
2060 => x"80deb805",
2061 => x"88110855",
2062 => x"5673762e",
2063 => x"82b33884",
2064 => x"1408fc06",
2065 => x"53767327",
2066 => x"8d388814",
2067 => x"08547376",
2068 => x"2e098106",
2069 => x"ea388c14",
2070 => x"08708c1a",
2071 => x"0c74881a",
2072 => x"0c788812",
2073 => x"0c56778c",
2074 => x"150c7a51",
2075 => x"ed933f8c",
2076 => x"3d0d0477",
2077 => x"08787131",
2078 => x"59770588",
2079 => x"19085457",
2080 => x"7280dec0",
2081 => x"2e80e038",
2082 => x"8c180870",
2083 => x"8c150c73",
2084 => x"88120c56",
2085 => x"fe893988",
2086 => x"15088c16",
2087 => x"08708c13",
2088 => x"0c578817",
2089 => x"0cfea339",
2090 => x"76832a70",
2091 => x"54558075",
2092 => x"24819838",
2093 => x"72822c81",
2094 => x"712b80de",
2095 => x"bc080780",
2096 => x"deb80b84",
2097 => x"050c5374",
2098 => x"10101080",
2099 => x"deb80588",
2100 => x"11085556",
2101 => x"758c190c",
2102 => x"7388190c",
2103 => x"7788170c",
2104 => x"778c150c",
2105 => x"ff843981",
2106 => x"5afdb439",
2107 => x"78177381",
2108 => x"06545772",
2109 => x"98387708",
2110 => x"78713159",
2111 => x"77058c19",
2112 => x"08881a08",
2113 => x"718c120c",
2114 => x"88120c57",
2115 => x"57768107",
2116 => x"84190c77",
2117 => x"80deb80b",
2118 => x"88050c80",
2119 => x"deb40877",
2120 => x"26fec738",
2121 => x"80deb008",
2122 => x"527a51fa",
2123 => x"fd3f7a51",
2124 => x"ebcf3ffe",
2125 => x"ba398178",
2126 => x"8c150c78",
2127 => x"88150c73",
2128 => x"8c1a0c73",
2129 => x"881a0c5a",
2130 => x"fd803983",
2131 => x"1570822c",
2132 => x"81712b80",
2133 => x"debc0807",
2134 => x"80deb80b",
2135 => x"84050c51",
2136 => x"53741010",
2137 => x"1080deb8",
2138 => x"05881108",
2139 => x"5556fee4",
2140 => x"39745380",
2141 => x"7524a738",
2142 => x"72822c81",
2143 => x"712b80de",
2144 => x"bc080780",
2145 => x"deb80b84",
2146 => x"050c5375",
2147 => x"8c190c73",
2148 => x"88190c77",
2149 => x"88170c77",
2150 => x"8c150cfd",
2151 => x"cd398315",
2152 => x"70822c81",
2153 => x"712b80de",
2154 => x"bc080780",
2155 => x"deb80b84",
2156 => x"050c5153",
2157 => x"d639f93d",
2158 => x"0d797b58",
2159 => x"53800b80",
2160 => x"d6fc0853",
2161 => x"5672722e",
2162 => x"80c03884",
2163 => x"dc135574",
2164 => x"762eb738",
2165 => x"88150884",
2166 => x"1608ff05",
2167 => x"54548073",
2168 => x"249d388c",
2169 => x"14227090",
2170 => x"2b70902c",
2171 => x"51535871",
2172 => x"80d83880",
2173 => x"dc14ff14",
2174 => x"54547280",
2175 => x"25e53874",
2176 => x"085574d0",
2177 => x"3880d6fc",
2178 => x"085284dc",
2179 => x"12557480",
2180 => x"2eb13888",
2181 => x"15088416",
2182 => x"08ff0554",
2183 => x"54807324",
2184 => x"9c388c14",
2185 => x"2270902b",
2186 => x"70902c51",
2187 => x"535871ad",
2188 => x"3880dc14",
2189 => x"ff145454",
2190 => x"728025e6",
2191 => x"38740855",
2192 => x"74d13875",
2193 => x"800c893d",
2194 => x"0d047351",
2195 => x"762d7580",
2196 => x"080780dc",
2197 => x"15ff1555",
2198 => x"5556ff9e",
2199 => x"39735176",
2200 => x"2d758008",
2201 => x"0780dc15",
2202 => x"ff155555",
2203 => x"56ca39ea",
2204 => x"3d0d688c",
2205 => x"1122700a",
2206 => x"100a8106",
2207 => x"57585674",
2208 => x"80e4388e",
2209 => x"16227090",
2210 => x"2b70902c",
2211 => x"51555880",
2212 => x"7424b138",
2213 => x"983dc405",
2214 => x"53735280",
2215 => x"d6fc0851",
2216 => x"86833f80",
2217 => x"0b800824",
2218 => x"97387983",
2219 => x"e0800654",
2220 => x"7380c080",
2221 => x"2e818f38",
2222 => x"73828080",
2223 => x"2e819138",
2224 => x"8c162257",
2225 => x"76908007",
2226 => x"54738c17",
2227 => x"23888052",
2228 => x"80d6fc08",
2229 => x"51d9d13f",
2230 => x"80089d38",
2231 => x"8c162282",
2232 => x"0754738c",
2233 => x"172380c3",
2234 => x"1670770c",
2235 => x"90170c81",
2236 => x"0b94170c",
2237 => x"983d0d04",
2238 => x"80d6fc08",
2239 => x"bd930bbc",
2240 => x"120c548c",
2241 => x"16228180",
2242 => x"0754738c",
2243 => x"17238008",
2244 => x"760c8008",
2245 => x"90170c88",
2246 => x"800b9417",
2247 => x"0c74802e",
2248 => x"d3388e16",
2249 => x"2270902b",
2250 => x"70902c53",
2251 => x"55588df3",
2252 => x"3f800880",
2253 => x"2effbd38",
2254 => x"8c162281",
2255 => x"0754738c",
2256 => x"1723983d",
2257 => x"0d04810b",
2258 => x"8c172258",
2259 => x"55fef539",
2260 => x"a8160880",
2261 => x"c9c92e09",
2262 => x"8106fee4",
2263 => x"388c1622",
2264 => x"88800754",
2265 => x"738c1723",
2266 => x"88800b80",
2267 => x"cc170cfe",
2268 => x"dc39fc3d",
2269 => x"0d767971",
2270 => x"028c059f",
2271 => x"05335755",
2272 => x"53558372",
2273 => x"278a3874",
2274 => x"83065170",
2275 => x"802ea238",
2276 => x"ff125271",
2277 => x"ff2e9338",
2278 => x"73737081",
2279 => x"055534ff",
2280 => x"125271ff",
2281 => x"2e098106",
2282 => x"ef387480",
2283 => x"0c863d0d",
2284 => x"04747488",
2285 => x"2b750770",
2286 => x"71902b07",
2287 => x"5154518f",
2288 => x"7227a538",
2289 => x"72717084",
2290 => x"05530c72",
2291 => x"71708405",
2292 => x"530c7271",
2293 => x"70840553",
2294 => x"0c727170",
2295 => x"8405530c",
2296 => x"f0125271",
2297 => x"8f26dd38",
2298 => x"83722790",
2299 => x"38727170",
2300 => x"8405530c",
2301 => x"fc125271",
2302 => x"8326f238",
2303 => x"7053ff90",
2304 => x"39f93d0d",
2305 => x"797c557b",
2306 => x"548e1122",
2307 => x"70902b70",
2308 => x"902c5557",
2309 => x"80d6fc08",
2310 => x"53585683",
2311 => x"f63f8008",
2312 => x"57800b80",
2313 => x"08249338",
2314 => x"80d01608",
2315 => x"80080580",
2316 => x"d0170c76",
2317 => x"800c893d",
2318 => x"0d048c16",
2319 => x"2283dfff",
2320 => x"0655748c",
2321 => x"17237680",
2322 => x"0c893d0d",
2323 => x"04fa3d0d",
2324 => x"788c1122",
2325 => x"70882a70",
2326 => x"81065157",
2327 => x"585674a9",
2328 => x"388c1622",
2329 => x"83dfff06",
2330 => x"55748c17",
2331 => x"237a5479",
2332 => x"538e1622",
2333 => x"70902b70",
2334 => x"902c5456",
2335 => x"80d6fc08",
2336 => x"525681b2",
2337 => x"3f883d0d",
2338 => x"04825480",
2339 => x"538e1622",
2340 => x"70902b70",
2341 => x"902c5456",
2342 => x"80d6fc08",
2343 => x"525782bb",
2344 => x"3f8c1622",
2345 => x"83dfff06",
2346 => x"55748c17",
2347 => x"237a5479",
2348 => x"538e1622",
2349 => x"70902b70",
2350 => x"902c5456",
2351 => x"80d6fc08",
2352 => x"525680f2",
2353 => x"3f883d0d",
2354 => x"04f93d0d",
2355 => x"797c557b",
2356 => x"548e1122",
2357 => x"70902b70",
2358 => x"902c5557",
2359 => x"80d6fc08",
2360 => x"53585681",
2361 => x"f63f8008",
2362 => x"578008ff",
2363 => x"2e99388c",
2364 => x"1622a080",
2365 => x"0755748c",
2366 => x"17238008",
2367 => x"80d0170c",
2368 => x"76800c89",
2369 => x"3d0d048c",
2370 => x"162283df",
2371 => x"ff065574",
2372 => x"8c172376",
2373 => x"800c893d",
2374 => x"0d047070",
2375 => x"70748e11",
2376 => x"2270902b",
2377 => x"70902c55",
2378 => x"51515380",
2379 => x"d6fc0851",
2380 => x"bd3f5050",
2381 => x"5004fb3d",
2382 => x"0d800b80",
2383 => x"e7800c7a",
2384 => x"53795278",
2385 => x"51839c3f",
2386 => x"80085580",
2387 => x"08ff2e88",
2388 => x"3874800c",
2389 => x"873d0d04",
2390 => x"80e78008",
2391 => x"5675802e",
2392 => x"f0387776",
2393 => x"710c5474",
2394 => x"800c873d",
2395 => x"0d047070",
2396 => x"7070800b",
2397 => x"80e7800c",
2398 => x"765185a4",
2399 => x"3f800853",
2400 => x"8008ff2e",
2401 => x"89387280",
2402 => x"0c505050",
2403 => x"500480e7",
2404 => x"80085473",
2405 => x"802eef38",
2406 => x"7574710c",
2407 => x"5272800c",
2408 => x"50505050",
2409 => x"04fc3d0d",
2410 => x"800b80e7",
2411 => x"800c7852",
2412 => x"775187d4",
2413 => x"3f800854",
2414 => x"8008ff2e",
2415 => x"88387380",
2416 => x"0c863d0d",
2417 => x"0480e780",
2418 => x"08557480",
2419 => x"2ef03876",
2420 => x"75710c53",
2421 => x"73800c86",
2422 => x"3d0d04fb",
2423 => x"3d0d800b",
2424 => x"80e7800c",
2425 => x"7a537952",
2426 => x"785185b0",
2427 => x"3f800855",
2428 => x"8008ff2e",
2429 => x"88387480",
2430 => x"0c873d0d",
2431 => x"0480e780",
2432 => x"08567580",
2433 => x"2ef03877",
2434 => x"76710c54",
2435 => x"74800c87",
2436 => x"3d0d04fb",
2437 => x"3d0d800b",
2438 => x"80e7800c",
2439 => x"7a537952",
2440 => x"785182b7",
2441 => x"3f800855",
2442 => x"8008ff2e",
2443 => x"88387480",
2444 => x"0c873d0d",
2445 => x"0480e780",
2446 => x"08567580",
2447 => x"2ef03877",
2448 => x"76710c54",
2449 => x"74800c87",
2450 => x"3d0d0481",
2451 => x"0b800c04",
2452 => x"7072812e",
2453 => x"8738800b",
2454 => x"800c5004",
2455 => x"735180fd",
2456 => x"3f707070",
2457 => x"80e78408",
2458 => x"51708a38",
2459 => x"80e78c70",
2460 => x"80e7840c",
2461 => x"51707512",
2462 => x"5252ff53",
2463 => x"7087fb80",
2464 => x"80268838",
2465 => x"7080e784",
2466 => x"0c715372",
2467 => x"800c5050",
2468 => x"50047070",
2469 => x"7070800b",
2470 => x"80d6f008",
2471 => x"54547281",
2472 => x"2e9e3873",
2473 => x"80e7880c",
2474 => x"ffbbbe3f",
2475 => x"ffbad13f",
2476 => x"80e6c052",
2477 => x"8151ffbe",
2478 => x"913f8008",
2479 => x"51879b3f",
2480 => x"7280e788",
2481 => x"0cffbba1",
2482 => x"3fffbab4",
2483 => x"3f80e6c0",
2484 => x"528151ff",
2485 => x"bdf43f80",
2486 => x"085186fe",
2487 => x"3f00ff39",
2488 => x"00ff39f5",
2489 => x"3d0d7e60",
2490 => x"80e78808",
2491 => x"705b585b",
2492 => x"5b7580c5",
2493 => x"38777a25",
2494 => x"a238771b",
2495 => x"70337081",
2496 => x"ff065858",
2497 => x"59758a2e",
2498 => x"99387681",
2499 => x"ff0651ff",
2500 => x"bab83f81",
2501 => x"18587978",
2502 => x"24e03879",
2503 => x"800c8d3d",
2504 => x"0d048d51",
2505 => x"ffbaa33f",
2506 => x"78337081",
2507 => x"ff065257",
2508 => x"ffba973f",
2509 => x"811858de",
2510 => x"3979557a",
2511 => x"547d5385",
2512 => x"528d3dfc",
2513 => x"0551ffb9",
2514 => x"e13f8008",
2515 => x"5686843f",
2516 => x"7b80080c",
2517 => x"75800c8d",
2518 => x"3d0d04f6",
2519 => x"3d0d7d7f",
2520 => x"80e78808",
2521 => x"705a585a",
2522 => x"5a7580c4",
2523 => x"38767925",
2524 => x"b238761a",
2525 => x"56ffb9b4",
2526 => x"3f800876",
2527 => x"34800b80",
2528 => x"0881ff06",
2529 => x"5758758a",
2530 => x"2ea23875",
2531 => x"8d327030",
2532 => x"7080257a",
2533 => x"07515156",
2534 => x"75b83881",
2535 => x"17577877",
2536 => x"24d03876",
2537 => x"5675800c",
2538 => x"8c3d0d04",
2539 => x"8158dc39",
2540 => x"78557954",
2541 => x"7c538452",
2542 => x"8c3dfc05",
2543 => x"51ffb8ea",
2544 => x"3f800856",
2545 => x"858d3f7a",
2546 => x"80080c75",
2547 => x"800c8c3d",
2548 => x"0d048117",
2549 => x"56cf39f9",
2550 => x"3d0d7957",
2551 => x"80e78808",
2552 => x"802ead38",
2553 => x"7651c8f8",
2554 => x"3f7b567a",
2555 => x"55800881",
2556 => x"05547653",
2557 => x"8252893d",
2558 => x"fc0551ff",
2559 => x"b8ac3f80",
2560 => x"085784cf",
2561 => x"3f778008",
2562 => x"0c76800c",
2563 => x"893d0d04",
2564 => x"84c13f85",
2565 => x"0b80080c",
2566 => x"ff0b800c",
2567 => x"893d0d04",
2568 => x"fb3d0d80",
2569 => x"e7880870",
2570 => x"56547388",
2571 => x"3874800c",
2572 => x"873d0d04",
2573 => x"77538352",
2574 => x"873dfc05",
2575 => x"51ffb7ea",
2576 => x"3f800854",
2577 => x"848d3f75",
2578 => x"80080c73",
2579 => x"800c873d",
2580 => x"0d04ff0b",
2581 => x"800c04fb",
2582 => x"3d0d7755",
2583 => x"80e78808",
2584 => x"802ea938",
2585 => x"7451c7f8",
2586 => x"3f800881",
2587 => x"05547453",
2588 => x"8752873d",
2589 => x"fc0551ff",
2590 => x"b7b03f80",
2591 => x"085583d3",
2592 => x"3f758008",
2593 => x"0c74800c",
2594 => x"873d0d04",
2595 => x"83c53f85",
2596 => x"0b80080c",
2597 => x"ff0b800c",
2598 => x"873d0d04",
2599 => x"fa3d0d80",
2600 => x"e7880880",
2601 => x"2ea3387a",
2602 => x"55795478",
2603 => x"53865288",
2604 => x"3dfc0551",
2605 => x"ffb6f33f",
2606 => x"80085683",
2607 => x"963f7680",
2608 => x"080c7580",
2609 => x"0c883d0d",
2610 => x"0483883f",
2611 => x"9d0b8008",
2612 => x"0cff0b80",
2613 => x"0c883d0d",
2614 => x"04fb3d0d",
2615 => x"77795656",
2616 => x"80705454",
2617 => x"7375259f",
2618 => x"38741010",
2619 => x"10f80552",
2620 => x"72167033",
2621 => x"70742b76",
2622 => x"078116f8",
2623 => x"16565656",
2624 => x"51517473",
2625 => x"24ea3873",
2626 => x"800c873d",
2627 => x"0d04fc3d",
2628 => x"0d767855",
2629 => x"55bc5380",
2630 => x"527351f4",
2631 => x"d53f8452",
2632 => x"7451ffb5",
2633 => x"3f800874",
2634 => x"23845284",
2635 => x"1551ffa9",
2636 => x"3f800882",
2637 => x"15238452",
2638 => x"881551ff",
2639 => x"9c3f8008",
2640 => x"84150c84",
2641 => x"528c1551",
2642 => x"ff8f3f80",
2643 => x"08881523",
2644 => x"84529015",
2645 => x"51ff823f",
2646 => x"80088a15",
2647 => x"23845294",
2648 => x"1551fef5",
2649 => x"3f80088c",
2650 => x"15238452",
2651 => x"981551fe",
2652 => x"e83f8008",
2653 => x"8e152388",
2654 => x"529c1551",
2655 => x"fedb3f80",
2656 => x"0890150c",
2657 => x"863d0d04",
2658 => x"e93d0d6a",
2659 => x"80e78808",
2660 => x"57577593",
2661 => x"3880c080",
2662 => x"0b84180c",
2663 => x"75ac180c",
2664 => x"75800c99",
2665 => x"3d0d0489",
2666 => x"3d70556a",
2667 => x"54558a52",
2668 => x"993dffbc",
2669 => x"0551ffb4",
2670 => x"f13f8008",
2671 => x"77537552",
2672 => x"56fecb3f",
2673 => x"818d3f77",
2674 => x"80080c75",
2675 => x"800c993d",
2676 => x"0d04e93d",
2677 => x"0d695780",
2678 => x"e7880880",
2679 => x"2eb63876",
2680 => x"51c4fd3f",
2681 => x"893d7056",
2682 => x"80088105",
2683 => x"55775456",
2684 => x"8f52993d",
2685 => x"ffbc0551",
2686 => x"ffb4af3f",
2687 => x"80086b53",
2688 => x"765257fe",
2689 => x"893f80cb",
2690 => x"3f778008",
2691 => x"0c76800c",
2692 => x"993d0d04",
2693 => x"be3f850b",
2694 => x"80080cff",
2695 => x"0b800c99",
2696 => x"3d0d04fc",
2697 => x"3d0d8154",
2698 => x"80e78808",
2699 => x"88387380",
2700 => x"0c863d0d",
2701 => x"04765397",
2702 => x"b952863d",
2703 => x"fc0551ff",
2704 => x"b3e83f80",
2705 => x"08548c3f",
2706 => x"7480080c",
2707 => x"73800c86",
2708 => x"3d0d0480",
2709 => x"d6fc0880",
2710 => x"0c04f73d",
2711 => x"0d7b80d6",
2712 => x"fc0882c8",
2713 => x"11085a54",
2714 => x"5a77802e",
2715 => x"80da3881",
2716 => x"88188419",
2717 => x"08ff0581",
2718 => x"712b5955",
2719 => x"59807424",
2720 => x"80ea3880",
2721 => x"7424b538",
2722 => x"73822b78",
2723 => x"11880556",
2724 => x"56818019",
2725 => x"08770653",
2726 => x"72802eb6",
2727 => x"38781670",
2728 => x"08535379",
2729 => x"51740853",
2730 => x"722dff14",
2731 => x"fc17fc17",
2732 => x"79812c5a",
2733 => x"57575473",
2734 => x"8025d638",
2735 => x"77085877",
2736 => x"ffad3880",
2737 => x"d6fc0853",
2738 => x"bc1308a5",
2739 => x"387951f8",
2740 => x"8c3f7408",
2741 => x"53722dff",
2742 => x"14fc17fc",
2743 => x"1779812c",
2744 => x"5a575754",
2745 => x"738025ff",
2746 => x"a838d139",
2747 => x"8057ff93",
2748 => x"397251bc",
2749 => x"13085372",
2750 => x"2d7951f7",
2751 => x"e03f7070",
2752 => x"80e6c80b",
2753 => x"fc057008",
2754 => x"525270ff",
2755 => x"2e913870",
2756 => x"2dfc1270",
2757 => x"08525270",
2758 => x"ff2e0981",
2759 => x"06f13850",
2760 => x"500404ff",
2761 => x"b4c73f04",
2762 => x"48656c6c",
2763 => x"6f20776f",
2764 => x"726c6420",
2765 => x"310a0000",
2766 => x"48656c6c",
2767 => x"6f20776f",
2768 => x"726c6420",
2769 => x"320a0000",
2770 => x"0a000000",
2771 => x"43000000",
2772 => x"64756d6d",
2773 => x"792e6578",
2774 => x"65000000",
2775 => x"00ffffff",
2776 => x"ff00ffff",
2777 => x"ffff00ff",
2778 => x"ffffff00",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00003350",
2783 => x"00002b80",
2784 => x"00000000",
2785 => x"00002de8",
2786 => x"00002e44",
2787 => x"00002ea0",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"00000000",
2792 => x"00000000",
2793 => x"00000000",
2794 => x"00000000",
2795 => x"00000000",
2796 => x"00000000",
2797 => x"00002b4c",
2798 => x"00000000",
2799 => x"00000000",
2800 => x"00000000",
2801 => x"00000000",
2802 => x"00000000",
2803 => x"00000000",
2804 => x"00000000",
2805 => x"00000000",
2806 => x"00000000",
2807 => x"00000000",
2808 => x"00000000",
2809 => x"00000000",
2810 => x"00000000",
2811 => x"00000000",
2812 => x"00000000",
2813 => x"00000000",
2814 => x"00000000",
2815 => x"00000000",
2816 => x"00000000",
2817 => x"00000000",
2818 => x"00000000",
2819 => x"00000000",
2820 => x"00000000",
2821 => x"00000000",
2822 => x"00000000",
2823 => x"00000000",
2824 => x"00000000",
2825 => x"00000000",
2826 => x"00000001",
2827 => x"330eabcd",
2828 => x"1234e66d",
2829 => x"deec0005",
2830 => x"000b0000",
2831 => x"00000000",
2832 => x"00000000",
2833 => x"00000000",
2834 => x"00000000",
2835 => x"00000000",
2836 => x"00000000",
2837 => x"00000000",
2838 => x"00000000",
2839 => x"00000000",
2840 => x"00000000",
2841 => x"00000000",
2842 => x"00000000",
2843 => x"00000000",
2844 => x"00000000",
2845 => x"00000000",
2846 => x"00000000",
2847 => x"00000000",
2848 => x"00000000",
2849 => x"00000000",
2850 => x"00000000",
2851 => x"00000000",
2852 => x"00000000",
2853 => x"00000000",
2854 => x"00000000",
2855 => x"00000000",
2856 => x"00000000",
2857 => x"00000000",
2858 => x"00000000",
2859 => x"00000000",
2860 => x"00000000",
2861 => x"00000000",
2862 => x"00000000",
2863 => x"00000000",
2864 => x"00000000",
2865 => x"00000000",
2866 => x"00000000",
2867 => x"00000000",
2868 => x"00000000",
2869 => x"00000000",
2870 => x"00000000",
2871 => x"00000000",
2872 => x"00000000",
2873 => x"00000000",
2874 => x"00000000",
2875 => x"00000000",
2876 => x"00000000",
2877 => x"00000000",
2878 => x"00000000",
2879 => x"00000000",
2880 => x"00000000",
2881 => x"00000000",
2882 => x"00000000",
2883 => x"00000000",
2884 => x"00000000",
2885 => x"00000000",
2886 => x"00000000",
2887 => x"00000000",
2888 => x"00000000",
2889 => x"00000000",
2890 => x"00000000",
2891 => x"00000000",
2892 => x"00000000",
2893 => x"00000000",
2894 => x"00000000",
2895 => x"00000000",
2896 => x"00000000",
2897 => x"00000000",
2898 => x"00000000",
2899 => x"00000000",
2900 => x"00000000",
2901 => x"00000000",
2902 => x"00000000",
2903 => x"00000000",
2904 => x"00000000",
2905 => x"00000000",
2906 => x"00000000",
2907 => x"00000000",
2908 => x"00000000",
2909 => x"00000000",
2910 => x"00000000",
2911 => x"00000000",
2912 => x"00000000",
2913 => x"00000000",
2914 => x"00000000",
2915 => x"00000000",
2916 => x"00000000",
2917 => x"00000000",
2918 => x"00000000",
2919 => x"00000000",
2920 => x"00000000",
2921 => x"00000000",
2922 => x"00000000",
2923 => x"00000000",
2924 => x"00000000",
2925 => x"00000000",
2926 => x"00000000",
2927 => x"00000000",
2928 => x"00000000",
2929 => x"00000000",
2930 => x"00000000",
2931 => x"00000000",
2932 => x"00000000",
2933 => x"00000000",
2934 => x"00000000",
2935 => x"00000000",
2936 => x"00000000",
2937 => x"00000000",
2938 => x"00000000",
2939 => x"00000000",
2940 => x"00000000",
2941 => x"00000000",
2942 => x"00000000",
2943 => x"00000000",
2944 => x"00000000",
2945 => x"00000000",
2946 => x"00000000",
2947 => x"00000000",
2948 => x"00000000",
2949 => x"00000000",
2950 => x"00000000",
2951 => x"00000000",
2952 => x"00000000",
2953 => x"00000000",
2954 => x"00000000",
2955 => x"00000000",
2956 => x"00000000",
2957 => x"00000000",
2958 => x"00000000",
2959 => x"00000000",
2960 => x"00000000",
2961 => x"00000000",
2962 => x"00000000",
2963 => x"00000000",
2964 => x"00000000",
2965 => x"00000000",
2966 => x"00000000",
2967 => x"00000000",
2968 => x"00000000",
2969 => x"00000000",
2970 => x"00000000",
2971 => x"00000000",
2972 => x"00000000",
2973 => x"00000000",
2974 => x"00000000",
2975 => x"00000000",
2976 => x"00000000",
2977 => x"00000000",
2978 => x"00000000",
2979 => x"00000000",
2980 => x"00000000",
2981 => x"00000000",
2982 => x"00000000",
2983 => x"00000000",
2984 => x"00000000",
2985 => x"00000000",
2986 => x"00000000",
2987 => x"00000000",
2988 => x"00000000",
2989 => x"00000000",
2990 => x"00000000",
2991 => x"00000000",
2992 => x"00000000",
2993 => x"00000000",
2994 => x"00000000",
2995 => x"00000000",
2996 => x"00000000",
2997 => x"00000000",
2998 => x"00000000",
2999 => x"00000000",
3000 => x"00000000",
3001 => x"00000000",
3002 => x"00000000",
3003 => x"00000000",
3004 => x"00000000",
3005 => x"00000000",
3006 => x"00000000",
3007 => x"00000000",
3008 => x"00000000",
3009 => x"00000000",
3010 => x"00000000",
3011 => x"00000000",
3012 => x"00000000",
3013 => x"00000000",
3014 => x"00000000",
3015 => x"00000000",
3016 => x"00000000",
3017 => x"00000000",
3018 => x"00000000",
3019 => x"ffffffff",
3020 => x"00000000",
3021 => x"00020000",
3022 => x"00000000",
3023 => x"00000000",
3024 => x"00002f38",
3025 => x"00002f38",
3026 => x"00002f40",
3027 => x"00002f40",
3028 => x"00002f48",
3029 => x"00002f48",
3030 => x"00002f50",
3031 => x"00002f50",
3032 => x"00002f58",
3033 => x"00002f58",
3034 => x"00002f60",
3035 => x"00002f60",
3036 => x"00002f68",
3037 => x"00002f68",
3038 => x"00002f70",
3039 => x"00002f70",
3040 => x"00002f78",
3041 => x"00002f78",
3042 => x"00002f80",
3043 => x"00002f80",
3044 => x"00002f88",
3045 => x"00002f88",
3046 => x"00002f90",
3047 => x"00002f90",
3048 => x"00002f98",
3049 => x"00002f98",
3050 => x"00002fa0",
3051 => x"00002fa0",
3052 => x"00002fa8",
3053 => x"00002fa8",
3054 => x"00002fb0",
3055 => x"00002fb0",
3056 => x"00002fb8",
3057 => x"00002fb8",
3058 => x"00002fc0",
3059 => x"00002fc0",
3060 => x"00002fc8",
3061 => x"00002fc8",
3062 => x"00002fd0",
3063 => x"00002fd0",
3064 => x"00002fd8",
3065 => x"00002fd8",
3066 => x"00002fe0",
3067 => x"00002fe0",
3068 => x"00002fe8",
3069 => x"00002fe8",
3070 => x"00002ff0",
3071 => x"00002ff0",
3072 => x"00002ff8",
3073 => x"00002ff8",
3074 => x"00003000",
3075 => x"00003000",
3076 => x"00003008",
3077 => x"00003008",
3078 => x"00003010",
3079 => x"00003010",
3080 => x"00003018",
3081 => x"00003018",
3082 => x"00003020",
3083 => x"00003020",
3084 => x"00003028",
3085 => x"00003028",
3086 => x"00003030",
3087 => x"00003030",
3088 => x"00003038",
3089 => x"00003038",
3090 => x"00003040",
3091 => x"00003040",
3092 => x"00003048",
3093 => x"00003048",
3094 => x"00003050",
3095 => x"00003050",
3096 => x"00003058",
3097 => x"00003058",
3098 => x"00003060",
3099 => x"00003060",
3100 => x"00003068",
3101 => x"00003068",
3102 => x"00003070",
3103 => x"00003070",
3104 => x"00003078",
3105 => x"00003078",
3106 => x"00003080",
3107 => x"00003080",
3108 => x"00003088",
3109 => x"00003088",
3110 => x"00003090",
3111 => x"00003090",
3112 => x"00003098",
3113 => x"00003098",
3114 => x"000030a0",
3115 => x"000030a0",
3116 => x"000030a8",
3117 => x"000030a8",
3118 => x"000030b0",
3119 => x"000030b0",
3120 => x"000030b8",
3121 => x"000030b8",
3122 => x"000030c0",
3123 => x"000030c0",
3124 => x"000030c8",
3125 => x"000030c8",
3126 => x"000030d0",
3127 => x"000030d0",
3128 => x"000030d8",
3129 => x"000030d8",
3130 => x"000030e0",
3131 => x"000030e0",
3132 => x"000030e8",
3133 => x"000030e8",
3134 => x"000030f0",
3135 => x"000030f0",
3136 => x"000030f8",
3137 => x"000030f8",
3138 => x"00003100",
3139 => x"00003100",
3140 => x"00003108",
3141 => x"00003108",
3142 => x"00003110",
3143 => x"00003110",
3144 => x"00003118",
3145 => x"00003118",
3146 => x"00003120",
3147 => x"00003120",
3148 => x"00003128",
3149 => x"00003128",
3150 => x"00003130",
3151 => x"00003130",
3152 => x"00003138",
3153 => x"00003138",
3154 => x"00003140",
3155 => x"00003140",
3156 => x"00003148",
3157 => x"00003148",
3158 => x"00003150",
3159 => x"00003150",
3160 => x"00003158",
3161 => x"00003158",
3162 => x"00003160",
3163 => x"00003160",
3164 => x"00003168",
3165 => x"00003168",
3166 => x"00003170",
3167 => x"00003170",
3168 => x"00003178",
3169 => x"00003178",
3170 => x"00003180",
3171 => x"00003180",
3172 => x"00003188",
3173 => x"00003188",
3174 => x"00003190",
3175 => x"00003190",
3176 => x"00003198",
3177 => x"00003198",
3178 => x"000031a0",
3179 => x"000031a0",
3180 => x"000031a8",
3181 => x"000031a8",
3182 => x"000031b0",
3183 => x"000031b0",
3184 => x"000031b8",
3185 => x"000031b8",
3186 => x"000031c0",
3187 => x"000031c0",
3188 => x"000031c8",
3189 => x"000031c8",
3190 => x"000031d0",
3191 => x"000031d0",
3192 => x"000031d8",
3193 => x"000031d8",
3194 => x"000031e0",
3195 => x"000031e0",
3196 => x"000031e8",
3197 => x"000031e8",
3198 => x"000031f0",
3199 => x"000031f0",
3200 => x"000031f8",
3201 => x"000031f8",
3202 => x"00003200",
3203 => x"00003200",
3204 => x"00003208",
3205 => x"00003208",
3206 => x"00003210",
3207 => x"00003210",
3208 => x"00003218",
3209 => x"00003218",
3210 => x"00003220",
3211 => x"00003220",
3212 => x"00003228",
3213 => x"00003228",
3214 => x"00003230",
3215 => x"00003230",
3216 => x"00003238",
3217 => x"00003238",
3218 => x"00003240",
3219 => x"00003240",
3220 => x"00003248",
3221 => x"00003248",
3222 => x"00003250",
3223 => x"00003250",
3224 => x"00003258",
3225 => x"00003258",
3226 => x"00003260",
3227 => x"00003260",
3228 => x"00003268",
3229 => x"00003268",
3230 => x"00003270",
3231 => x"00003270",
3232 => x"00003278",
3233 => x"00003278",
3234 => x"00003280",
3235 => x"00003280",
3236 => x"00003288",
3237 => x"00003288",
3238 => x"00003290",
3239 => x"00003290",
3240 => x"00003298",
3241 => x"00003298",
3242 => x"000032a0",
3243 => x"000032a0",
3244 => x"000032a8",
3245 => x"000032a8",
3246 => x"000032b0",
3247 => x"000032b0",
3248 => x"000032b8",
3249 => x"000032b8",
3250 => x"000032c0",
3251 => x"000032c0",
3252 => x"000032c8",
3253 => x"000032c8",
3254 => x"000032d0",
3255 => x"000032d0",
3256 => x"000032d8",
3257 => x"000032d8",
3258 => x"000032e0",
3259 => x"000032e0",
3260 => x"000032e8",
3261 => x"000032e8",
3262 => x"000032f0",
3263 => x"000032f0",
3264 => x"000032f8",
3265 => x"000032f8",
3266 => x"00003300",
3267 => x"00003300",
3268 => x"00003308",
3269 => x"00003308",
3270 => x"00003310",
3271 => x"00003310",
3272 => x"00003318",
3273 => x"00003318",
3274 => x"00003320",
3275 => x"00003320",
3276 => x"00003328",
3277 => x"00003328",
3278 => x"00003330",
3279 => x"00003330",
3280 => x"00002b50",
3281 => x"ffffffff",
3282 => x"00000000",
3283 => x"ffffffff",
3284 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') then
			ram(conv_integer(memAAddr)) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(conv_integer(memAAddr));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(conv_integer(memBAddr)) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(conv_integer(memBAddr));
		end if;
	end if;
end process;




end dualport_ram_arch;
