-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0bb5",
     1 => x"a7040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0bb8",
     9 => x"8c040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0bb7",
    73 => x"c0040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0bb7a3",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80f5",
   162 => x"d8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"b7a60400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0bb7",
   169 => x"f4040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0bb7",
   177 => x"dc040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80f5e80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053351",
   258 => x"b5cc3f71",
   259 => x"b00c833d",
   260 => x"0d04fa3d",
   261 => x"0d8a51b0",
   262 => x"993f8b9a",
   263 => x"3fff54a5",
   264 => x"bd530b0b",
   265 => x"80e0dc52",
   266 => x"0b0b80e0",
   267 => x"ec518b9f",
   268 => x"3fff54a5",
   269 => x"d4530b0b",
   270 => x"80e0f452",
   271 => x"0b0b80e1",
   272 => x"90518b8b",
   273 => x"3f86548e",
   274 => x"e5530b0b",
   275 => x"80e19852",
   276 => x"0b0b80e1",
   277 => x"a8518af7",
   278 => x"3f8754ad",
   279 => x"e5530b0b",
   280 => x"80e1b052",
   281 => x"0b0b80ec",
   282 => x"9c518ae3",
   283 => x"3f8854af",
   284 => x"cd530b0b",
   285 => x"80e1c852",
   286 => x"0b0b80e1",
   287 => x"c0518acf",
   288 => x"3f8954b2",
   289 => x"b4530b0b",
   290 => x"80e1d452",
   291 => x"0b0b80e1",
   292 => x"f4518abb",
   293 => x"3fff54b3",
   294 => x"a2530b0b",
   295 => x"80e1fc52",
   296 => x"0b0b80e2",
   297 => x"a4518aa7",
   298 => x"3fff54b3",
   299 => x"fe530b0b",
   300 => x"80e2ac52",
   301 => x"0b0b80e2",
   302 => x"c8518a93",
   303 => x"3fff5490",
   304 => x"c1530b0b",
   305 => x"80e2d052",
   306 => x"0b0b80e2",
   307 => x"f85189ff",
   308 => x"3fff5490",
   309 => x"d6530b0b",
   310 => x"80e38052",
   311 => x"0b0b80e3",
   312 => x"9c5189eb",
   313 => x"3f8b54b2",
   314 => x"f7530b0b",
   315 => x"80e3a452",
   316 => x"0b0b80e3",
   317 => x"bc5189d7",
   318 => x"3f8c54b3",
   319 => x"90530b0b",
   320 => x"80e3c452",
   321 => x"0b0b80e3",
   322 => x"e05189c3",
   323 => x"3f8d54b0",
   324 => x"c3530b0b",
   325 => x"80e3e852",
   326 => x"0b0b80e4",
   327 => x"805189af",
   328 => x"3f8e54b1",
   329 => x"df530b0b",
   330 => x"80e48852",
   331 => x"0b0b80e4",
   332 => x"a451899b",
   333 => x"3fff548f",
   334 => x"be530b0b",
   335 => x"80e4ac52",
   336 => x"0b0b80e4",
   337 => x"d0518987",
   338 => x"3f8f548e",
   339 => x"fe530b0b",
   340 => x"80e4d852",
   341 => x"0b0b80e5",
   342 => x"805188f3",
   343 => x"3fff54ac",
   344 => x"c6530b0b",
   345 => x"80e58852",
   346 => x"0b0b80e5",
   347 => x"9c5188df",
   348 => x"3fff5490",
   349 => x"eb530b0b",
   350 => x"80e5a452",
   351 => x"0b0b80e5",
   352 => x"bc5188cb",
   353 => x"3fff54ad",
   354 => x"b9530b0b",
   355 => x"80e5c452",
   356 => x"0b0b80e5",
   357 => x"d45188b7",
   358 => x"3f82548e",
   359 => x"b1530b0b",
   360 => x"80f3b052",
   361 => x"0b0b80e0",
   362 => x"d45188a3",
   363 => x"3f8f8e3f",
   364 => x"898e3f81",
   365 => x"0b819dc0",
   366 => x"348185d0",
   367 => x"337081ff",
   368 => x"06565674",
   369 => x"81ea38b1",
   370 => x"d83fb008",
   371 => x"81d33888",
   372 => x"fd3f80f5",
   373 => x"f4087008",
   374 => x"70842a81",
   375 => x"06515657",
   376 => x"74802e80",
   377 => x"f238f881",
   378 => x"c08e8056",
   379 => x"8185cc08",
   380 => x"802e8183",
   381 => x"387581ff",
   382 => x"0684180c",
   383 => x"80f5c833",
   384 => x"7081ff06",
   385 => x"51557480",
   386 => x"2e80c138",
   387 => x"759f2a76",
   388 => x"10075681",
   389 => x"85d03370",
   390 => x"81ff0651",
   391 => x"5574802e",
   392 => x"d438800b",
   393 => x"8185d034",
   394 => x"8fd43f80",
   395 => x"f5c43357",
   396 => x"76a53880",
   397 => x"f5f40876",
   398 => x"81ff0684",
   399 => x"120c80f5",
   400 => x"c8337081",
   401 => x"ff065156",
   402 => x"5774c138",
   403 => x"75812a76",
   404 => x"9f2b0756",
   405 => x"ffbd3981",
   406 => x"9dc03356",
   407 => x"75feda38",
   408 => x"883d0d04",
   409 => x"75812a76",
   410 => x"9f2b0756",
   411 => x"80fd51af",
   412 => x"ce3f80f5",
   413 => x"f4085775",
   414 => x"81ff0684",
   415 => x"180c80f5",
   416 => x"c8337081",
   417 => x"ff065855",
   418 => x"76802ed8",
   419 => x"38759f2a",
   420 => x"76100756",
   421 => x"80fd51af",
   422 => x"a63f80f5",
   423 => x"f40857d7",
   424 => x"39b0913f",
   425 => x"b00881ff",
   426 => x"065187f3",
   427 => x"3ffea039",
   428 => x"800b8185",
   429 => x"d0348ec6",
   430 => x"3fafe63f",
   431 => x"b008802e",
   432 => x"fe8d38dd",
   433 => x"39803d0d",
   434 => x"0b0b80e5",
   435 => x"d851aafc",
   436 => x"3f0b0b80",
   437 => x"e5dc51aa",
   438 => x"f33f8185",
   439 => x"cc08802e",
   440 => x"8e380b0b",
   441 => x"80e5f851",
   442 => x"aae23f82",
   443 => x"3d0d048a",
   444 => x"51aabf3f",
   445 => x"0b0b80e6",
   446 => x"8451aad0",
   447 => x"3f0b0b80",
   448 => x"e69c51aa",
   449 => x"c73f810a",
   450 => x"51aac13f",
   451 => x"0b0b80e6",
   452 => x"b051aab8",
   453 => x"3f0b0b80",
   454 => x"e6d851aa",
   455 => x"af3f80e4",
   456 => x"51abff3f",
   457 => x"0b0b80e6",
   458 => x"ec51aaa0",
   459 => x"3f823d0d",
   460 => x"04ff923f",
   461 => x"8c873f80",
   462 => x"0bb00c04",
   463 => x"fe3d0d80",
   464 => x"f5f80898",
   465 => x"11087084",
   466 => x"2a708106",
   467 => x"51535353",
   468 => x"70802e8d",
   469 => x"3871ef06",
   470 => x"98140c81",
   471 => x"0b8185d0",
   472 => x"34843d0d",
   473 => x"04803d0d",
   474 => x"0b0b80e6",
   475 => x"8451a9dc",
   476 => x"3f8a51a9",
   477 => x"bd3f800b",
   478 => x"b00c823d",
   479 => x"0d04f93d",
   480 => x"0d81518a",
   481 => x"863fb008",
   482 => x"55825189",
   483 => x"fe3f74b0",
   484 => x"08075399",
   485 => x"cc57fce2",
   486 => x"97f68058",
   487 => x"72802e90",
   488 => x"38747554",
   489 => x"57805480",
   490 => x"770774b0",
   491 => x"08075957",
   492 => x"76517752",
   493 => x"97943f72",
   494 => x"b00c893d",
   495 => x"0d04fa3d",
   496 => x"0d815188",
   497 => x"943fb008",
   498 => x"81ff0656",
   499 => x"82518889",
   500 => x"3f75802e",
   501 => x"80e438b0",
   502 => x"08832b86",
   503 => x"8fc09082",
   504 => x"0757a3ac",
   505 => x"3fa4973f",
   506 => x"76538252",
   507 => x"8051a0a3",
   508 => x"3f80f5d4",
   509 => x"0855800b",
   510 => x"90160c82",
   511 => x"750c80f5",
   512 => x"f4088411",
   513 => x"0870810a",
   514 => x"0784130c",
   515 => x"55558a51",
   516 => x"ac873f80",
   517 => x"f5f40884",
   518 => x"110870fe",
   519 => x"0a068413",
   520 => x"0c555594",
   521 => x"51abf23f",
   522 => x"9dbb3f9f",
   523 => x"a03fff16",
   524 => x"7081ff06",
   525 => x"575475ff",
   526 => x"a93876b0",
   527 => x"0c883d0d",
   528 => x"04803d0d",
   529 => x"81518791",
   530 => x"3fb00881",
   531 => x"ff0651a3",
   532 => x"e33f823d",
   533 => x"0d04803d",
   534 => x"0d815186",
   535 => x"fc3fb008",
   536 => x"81ff0651",
   537 => x"a4963f82",
   538 => x"3d0d04fe",
   539 => x"3d0d8151",
   540 => x"86e73f80",
   541 => x"f5f40884",
   542 => x"11087081",
   543 => x"0a078413",
   544 => x"0c5353b0",
   545 => x"0851ab91",
   546 => x"3f80f5f4",
   547 => x"08841108",
   548 => x"70fe0a06",
   549 => x"7084140c",
   550 => x"b00c5353",
   551 => x"843d0d04",
   552 => x"fc3d0d80",
   553 => x"f5f40870",
   554 => x"08810a06",
   555 => x"8185cc0c",
   556 => x"54abb03f",
   557 => x"abd43f8b",
   558 => x"a53f93ec",
   559 => x"3f80f5f8",
   560 => x"08981108",
   561 => x"70880798",
   562 => x"130c5555",
   563 => x"8185cc08",
   564 => x"81803888",
   565 => x"800b819e",
   566 => x"c80cfbe9",
   567 => x"3f8185cc",
   568 => x"08802e80",
   569 => x"fe388653",
   570 => x"82528051",
   571 => x"9ea53f80",
   572 => x"f5d40855",
   573 => x"80e40b90",
   574 => x"160c8275",
   575 => x"0cb251aa",
   576 => x"983f80f5",
   577 => x"f4088411",
   578 => x"0870810a",
   579 => x"0784130c",
   580 => x"55558051",
   581 => x"aa833f80",
   582 => x"f5f40884",
   583 => x"110870fe",
   584 => x"0a068413",
   585 => x"0c555580",
   586 => x"f5d40855",
   587 => x"74085473",
   588 => x"fb380b0b",
   589 => x"80e6f451",
   590 => x"a6923f80",
   591 => x"f5d4089c",
   592 => x"11085255",
   593 => x"a7dc3f8a",
   594 => x"51a5e73f",
   595 => x"9df53fac",
   596 => x"9f3fb89c",
   597 => x"0b819ec8",
   598 => x"0cfaea3f",
   599 => x"8185cc08",
   600 => x"ff8438bd",
   601 => x"d60b819e",
   602 => x"c80cf5a6",
   603 => x"3f865382",
   604 => x"5280519d",
   605 => x"9e3f80f5",
   606 => x"d4085580",
   607 => x"e40b9016",
   608 => x"0c82750c",
   609 => x"b251a991",
   610 => x"3f80f5f4",
   611 => x"08841108",
   612 => x"70810a07",
   613 => x"84130c55",
   614 => x"558051a8",
   615 => x"fc3f80f5",
   616 => x"f4088411",
   617 => x"0870fe0a",
   618 => x"0684130c",
   619 => x"555580f5",
   620 => x"d40855fe",
   621 => x"f739800b",
   622 => x"819db834",
   623 => x"800b819d",
   624 => x"b434800b",
   625 => x"819dbc0c",
   626 => x"ff0b819d",
   627 => x"ec3404fb",
   628 => x"3d0d7a98",
   629 => x"2b70982c",
   630 => x"819db433",
   631 => x"52565372",
   632 => x"a72680d1",
   633 => x"38775272",
   634 => x"10101073",
   635 => x"10058185",
   636 => x"d40551b0",
   637 => x"963f7852",
   638 => x"819db433",
   639 => x"70902971",
   640 => x"31701010",
   641 => x"8188e405",
   642 => x"535754af",
   643 => x"fe3f819d",
   644 => x"b4337081",
   645 => x"ff065456",
   646 => x"74819dc4",
   647 => x"14347210",
   648 => x"10819bc4",
   649 => x"057a710c",
   650 => x"55811654",
   651 => x"73819db4",
   652 => x"34873d0d",
   653 => x"0480e780",
   654 => x"51a4913f",
   655 => x"873d0d04",
   656 => x"803d0d80",
   657 => x"e79c51a4",
   658 => x"833f823d",
   659 => x"0d04fc3d",
   660 => x"0d819dbc",
   661 => x"08537285",
   662 => x"38863d0d",
   663 => x"04722db0",
   664 => x"0854800b",
   665 => x"819dbc0c",
   666 => x"80e7b451",
   667 => x"a3de3f81",
   668 => x"9dec3370",
   669 => x"982b7098",
   670 => x"2c545455",
   671 => x"a051a3ef",
   672 => x"3f80e7c0",
   673 => x"51a3c53f",
   674 => x"7352a051",
   675 => x"a3e13f8a",
   676 => x"51a39f3f",
   677 => x"80e79c51",
   678 => x"a3b23f86",
   679 => x"3d0d04fa",
   680 => x"3d0d02a3",
   681 => x"05335675",
   682 => x"8d2e80f4",
   683 => x"38758832",
   684 => x"70307780",
   685 => x"ff327030",
   686 => x"72802571",
   687 => x"80250754",
   688 => x"51565855",
   689 => x"7495389f",
   690 => x"76278c38",
   691 => x"819db833",
   692 => x"5580ce75",
   693 => x"27ae3888",
   694 => x"3d0d0481",
   695 => x"9db83356",
   696 => x"75802ef3",
   697 => x"388851a2",
   698 => x"c93fa051",
   699 => x"a2c43f88",
   700 => x"51a2bf3f",
   701 => x"819db833",
   702 => x"ff055776",
   703 => x"819db834",
   704 => x"883d0d04",
   705 => x"7551a2aa",
   706 => x"3f819db8",
   707 => x"33811155",
   708 => x"5773819d",
   709 => x"b8347581",
   710 => x"9ce41834",
   711 => x"883d0d04",
   712 => x"8a51a28e",
   713 => x"3f819db8",
   714 => x"33811156",
   715 => x"5474819d",
   716 => x"b834800b",
   717 => x"819ce415",
   718 => x"34805680",
   719 => x"0b819ce4",
   720 => x"17335654",
   721 => x"74a02e83",
   722 => x"38815474",
   723 => x"802e9038",
   724 => x"73802e8b",
   725 => x"38811670",
   726 => x"81ff0657",
   727 => x"57dd3975",
   728 => x"802e80c5",
   729 => x"38800b81",
   730 => x"9db43355",
   731 => x"55747427",
   732 => x"ab387357",
   733 => x"74101010",
   734 => x"75100576",
   735 => x"54819ce4",
   736 => x"538185d4",
   737 => x"0551aecf",
   738 => x"3fb00880",
   739 => x"2eac3881",
   740 => x"157081ff",
   741 => x"06565476",
   742 => x"7526d938",
   743 => x"80e7a051",
   744 => x"a1aa3fff",
   745 => x"0b819dec",
   746 => x"3480e79c",
   747 => x"51a19d3f",
   748 => x"800b819d",
   749 => x"b834883d",
   750 => x"0d047410",
   751 => x"10819bc4",
   752 => x"05700881",
   753 => x"9dbc0c56",
   754 => x"819dc415",
   755 => x"33819dec",
   756 => x"34800b81",
   757 => x"9db834de",
   758 => x"39f73d0d",
   759 => x"02af0533",
   760 => x"59800b81",
   761 => x"9ce43381",
   762 => x"9ce45955",
   763 => x"5673a02e",
   764 => x"09810696",
   765 => x"38811670",
   766 => x"81ff0681",
   767 => x"9ce41170",
   768 => x"33535957",
   769 => x"5473a02e",
   770 => x"ec388058",
   771 => x"77792780",
   772 => x"ea388077",
   773 => x"33565474",
   774 => x"742e8338",
   775 => x"815474a0",
   776 => x"2e9a3873",
   777 => x"80c53874",
   778 => x"a02e9138",
   779 => x"81187081",
   780 => x"ff065955",
   781 => x"787826da",
   782 => x"3880c039",
   783 => x"81167081",
   784 => x"ff06819c",
   785 => x"e4117033",
   786 => x"57525757",
   787 => x"73a02e09",
   788 => x"8106d938",
   789 => x"81167081",
   790 => x"ff06819c",
   791 => x"e4117033",
   792 => x"57525757",
   793 => x"73a02ed4",
   794 => x"38c23981",
   795 => x"167081ff",
   796 => x"06819ce4",
   797 => x"11595755",
   798 => x"ff983980",
   799 => x"538b3dfc",
   800 => x"05527651",
   801 => x"b1963f8b",
   802 => x"3d0d04f7",
   803 => x"3d0d02af",
   804 => x"05335980",
   805 => x"0b819ce4",
   806 => x"33819ce4",
   807 => x"59555673",
   808 => x"a02e0981",
   809 => x"06963881",
   810 => x"167081ff",
   811 => x"06819ce4",
   812 => x"11703353",
   813 => x"59575473",
   814 => x"a02eec38",
   815 => x"80587779",
   816 => x"2780ea38",
   817 => x"80773356",
   818 => x"5474742e",
   819 => x"83388154",
   820 => x"74a02e9a",
   821 => x"387380c5",
   822 => x"3874a02e",
   823 => x"91388118",
   824 => x"7081ff06",
   825 => x"59557878",
   826 => x"26da3880",
   827 => x"c0398116",
   828 => x"7081ff06",
   829 => x"819ce411",
   830 => x"70335752",
   831 => x"575773a0",
   832 => x"2e098106",
   833 => x"d9388116",
   834 => x"7081ff06",
   835 => x"819ce411",
   836 => x"70335752",
   837 => x"575773a0",
   838 => x"2ed438c2",
   839 => x"39811670",
   840 => x"81ff0681",
   841 => x"9ce41159",
   842 => x"5755ff98",
   843 => x"3990538b",
   844 => x"3dfc0552",
   845 => x"7651b381",
   846 => x"3f8b3d0d",
   847 => x"04fb3d0d",
   848 => x"8a519dee",
   849 => x"3f80e7cc",
   850 => x"519e813f",
   851 => x"800b819d",
   852 => x"b4335454",
   853 => x"73732781",
   854 => x"963880f2",
   855 => x"90519dec",
   856 => x"3f819dc4",
   857 => x"14337098",
   858 => x"2b70982c",
   859 => x"545455a0",
   860 => x"519dfc3f",
   861 => x"80f3a451",
   862 => x"9dd23f73",
   863 => x"10101074",
   864 => x"10058185",
   865 => x"d4057052",
   866 => x"559dc13f",
   867 => x"73842b70",
   868 => x"7531822b",
   869 => x"8188e411",
   870 => x"33515456",
   871 => x"72802eb7",
   872 => x"387451a9",
   873 => x"d33fb008",
   874 => x"81ff0653",
   875 => x"72892693",
   876 => x"38a0519c",
   877 => x"fd3f8113",
   878 => x"7081ff06",
   879 => x"51538973",
   880 => x"27ef3880",
   881 => x"e7e4519d",
   882 => x"833f7574",
   883 => x"31822b81",
   884 => x"88e40551",
   885 => x"9cf63f8a",
   886 => x"519cd73f",
   887 => x"81147081",
   888 => x"ff06819d",
   889 => x"b4335555",
   890 => x"56727426",
   891 => x"feec388a",
   892 => x"519cbf3f",
   893 => x"819db433",
   894 => x"b00c873d",
   895 => x"0d04fe3d",
   896 => x"0d819ec0",
   897 => x"22ff0551",
   898 => x"70819ec0",
   899 => x"237083ff",
   900 => x"ff065170",
   901 => x"80c43881",
   902 => x"9ec43351",
   903 => x"7081ff2e",
   904 => x"b9387010",
   905 => x"1010819d",
   906 => x"f0055271",
   907 => x"33819ec4",
   908 => x"34fe7234",
   909 => x"819ec433",
   910 => x"70101010",
   911 => x"819df005",
   912 => x"52538211",
   913 => x"22819ec0",
   914 => x"23841208",
   915 => x"53722d81",
   916 => x"9ec02251",
   917 => x"70802eff",
   918 => x"be38843d",
   919 => x"0d04ff3d",
   920 => x"0d8a5271",
   921 => x"10101081",
   922 => x"9de80551",
   923 => x"fe7134ff",
   924 => x"127081ff",
   925 => x"06535171",
   926 => x"ea38ff0b",
   927 => x"819ec434",
   928 => x"833d0d04",
   929 => x"fe3d0d02",
   930 => x"93053302",
   931 => x"84059705",
   932 => x"33545271",
   933 => x"842e80d1",
   934 => x"38718424",
   935 => x"91387181",
   936 => x"2eac3880",
   937 => x"e7e8519b",
   938 => x"a33f843d",
   939 => x"0d047180",
   940 => x"d52e0981",
   941 => x"06ed3880",
   942 => x"e7f4519b",
   943 => x"8f3f728c",
   944 => x"26b33872",
   945 => x"101080ec",
   946 => x"e8055271",
   947 => x"080480e8",
   948 => x"80519af8",
   949 => x"3ffa1352",
   950 => x"7180db26",
   951 => x"98387110",
   952 => x"1080ed9c",
   953 => x"05527108",
   954 => x"0480e88c",
   955 => x"519add3f",
   956 => x"728f2e8c",
   957 => x"3880e898",
   958 => x"519ad13f",
   959 => x"843d0d04",
   960 => x"80e8a851",
   961 => x"9ac63f84",
   962 => x"3d0d0480",
   963 => x"e8c0519a",
   964 => x"bb3f843d",
   965 => x"0d0480e8",
   966 => x"d0519ab0",
   967 => x"3f843d0d",
   968 => x"0480e8e8",
   969 => x"519aa53f",
   970 => x"843d0d04",
   971 => x"80e8f851",
   972 => x"9a9a3f84",
   973 => x"3d0d0480",
   974 => x"e998519a",
   975 => x"8f3f843d",
   976 => x"0d0480e9",
   977 => x"b4519a84",
   978 => x"3f843d0d",
   979 => x"0480e9d0",
   980 => x"5199f93f",
   981 => x"843d0d04",
   982 => x"80e9e451",
   983 => x"99ee3f84",
   984 => x"3d0d0480",
   985 => x"ea805199",
   986 => x"e33f843d",
   987 => x"0d0480ea",
   988 => x"905199d8",
   989 => x"3f843d0d",
   990 => x"0480eaa0",
   991 => x"5199cd3f",
   992 => x"843d0d04",
   993 => x"80eac051",
   994 => x"99c23f84",
   995 => x"3d0d0480",
   996 => x"ead45199",
   997 => x"b73f843d",
   998 => x"0d0480ea",
   999 => x"f05199ac",
  1000 => x"3f843d0d",
  1001 => x"0480eb88",
  1002 => x"5199a13f",
  1003 => x"843d0d04",
  1004 => x"80eb9c51",
  1005 => x"99963f84",
  1006 => x"3d0d0480",
  1007 => x"ebac5199",
  1008 => x"8b3f843d",
  1009 => x"0d0480eb",
  1010 => x"c0519980",
  1011 => x"3f843d0d",
  1012 => x"0480ebd0",
  1013 => x"5198f53f",
  1014 => x"843d0d04",
  1015 => x"80ebe851",
  1016 => x"98ea3f84",
  1017 => x"3d0d0480",
  1018 => x"ebfc5198",
  1019 => x"df3f843d",
  1020 => x"0d0480ec",
  1021 => x"8c5198d4",
  1022 => x"3f843d0d",
  1023 => x"04f73d0d",
  1024 => x"02b30533",
  1025 => x"7c7008c0",
  1026 => x"80800659",
  1027 => x"545a8056",
  1028 => x"75832b77",
  1029 => x"07bfe080",
  1030 => x"07707084",
  1031 => x"05520871",
  1032 => x"088c2abf",
  1033 => x"fe800679",
  1034 => x"0771982a",
  1035 => x"728c2a9f",
  1036 => x"ff067385",
  1037 => x"2a708f06",
  1038 => x"759f0656",
  1039 => x"51585d58",
  1040 => x"52555874",
  1041 => x"8d388116",
  1042 => x"568f7627",
  1043 => x"c3388b3d",
  1044 => x"0d0480ec",
  1045 => x"a45197f4",
  1046 => x"3f755199",
  1047 => x"c53f8452",
  1048 => x"b008519b",
  1049 => x"863f80ec",
  1050 => x"b05197e0",
  1051 => x"3f745288",
  1052 => x"5197fc3f",
  1053 => x"8452b008",
  1054 => x"519af03f",
  1055 => x"80ecb851",
  1056 => x"97ca3f78",
  1057 => x"52905197",
  1058 => x"e63f8652",
  1059 => x"b008519a",
  1060 => x"da3f80ec",
  1061 => x"c05197b4",
  1062 => x"3f725199",
  1063 => x"853f8452",
  1064 => x"b008519a",
  1065 => x"c63f80ec",
  1066 => x"c85197a0",
  1067 => x"3f735198",
  1068 => x"f13f8452",
  1069 => x"b008519a",
  1070 => x"b23f80ec",
  1071 => x"d051978c",
  1072 => x"3f7752a0",
  1073 => x"5197a83f",
  1074 => x"8a52b008",
  1075 => x"519a9c3f",
  1076 => x"7992388a",
  1077 => x"5196db3f",
  1078 => x"8116568f",
  1079 => x"7627feb0",
  1080 => x"38feeb39",
  1081 => x"7881ff06",
  1082 => x"527451fb",
  1083 => x"973f8a51",
  1084 => x"96c03fe4",
  1085 => x"39f83d0d",
  1086 => x"02ab0533",
  1087 => x"59805675",
  1088 => x"852be090",
  1089 => x"11e08012",
  1090 => x"0870982a",
  1091 => x"718c2a9f",
  1092 => x"ff067285",
  1093 => x"2a708f06",
  1094 => x"749f0655",
  1095 => x"51585b53",
  1096 => x"56595574",
  1097 => x"802e81a1",
  1098 => x"3875bf26",
  1099 => x"81a93880",
  1100 => x"ecd85196",
  1101 => x"973f7551",
  1102 => x"97e83f86",
  1103 => x"52b00851",
  1104 => x"99a93f80",
  1105 => x"ecb05196",
  1106 => x"833f7452",
  1107 => x"8851969f",
  1108 => x"3f8452b0",
  1109 => x"08519993",
  1110 => x"3f80ecb8",
  1111 => x"5195ed3f",
  1112 => x"76529051",
  1113 => x"96893f86",
  1114 => x"52b00851",
  1115 => x"98fd3f80",
  1116 => x"ecc05195",
  1117 => x"d73f7251",
  1118 => x"97a83f84",
  1119 => x"52b00851",
  1120 => x"98e93f80",
  1121 => x"ecc85195",
  1122 => x"c33f7351",
  1123 => x"97943f84",
  1124 => x"52b00851",
  1125 => x"98d53f80",
  1126 => x"ecd05195",
  1127 => x"af3f7708",
  1128 => x"c0808006",
  1129 => x"52a05195",
  1130 => x"c63f8a52",
  1131 => x"b0085198",
  1132 => x"ba3f7881",
  1133 => x"ac388a51",
  1134 => x"94f83f80",
  1135 => x"5374812e",
  1136 => x"81d93876",
  1137 => x"862e81b5",
  1138 => x"38811656",
  1139 => x"80ff7627",
  1140 => x"fead388a",
  1141 => x"3d0d0480",
  1142 => x"ece05194",
  1143 => x"ef3fc016",
  1144 => x"5196bf3f",
  1145 => x"8652b008",
  1146 => x"5198803f",
  1147 => x"80ecb051",
  1148 => x"94da3f74",
  1149 => x"52885194",
  1150 => x"f63f8452",
  1151 => x"b0085197",
  1152 => x"ea3f80ec",
  1153 => x"b85194c4",
  1154 => x"3f765290",
  1155 => x"5194e03f",
  1156 => x"8652b008",
  1157 => x"5197d43f",
  1158 => x"80ecc051",
  1159 => x"94ae3f72",
  1160 => x"5195ff3f",
  1161 => x"8452b008",
  1162 => x"5197c03f",
  1163 => x"80ecc851",
  1164 => x"949a3f73",
  1165 => x"5195eb3f",
  1166 => x"8452b008",
  1167 => x"5197ac3f",
  1168 => x"80ecd051",
  1169 => x"94863f77",
  1170 => x"08c08080",
  1171 => x"0652a051",
  1172 => x"949d3f8a",
  1173 => x"52b00851",
  1174 => x"97913f78",
  1175 => x"802efed6",
  1176 => x"387681ff",
  1177 => x"06527451",
  1178 => x"f89a3f8a",
  1179 => x"5193c33f",
  1180 => x"80537481",
  1181 => x"2e098106",
  1182 => x"fec9389f",
  1183 => x"39728106",
  1184 => x"5776802e",
  1185 => x"fec33878",
  1186 => x"527751fa",
  1187 => x"f03f8116",
  1188 => x"5680ff76",
  1189 => x"27fce838",
  1190 => x"feb93974",
  1191 => x"5376862e",
  1192 => x"098106fe",
  1193 => x"a438d639",
  1194 => x"803d0d80",
  1195 => x"f5f00851",
  1196 => x"b1710c81",
  1197 => x"800b8412",
  1198 => x"0c823d0d",
  1199 => x"04803d0d",
  1200 => x"80f68008",
  1201 => x"51f8bb95",
  1202 => x"86a1710c",
  1203 => x"810bb00c",
  1204 => x"823d0d04",
  1205 => x"803d0d81",
  1206 => x"51f1fe3f",
  1207 => x"b00881ff",
  1208 => x"0651fc91",
  1209 => x"3f800bb0",
  1210 => x"0c823d0d",
  1211 => x"04ff3d0d",
  1212 => x"80f5cc08",
  1213 => x"a0110870",
  1214 => x"80ff0a06",
  1215 => x"a0130c52",
  1216 => x"52bbc880",
  1217 => x"800ba013",
  1218 => x"0c833d0d",
  1219 => x"04ff3d0d",
  1220 => x"028f0533",
  1221 => x"70982b80",
  1222 => x"f5cc0852",
  1223 => x"b0120c51",
  1224 => x"833d0d04",
  1225 => x"ff3d0d80",
  1226 => x"f5cc0852",
  1227 => x"a4120870",
  1228 => x"892a7081",
  1229 => x"06515151",
  1230 => x"70802ef0",
  1231 => x"38b41208",
  1232 => x"70902ab0",
  1233 => x"0c51833d",
  1234 => x"0d04f83d",
  1235 => x"0d7a7c57",
  1236 => x"55ff9a3f",
  1237 => x"80f5f408",
  1238 => x"84110882",
  1239 => x"80800784",
  1240 => x"120c8411",
  1241 => x"08fdffff",
  1242 => x"0684120c",
  1243 => x"84110881",
  1244 => x"80800784",
  1245 => x"120c8411",
  1246 => x"08feffff",
  1247 => x"0684120c",
  1248 => x"53900b89",
  1249 => x"3d349402",
  1250 => x"84059d05",
  1251 => x"34800284",
  1252 => x"059e0534",
  1253 => x"80e10284",
  1254 => x"059f0534",
  1255 => x"883d80f5",
  1256 => x"cc085457",
  1257 => x"a4130870",
  1258 => x"882a8106",
  1259 => x"51527180",
  1260 => x"2ef23887",
  1261 => x"51fed63f",
  1262 => x"800b80f0",
  1263 => x"93335353",
  1264 => x"72722799",
  1265 => x"38715476",
  1266 => x"13703352",
  1267 => x"52febe3f",
  1268 => x"81137081",
  1269 => x"ff065452",
  1270 => x"737326eb",
  1271 => x"38fec53f",
  1272 => x"800b80f0",
  1273 => x"93335353",
  1274 => x"72722793",
  1275 => x"387154fe",
  1276 => x"b33f8113",
  1277 => x"7081ff06",
  1278 => x"54527373",
  1279 => x"26f13874",
  1280 => x"882a5473",
  1281 => x"893d3474",
  1282 => x"0284059d",
  1283 => x"05347488",
  1284 => x"2b76982a",
  1285 => x"07527102",
  1286 => x"84059e05",
  1287 => x"3474902b",
  1288 => x"76902a07",
  1289 => x"54730284",
  1290 => x"059f0534",
  1291 => x"74982b76",
  1292 => x"882a0753",
  1293 => x"728a3d34",
  1294 => x"75028405",
  1295 => x"a1053480",
  1296 => x"f5cc0853",
  1297 => x"a4130870",
  1298 => x"882a8106",
  1299 => x"56527480",
  1300 => x"2ef23882",
  1301 => x"51fdb63f",
  1302 => x"800b80f0",
  1303 => x"8e335353",
  1304 => x"72722799",
  1305 => x"38715476",
  1306 => x"13703352",
  1307 => x"56fd9e3f",
  1308 => x"81137081",
  1309 => x"ff065455",
  1310 => x"737326eb",
  1311 => x"38fda53f",
  1312 => x"800b80f0",
  1313 => x"8e335353",
  1314 => x"72722793",
  1315 => x"387154fd",
  1316 => x"933f8113",
  1317 => x"7081ff06",
  1318 => x"54527373",
  1319 => x"26f1388a",
  1320 => x"0b893d34",
  1321 => x"ff8c0284",
  1322 => x"059d0534",
  1323 => x"80f5cc08",
  1324 => x"53a41308",
  1325 => x"70882a81",
  1326 => x"06555673",
  1327 => x"802ef238",
  1328 => x"8851fcc9",
  1329 => x"3f800b80",
  1330 => x"f0943353",
  1331 => x"53727227",
  1332 => x"99387154",
  1333 => x"76137033",
  1334 => x"5255fcb1",
  1335 => x"3f811370",
  1336 => x"81ff0654",
  1337 => x"52737326",
  1338 => x"eb38fcb8",
  1339 => x"3f800b80",
  1340 => x"f0943353",
  1341 => x"53727227",
  1342 => x"93387154",
  1343 => x"fca63f81",
  1344 => x"137081ff",
  1345 => x"06545673",
  1346 => x"7326f138",
  1347 => x"8a0b893d",
  1348 => x"34ff8c02",
  1349 => x"84059d05",
  1350 => x"3480f5cc",
  1351 => x"0853a413",
  1352 => x"0870882a",
  1353 => x"81065555",
  1354 => x"73802ef2",
  1355 => x"388951fb",
  1356 => x"dc3f800b",
  1357 => x"80f09533",
  1358 => x"53537272",
  1359 => x"27993871",
  1360 => x"54761370",
  1361 => x"335252fb",
  1362 => x"c43f8113",
  1363 => x"7081ff06",
  1364 => x"54567373",
  1365 => x"26eb38fb",
  1366 => x"cb3f800b",
  1367 => x"80f09533",
  1368 => x"53537272",
  1369 => x"27933871",
  1370 => x"54fbb93f",
  1371 => x"81137081",
  1372 => x"ff065457",
  1373 => x"737326f1",
  1374 => x"3880f5f4",
  1375 => x"08841108",
  1376 => x"80c08007",
  1377 => x"84120c84",
  1378 => x"1108ffbf",
  1379 => x"ff068412",
  1380 => x"0c54800b",
  1381 => x"b00c8a3d",
  1382 => x"0d04f83d",
  1383 => x"0d02ab05",
  1384 => x"33893d80",
  1385 => x"f5cc0856",
  1386 => x"5856a414",
  1387 => x"0870882a",
  1388 => x"81065153",
  1389 => x"72802ef2",
  1390 => x"38758180",
  1391 => x"0751facd",
  1392 => x"3f800b80",
  1393 => x"f08c1733",
  1394 => x"54547373",
  1395 => x"27953872",
  1396 => x"558051fa",
  1397 => x"b83f8114",
  1398 => x"7081ff06",
  1399 => x"55537474",
  1400 => x"26ef38fa",
  1401 => x"bf3f800b",
  1402 => x"80f08c17",
  1403 => x"337081ff",
  1404 => x"06555754",
  1405 => x"7373279a",
  1406 => x"38725576",
  1407 => x"1453faa4",
  1408 => x"3fb00873",
  1409 => x"34811470",
  1410 => x"81ff0655",
  1411 => x"53747426",
  1412 => x"ea387581",
  1413 => x"ff0680f2",
  1414 => x"9052558c",
  1415 => x"af3f8054",
  1416 => x"73752799",
  1417 => x"38731770",
  1418 => x"33535388",
  1419 => x"518cc03f",
  1420 => x"81147081",
  1421 => x"ff065556",
  1422 => x"747426e9",
  1423 => x"388a518b",
  1424 => x"f13f8a3d",
  1425 => x"0d04fe3d",
  1426 => x"0d80f5f4",
  1427 => x"08841108",
  1428 => x"70818080",
  1429 => x"0784130c",
  1430 => x"54841108",
  1431 => x"70feffff",
  1432 => x"0684130c",
  1433 => x"5452f985",
  1434 => x"3f80f098",
  1435 => x"518bdd3f",
  1436 => x"8751fea6",
  1437 => x"3f80f0a8",
  1438 => x"518bd13f",
  1439 => x"8251fe9a",
  1440 => x"3f80f0b8",
  1441 => x"518bc53f",
  1442 => x"8551fe8e",
  1443 => x"3f80f0c8",
  1444 => x"518bb93f",
  1445 => x"8651fe82",
  1446 => x"3f80f0d8",
  1447 => x"518bad3f",
  1448 => x"8851fdf6",
  1449 => x"3f80f0e8",
  1450 => x"518ba13f",
  1451 => x"8951fdea",
  1452 => x"3f800bb0",
  1453 => x"0c843d0d",
  1454 => x"04fe3d0d",
  1455 => x"80f5f408",
  1456 => x"84110882",
  1457 => x"0a078412",
  1458 => x"0c700870",
  1459 => x"902a8413",
  1460 => x"0870fd0a",
  1461 => x"0684150c",
  1462 => x"5481ffff",
  1463 => x"06b00c53",
  1464 => x"53843d0d",
  1465 => x"04ff3d0d",
  1466 => x"80f5d408",
  1467 => x"70087081",
  1468 => x"ff065151",
  1469 => x"52718926",
  1470 => x"8c387110",
  1471 => x"1080f2dc",
  1472 => x"05527108",
  1473 => x"0480f0f8",
  1474 => x"518ac13f",
  1475 => x"8a518aa2",
  1476 => x"3f800bb0",
  1477 => x"0c833d0d",
  1478 => x"0480e2f8",
  1479 => x"518aad3f",
  1480 => x"8a518a8e",
  1481 => x"3f800bb0",
  1482 => x"0c833d0d",
  1483 => x"0480f180",
  1484 => x"518a993f",
  1485 => x"8a5189fa",
  1486 => x"3f800bb0",
  1487 => x"0c833d0d",
  1488 => x"0480f188",
  1489 => x"518a853f",
  1490 => x"8a5189e6",
  1491 => x"3f800bb0",
  1492 => x"0c833d0d",
  1493 => x"0480f194",
  1494 => x"5189f13f",
  1495 => x"8a5189d2",
  1496 => x"3f800bb0",
  1497 => x"0c833d0d",
  1498 => x"0480f19c",
  1499 => x"5189dd3f",
  1500 => x"8a5189be",
  1501 => x"3f800bb0",
  1502 => x"0c833d0d",
  1503 => x"0480f1a4",
  1504 => x"5189c93f",
  1505 => x"8a5189aa",
  1506 => x"3f800bb0",
  1507 => x"0c833d0d",
  1508 => x"0480f1ac",
  1509 => x"5189b53f",
  1510 => x"8a518996",
  1511 => x"3f800bb0",
  1512 => x"0c833d0d",
  1513 => x"0480f1b4",
  1514 => x"5189a13f",
  1515 => x"8a518982",
  1516 => x"3f800bb0",
  1517 => x"0c833d0d",
  1518 => x"0480f1bc",
  1519 => x"51898d3f",
  1520 => x"8a5188ee",
  1521 => x"3f800bb0",
  1522 => x"0c833d0d",
  1523 => x"04fe3d0d",
  1524 => x"80f5d408",
  1525 => x"84110880",
  1526 => x"f1c45354",
  1527 => x"5288ed3f",
  1528 => x"72822a81",
  1529 => x"06518aba",
  1530 => x"3f80f1d4",
  1531 => x"5188dd3f",
  1532 => x"72812a81",
  1533 => x"06518aaa",
  1534 => x"3f80f1e8",
  1535 => x"5188cd3f",
  1536 => x"72810651",
  1537 => x"8a9c3f8a",
  1538 => x"5188a73f",
  1539 => x"72b00c84",
  1540 => x"3d0d04fe",
  1541 => x"3d0d0293",
  1542 => x"05330284",
  1543 => x"05970533",
  1544 => x"80f5d408",
  1545 => x"55535180",
  1546 => x"730c7688",
  1547 => x"140c7083",
  1548 => x"2b72078c",
  1549 => x"140c7208",
  1550 => x"5170fb38",
  1551 => x"70b00c84",
  1552 => x"3d0d04fe",
  1553 => x"3d0d80f1",
  1554 => x"fc518880",
  1555 => x"3f80f5d4",
  1556 => x"08a41108",
  1557 => x"53538451",
  1558 => x"88953f80",
  1559 => x"f5d408a0",
  1560 => x"11085353",
  1561 => x"a0518887",
  1562 => x"3f80f294",
  1563 => x"5187dd3f",
  1564 => x"80f5d408",
  1565 => x"ac110853",
  1566 => x"53845187",
  1567 => x"f23f80f5",
  1568 => x"d408a811",
  1569 => x"085353a0",
  1570 => x"5187e43f",
  1571 => x"80f2ac51",
  1572 => x"87ba3f80",
  1573 => x"f5d40898",
  1574 => x"11085353",
  1575 => x"845187cf",
  1576 => x"3f80f5d4",
  1577 => x"08941108",
  1578 => x"5353a051",
  1579 => x"87c13f80",
  1580 => x"f2c45187",
  1581 => x"973f80f5",
  1582 => x"d408b411",
  1583 => x"08535384",
  1584 => x"5187ac3f",
  1585 => x"80f5d408",
  1586 => x"b0110853",
  1587 => x"53a05187",
  1588 => x"9e3f8a51",
  1589 => x"86dc3f80",
  1590 => x"0bb00c84",
  1591 => x"3d0d04fc",
  1592 => x"3d0d80f5",
  1593 => x"d4089c11",
  1594 => x"087081ff",
  1595 => x"0680e6f4",
  1596 => x"54575353",
  1597 => x"86d63f74",
  1598 => x"5188a73f",
  1599 => x"8a5186b2",
  1600 => x"3f800bff",
  1601 => x"16555372",
  1602 => x"7425a238",
  1603 => x"72101080",
  1604 => x"f5d00805",
  1605 => x"70085252",
  1606 => x"88883f8a",
  1607 => x"5186933f",
  1608 => x"81137081",
  1609 => x"ff065452",
  1610 => x"737324e0",
  1611 => x"3874b00c",
  1612 => x"863d0d04",
  1613 => x"fc3d0d81",
  1614 => x"51e59e3f",
  1615 => x"b00881ff",
  1616 => x"06528251",
  1617 => x"e6c53fb0",
  1618 => x"0881ff06",
  1619 => x"538351e6",
  1620 => x"ba3fb008",
  1621 => x"80f5d408",
  1622 => x"55558074",
  1623 => x"0cb00888",
  1624 => x"150c7183",
  1625 => x"2b73078c",
  1626 => x"150c7308",
  1627 => x"5271fb38",
  1628 => x"74b00c86",
  1629 => x"3d0d04ff",
  1630 => x"3d0d8151",
  1631 => x"e4db3f80",
  1632 => x"f5d408b0",
  1633 => x"0890120c",
  1634 => x"5282720c",
  1635 => x"833d0d04",
  1636 => x"803d0d80",
  1637 => x"f5d40851",
  1638 => x"80710c70",
  1639 => x"b00c823d",
  1640 => x"0d04fb3d",
  1641 => x"0d8151e4",
  1642 => x"b03fb008",
  1643 => x"81ff0656",
  1644 => x"800b80f5",
  1645 => x"d4085555",
  1646 => x"80740c86",
  1647 => x"8fdff7fa",
  1648 => x"0b88150c",
  1649 => x"74832b8c",
  1650 => x"150c7308",
  1651 => x"5372fb38",
  1652 => x"81157081",
  1653 => x"ff065652",
  1654 => x"a27527dc",
  1655 => x"3872740c",
  1656 => x"868fdff7",
  1657 => x"fa0b8815",
  1658 => x"0c75832b",
  1659 => x"82078c15",
  1660 => x"0c730852",
  1661 => x"71fb3871",
  1662 => x"b00c873d",
  1663 => x"0d04fd3d",
  1664 => x"0d800b80",
  1665 => x"f5d40854",
  1666 => x"5480730c",
  1667 => x"880a0b88",
  1668 => x"140c7383",
  1669 => x"2b81078c",
  1670 => x"140c7208",
  1671 => x"5271fb38",
  1672 => x"81147081",
  1673 => x"ff065551",
  1674 => x"a27427dd",
  1675 => x"3871b00c",
  1676 => x"853d0d04",
  1677 => x"ff3d0d02",
  1678 => x"8f053351",
  1679 => x"709f269d",
  1680 => x"3880f5d4",
  1681 => x"0881722b",
  1682 => x"b0120c52",
  1683 => x"800bb413",
  1684 => x"0c89720c",
  1685 => x"b01208b0",
  1686 => x"0c833d0d",
  1687 => x"0480f5d4",
  1688 => x"0852800b",
  1689 => x"b0130ce0",
  1690 => x"1181712b",
  1691 => x"b4140c51",
  1692 => x"89720cb0",
  1693 => x"1208b00c",
  1694 => x"833d0d04",
  1695 => x"ff3d0d02",
  1696 => x"8f053380",
  1697 => x"f5d40853",
  1698 => x"5180720c",
  1699 => x"810b8813",
  1700 => x"0c70832b",
  1701 => x"82078c13",
  1702 => x"0c710851",
  1703 => x"70fb3881",
  1704 => x"0bb00c83",
  1705 => x"3d0d04db",
  1706 => x"f73f04fb",
  1707 => x"3d0d7779",
  1708 => x"55558056",
  1709 => x"757524ab",
  1710 => x"38807424",
  1711 => x"9d388053",
  1712 => x"73527451",
  1713 => x"80e13fb0",
  1714 => x"08547580",
  1715 => x"2e8538b0",
  1716 => x"08305473",
  1717 => x"b00c873d",
  1718 => x"0d047330",
  1719 => x"76813257",
  1720 => x"54dc3974",
  1721 => x"30558156",
  1722 => x"738025d2",
  1723 => x"38ec39fa",
  1724 => x"3d0d787a",
  1725 => x"57558057",
  1726 => x"767524a4",
  1727 => x"38759f2c",
  1728 => x"54815375",
  1729 => x"74327431",
  1730 => x"5274519b",
  1731 => x"3fb00854",
  1732 => x"76802e85",
  1733 => x"38b00830",
  1734 => x"5473b00c",
  1735 => x"883d0d04",
  1736 => x"74305581",
  1737 => x"57d739fc",
  1738 => x"3d0d7678",
  1739 => x"53548153",
  1740 => x"80747326",
  1741 => x"52557280",
  1742 => x"2e983870",
  1743 => x"802ea938",
  1744 => x"807224a4",
  1745 => x"38711073",
  1746 => x"10757226",
  1747 => x"53545272",
  1748 => x"ea387351",
  1749 => x"78833874",
  1750 => x"5170b00c",
  1751 => x"863d0d04",
  1752 => x"72812a72",
  1753 => x"812a5353",
  1754 => x"72802ee6",
  1755 => x"38717426",
  1756 => x"ef387372",
  1757 => x"31757407",
  1758 => x"74812a74",
  1759 => x"812a5555",
  1760 => x"5654e539",
  1761 => x"10101010",
  1762 => x"10101010",
  1763 => x"10101010",
  1764 => x"10101010",
  1765 => x"10101010",
  1766 => x"10101010",
  1767 => x"10101010",
  1768 => x"10101053",
  1769 => x"51047381",
  1770 => x"ff067383",
  1771 => x"06098105",
  1772 => x"83051010",
  1773 => x"102b0772",
  1774 => x"fc060c51",
  1775 => x"51043c04",
  1776 => x"72728072",
  1777 => x"8106ff05",
  1778 => x"09720605",
  1779 => x"71105272",
  1780 => x"0a100a53",
  1781 => x"72ed3851",
  1782 => x"51535104",
  1783 => x"b008b408",
  1784 => x"b8087575",
  1785 => x"b5ef2d50",
  1786 => x"50b00856",
  1787 => x"b80cb40c",
  1788 => x"b00c5104",
  1789 => x"b008b408",
  1790 => x"b8087575",
  1791 => x"b5ab2d50",
  1792 => x"50b00856",
  1793 => x"b80cb40c",
  1794 => x"b00c5104",
  1795 => x"b008b408",
  1796 => x"b8088ebc",
  1797 => x"2db80cb4",
  1798 => x"0cb00c04",
  1799 => x"ff3d0d02",
  1800 => x"8f053380",
  1801 => x"f6840852",
  1802 => x"710c800b",
  1803 => x"b00c833d",
  1804 => x"0d04ff3d",
  1805 => x"0d028f05",
  1806 => x"3351819e",
  1807 => x"c8085271",
  1808 => x"2db00881",
  1809 => x"ff06b00c",
  1810 => x"833d0d04",
  1811 => x"fe3d0d74",
  1812 => x"70335353",
  1813 => x"71802e93",
  1814 => x"38811372",
  1815 => x"52819ec8",
  1816 => x"08535371",
  1817 => x"2d723352",
  1818 => x"71ef3884",
  1819 => x"3d0d04f4",
  1820 => x"3d0d7f02",
  1821 => x"8405bb05",
  1822 => x"33555788",
  1823 => x"0b8c3d5b",
  1824 => x"59895380",
  1825 => x"f3a85279",
  1826 => x"5185f23f",
  1827 => x"73842e80",
  1828 => x"fa387388",
  1829 => x"2e80ff38",
  1830 => x"78567390",
  1831 => x"2e80fd38",
  1832 => x"02a70558",
  1833 => x"768f0654",
  1834 => x"73892680",
  1835 => x"c2387518",
  1836 => x"b0155555",
  1837 => x"73753476",
  1838 => x"842aff17",
  1839 => x"7081ff06",
  1840 => x"58555775",
  1841 => x"df38781a",
  1842 => x"55757534",
  1843 => x"79703355",
  1844 => x"5573802e",
  1845 => x"93388115",
  1846 => x"7452819e",
  1847 => x"c8085755",
  1848 => x"752d7433",
  1849 => x"5473ef38",
  1850 => x"78b00c8e",
  1851 => x"3d0d0475",
  1852 => x"18b71555",
  1853 => x"55737534",
  1854 => x"76842aff",
  1855 => x"177081ff",
  1856 => x"06585557",
  1857 => x"75ff9d38",
  1858 => x"ffbc3981",
  1859 => x"70575902",
  1860 => x"a70558ff",
  1861 => x"8f398270",
  1862 => x"5759f439",
  1863 => x"84705759",
  1864 => x"ee39f13d",
  1865 => x"0d618d3d",
  1866 => x"705b5c5a",
  1867 => x"807a5657",
  1868 => x"767a2481",
  1869 => x"85387817",
  1870 => x"548a5274",
  1871 => x"51848c3f",
  1872 => x"b008b005",
  1873 => x"53727434",
  1874 => x"8117578a",
  1875 => x"52745183",
  1876 => x"d53fb008",
  1877 => x"55b008de",
  1878 => x"38b00877",
  1879 => x"9f2a1870",
  1880 => x"812c5a56",
  1881 => x"56807825",
  1882 => x"9e387817",
  1883 => x"ff055575",
  1884 => x"19703355",
  1885 => x"53743373",
  1886 => x"34737534",
  1887 => x"8116ff16",
  1888 => x"56567776",
  1889 => x"24e93876",
  1890 => x"19588078",
  1891 => x"34807a24",
  1892 => x"177081ff",
  1893 => x"067c7033",
  1894 => x"56575556",
  1895 => x"72802e93",
  1896 => x"38811573",
  1897 => x"52819ec8",
  1898 => x"08585576",
  1899 => x"2d743353",
  1900 => x"72ef3873",
  1901 => x"b00c913d",
  1902 => x"0d04ad7b",
  1903 => x"3402ad05",
  1904 => x"7a307119",
  1905 => x"5656598a",
  1906 => x"52745182",
  1907 => x"fe3fb008",
  1908 => x"b0055372",
  1909 => x"74348117",
  1910 => x"578a5274",
  1911 => x"5182c73f",
  1912 => x"b00855b0",
  1913 => x"08fecf38",
  1914 => x"feef39fd",
  1915 => x"3d0d0297",
  1916 => x"05330284",
  1917 => x"059b0533",
  1918 => x"55537274",
  1919 => x"279738a0",
  1920 => x"51819ec8",
  1921 => x"0852712d",
  1922 => x"81137081",
  1923 => x"ff065452",
  1924 => x"737326eb",
  1925 => x"38853d0d",
  1926 => x"04ff3d0d",
  1927 => x"80f5f808",
  1928 => x"74101570",
  1929 => x"822b9413",
  1930 => x"0c525285",
  1931 => x"0b98130c",
  1932 => x"98120870",
  1933 => x"81065151",
  1934 => x"70f63883",
  1935 => x"3d0d04fd",
  1936 => x"3d0d80f5",
  1937 => x"f8087680",
  1938 => x"e1d42994",
  1939 => x"120c5485",
  1940 => x"0b98150c",
  1941 => x"98140870",
  1942 => x"81065153",
  1943 => x"72f63885",
  1944 => x"3d0d0480",
  1945 => x"3d0d80f5",
  1946 => x"f8085187",
  1947 => x"0b84120c",
  1948 => x"ff0ba412",
  1949 => x"0ca70ba8",
  1950 => x"120c80e1",
  1951 => x"d40b9412",
  1952 => x"0c870b98",
  1953 => x"120c823d",
  1954 => x"0d04803d",
  1955 => x"0d80f5fc",
  1956 => x"085180ec",
  1957 => x"0b8c120c",
  1958 => x"830b8812",
  1959 => x"0c823d0d",
  1960 => x"04803d0d",
  1961 => x"80f5fc08",
  1962 => x"84110881",
  1963 => x"06b00c51",
  1964 => x"823d0d04",
  1965 => x"ff3d0d80",
  1966 => x"f5fc0852",
  1967 => x"84120870",
  1968 => x"81065151",
  1969 => x"70802ef4",
  1970 => x"38710870",
  1971 => x"81ff06b0",
  1972 => x"0c51833d",
  1973 => x"0d04fe3d",
  1974 => x"0d029305",
  1975 => x"3353728a",
  1976 => x"2e9c3880",
  1977 => x"f5fc0852",
  1978 => x"84120870",
  1979 => x"892a7081",
  1980 => x"06515151",
  1981 => x"70f23872",
  1982 => x"720c843d",
  1983 => x"0d0480f5",
  1984 => x"fc085284",
  1985 => x"12087089",
  1986 => x"2a708106",
  1987 => x"51515170",
  1988 => x"f2388d72",
  1989 => x"0c841208",
  1990 => x"70892a70",
  1991 => x"81065151",
  1992 => x"5170c538",
  1993 => x"d239bc08",
  1994 => x"02bc0cfd",
  1995 => x"3d0d8053",
  1996 => x"bc088c05",
  1997 => x"0852bc08",
  1998 => x"88050851",
  1999 => x"f7e93fb0",
  2000 => x"0870b00c",
  2001 => x"54853d0d",
  2002 => x"bc0c04bc",
  2003 => x"0802bc0c",
  2004 => x"fd3d0d81",
  2005 => x"53bc088c",
  2006 => x"050852bc",
  2007 => x"08880508",
  2008 => x"51f7c43f",
  2009 => x"b00870b0",
  2010 => x"0c54853d",
  2011 => x"0dbc0c04",
  2012 => x"803d0d86",
  2013 => x"5184963f",
  2014 => x"8151a1d3",
  2015 => x"3ffc3d0d",
  2016 => x"7670797b",
  2017 => x"55555555",
  2018 => x"8f72278c",
  2019 => x"38727507",
  2020 => x"83065170",
  2021 => x"802ea738",
  2022 => x"ff125271",
  2023 => x"ff2e9838",
  2024 => x"72708105",
  2025 => x"54337470",
  2026 => x"81055634",
  2027 => x"ff125271",
  2028 => x"ff2e0981",
  2029 => x"06ea3874",
  2030 => x"b00c863d",
  2031 => x"0d047451",
  2032 => x"72708405",
  2033 => x"54087170",
  2034 => x"8405530c",
  2035 => x"72708405",
  2036 => x"54087170",
  2037 => x"8405530c",
  2038 => x"72708405",
  2039 => x"54087170",
  2040 => x"8405530c",
  2041 => x"72708405",
  2042 => x"54087170",
  2043 => x"8405530c",
  2044 => x"f0125271",
  2045 => x"8f26c938",
  2046 => x"83722795",
  2047 => x"38727084",
  2048 => x"05540871",
  2049 => x"70840553",
  2050 => x"0cfc1252",
  2051 => x"718326ed",
  2052 => x"387054ff",
  2053 => x"8339fd3d",
  2054 => x"0d755384",
  2055 => x"d8130880",
  2056 => x"2e8a3880",
  2057 => x"5372b00c",
  2058 => x"853d0d04",
  2059 => x"81805272",
  2060 => x"518d9b3f",
  2061 => x"b00884d8",
  2062 => x"140cff53",
  2063 => x"b008802e",
  2064 => x"e438b008",
  2065 => x"549f5380",
  2066 => x"74708405",
  2067 => x"560cff13",
  2068 => x"53807324",
  2069 => x"ce388074",
  2070 => x"70840556",
  2071 => x"0cff1353",
  2072 => x"728025e3",
  2073 => x"38ffbc39",
  2074 => x"fd3d0d75",
  2075 => x"7755539f",
  2076 => x"74278d38",
  2077 => x"96730cff",
  2078 => x"5271b00c",
  2079 => x"853d0d04",
  2080 => x"84d81308",
  2081 => x"5271802e",
  2082 => x"93387310",
  2083 => x"10127008",
  2084 => x"79720c51",
  2085 => x"5271b00c",
  2086 => x"853d0d04",
  2087 => x"7251fef6",
  2088 => x"3fff52b0",
  2089 => x"08d33884",
  2090 => x"d8130874",
  2091 => x"10101170",
  2092 => x"087a720c",
  2093 => x"515152dd",
  2094 => x"39f93d0d",
  2095 => x"797b5856",
  2096 => x"769f2680",
  2097 => x"e83884d8",
  2098 => x"16085473",
  2099 => x"802eaa38",
  2100 => x"76101014",
  2101 => x"70085555",
  2102 => x"73802eba",
  2103 => x"38805873",
  2104 => x"812e8f38",
  2105 => x"73ff2ea3",
  2106 => x"3880750c",
  2107 => x"7651732d",
  2108 => x"805877b0",
  2109 => x"0c893d0d",
  2110 => x"047551fe",
  2111 => x"993fff58",
  2112 => x"b008ef38",
  2113 => x"84d81608",
  2114 => x"54c63996",
  2115 => x"760c810b",
  2116 => x"b00c893d",
  2117 => x"0d047551",
  2118 => x"81ed3f76",
  2119 => x"53b00852",
  2120 => x"755181ad",
  2121 => x"3fb008b0",
  2122 => x"0c893d0d",
  2123 => x"0496760c",
  2124 => x"ff0bb00c",
  2125 => x"893d0d04",
  2126 => x"fc3d0d76",
  2127 => x"785653ff",
  2128 => x"54749f26",
  2129 => x"b13884d8",
  2130 => x"13085271",
  2131 => x"802eae38",
  2132 => x"74101012",
  2133 => x"70085353",
  2134 => x"81547180",
  2135 => x"2e983882",
  2136 => x"5471ff2e",
  2137 => x"91388354",
  2138 => x"71812e8a",
  2139 => x"3880730c",
  2140 => x"7451712d",
  2141 => x"805473b0",
  2142 => x"0c863d0d",
  2143 => x"047251fd",
  2144 => x"953fb008",
  2145 => x"f13884d8",
  2146 => x"130852c4",
  2147 => x"39ff3d0d",
  2148 => x"735280f6",
  2149 => x"880851fe",
  2150 => x"a03f833d",
  2151 => x"0d04fe3d",
  2152 => x"0d755374",
  2153 => x"5280f688",
  2154 => x"0851fdbc",
  2155 => x"3f843d0d",
  2156 => x"04803d0d",
  2157 => x"80f68808",
  2158 => x"51fcdb3f",
  2159 => x"823d0d04",
  2160 => x"ff3d0d73",
  2161 => x"5280f688",
  2162 => x"0851feec",
  2163 => x"3f833d0d",
  2164 => x"04fc3d0d",
  2165 => x"800b819e",
  2166 => x"d00c7852",
  2167 => x"77519caa",
  2168 => x"3fb00854",
  2169 => x"b008ff2e",
  2170 => x"883873b0",
  2171 => x"0c863d0d",
  2172 => x"04819ed0",
  2173 => x"08557480",
  2174 => x"2ef03876",
  2175 => x"75710c53",
  2176 => x"73b00c86",
  2177 => x"3d0d049b",
  2178 => x"fc3f04fc",
  2179 => x"3d0d7670",
  2180 => x"79707307",
  2181 => x"83065454",
  2182 => x"54557080",
  2183 => x"c3387170",
  2184 => x"08700970",
  2185 => x"f7fbfdff",
  2186 => x"130670f8",
  2187 => x"84828180",
  2188 => x"06515153",
  2189 => x"535470a6",
  2190 => x"38841472",
  2191 => x"74708405",
  2192 => x"560c7008",
  2193 => x"700970f7",
  2194 => x"fbfdff13",
  2195 => x"0670f884",
  2196 => x"82818006",
  2197 => x"51515353",
  2198 => x"5470802e",
  2199 => x"dc387352",
  2200 => x"71708105",
  2201 => x"53335170",
  2202 => x"73708105",
  2203 => x"553470f0",
  2204 => x"3874b00c",
  2205 => x"863d0d04",
  2206 => x"fd3d0d75",
  2207 => x"70718306",
  2208 => x"53555270",
  2209 => x"b8387170",
  2210 => x"087009f7",
  2211 => x"fbfdff12",
  2212 => x"0670f884",
  2213 => x"82818006",
  2214 => x"51515253",
  2215 => x"709d3884",
  2216 => x"13700870",
  2217 => x"09f7fbfd",
  2218 => x"ff120670",
  2219 => x"f8848281",
  2220 => x"80065151",
  2221 => x"52537080",
  2222 => x"2ee53872",
  2223 => x"52713351",
  2224 => x"70802e8a",
  2225 => x"38811270",
  2226 => x"33525270",
  2227 => x"f8387174",
  2228 => x"31b00c85",
  2229 => x"3d0d04fa",
  2230 => x"3d0d787a",
  2231 => x"7c705455",
  2232 => x"55527280",
  2233 => x"2e80d938",
  2234 => x"71740783",
  2235 => x"06517080",
  2236 => x"2e80d438",
  2237 => x"ff135372",
  2238 => x"ff2eb138",
  2239 => x"71337433",
  2240 => x"56517471",
  2241 => x"2e098106",
  2242 => x"a9387280",
  2243 => x"2e818738",
  2244 => x"7081ff06",
  2245 => x"5170802e",
  2246 => x"80fc3881",
  2247 => x"128115ff",
  2248 => x"15555552",
  2249 => x"72ff2e09",
  2250 => x"8106d138",
  2251 => x"71337433",
  2252 => x"56517081",
  2253 => x"ff067581",
  2254 => x"ff067171",
  2255 => x"31515252",
  2256 => x"70b00c88",
  2257 => x"3d0d0471",
  2258 => x"74575583",
  2259 => x"73278838",
  2260 => x"71087408",
  2261 => x"2e883874",
  2262 => x"765552ff",
  2263 => x"9739fc13",
  2264 => x"5372802e",
  2265 => x"b1387408",
  2266 => x"7009f7fb",
  2267 => x"fdff1206",
  2268 => x"70f88482",
  2269 => x"81800651",
  2270 => x"5151709a",
  2271 => x"38841584",
  2272 => x"17575583",
  2273 => x"7327d038",
  2274 => x"74087608",
  2275 => x"2ed03874",
  2276 => x"765552fe",
  2277 => x"df39800b",
  2278 => x"b00c883d",
  2279 => x"0d04f33d",
  2280 => x"0d606264",
  2281 => x"725a5a5e",
  2282 => x"5e805c76",
  2283 => x"70810558",
  2284 => x"3380f3bd",
  2285 => x"11337083",
  2286 => x"2a708106",
  2287 => x"51555556",
  2288 => x"72e93875",
  2289 => x"ad2e8288",
  2290 => x"3875ab2e",
  2291 => x"82843877",
  2292 => x"30707907",
  2293 => x"80257990",
  2294 => x"32703070",
  2295 => x"72078025",
  2296 => x"73075357",
  2297 => x"57515372",
  2298 => x"802e8738",
  2299 => x"75b02e81",
  2300 => x"eb38778a",
  2301 => x"38885875",
  2302 => x"b02e8338",
  2303 => x"8a58810a",
  2304 => x"5a7b8438",
  2305 => x"fe0a5a77",
  2306 => x"527951f6",
  2307 => x"be3fb008",
  2308 => x"78537a52",
  2309 => x"5bf68f3f",
  2310 => x"b0085a80",
  2311 => x"7080f3bd",
  2312 => x"18337082",
  2313 => x"2a708106",
  2314 => x"5156565a",
  2315 => x"5572802e",
  2316 => x"80c138d0",
  2317 => x"16567578",
  2318 => x"2580d738",
  2319 => x"80792475",
  2320 => x"7b260753",
  2321 => x"72933874",
  2322 => x"7a2e80eb",
  2323 => x"387a7625",
  2324 => x"80ed3872",
  2325 => x"802e80e7",
  2326 => x"38ff7770",
  2327 => x"81055933",
  2328 => x"575980f3",
  2329 => x"bd163370",
  2330 => x"822a7081",
  2331 => x"06515454",
  2332 => x"72c13873",
  2333 => x"83065372",
  2334 => x"802e9738",
  2335 => x"738106c9",
  2336 => x"17555372",
  2337 => x"8538ffa9",
  2338 => x"16547356",
  2339 => x"777624ff",
  2340 => x"ab388079",
  2341 => x"2480f038",
  2342 => x"7b802e84",
  2343 => x"38743055",
  2344 => x"7c802e8c",
  2345 => x"38ff1753",
  2346 => x"7883387d",
  2347 => x"53727d0c",
  2348 => x"74b00c8f",
  2349 => x"3d0d0481",
  2350 => x"53757b24",
  2351 => x"ff953881",
  2352 => x"75792917",
  2353 => x"78708105",
  2354 => x"5a335856",
  2355 => x"59ff9339",
  2356 => x"815c7670",
  2357 => x"81055833",
  2358 => x"56fdf439",
  2359 => x"80773354",
  2360 => x"547280f8",
  2361 => x"2eb23872",
  2362 => x"80d83270",
  2363 => x"30708025",
  2364 => x"76075151",
  2365 => x"5372802e",
  2366 => x"fdf83881",
  2367 => x"17338218",
  2368 => x"58569058",
  2369 => x"fdf83981",
  2370 => x"0a557b84",
  2371 => x"38fe0a55",
  2372 => x"7f53a273",
  2373 => x"0cff8939",
  2374 => x"8154cc39",
  2375 => x"fd3d0d77",
  2376 => x"54765375",
  2377 => x"5280f688",
  2378 => x"0851fcf2",
  2379 => x"3f853d0d",
  2380 => x"04f33d0d",
  2381 => x"60626472",
  2382 => x"5a5a5d5d",
  2383 => x"805e7670",
  2384 => x"81055833",
  2385 => x"80f3bd11",
  2386 => x"3370832a",
  2387 => x"70810651",
  2388 => x"55555672",
  2389 => x"e93875ad",
  2390 => x"2e81ff38",
  2391 => x"75ab2e81",
  2392 => x"fb387730",
  2393 => x"70790780",
  2394 => x"25799032",
  2395 => x"70307072",
  2396 => x"07802573",
  2397 => x"07535757",
  2398 => x"51537280",
  2399 => x"2e873875",
  2400 => x"b02e81e2",
  2401 => x"38778a38",
  2402 => x"885875b0",
  2403 => x"2e83388a",
  2404 => x"587752ff",
  2405 => x"51f38f3f",
  2406 => x"b0087853",
  2407 => x"5aff51f3",
  2408 => x"aa3fb008",
  2409 => x"5b80705a",
  2410 => x"5580f3bd",
  2411 => x"16337082",
  2412 => x"2a708106",
  2413 => x"51545472",
  2414 => x"802e80c1",
  2415 => x"38d01656",
  2416 => x"75782580",
  2417 => x"d7388079",
  2418 => x"24757b26",
  2419 => x"07537293",
  2420 => x"38747a2e",
  2421 => x"80eb387a",
  2422 => x"762580ed",
  2423 => x"3872802e",
  2424 => x"80e738ff",
  2425 => x"77708105",
  2426 => x"59335759",
  2427 => x"80f3bd16",
  2428 => x"3370822a",
  2429 => x"70810651",
  2430 => x"545472c1",
  2431 => x"38738306",
  2432 => x"5372802e",
  2433 => x"97387381",
  2434 => x"06c91755",
  2435 => x"53728538",
  2436 => x"ffa91654",
  2437 => x"73567776",
  2438 => x"24ffab38",
  2439 => x"80792481",
  2440 => x"89387d80",
  2441 => x"2e843874",
  2442 => x"30557b80",
  2443 => x"2e8c38ff",
  2444 => x"17537883",
  2445 => x"387c5372",
  2446 => x"7c0c74b0",
  2447 => x"0c8f3d0d",
  2448 => x"04815375",
  2449 => x"7b24ff95",
  2450 => x"38817579",
  2451 => x"29177870",
  2452 => x"81055a33",
  2453 => x"585659ff",
  2454 => x"9339815e",
  2455 => x"76708105",
  2456 => x"583356fd",
  2457 => x"fd398077",
  2458 => x"33545472",
  2459 => x"80f82e80",
  2460 => x"c3387280",
  2461 => x"d8327030",
  2462 => x"70802576",
  2463 => x"07515153",
  2464 => x"72802efe",
  2465 => x"80388117",
  2466 => x"33821858",
  2467 => x"56907053",
  2468 => x"58ff51f1",
  2469 => x"913fb008",
  2470 => x"78535aff",
  2471 => x"51f1ac3f",
  2472 => x"b0085b80",
  2473 => x"705a55fe",
  2474 => x"8039ff60",
  2475 => x"5455a273",
  2476 => x"0cfef739",
  2477 => x"8154ffba",
  2478 => x"39fd3d0d",
  2479 => x"77547653",
  2480 => x"755280f6",
  2481 => x"880851fc",
  2482 => x"e83f853d",
  2483 => x"0d04f33d",
  2484 => x"0d7f618b",
  2485 => x"1170f806",
  2486 => x"5c55555e",
  2487 => x"72962683",
  2488 => x"38905980",
  2489 => x"7924747a",
  2490 => x"26075380",
  2491 => x"5472742e",
  2492 => x"09810680",
  2493 => x"cb387d51",
  2494 => x"8bca3f78",
  2495 => x"83f72680",
  2496 => x"c6387883",
  2497 => x"2a701010",
  2498 => x"1080fdc4",
  2499 => x"058c1108",
  2500 => x"59595a76",
  2501 => x"782e83b0",
  2502 => x"38841708",
  2503 => x"fc06568c",
  2504 => x"17088818",
  2505 => x"08718c12",
  2506 => x"0c88120c",
  2507 => x"58751784",
  2508 => x"11088107",
  2509 => x"84120c53",
  2510 => x"7d518b89",
  2511 => x"3f881754",
  2512 => x"73b00c8f",
  2513 => x"3d0d0478",
  2514 => x"892a7983",
  2515 => x"2a5b5372",
  2516 => x"802ebf38",
  2517 => x"78862ab8",
  2518 => x"055a8473",
  2519 => x"27b43880",
  2520 => x"db135a94",
  2521 => x"7327ab38",
  2522 => x"788c2a80",
  2523 => x"ee055a80",
  2524 => x"d473279e",
  2525 => x"38788f2a",
  2526 => x"80f7055a",
  2527 => x"82d47327",
  2528 => x"91387892",
  2529 => x"2a80fc05",
  2530 => x"5a8ad473",
  2531 => x"27843880",
  2532 => x"fe5a7910",
  2533 => x"101080fd",
  2534 => x"c4058c11",
  2535 => x"08585576",
  2536 => x"752ea338",
  2537 => x"841708fc",
  2538 => x"06707a31",
  2539 => x"5556738f",
  2540 => x"2488d538",
  2541 => x"738025fe",
  2542 => x"e6388c17",
  2543 => x"08577675",
  2544 => x"2e098106",
  2545 => x"df38811a",
  2546 => x"5a80fdd4",
  2547 => x"08577680",
  2548 => x"fdcc2e82",
  2549 => x"c0388417",
  2550 => x"08fc0670",
  2551 => x"7a315556",
  2552 => x"738f2481",
  2553 => x"f93880fd",
  2554 => x"cc0b80fd",
  2555 => x"d80c80fd",
  2556 => x"cc0b80fd",
  2557 => x"d40c7380",
  2558 => x"25feb238",
  2559 => x"83ff7627",
  2560 => x"83df3875",
  2561 => x"892a7683",
  2562 => x"2a555372",
  2563 => x"802ebf38",
  2564 => x"75862ab8",
  2565 => x"05548473",
  2566 => x"27b43880",
  2567 => x"db135494",
  2568 => x"7327ab38",
  2569 => x"758c2a80",
  2570 => x"ee055480",
  2571 => x"d473279e",
  2572 => x"38758f2a",
  2573 => x"80f70554",
  2574 => x"82d47327",
  2575 => x"91387592",
  2576 => x"2a80fc05",
  2577 => x"548ad473",
  2578 => x"27843880",
  2579 => x"fe547310",
  2580 => x"101080fd",
  2581 => x"c4058811",
  2582 => x"08565874",
  2583 => x"782e86cf",
  2584 => x"38841508",
  2585 => x"fc065375",
  2586 => x"73278d38",
  2587 => x"88150855",
  2588 => x"74782e09",
  2589 => x"8106ea38",
  2590 => x"8c150880",
  2591 => x"fdc40b84",
  2592 => x"0508718c",
  2593 => x"1a0c7688",
  2594 => x"1a0c7888",
  2595 => x"130c788c",
  2596 => x"180c5d58",
  2597 => x"7953807a",
  2598 => x"2483e638",
  2599 => x"72822c81",
  2600 => x"712b5c53",
  2601 => x"7a7c2681",
  2602 => x"98387b7b",
  2603 => x"06537282",
  2604 => x"f13879fc",
  2605 => x"0684055a",
  2606 => x"7a10707d",
  2607 => x"06545b72",
  2608 => x"82e03884",
  2609 => x"1a5af139",
  2610 => x"88178c11",
  2611 => x"08585876",
  2612 => x"782e0981",
  2613 => x"06fcc238",
  2614 => x"821a5afd",
  2615 => x"ec397817",
  2616 => x"79810784",
  2617 => x"190c7080",
  2618 => x"fdd80c70",
  2619 => x"80fdd40c",
  2620 => x"80fdcc0b",
  2621 => x"8c120c8c",
  2622 => x"11088812",
  2623 => x"0c748107",
  2624 => x"84120c74",
  2625 => x"1175710c",
  2626 => x"51537d51",
  2627 => x"87b73f88",
  2628 => x"1754fcac",
  2629 => x"3980fdc4",
  2630 => x"0b840508",
  2631 => x"7a545c79",
  2632 => x"8025fef8",
  2633 => x"3882da39",
  2634 => x"7a097c06",
  2635 => x"7080fdc4",
  2636 => x"0b84050c",
  2637 => x"5c7a105b",
  2638 => x"7a7c2685",
  2639 => x"387a85b8",
  2640 => x"3880fdc4",
  2641 => x"0b880508",
  2642 => x"70841208",
  2643 => x"fc06707c",
  2644 => x"317c7226",
  2645 => x"8f722507",
  2646 => x"57575c5d",
  2647 => x"5572802e",
  2648 => x"80db3879",
  2649 => x"7a1680fd",
  2650 => x"bc081b90",
  2651 => x"115a5557",
  2652 => x"5b80fdb8",
  2653 => x"08ff2e88",
  2654 => x"38a08f13",
  2655 => x"e0800657",
  2656 => x"76527d51",
  2657 => x"86c03fb0",
  2658 => x"0854b008",
  2659 => x"ff2e9038",
  2660 => x"b0087627",
  2661 => x"82993874",
  2662 => x"80fdc42e",
  2663 => x"82913880",
  2664 => x"fdc40b88",
  2665 => x"05085584",
  2666 => x"1508fc06",
  2667 => x"707a317a",
  2668 => x"72268f72",
  2669 => x"25075255",
  2670 => x"537283e6",
  2671 => x"38747981",
  2672 => x"0784170c",
  2673 => x"79167080",
  2674 => x"fdc40b88",
  2675 => x"050c7581",
  2676 => x"0784120c",
  2677 => x"547e5257",
  2678 => x"85eb3f88",
  2679 => x"1754fae0",
  2680 => x"3975832a",
  2681 => x"70545480",
  2682 => x"7424819b",
  2683 => x"3872822c",
  2684 => x"81712b80",
  2685 => x"fdc80807",
  2686 => x"7080fdc4",
  2687 => x"0b84050c",
  2688 => x"75101010",
  2689 => x"80fdc405",
  2690 => x"88110858",
  2691 => x"5a5d5377",
  2692 => x"8c180c74",
  2693 => x"88180c76",
  2694 => x"88190c76",
  2695 => x"8c160cfc",
  2696 => x"f339797a",
  2697 => x"10101080",
  2698 => x"fdc40570",
  2699 => x"57595d8c",
  2700 => x"15085776",
  2701 => x"752ea338",
  2702 => x"841708fc",
  2703 => x"06707a31",
  2704 => x"5556738f",
  2705 => x"2483ca38",
  2706 => x"73802584",
  2707 => x"81388c17",
  2708 => x"08577675",
  2709 => x"2e098106",
  2710 => x"df388815",
  2711 => x"811b7083",
  2712 => x"06555b55",
  2713 => x"72c9387c",
  2714 => x"83065372",
  2715 => x"802efdb8",
  2716 => x"38ff1df8",
  2717 => x"19595d88",
  2718 => x"1808782e",
  2719 => x"ea38fdb5",
  2720 => x"39831a53",
  2721 => x"fc963983",
  2722 => x"1470822c",
  2723 => x"81712b80",
  2724 => x"fdc80807",
  2725 => x"7080fdc4",
  2726 => x"0b84050c",
  2727 => x"76101010",
  2728 => x"80fdc405",
  2729 => x"88110859",
  2730 => x"5b5e5153",
  2731 => x"fee13980",
  2732 => x"fd880817",
  2733 => x"58b00876",
  2734 => x"2e818d38",
  2735 => x"80fdb808",
  2736 => x"ff2e83ec",
  2737 => x"38737631",
  2738 => x"1880fd88",
  2739 => x"0c738706",
  2740 => x"70575372",
  2741 => x"802e8838",
  2742 => x"88733170",
  2743 => x"15555676",
  2744 => x"149fff06",
  2745 => x"a0807131",
  2746 => x"1770547f",
  2747 => x"53575383",
  2748 => x"d53fb008",
  2749 => x"53b008ff",
  2750 => x"2e81a038",
  2751 => x"80fd8808",
  2752 => x"167080fd",
  2753 => x"880c7475",
  2754 => x"80fdc40b",
  2755 => x"88050c74",
  2756 => x"76311870",
  2757 => x"81075155",
  2758 => x"56587b80",
  2759 => x"fdc42e83",
  2760 => x"9c38798f",
  2761 => x"2682cb38",
  2762 => x"810b8415",
  2763 => x"0c841508",
  2764 => x"fc06707a",
  2765 => x"317a7226",
  2766 => x"8f722507",
  2767 => x"52555372",
  2768 => x"802efcf9",
  2769 => x"3880db39",
  2770 => x"b0089fff",
  2771 => x"065372fe",
  2772 => x"eb387780",
  2773 => x"fd880c80",
  2774 => x"fdc40b88",
  2775 => x"05087b18",
  2776 => x"81078412",
  2777 => x"0c5580fd",
  2778 => x"b4087827",
  2779 => x"86387780",
  2780 => x"fdb40c80",
  2781 => x"fdb00878",
  2782 => x"27fcac38",
  2783 => x"7780fdb0",
  2784 => x"0c841508",
  2785 => x"fc06707a",
  2786 => x"317a7226",
  2787 => x"8f722507",
  2788 => x"52555372",
  2789 => x"802efca5",
  2790 => x"38883980",
  2791 => x"745456fe",
  2792 => x"db397d51",
  2793 => x"829f3f80",
  2794 => x"0bb00c8f",
  2795 => x"3d0d0473",
  2796 => x"53807424",
  2797 => x"a9387282",
  2798 => x"2c81712b",
  2799 => x"80fdc808",
  2800 => x"077080fd",
  2801 => x"c40b8405",
  2802 => x"0c5d5377",
  2803 => x"8c180c74",
  2804 => x"88180c76",
  2805 => x"88190c76",
  2806 => x"8c160cf9",
  2807 => x"b7398314",
  2808 => x"70822c81",
  2809 => x"712b80fd",
  2810 => x"c8080770",
  2811 => x"80fdc40b",
  2812 => x"84050c5e",
  2813 => x"5153d439",
  2814 => x"7b7b0653",
  2815 => x"72fca338",
  2816 => x"841a7b10",
  2817 => x"5c5af139",
  2818 => x"ff1a8111",
  2819 => x"515af7b9",
  2820 => x"39781779",
  2821 => x"81078419",
  2822 => x"0c8c1808",
  2823 => x"88190871",
  2824 => x"8c120c88",
  2825 => x"120c5970",
  2826 => x"80fdd80c",
  2827 => x"7080fdd4",
  2828 => x"0c80fdcc",
  2829 => x"0b8c120c",
  2830 => x"8c110888",
  2831 => x"120c7481",
  2832 => x"0784120c",
  2833 => x"74117571",
  2834 => x"0c5153f9",
  2835 => x"bd397517",
  2836 => x"84110881",
  2837 => x"0784120c",
  2838 => x"538c1708",
  2839 => x"88180871",
  2840 => x"8c120c88",
  2841 => x"120c587d",
  2842 => x"5180da3f",
  2843 => x"881754f5",
  2844 => x"cf397284",
  2845 => x"150cf41a",
  2846 => x"f8067084",
  2847 => x"1e088106",
  2848 => x"07841e0c",
  2849 => x"701d545b",
  2850 => x"850b8414",
  2851 => x"0c850b88",
  2852 => x"140c8f7b",
  2853 => x"27fdcf38",
  2854 => x"881c527d",
  2855 => x"5182903f",
  2856 => x"80fdc40b",
  2857 => x"88050880",
  2858 => x"fd880859",
  2859 => x"55fdb739",
  2860 => x"7780fd88",
  2861 => x"0c7380fd",
  2862 => x"b80cfc91",
  2863 => x"39728415",
  2864 => x"0cfda339",
  2865 => x"0404fd3d",
  2866 => x"0d800b81",
  2867 => x"9ed00c76",
  2868 => x"5186cb3f",
  2869 => x"b00853b0",
  2870 => x"08ff2e88",
  2871 => x"3872b00c",
  2872 => x"853d0d04",
  2873 => x"819ed008",
  2874 => x"5473802e",
  2875 => x"f0387574",
  2876 => x"710c5272",
  2877 => x"b00c853d",
  2878 => x"0d04fb3d",
  2879 => x"0d777052",
  2880 => x"56c23f80",
  2881 => x"fdc40b88",
  2882 => x"05088411",
  2883 => x"08fc0670",
  2884 => x"7b319fef",
  2885 => x"05e08006",
  2886 => x"e0800556",
  2887 => x"5653a080",
  2888 => x"74249438",
  2889 => x"80527551",
  2890 => x"ff9c3f80",
  2891 => x"fdcc0815",
  2892 => x"5372b008",
  2893 => x"2e8f3875",
  2894 => x"51ff8a3f",
  2895 => x"805372b0",
  2896 => x"0c873d0d",
  2897 => x"04733052",
  2898 => x"7551fefa",
  2899 => x"3fb008ff",
  2900 => x"2ea83880",
  2901 => x"fdc40b88",
  2902 => x"05087575",
  2903 => x"31810784",
  2904 => x"120c5380",
  2905 => x"fd880874",
  2906 => x"3180fd88",
  2907 => x"0c7551fe",
  2908 => x"d43f810b",
  2909 => x"b00c873d",
  2910 => x"0d048052",
  2911 => x"7551fec6",
  2912 => x"3f80fdc4",
  2913 => x"0b880508",
  2914 => x"b0087131",
  2915 => x"56538f75",
  2916 => x"25ffa438",
  2917 => x"b00880fd",
  2918 => x"b8083180",
  2919 => x"fd880c74",
  2920 => x"81078414",
  2921 => x"0c7551fe",
  2922 => x"9c3f8053",
  2923 => x"ff9039f6",
  2924 => x"3d0d7c7e",
  2925 => x"545b7280",
  2926 => x"2e828338",
  2927 => x"7a51fe84",
  2928 => x"3ff81384",
  2929 => x"110870fe",
  2930 => x"06701384",
  2931 => x"1108fc06",
  2932 => x"5d585954",
  2933 => x"5880fdcc",
  2934 => x"08752e82",
  2935 => x"de387884",
  2936 => x"160c8073",
  2937 => x"8106545a",
  2938 => x"727a2e81",
  2939 => x"d5387815",
  2940 => x"84110881",
  2941 => x"06515372",
  2942 => x"a0387817",
  2943 => x"577981e6",
  2944 => x"38881508",
  2945 => x"537280fd",
  2946 => x"cc2e82f9",
  2947 => x"388c1508",
  2948 => x"708c150c",
  2949 => x"7388120c",
  2950 => x"56768107",
  2951 => x"84190c76",
  2952 => x"1877710c",
  2953 => x"53798191",
  2954 => x"3883ff77",
  2955 => x"2781c838",
  2956 => x"76892a77",
  2957 => x"832a5653",
  2958 => x"72802ebf",
  2959 => x"3876862a",
  2960 => x"b8055584",
  2961 => x"7327b438",
  2962 => x"80db1355",
  2963 => x"947327ab",
  2964 => x"38768c2a",
  2965 => x"80ee0555",
  2966 => x"80d47327",
  2967 => x"9e38768f",
  2968 => x"2a80f705",
  2969 => x"5582d473",
  2970 => x"27913876",
  2971 => x"922a80fc",
  2972 => x"05558ad4",
  2973 => x"73278438",
  2974 => x"80fe5574",
  2975 => x"10101080",
  2976 => x"fdc40588",
  2977 => x"11085556",
  2978 => x"73762e82",
  2979 => x"b3388414",
  2980 => x"08fc0653",
  2981 => x"7673278d",
  2982 => x"38881408",
  2983 => x"5473762e",
  2984 => x"098106ea",
  2985 => x"388c1408",
  2986 => x"708c1a0c",
  2987 => x"74881a0c",
  2988 => x"7888120c",
  2989 => x"56778c15",
  2990 => x"0c7a51fc",
  2991 => x"883f8c3d",
  2992 => x"0d047708",
  2993 => x"78713159",
  2994 => x"77058819",
  2995 => x"08545772",
  2996 => x"80fdcc2e",
  2997 => x"80e0388c",
  2998 => x"1808708c",
  2999 => x"150c7388",
  3000 => x"120c56fe",
  3001 => x"89398815",
  3002 => x"088c1608",
  3003 => x"708c130c",
  3004 => x"5788170c",
  3005 => x"fea33976",
  3006 => x"832a7054",
  3007 => x"55807524",
  3008 => x"81983872",
  3009 => x"822c8171",
  3010 => x"2b80fdc8",
  3011 => x"080780fd",
  3012 => x"c40b8405",
  3013 => x"0c537410",
  3014 => x"101080fd",
  3015 => x"c4058811",
  3016 => x"08555675",
  3017 => x"8c190c73",
  3018 => x"88190c77",
  3019 => x"88170c77",
  3020 => x"8c150cff",
  3021 => x"8439815a",
  3022 => x"fdb43978",
  3023 => x"17738106",
  3024 => x"54577298",
  3025 => x"38770878",
  3026 => x"71315977",
  3027 => x"058c1908",
  3028 => x"881a0871",
  3029 => x"8c120c88",
  3030 => x"120c5757",
  3031 => x"76810784",
  3032 => x"190c7780",
  3033 => x"fdc40b88",
  3034 => x"050c80fd",
  3035 => x"c0087726",
  3036 => x"fec73880",
  3037 => x"fdbc0852",
  3038 => x"7a51fafe",
  3039 => x"3f7a51fa",
  3040 => x"c43ffeba",
  3041 => x"3981788c",
  3042 => x"150c7888",
  3043 => x"150c738c",
  3044 => x"1a0c7388",
  3045 => x"1a0c5afd",
  3046 => x"80398315",
  3047 => x"70822c81",
  3048 => x"712b80fd",
  3049 => x"c8080780",
  3050 => x"fdc40b84",
  3051 => x"050c5153",
  3052 => x"74101010",
  3053 => x"80fdc405",
  3054 => x"88110855",
  3055 => x"56fee439",
  3056 => x"74538075",
  3057 => x"24a73872",
  3058 => x"822c8171",
  3059 => x"2b80fdc8",
  3060 => x"080780fd",
  3061 => x"c40b8405",
  3062 => x"0c53758c",
  3063 => x"190c7388",
  3064 => x"190c7788",
  3065 => x"170c778c",
  3066 => x"150cfdcd",
  3067 => x"39831570",
  3068 => x"822c8171",
  3069 => x"2b80fdc8",
  3070 => x"080780fd",
  3071 => x"c40b8405",
  3072 => x"0c5153d6",
  3073 => x"39810bb0",
  3074 => x"0c04803d",
  3075 => x"0d72812e",
  3076 => x"8938800b",
  3077 => x"b00c823d",
  3078 => x"0d047351",
  3079 => x"b23ffe3d",
  3080 => x"0d819ecc",
  3081 => x"0851708a",
  3082 => x"38819ed4",
  3083 => x"70819ecc",
  3084 => x"0c517075",
  3085 => x"125252ff",
  3086 => x"537087fb",
  3087 => x"80802688",
  3088 => x"3870819e",
  3089 => x"cc0c7153",
  3090 => x"72b00c84",
  3091 => x"3d0d0400",
  3092 => x"ff390000",
  3093 => x"68656c70",
  3094 => x"00000000",
  3095 => x"73797374",
  3096 => x"656d2072",
  3097 => x"65736574",
  3098 => x"00000000",
  3099 => x"72657365",
  3100 => x"74000000",
  3101 => x"73686f77",
  3102 => x"20737973",
  3103 => x"74656d20",
  3104 => x"696e666f",
  3105 => x"203c7665",
  3106 => x"72626f73",
  3107 => x"653e0000",
  3108 => x"73797369",
  3109 => x"6e666f00",
  3110 => x"7265706f",
  3111 => x"72742076",
  3112 => x"65727369",
  3113 => x"6f6e0000",
  3114 => x"76657273",
  3115 => x"696f6e00",
  3116 => x"72656e61",
  3117 => x"20636f6e",
  3118 => x"74726f6c",
  3119 => x"6c657220",
  3120 => x"73746174",
  3121 => x"75730000",
  3122 => x"72656e61",
  3123 => x"20737461",
  3124 => x"74757300",
  3125 => x"3c636861",
  3126 => x"6e6e656c",
  3127 => x"3e203c68",
  3128 => x"6967683e",
  3129 => x"203c6c6f",
  3130 => x"775f636f",
  3131 => x"6e666967",
  3132 => x"3e000000",
  3133 => x"636f6e66",
  3134 => x"69670000",
  3135 => x"3c636861",
  3136 => x"6e6e656c",
  3137 => x"3e204543",
  3138 => x"414c2c20",
  3139 => x"64656d6f",
  3140 => x"20636f6e",
  3141 => x"66696720",
  3142 => x"666f7220",
  3143 => x"52454e41",
  3144 => x"00000000",
  3145 => x"64656d6f",
  3146 => x"00000000",
  3147 => x"73657420",
  3148 => x"52454e41",
  3149 => x"20746f20",
  3150 => x"706f7765",
  3151 => x"7220646f",
  3152 => x"776e206d",
  3153 => x"6f646500",
  3154 => x"706f6666",
  3155 => x"00000000",
  3156 => x"3c636861",
  3157 => x"6e6e656c",
  3158 => x"3e207365",
  3159 => x"74206120",
  3160 => x"72656e61",
  3161 => x"20746f20",
  3162 => x"666f6c6c",
  3163 => x"6f776572",
  3164 => x"206d6f64",
  3165 => x"65000000",
  3166 => x"666f6c6c",
  3167 => x"6f770000",
  3168 => x"3c636861",
  3169 => x"6e6e656c",
  3170 => x"3e20636f",
  3171 => x"6e666967",
  3172 => x"20746f20",
  3173 => x"4543414c",
  3174 => x"00000000",
  3175 => x"6563616c",
  3176 => x"00000000",
  3177 => x"3c74696d",
  3178 => x"653e2061",
  3179 => x"63746976",
  3180 => x"61746520",
  3181 => x"52454e41",
  3182 => x"00000000",
  3183 => x"61637175",
  3184 => x"69726500",
  3185 => x"73657420",
  3186 => x"52454e41",
  3187 => x"20636f6e",
  3188 => x"74726f6c",
  3189 => x"6c657220",
  3190 => x"746f2049",
  3191 => x"444c4500",
  3192 => x"73746f70",
  3193 => x"00000000",
  3194 => x"7072696e",
  3195 => x"74207472",
  3196 => x"69676765",
  3197 => x"72206368",
  3198 => x"61696e73",
  3199 => x"00000000",
  3200 => x"63686169",
  3201 => x"6e730000",
  3202 => x"7072696e",
  3203 => x"74207361",
  3204 => x"6d706c65",
  3205 => x"64205245",
  3206 => x"4e412074",
  3207 => x"6f6b656e",
  3208 => x"73000000",
  3209 => x"746f6b65",
  3210 => x"6e000000",
  3211 => x"3c636f75",
  3212 => x"6e743e20",
  3213 => x"3c74696d",
  3214 => x"653e2074",
  3215 => x"726f7562",
  3216 => x"6c657365",
  3217 => x"61726368",
  3218 => x"2052454e",
  3219 => x"41000000",
  3220 => x"74726f75",
  3221 => x"626c6500",
  3222 => x"696e6974",
  3223 => x"616c697a",
  3224 => x"65204444",
  3225 => x"53206368",
  3226 => x"6970203c",
  3227 => x"66726571",
  3228 => x"2074756e",
  3229 => x"696e6720",
  3230 => x"776f7264",
  3231 => x"3e000000",
  3232 => x"64647369",
  3233 => x"6e697400",
  3234 => x"72656164",
  3235 => x"20646473",
  3236 => x"20726567",
  3237 => x"69737465",
  3238 => x"72730000",
  3239 => x"64647369",
  3240 => x"6e666f00",
  3241 => x"67656e65",
  3242 => x"72617465",
  3243 => x"20746573",
  3244 => x"7420696d",
  3245 => x"70756c73",
  3246 => x"65000000",
  3247 => x"74657374",
  3248 => x"67656e00",
  3249 => x"72656164",
  3250 => x"20616463",
  3251 => x"2076616c",
  3252 => x"75650000",
  3253 => x"61646300",
  3254 => x"0a0a0000",
  3255 => x"72656e61",
  3256 => x"33202d20",
  3257 => x"72656164",
  3258 => x"206f7574",
  3259 => x"20656c65",
  3260 => x"6374726f",
  3261 => x"6e696300",
  3262 => x"20286f6e",
  3263 => x"2073696d",
  3264 => x"290a0000",
  3265 => x"56312e30",
  3266 => x"2d31322e",
  3267 => x"32303131",
  3268 => x"5f524f45",
  3269 => x"5f5a5055",
  3270 => x"00000000",
  3271 => x"0a485720",
  3272 => x"73796e74",
  3273 => x"68657369",
  3274 => x"7a65643a",
  3275 => x"20000000",
  3276 => x"0a535720",
  3277 => x"636f6d70",
  3278 => x"696c6564",
  3279 => x"2020203a",
  3280 => x"20466562",
  3281 => x"20313020",
  3282 => x"32303132",
  3283 => x"20203039",
  3284 => x"3a34353a",
  3285 => x"34340000",
  3286 => x"0a737973",
  3287 => x"74656d20",
  3288 => x"636c6f63",
  3289 => x"6b20203a",
  3290 => x"20000000",
  3291 => x"204d487a",
  3292 => x"0a000000",
  3293 => x"746f6b65",
  3294 => x"6e733a20",
  3295 => x"00000000",
  3296 => x"4552524f",
  3297 => x"523a2074",
  3298 => x"6f6f206d",
  3299 => x"75636820",
  3300 => x"636f6d6d",
  3301 => x"616e6473",
  3302 => x"2e0a0000",
  3303 => x"3e200000",
  3304 => x"636f6d6d",
  3305 => x"616e6420",
  3306 => x"6e6f7420",
  3307 => x"666f756e",
  3308 => x"642e0a00",
  3309 => x"66756e63",
  3310 => x"3a203078",
  3311 => x"00000000",
  3312 => x"20207265",
  3313 => x"743a2030",
  3314 => x"78000000",
  3315 => x"73757070",
  3316 => x"6f727465",
  3317 => x"6420636f",
  3318 => x"6d6d616e",
  3319 => x"64733a0a",
  3320 => x"0a000000",
  3321 => x"202d2000",
  3322 => x"76656e64",
  3323 => x"6f723f20",
  3324 => x"20000000",
  3325 => x"485a4452",
  3326 => x"20202020",
  3327 => x"20000000",
  3328 => x"67616973",
  3329 => x"6c657220",
  3330 => x"20000000",
  3331 => x"45534120",
  3332 => x"20202020",
  3333 => x"20000000",
  3334 => x"756e6b6e",
  3335 => x"6f776e20",
  3336 => x"64657669",
  3337 => x"63650000",
  3338 => x"4c656f6e",
  3339 => x"32204d65",
  3340 => x"6d6f7279",
  3341 => x"20436f6e",
  3342 => x"74726f6c",
  3343 => x"6c657200",
  3344 => x"56474120",
  3345 => x"636f6e74",
  3346 => x"726f6c6c",
  3347 => x"65720000",
  3348 => x"53504920",
  3349 => x"4d656d6f",
  3350 => x"72792043",
  3351 => x"6f6e7472",
  3352 => x"6f6c6c65",
  3353 => x"72000000",
  3354 => x"53504920",
  3355 => x"436f6e74",
  3356 => x"726f6c6c",
  3357 => x"65720000",
  3358 => x"414d4241",
  3359 => x"20577261",
  3360 => x"70706572",
  3361 => x"20666f72",
  3362 => x"204f4320",
  3363 => x"4932432d",
  3364 => x"6d617374",
  3365 => x"65720000",
  3366 => x"47522031",
  3367 => x"302f3130",
  3368 => x"30204d62",
  3369 => x"69742045",
  3370 => x"74686572",
  3371 => x"6e657420",
  3372 => x"4d414300",
  3373 => x"47656e65",
  3374 => x"72616c20",
  3375 => x"50757270",
  3376 => x"6f736520",
  3377 => x"492f4f20",
  3378 => x"706f7274",
  3379 => x"00000000",
  3380 => x"4d6f6475",
  3381 => x"6c617220",
  3382 => x"54696d65",
  3383 => x"7220556e",
  3384 => x"69740000",
  3385 => x"4475616c",
  3386 => x"2d706f72",
  3387 => x"74204148",
  3388 => x"42205352",
  3389 => x"414d206d",
  3390 => x"6f64756c",
  3391 => x"65000000",
  3392 => x"47656e65",
  3393 => x"72696320",
  3394 => x"55415254",
  3395 => x"00000000",
  3396 => x"4148422f",
  3397 => x"41504220",
  3398 => x"42726964",
  3399 => x"67650000",
  3400 => x"64696666",
  3401 => x"6572656e",
  3402 => x"7469616c",
  3403 => x"20637572",
  3404 => x"72656e74",
  3405 => x"206d6f6e",
  3406 => x"69746f72",
  3407 => x"00000000",
  3408 => x"64656275",
  3409 => x"67207472",
  3410 => x"61636572",
  3411 => x"206d656d",
  3412 => x"6f727900",
  3413 => x"4541444f",
  3414 => x"47533130",
  3415 => x"32206469",
  3416 => x"73706c61",
  3417 => x"79206472",
  3418 => x"69766572",
  3419 => x"00000000",
  3420 => x"64656275",
  3421 => x"67206275",
  3422 => x"66666572",
  3423 => x"20636f6e",
  3424 => x"74726f6c",
  3425 => x"00000000",
  3426 => x"52454e41",
  3427 => x"3320636f",
  3428 => x"6e74726f",
  3429 => x"6c6c6572",
  3430 => x"00000000",
  3431 => x"53465020",
  3432 => x"636f6e74",
  3433 => x"726f6c6c",
  3434 => x"65720000",
  3435 => x"5a505520",
  3436 => x"4d656d6f",
  3437 => x"72792077",
  3438 => x"72617070",
  3439 => x"65720000",
  3440 => x"5a505520",
  3441 => x"41484220",
  3442 => x"57726170",
  3443 => x"70657200",
  3444 => x"6265616d",
  3445 => x"20706f73",
  3446 => x"6974696f",
  3447 => x"6e206d6f",
  3448 => x"6e69746f",
  3449 => x"72000000",
  3450 => x"74726967",
  3451 => x"67657220",
  3452 => x"67656e65",
  3453 => x"7261746f",
  3454 => x"72000000",
  3455 => x"64656275",
  3456 => x"6720636f",
  3457 => x"6e736f6c",
  3458 => x"65000000",
  3459 => x"44434d20",
  3460 => x"70686173",
  3461 => x"65207368",
  3462 => x"69667420",
  3463 => x"636f6e74",
  3464 => x"726f6c00",
  3465 => x"20206170",
  3466 => x"62736c76",
  3467 => x"00000000",
  3468 => x"76656e64",
  3469 => x"20307800",
  3470 => x"64657620",
  3471 => x"30780000",
  3472 => x"76657220",
  3473 => x"00000000",
  3474 => x"69727120",
  3475 => x"00000000",
  3476 => x"61646472",
  3477 => x"20307800",
  3478 => x"6168626d",
  3479 => x"73740000",
  3480 => x"61686273",
  3481 => x"6c760000",
  3482 => x"00000ef5",
  3483 => x"00000fc6",
  3484 => x"00000fbb",
  3485 => x"00000ff2",
  3486 => x"00000fe7",
  3487 => x"00000fdc",
  3488 => x"00000fd1",
  3489 => x"00000f9a",
  3490 => x"00000f8f",
  3491 => x"00000f84",
  3492 => x"00000f79",
  3493 => x"00000fb0",
  3494 => x"00000fa5",
  3495 => x"00000f6e",
  3496 => x"00000ef5",
  3497 => x"00000ef5",
  3498 => x"00000ef5",
  3499 => x"00000ef5",
  3500 => x"00000ef5",
  3501 => x"00000f63",
  3502 => x"00000ef5",
  3503 => x"00000ef5",
  3504 => x"00000f58",
  3505 => x"00000ef5",
  3506 => x"00000f4d",
  3507 => x"00000ef5",
  3508 => x"00000ef5",
  3509 => x"00000ef5",
  3510 => x"00000ef5",
  3511 => x"00000ef5",
  3512 => x"00000ef5",
  3513 => x"00000ef5",
  3514 => x"00000ef5",
  3515 => x"00000f42",
  3516 => x"00000ef5",
  3517 => x"00000ef5",
  3518 => x"00000f37",
  3519 => x"00000ef5",
  3520 => x"00000ef5",
  3521 => x"00000ef5",
  3522 => x"00000ef5",
  3523 => x"00000ef5",
  3524 => x"00000ef5",
  3525 => x"00000ef5",
  3526 => x"00000ef5",
  3527 => x"00000ef5",
  3528 => x"00000ef5",
  3529 => x"00000f2c",
  3530 => x"00000ef5",
  3531 => x"00000ef5",
  3532 => x"00000ef5",
  3533 => x"00000ef5",
  3534 => x"00000f21",
  3535 => x"00000ef5",
  3536 => x"00000ef5",
  3537 => x"00000ef5",
  3538 => x"00000ef5",
  3539 => x"00000ef5",
  3540 => x"00000ef5",
  3541 => x"00000ef5",
  3542 => x"00000ef5",
  3543 => x"00000ef5",
  3544 => x"00000ef5",
  3545 => x"00000ef5",
  3546 => x"00000ef5",
  3547 => x"00000ef5",
  3548 => x"00000ef5",
  3549 => x"00000ef5",
  3550 => x"00000ef5",
  3551 => x"00000ef5",
  3552 => x"00000ef5",
  3553 => x"00000ef5",
  3554 => x"00000ef5",
  3555 => x"00000ef5",
  3556 => x"00000ef5",
  3557 => x"00000ef5",
  3558 => x"00000f16",
  3559 => x"00000ef5",
  3560 => x"00000ef5",
  3561 => x"00000ef5",
  3562 => x"00000ef5",
  3563 => x"00000ef5",
  3564 => x"00000ef5",
  3565 => x"00000ef5",
  3566 => x"00000ef5",
  3567 => x"00000ef5",
  3568 => x"00000ef5",
  3569 => x"00000ef5",
  3570 => x"00000ef5",
  3571 => x"00000ef5",
  3572 => x"00000ef5",
  3573 => x"00000ef5",
  3574 => x"00000ef5",
  3575 => x"00000ef5",
  3576 => x"00000ef5",
  3577 => x"00000ef5",
  3578 => x"00000ef5",
  3579 => x"00000ef5",
  3580 => x"00000ef5",
  3581 => x"00000ef5",
  3582 => x"00000ef5",
  3583 => x"00000ef5",
  3584 => x"00000ef5",
  3585 => x"00000ef5",
  3586 => x"00000f0b",
  3587 => x"02020606",
  3588 => x"06040304",
  3589 => x"02020102",
  3590 => x"636f6e74",
  3591 => x"726f6c20",
  3592 => x"2020203a",
  3593 => x"20000000",
  3594 => x"66726571",
  3595 => x"75656e63",
  3596 => x"7920203a",
  3597 => x"20000000",
  3598 => x"75706461",
  3599 => x"74652063",
  3600 => x"6c6b203a",
  3601 => x"20000000",
  3602 => x"72616d70",
  3603 => x"20726174",
  3604 => x"6520203a",
  3605 => x"20000000",
  3606 => x"49206d75",
  3607 => x"6c742072",
  3608 => x"6567203a",
  3609 => x"20000000",
  3610 => x"51206d75",
  3611 => x"6c742072",
  3612 => x"6567203a",
  3613 => x"20000000",
  3614 => x"554e4b4e",
  3615 => x"4f574e00",
  3616 => x"69646c65",
  3617 => x"00000000",
  3618 => x"636f6e66",
  3619 => x"69677572",
  3620 => x"65000000",
  3621 => x"64657465",
  3622 => x"63740000",
  3623 => x"61717569",
  3624 => x"72650000",
  3625 => x"616e616c",
  3626 => x"797a6500",
  3627 => x"64657369",
  3628 => x"72650000",
  3629 => x"72656164",
  3630 => x"6f757400",
  3631 => x"72656164",
  3632 => x"6c616700",
  3633 => x"66617374",
  3634 => x"20747269",
  3635 => x"67676572",
  3636 => x"203a2000",
  3637 => x"0a736c6f",
  3638 => x"77207472",
  3639 => x"69676765",
  3640 => x"72203a20",
  3641 => x"00000000",
  3642 => x"0a6f7665",
  3643 => x"72666c6f",
  3644 => x"77202020",
  3645 => x"20203a20",
  3646 => x"00000000",
  3647 => x"66617374",
  3648 => x"20747269",
  3649 => x"67676572",
  3650 => x"20636861",
  3651 => x"696e3a20",
  3652 => x"30780000",
  3653 => x"0a736c6f",
  3654 => x"77207472",
  3655 => x"69676765",
  3656 => x"72206368",
  3657 => x"61696e3a",
  3658 => x"20307800",
  3659 => x"0a636861",
  3660 => x"6e6e656c",
  3661 => x"206d6173",
  3662 => x"6b202861",
  3663 => x"6e64293a",
  3664 => x"20307800",
  3665 => x"0a666f72",
  3666 => x"6365206d",
  3667 => x"61736b20",
  3668 => x"286f7229",
  3669 => x"3a202020",
  3670 => x"20307800",
  3671 => x"0000172d",
  3672 => x"00001741",
  3673 => x"00001705",
  3674 => x"00001755",
  3675 => x"00001769",
  3676 => x"0000177d",
  3677 => x"00001791",
  3678 => x"000017a5",
  3679 => x"000017b9",
  3680 => x"00001719",
  3681 => x"30622020",
  3682 => x"20202020",
  3683 => x"20202020",
  3684 => x"20202020",
  3685 => x"20202020",
  3686 => x"20202020",
  3687 => x"20202020",
  3688 => x"20202020",
  3689 => x"20200000",
  3690 => x"20202020",
  3691 => x"20202020",
  3692 => x"00000000",
  3693 => x"79657300",
  3694 => x"6e6f0000",
  3695 => x"00202020",
  3696 => x"20202020",
  3697 => x"20202828",
  3698 => x"28282820",
  3699 => x"20202020",
  3700 => x"20202020",
  3701 => x"20202020",
  3702 => x"20202020",
  3703 => x"20881010",
  3704 => x"10101010",
  3705 => x"10101010",
  3706 => x"10101010",
  3707 => x"10040404",
  3708 => x"04040404",
  3709 => x"04040410",
  3710 => x"10101010",
  3711 => x"10104141",
  3712 => x"41414141",
  3713 => x"01010101",
  3714 => x"01010101",
  3715 => x"01010101",
  3716 => x"01010101",
  3717 => x"01010101",
  3718 => x"10101010",
  3719 => x"10104242",
  3720 => x"42424242",
  3721 => x"02020202",
  3722 => x"02020202",
  3723 => x"02020202",
  3724 => x"02020202",
  3725 => x"02020202",
  3726 => x"10101010",
  3727 => x"20000000",
  3728 => x"00000000",
  3729 => x"00000000",
  3730 => x"00000000",
  3731 => x"00000000",
  3732 => x"00000000",
  3733 => x"00000000",
  3734 => x"00000000",
  3735 => x"00000000",
  3736 => x"00000000",
  3737 => x"00000000",
  3738 => x"00000000",
  3739 => x"00000000",
  3740 => x"00000000",
  3741 => x"00000000",
  3742 => x"00000000",
  3743 => x"00000000",
  3744 => x"00000000",
  3745 => x"00000000",
  3746 => x"00000000",
  3747 => x"00000000",
  3748 => x"00000000",
  3749 => x"00000000",
  3750 => x"00000000",
  3751 => x"00000000",
  3752 => x"00000000",
  3753 => x"00000000",
  3754 => x"00000000",
  3755 => x"00000000",
  3756 => x"00000000",
  3757 => x"00000000",
  3758 => x"00000000",
  3759 => x"00000000",
  3760 => x"43000000",
  3761 => x"00000000",
  3762 => x"00000000",
  3763 => x"80000b00",
  3764 => x"10000000",
  3765 => x"80000d00",
  3766 => x"00ffffff",
  3767 => x"ff00ffff",
  3768 => x"ffff00ff",
  3769 => x"ffffff00",
  3770 => x"00000000",
  3771 => x"00000000",
  3772 => x"80000a00",
  3773 => x"80000400",
  3774 => x"80000200",
  3775 => x"80000100",
  3776 => x"80000004",
  3777 => x"80000000",
  3778 => x"00003b0c",
  3779 => x"00000000",
  3780 => x"00003d74",
  3781 => x"00003dd0",
  3782 => x"00003e2c",
  3783 => x"00000000",
  3784 => x"00000000",
  3785 => x"00000000",
  3786 => x"00000000",
  3787 => x"00000000",
  3788 => x"00000000",
  3789 => x"00000000",
  3790 => x"00000000",
  3791 => x"00000000",
  3792 => x"00003ac0",
  3793 => x"00000000",
  3794 => x"00000000",
  3795 => x"00000000",
  3796 => x"00000000",
  3797 => x"00000000",
  3798 => x"00000000",
  3799 => x"00000000",
  3800 => x"00000000",
  3801 => x"00000000",
  3802 => x"00000000",
  3803 => x"00000000",
  3804 => x"00000000",
  3805 => x"00000000",
  3806 => x"00000000",
  3807 => x"00000000",
  3808 => x"00000000",
  3809 => x"00000000",
  3810 => x"00000000",
  3811 => x"00000000",
  3812 => x"00000000",
  3813 => x"00000000",
  3814 => x"00000000",
  3815 => x"00000000",
  3816 => x"00000000",
  3817 => x"00000000",
  3818 => x"00000000",
  3819 => x"00000000",
  3820 => x"00000000",
  3821 => x"00000001",
  3822 => x"330eabcd",
  3823 => x"1234e66d",
  3824 => x"deec0005",
  3825 => x"000b0000",
  3826 => x"00000000",
  3827 => x"00000000",
  3828 => x"00000000",
  3829 => x"00000000",
  3830 => x"00000000",
  3831 => x"00000000",
  3832 => x"00000000",
  3833 => x"00000000",
  3834 => x"00000000",
  3835 => x"00000000",
  3836 => x"00000000",
  3837 => x"00000000",
  3838 => x"00000000",
  3839 => x"00000000",
  3840 => x"00000000",
  3841 => x"00000000",
  3842 => x"00000000",
  3843 => x"00000000",
  3844 => x"00000000",
  3845 => x"00000000",
  3846 => x"00000000",
  3847 => x"00000000",
  3848 => x"00000000",
  3849 => x"00000000",
  3850 => x"00000000",
  3851 => x"00000000",
  3852 => x"00000000",
  3853 => x"00000000",
  3854 => x"00000000",
  3855 => x"00000000",
  3856 => x"00000000",
  3857 => x"00000000",
  3858 => x"00000000",
  3859 => x"00000000",
  3860 => x"00000000",
  3861 => x"00000000",
  3862 => x"00000000",
  3863 => x"00000000",
  3864 => x"00000000",
  3865 => x"00000000",
  3866 => x"00000000",
  3867 => x"00000000",
  3868 => x"00000000",
  3869 => x"00000000",
  3870 => x"00000000",
  3871 => x"00000000",
  3872 => x"00000000",
  3873 => x"00000000",
  3874 => x"00000000",
  3875 => x"00000000",
  3876 => x"00000000",
  3877 => x"00000000",
  3878 => x"00000000",
  3879 => x"00000000",
  3880 => x"00000000",
  3881 => x"00000000",
  3882 => x"00000000",
  3883 => x"00000000",
  3884 => x"00000000",
  3885 => x"00000000",
  3886 => x"00000000",
  3887 => x"00000000",
  3888 => x"00000000",
  3889 => x"00000000",
  3890 => x"00000000",
  3891 => x"00000000",
  3892 => x"00000000",
  3893 => x"00000000",
  3894 => x"00000000",
  3895 => x"00000000",
  3896 => x"00000000",
  3897 => x"00000000",
  3898 => x"00000000",
  3899 => x"00000000",
  3900 => x"00000000",
  3901 => x"00000000",
  3902 => x"00000000",
  3903 => x"00000000",
  3904 => x"00000000",
  3905 => x"00000000",
  3906 => x"00000000",
  3907 => x"00000000",
  3908 => x"00000000",
  3909 => x"00000000",
  3910 => x"00000000",
  3911 => x"00000000",
  3912 => x"00000000",
  3913 => x"00000000",
  3914 => x"00000000",
  3915 => x"00000000",
  3916 => x"00000000",
  3917 => x"00000000",
  3918 => x"00000000",
  3919 => x"00000000",
  3920 => x"00000000",
  3921 => x"00000000",
  3922 => x"00000000",
  3923 => x"00000000",
  3924 => x"00000000",
  3925 => x"00000000",
  3926 => x"00000000",
  3927 => x"00000000",
  3928 => x"00000000",
  3929 => x"00000000",
  3930 => x"00000000",
  3931 => x"00000000",
  3932 => x"00000000",
  3933 => x"00000000",
  3934 => x"00000000",
  3935 => x"00000000",
  3936 => x"00000000",
  3937 => x"00000000",
  3938 => x"00000000",
  3939 => x"00000000",
  3940 => x"00000000",
  3941 => x"00000000",
  3942 => x"00000000",
  3943 => x"00000000",
  3944 => x"00000000",
  3945 => x"00000000",
  3946 => x"00000000",
  3947 => x"00000000",
  3948 => x"00000000",
  3949 => x"00000000",
  3950 => x"00000000",
  3951 => x"00000000",
  3952 => x"00000000",
  3953 => x"00000000",
  3954 => x"00000000",
  3955 => x"00000000",
  3956 => x"00000000",
  3957 => x"00000000",
  3958 => x"00000000",
  3959 => x"00000000",
  3960 => x"00000000",
  3961 => x"00000000",
  3962 => x"00000000",
  3963 => x"00000000",
  3964 => x"00000000",
  3965 => x"00000000",
  3966 => x"00000000",
  3967 => x"00000000",
  3968 => x"00000000",
  3969 => x"00000000",
  3970 => x"00000000",
  3971 => x"00000000",
  3972 => x"00000000",
  3973 => x"00000000",
  3974 => x"00000000",
  3975 => x"00000000",
  3976 => x"00000000",
  3977 => x"00000000",
  3978 => x"00000000",
  3979 => x"00000000",
  3980 => x"00000000",
  3981 => x"00000000",
  3982 => x"00000000",
  3983 => x"00000000",
  3984 => x"00000000",
  3985 => x"00000000",
  3986 => x"00000000",
  3987 => x"00000000",
  3988 => x"00000000",
  3989 => x"00000000",
  3990 => x"00000000",
  3991 => x"00000000",
  3992 => x"00000000",
  3993 => x"00000000",
  3994 => x"00000000",
  3995 => x"00000000",
  3996 => x"00000000",
  3997 => x"00000000",
  3998 => x"00000000",
  3999 => x"00000000",
  4000 => x"00000000",
  4001 => x"00000000",
  4002 => x"00000000",
  4003 => x"00000000",
  4004 => x"00000000",
  4005 => x"00000000",
  4006 => x"00000000",
  4007 => x"00000000",
  4008 => x"00000000",
  4009 => x"00000000",
  4010 => x"00000000",
  4011 => x"00000000",
  4012 => x"00000000",
  4013 => x"00000000",
  4014 => x"ffffffff",
  4015 => x"00000000",
  4016 => x"00020000",
  4017 => x"00000000",
  4018 => x"00000000",
  4019 => x"00003ec4",
  4020 => x"00003ec4",
  4021 => x"00003ecc",
  4022 => x"00003ecc",
  4023 => x"00003ed4",
  4024 => x"00003ed4",
  4025 => x"00003edc",
  4026 => x"00003edc",
  4027 => x"00003ee4",
  4028 => x"00003ee4",
  4029 => x"00003eec",
  4030 => x"00003eec",
  4031 => x"00003ef4",
  4032 => x"00003ef4",
  4033 => x"00003efc",
  4034 => x"00003efc",
  4035 => x"00003f04",
  4036 => x"00003f04",
  4037 => x"00003f0c",
  4038 => x"00003f0c",
  4039 => x"00003f14",
  4040 => x"00003f14",
  4041 => x"00003f1c",
  4042 => x"00003f1c",
  4043 => x"00003f24",
  4044 => x"00003f24",
  4045 => x"00003f2c",
  4046 => x"00003f2c",
  4047 => x"00003f34",
  4048 => x"00003f34",
  4049 => x"00003f3c",
  4050 => x"00003f3c",
  4051 => x"00003f44",
  4052 => x"00003f44",
  4053 => x"00003f4c",
  4054 => x"00003f4c",
  4055 => x"00003f54",
  4056 => x"00003f54",
  4057 => x"00003f5c",
  4058 => x"00003f5c",
  4059 => x"00003f64",
  4060 => x"00003f64",
  4061 => x"00003f6c",
  4062 => x"00003f6c",
  4063 => x"00003f74",
  4064 => x"00003f74",
  4065 => x"00003f7c",
  4066 => x"00003f7c",
  4067 => x"00003f84",
  4068 => x"00003f84",
  4069 => x"00003f8c",
  4070 => x"00003f8c",
  4071 => x"00003f94",
  4072 => x"00003f94",
  4073 => x"00003f9c",
  4074 => x"00003f9c",
  4075 => x"00003fa4",
  4076 => x"00003fa4",
  4077 => x"00003fac",
  4078 => x"00003fac",
  4079 => x"00003fb4",
  4080 => x"00003fb4",
  4081 => x"00003fbc",
  4082 => x"00003fbc",
  4083 => x"00003fc4",
  4084 => x"00003fc4",
  4085 => x"00003fcc",
  4086 => x"00003fcc",
  4087 => x"00003fd4",
  4088 => x"00003fd4",
  4089 => x"00003fdc",
  4090 => x"00003fdc",
  4091 => x"00003fe4",
  4092 => x"00003fe4",
  4093 => x"00003fec",
  4094 => x"00003fec",
  4095 => x"00003ff4",
  4096 => x"00003ff4",
  4097 => x"00003ffc",
  4098 => x"00003ffc",
  4099 => x"00004004",
  4100 => x"00004004",
  4101 => x"0000400c",
  4102 => x"0000400c",
  4103 => x"00004014",
  4104 => x"00004014",
  4105 => x"0000401c",
  4106 => x"0000401c",
  4107 => x"00004024",
  4108 => x"00004024",
  4109 => x"0000402c",
  4110 => x"0000402c",
  4111 => x"00004034",
  4112 => x"00004034",
  4113 => x"0000403c",
  4114 => x"0000403c",
  4115 => x"00004044",
  4116 => x"00004044",
  4117 => x"0000404c",
  4118 => x"0000404c",
  4119 => x"00004054",
  4120 => x"00004054",
  4121 => x"0000405c",
  4122 => x"0000405c",
  4123 => x"00004064",
  4124 => x"00004064",
  4125 => x"0000406c",
  4126 => x"0000406c",
  4127 => x"00004074",
  4128 => x"00004074",
  4129 => x"0000407c",
  4130 => x"0000407c",
  4131 => x"00004084",
  4132 => x"00004084",
  4133 => x"0000408c",
  4134 => x"0000408c",
  4135 => x"00004094",
  4136 => x"00004094",
  4137 => x"0000409c",
  4138 => x"0000409c",
  4139 => x"000040a4",
  4140 => x"000040a4",
  4141 => x"000040ac",
  4142 => x"000040ac",
  4143 => x"000040b4",
  4144 => x"000040b4",
  4145 => x"000040bc",
  4146 => x"000040bc",
  4147 => x"000040c4",
  4148 => x"000040c4",
  4149 => x"000040cc",
  4150 => x"000040cc",
  4151 => x"000040d4",
  4152 => x"000040d4",
  4153 => x"000040dc",
  4154 => x"000040dc",
  4155 => x"000040e4",
  4156 => x"000040e4",
  4157 => x"000040ec",
  4158 => x"000040ec",
  4159 => x"000040f4",
  4160 => x"000040f4",
  4161 => x"000040fc",
  4162 => x"000040fc",
  4163 => x"00004104",
  4164 => x"00004104",
  4165 => x"0000410c",
  4166 => x"0000410c",
  4167 => x"00004114",
  4168 => x"00004114",
  4169 => x"0000411c",
  4170 => x"0000411c",
  4171 => x"00004124",
  4172 => x"00004124",
  4173 => x"0000412c",
  4174 => x"0000412c",
  4175 => x"00004134",
  4176 => x"00004134",
  4177 => x"0000413c",
  4178 => x"0000413c",
  4179 => x"00004144",
  4180 => x"00004144",
  4181 => x"0000414c",
  4182 => x"0000414c",
  4183 => x"00004154",
  4184 => x"00004154",
  4185 => x"0000415c",
  4186 => x"0000415c",
  4187 => x"00004164",
  4188 => x"00004164",
  4189 => x"0000416c",
  4190 => x"0000416c",
  4191 => x"00004174",
  4192 => x"00004174",
  4193 => x"0000417c",
  4194 => x"0000417c",
  4195 => x"00004184",
  4196 => x"00004184",
  4197 => x"0000418c",
  4198 => x"0000418c",
  4199 => x"00004194",
  4200 => x"00004194",
  4201 => x"0000419c",
  4202 => x"0000419c",
  4203 => x"000041a4",
  4204 => x"000041a4",
  4205 => x"000041ac",
  4206 => x"000041ac",
  4207 => x"000041b4",
  4208 => x"000041b4",
  4209 => x"000041bc",
  4210 => x"000041bc",
  4211 => x"000041c4",
  4212 => x"000041c4",
  4213 => x"000041cc",
  4214 => x"000041cc",
  4215 => x"000041d4",
  4216 => x"000041d4",
  4217 => x"000041dc",
  4218 => x"000041dc",
  4219 => x"000041e4",
  4220 => x"000041e4",
  4221 => x"000041ec",
  4222 => x"000041ec",
  4223 => x"000041f4",
  4224 => x"000041f4",
  4225 => x"000041fc",
  4226 => x"000041fc",
  4227 => x"00004204",
  4228 => x"00004204",
  4229 => x"0000420c",
  4230 => x"0000420c",
  4231 => x"00004214",
  4232 => x"00004214",
  4233 => x"0000421c",
  4234 => x"0000421c",
  4235 => x"00004224",
  4236 => x"00004224",
  4237 => x"0000422c",
  4238 => x"0000422c",
  4239 => x"00004234",
  4240 => x"00004234",
  4241 => x"0000423c",
  4242 => x"0000423c",
  4243 => x"00004244",
  4244 => x"00004244",
  4245 => x"0000424c",
  4246 => x"0000424c",
  4247 => x"00004254",
  4248 => x"00004254",
  4249 => x"0000425c",
  4250 => x"0000425c",
  4251 => x"00004264",
  4252 => x"00004264",
  4253 => x"0000426c",
  4254 => x"0000426c",
  4255 => x"00004274",
  4256 => x"00004274",
  4257 => x"0000427c",
  4258 => x"0000427c",
  4259 => x"00004284",
  4260 => x"00004284",
  4261 => x"0000428c",
  4262 => x"0000428c",
  4263 => x"00004294",
  4264 => x"00004294",
  4265 => x"0000429c",
  4266 => x"0000429c",
  4267 => x"000042a4",
  4268 => x"000042a4",
  4269 => x"000042ac",
  4270 => x"000042ac",
  4271 => x"000042b4",
  4272 => x"000042b4",
  4273 => x"000042bc",
  4274 => x"000042bc",
	--others => x"00dead00" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
