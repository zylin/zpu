-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b80e1",
     1 => x"d7040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b80e4",
     9 => x"be040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b80e3",
    73 => x"f0040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b80e3d3",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b81b1",
   162 => x"f8738306",
   163 => x"10100508",
   164 => x"060b0b80",
   165 => x"e3d60400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b80e4",
   169 => x"a5040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b80e4",
   177 => x"8c040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"81b2880c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053370",
   258 => x"525280e1",
   259 => x"bb3f7151",
   260 => x"80e2a93f",
   261 => x"71b00c83",
   262 => x"3d0d04fd",
   263 => x"3d0d8a51",
   264 => x"80dcc13f",
   265 => x"aaad3f97",
   266 => x"8a538193",
   267 => x"e4528193",
   268 => x"f851aab2",
   269 => x"3fa49253",
   270 => x"8193fc52",
   271 => x"8194a051",
   272 => x"aaa43fa7",
   273 => x"ab538194",
   274 => x"a8528194",
   275 => x"b851aa96",
   276 => x"3fa09d53",
   277 => x"8194c052",
   278 => x"8195b851",
   279 => x"aa883fa2",
   280 => x"87538194",
   281 => x"dc528194",
   282 => x"fc51a9fa",
   283 => x"3fa2ed53",
   284 => x"81958452",
   285 => x"8195a451",
   286 => x"a9ec3f9f",
   287 => x"e9538195",
   288 => x"ac528195",
   289 => x"c051a9de",
   290 => x"3fa5b153",
   291 => x"8195c852",
   292 => x"8195e451",
   293 => x"a9d03fa7",
   294 => x"c2538195",
   295 => x"ec528196",
   296 => x"9051a9c2",
   297 => x"3fa88353",
   298 => x"81969852",
   299 => x"8196c051",
   300 => x"a9b43fa9",
   301 => x"ab538196",
   302 => x"c8528196",
   303 => x"e851a9a6",
   304 => x"3fa79253",
   305 => x"8196ec52",
   306 => x"81978851",
   307 => x"a9983faa",
   308 => x"86538197",
   309 => x"90528197",
   310 => x"a051a98a",
   311 => x"3facd253",
   312 => x"8197a452",
   313 => x"8197c051",
   314 => x"a8fc3fa6",
   315 => x"d8538197",
   316 => x"c8528197",
   317 => x"e051a8ee",
   318 => x"3facda53",
   319 => x"8197e852",
   320 => x"8197fc51",
   321 => x"a8e03f8d",
   322 => x"f9538198",
   323 => x"84528198",
   324 => x"9851a8d2",
   325 => x"3f918353",
   326 => x"81989c52",
   327 => x"8198c451",
   328 => x"a8c43fa6",
   329 => x"f4538198",
   330 => x"cc528198",
   331 => x"ec51a8b6",
   332 => x"3f96a753",
   333 => x"8198f452",
   334 => x"81998851",
   335 => x"a8a83f8b",
   336 => x"fd538199",
   337 => x"90528199",
   338 => x"9c51a89a",
   339 => x"3f8da253",
   340 => x"8199a052",
   341 => x"8199c851",
   342 => x"a88c3f8b",
   343 => x"fd538199",
   344 => x"d05281a0",
   345 => x"f451a7fe",
   346 => x"3f8de853",
   347 => x"8199e052",
   348 => x"8199f051",
   349 => x"a7f03f8b",
   350 => x"f253819a",
   351 => x"84528193",
   352 => x"d451a7e2",
   353 => x"3fb9bd53",
   354 => x"819a8452",
   355 => x"8193dc51",
   356 => x"a7d43fae",
   357 => x"a83fa89a",
   358 => x"3f810b81",
   359 => x"d5983481",
   360 => x"c1f83370",
   361 => x"81ff0651",
   362 => x"5473b238",
   363 => x"80ddc13f",
   364 => x"b0089038",
   365 => x"a88a3f81",
   366 => x"d5983354",
   367 => x"73e13885",
   368 => x"3d0d0480",
   369 => x"ddbd3fb0",
   370 => x"0881ff06",
   371 => x"51a8df3f",
   372 => x"a7ee3f81",
   373 => x"d5983354",
   374 => x"73c538e3",
   375 => x"39800b81",
   376 => x"c1f834ae",
   377 => x"f83f80dd",
   378 => x"873fb008",
   379 => x"802ec538",
   380 => x"d239800b",
   381 => x"81d59834",
   382 => x"800bb00c",
   383 => x"04fb3d0d",
   384 => x"8151ac86",
   385 => x"3fb00853",
   386 => x"8251abfe",
   387 => x"3fb00856",
   388 => x"b0088338",
   389 => x"905672fc",
   390 => x"06547581",
   391 => x"2e80fb38",
   392 => x"80557476",
   393 => x"27ad3874",
   394 => x"83065372",
   395 => x"802eb238",
   396 => x"81a5f051",
   397 => x"80d8c73f",
   398 => x"73708405",
   399 => x"550852a0",
   400 => x"5180d8dd",
   401 => x"3fa05180",
   402 => x"d89a3f81",
   403 => x"15557575",
   404 => x"26d5388a",
   405 => x"5180d88c",
   406 => x"3f800bb0",
   407 => x"0c873d0d",
   408 => x"048199f8",
   409 => x"5180d896",
   410 => x"3f7352a0",
   411 => x"5180d8b1",
   412 => x"3f81a0e0",
   413 => x"5180d886",
   414 => x"3f81a5f0",
   415 => x"5180d7fe",
   416 => x"3f737084",
   417 => x"05550852",
   418 => x"a05180d8",
   419 => x"943fa051",
   420 => x"80d7d13f",
   421 => x"811555ff",
   422 => x"b5397308",
   423 => x"b00c873d",
   424 => x"0d04fc3d",
   425 => x"0d8151aa",
   426 => x"e13fb008",
   427 => x"528251a9",
   428 => x"a73fb008",
   429 => x"81ff0672",
   430 => x"56538354",
   431 => x"72802ea1",
   432 => x"387351aa",
   433 => x"c53f8114",
   434 => x"7081ff06",
   435 => x"ff157081",
   436 => x"ff06b008",
   437 => x"79708405",
   438 => x"5b0c5652",
   439 => x"555272e1",
   440 => x"3872b00c",
   441 => x"863d0d04",
   442 => x"803d0d8c",
   443 => x"5180d6f4",
   444 => x"3f800bb0",
   445 => x"0c823d0d",
   446 => x"04fb3d0d",
   447 => x"800b8199",
   448 => x"fc525680",
   449 => x"d6f83f75",
   450 => x"55741081",
   451 => x"fe065381",
   452 => x"d05281b2",
   453 => x"900851bd",
   454 => x"983fb008",
   455 => x"982b5480",
   456 => x"7424a238",
   457 => x"819a8851",
   458 => x"80d6d33f",
   459 => x"74528851",
   460 => x"80d6ee3f",
   461 => x"819a9451",
   462 => x"80d6c33f",
   463 => x"81167083",
   464 => x"ffff0657",
   465 => x"54811570",
   466 => x"81ff0670",
   467 => x"982b5256",
   468 => x"54738025",
   469 => x"ffb33875",
   470 => x"b00c873d",
   471 => x"0d04f33d",
   472 => x"0d7f0284",
   473 => x"0580c305",
   474 => x"33028805",
   475 => x"80c60522",
   476 => x"819aa454",
   477 => x"5b555880",
   478 => x"d6843f78",
   479 => x"5180d7c8",
   480 => x"3f819ab0",
   481 => x"5180d5f6",
   482 => x"3f735288",
   483 => x"5180d691",
   484 => x"3f819acc",
   485 => x"5180d5e6",
   486 => x"3f805776",
   487 => x"7927819c",
   488 => x"3873108e",
   489 => x"3d5d5a79",
   490 => x"81ff0653",
   491 => x"81905277",
   492 => x"51bbfe3f",
   493 => x"76882a53",
   494 => x"90527751",
   495 => x"bbf33f76",
   496 => x"81ff0653",
   497 => x"90527751",
   498 => x"bbe73f81",
   499 => x"1a7081ff",
   500 => x"06545581",
   501 => x"90527751",
   502 => x"bbd73f80",
   503 => x"5380e052",
   504 => x"7751bbcd",
   505 => x"3fb00898",
   506 => x"2b548074",
   507 => x"248a3888",
   508 => x"18087081",
   509 => x"ff065c56",
   510 => x"7a81ff06",
   511 => x"81a5f052",
   512 => x"5680d4fa",
   513 => x"3f755288",
   514 => x"5180d595",
   515 => x"3f819dec",
   516 => x"5180d4ea",
   517 => x"3fe01654",
   518 => x"80df7427",
   519 => x"b6387687",
   520 => x"06701d57",
   521 => x"55a07634",
   522 => x"74872eb9",
   523 => x"38811770",
   524 => x"83ffff06",
   525 => x"58557877",
   526 => x"26feec38",
   527 => x"80e00b8c",
   528 => x"190c8c18",
   529 => x"0870812a",
   530 => x"8106585a",
   531 => x"76f4388f",
   532 => x"3d0d0476",
   533 => x"8706701d",
   534 => x"55557574",
   535 => x"3474872e",
   536 => x"098106c9",
   537 => x"387b5180",
   538 => x"d4943f8a",
   539 => x"5180d3f4",
   540 => x"3f811770",
   541 => x"83ffff06",
   542 => x"58557877",
   543 => x"26fea838",
   544 => x"ffba39fb",
   545 => x"3d0d8151",
   546 => x"a5ce3fb0",
   547 => x"0881ff06",
   548 => x"548251a6",
   549 => x"f53fb008",
   550 => x"81ff0656",
   551 => x"8351a5b8",
   552 => x"3fb00883",
   553 => x"ffff0655",
   554 => x"739c3881",
   555 => x"b2900854",
   556 => x"74843881",
   557 => x"80557453",
   558 => x"75527351",
   559 => x"fda03f74",
   560 => x"b00c873d",
   561 => x"0d0481b2",
   562 => x"940854e4",
   563 => x"39f83d0d",
   564 => x"02aa0522",
   565 => x"81b1ec33",
   566 => x"81f70658",
   567 => x"587681b1",
   568 => x"ec3481b2",
   569 => x"90085580",
   570 => x"c0538190",
   571 => x"527451b9",
   572 => x"c03f7451",
   573 => x"b9ed3fb0",
   574 => x"0881ff06",
   575 => x"5473802e",
   576 => x"83fc3876",
   577 => x"5380d052",
   578 => x"7451b9a5",
   579 => x"3f80598f",
   580 => x"5781b1ec",
   581 => x"3381fe06",
   582 => x"547381b1",
   583 => x"ec3481b2",
   584 => x"90087457",
   585 => x"5580c053",
   586 => x"81905274",
   587 => x"51b9823f",
   588 => x"7451b9af",
   589 => x"3fb00881",
   590 => x"ff065473",
   591 => x"802e83b3",
   592 => x"38755380",
   593 => x"d0527451",
   594 => x"b8e73f77",
   595 => x"772c8106",
   596 => x"5574802e",
   597 => x"83923881",
   598 => x"b1ec3382",
   599 => x"07547381",
   600 => x"b1ec3481",
   601 => x"b2900874",
   602 => x"575580c0",
   603 => x"53819052",
   604 => x"7451b8bd",
   605 => x"3f7451b8",
   606 => x"ea3fb008",
   607 => x"81ff0654",
   608 => x"73802e82",
   609 => x"d8387553",
   610 => x"80d05274",
   611 => x"51b8a23f",
   612 => x"81b29008",
   613 => x"5580c153",
   614 => x"81905274",
   615 => x"51b8923f",
   616 => x"7451b8bf",
   617 => x"3fb00881",
   618 => x"ff065675",
   619 => x"802e8281",
   620 => x"38805380",
   621 => x"e0527451",
   622 => x"b7f73f74",
   623 => x"51b8a43f",
   624 => x"b00881ff",
   625 => x"06547380",
   626 => x"2e81e638",
   627 => x"88150870",
   628 => x"902b7090",
   629 => x"2c565656",
   630 => x"73822a81",
   631 => x"06547380",
   632 => x"2e8d3881",
   633 => x"772b7907",
   634 => x"7083ffff",
   635 => x"065a5681",
   636 => x"b1ec3381",
   637 => x"07547381",
   638 => x"b1ec3481",
   639 => x"b2900874",
   640 => x"575580c0",
   641 => x"53819052",
   642 => x"7451b7a5",
   643 => x"3f7451b7",
   644 => x"d23fb008",
   645 => x"81ff0654",
   646 => x"73802e81",
   647 => x"a1387553",
   648 => x"80d05274",
   649 => x"51b78a3f",
   650 => x"7681800a",
   651 => x"2981ff0a",
   652 => x"0570982c",
   653 => x"58567680",
   654 => x"25fdd638",
   655 => x"81b1ec33",
   656 => x"82075776",
   657 => x"81b1ec34",
   658 => x"81b29008",
   659 => x"5580c053",
   660 => x"81905274",
   661 => x"51b6da3f",
   662 => x"7451b787",
   663 => x"3fb00881",
   664 => x"ff065877",
   665 => x"802e81b4",
   666 => x"38765380",
   667 => x"d0527451",
   668 => x"b6bf3f81",
   669 => x"b1ec3388",
   670 => x"07577681",
   671 => x"b1ec3481",
   672 => x"b2900855",
   673 => x"80c05381",
   674 => x"90527451",
   675 => x"b6a33f74",
   676 => x"51b6d03f",
   677 => x"b00881ff",
   678 => x"06587780",
   679 => x"2e80ee38",
   680 => x"765380d0",
   681 => x"527451b6",
   682 => x"883f78b0",
   683 => x"0c8a3d0d",
   684 => x"04819ad0",
   685 => x"5180cfc6",
   686 => x"3fff54fe",
   687 => x"9b39819a",
   688 => x"d05180cf",
   689 => x"b93f7681",
   690 => x"800a2981",
   691 => x"ff0a0570",
   692 => x"982c5856",
   693 => x"768025fc",
   694 => x"b838fee0",
   695 => x"39819ad0",
   696 => x"5180cf9a",
   697 => x"3ffda939",
   698 => x"81b1ec33",
   699 => x"81fd0654",
   700 => x"fcec3981",
   701 => x"9ad05180",
   702 => x"cf843ffc",
   703 => x"ce39819a",
   704 => x"d05180ce",
   705 => x"f93f8059",
   706 => x"8f57fc85",
   707 => x"39819ad0",
   708 => x"5180ceea",
   709 => x"3f78b00c",
   710 => x"8a3d0d04",
   711 => x"819ad051",
   712 => x"80cedb3f",
   713 => x"fecd39ff",
   714 => x"3d0d8151",
   715 => x"a0aa3fb0",
   716 => x"0881ff06",
   717 => x"52818051",
   718 => x"fb933f82",
   719 => x"8051fb8d",
   720 => x"3f848351",
   721 => x"fb873f86",
   722 => x"f151fb81",
   723 => x"3f71832b",
   724 => x"88830751",
   725 => x"faf73f80",
   726 => x"0bb00c83",
   727 => x"3d0d04fe",
   728 => x"3d0d0293",
   729 => x"05330284",
   730 => x"05970533",
   731 => x"54527173",
   732 => x"279438a0",
   733 => x"5180cdec",
   734 => x"3f811270",
   735 => x"81ff0651",
   736 => x"52727226",
   737 => x"ee38843d",
   738 => x"0d04fd3d",
   739 => x"0d819b88",
   740 => x"5180cdea",
   741 => x"3f819ba8",
   742 => x"5180cde2",
   743 => x"3f819bf0",
   744 => x"5180cdda",
   745 => x"3f819cb8",
   746 => x"5180cdd2",
   747 => x"3f81b1e4",
   748 => x"08700852",
   749 => x"5380cf90",
   750 => x"3fb00881",
   751 => x"ff065372",
   752 => x"8c279438",
   753 => x"a05180cd",
   754 => x"9b3f8113",
   755 => x"7081ff06",
   756 => x"54548c73",
   757 => x"26ee3881",
   758 => x"b1e40884",
   759 => x"11085253",
   760 => x"80cee53f",
   761 => x"b00881ff",
   762 => x"0653728c",
   763 => x"279438a0",
   764 => x"5180ccf0",
   765 => x"3f811370",
   766 => x"81ff0654",
   767 => x"548c7326",
   768 => x"ee3881b1",
   769 => x"e4088811",
   770 => x"08525380",
   771 => x"ceba3fb0",
   772 => x"0881ff06",
   773 => x"53728c27",
   774 => x"9438a051",
   775 => x"80ccc53f",
   776 => x"81137081",
   777 => x"ff065454",
   778 => x"8c7326ee",
   779 => x"3881b1e4",
   780 => x"088c1108",
   781 => x"525380ce",
   782 => x"8f3fb008",
   783 => x"81ff0653",
   784 => x"728c2794",
   785 => x"38a05180",
   786 => x"cc9a3f81",
   787 => x"137081ff",
   788 => x"0654548c",
   789 => x"7326ee38",
   790 => x"819cd451",
   791 => x"80cc9f3f",
   792 => x"81b1e408",
   793 => x"90110852",
   794 => x"5380cddc",
   795 => x"3fb00881",
   796 => x"ff065372",
   797 => x"8c279438",
   798 => x"a05180cb",
   799 => x"e73f8113",
   800 => x"7081ff06",
   801 => x"54548c73",
   802 => x"26ee3881",
   803 => x"b1e40894",
   804 => x"11085253",
   805 => x"80cdb13f",
   806 => x"b00881ff",
   807 => x"0653728c",
   808 => x"279438a0",
   809 => x"5180cbbc",
   810 => x"3f811370",
   811 => x"81ff0654",
   812 => x"548c7326",
   813 => x"ee3881b1",
   814 => x"e4089811",
   815 => x"08525380",
   816 => x"cd863fb0",
   817 => x"0881ff06",
   818 => x"53728c27",
   819 => x"9438a051",
   820 => x"80cb913f",
   821 => x"81137081",
   822 => x"ff065454",
   823 => x"8c7326ee",
   824 => x"3881b1e4",
   825 => x"089c1108",
   826 => x"525380cc",
   827 => x"db3fb008",
   828 => x"81ff0653",
   829 => x"728c2794",
   830 => x"38a05180",
   831 => x"cae63f81",
   832 => x"137081ff",
   833 => x"0654548c",
   834 => x"7326ee38",
   835 => x"819cf051",
   836 => x"80caeb3f",
   837 => x"81b1e408",
   838 => x"54810bb0",
   839 => x"150cb014",
   840 => x"08537280",
   841 => x"25f838a0",
   842 => x"14085180",
   843 => x"cc9a3fb0",
   844 => x"0881ff06",
   845 => x"53728c27",
   846 => x"9438a051",
   847 => x"80caa53f",
   848 => x"81137081",
   849 => x"ff065454",
   850 => x"8c7326ee",
   851 => x"3881b1e4",
   852 => x"08a41108",
   853 => x"525380cb",
   854 => x"ef3fb008",
   855 => x"81ff0653",
   856 => x"728c2794",
   857 => x"38a05180",
   858 => x"c9fa3f81",
   859 => x"137081ff",
   860 => x"0654548c",
   861 => x"7326ee38",
   862 => x"81b1e408",
   863 => x"a8110852",
   864 => x"5380cbc4",
   865 => x"3fb00881",
   866 => x"ff065372",
   867 => x"8c279438",
   868 => x"a05180c9",
   869 => x"cf3f8113",
   870 => x"7081ff06",
   871 => x"54548c73",
   872 => x"26ee3881",
   873 => x"b1e408ac",
   874 => x"11085253",
   875 => x"80cb993f",
   876 => x"b00881ff",
   877 => x"0653728c",
   878 => x"279438a0",
   879 => x"5180c9a4",
   880 => x"3f811370",
   881 => x"81ff0654",
   882 => x"548c7326",
   883 => x"ee38819d",
   884 => x"8c5180c9",
   885 => x"a93f81b1",
   886 => x"e408b011",
   887 => x"08fe0a06",
   888 => x"525480ca",
   889 => x"e33f81b1",
   890 => x"e4085480",
   891 => x"0bb0150c",
   892 => x"819da051",
   893 => x"80c9873f",
   894 => x"819db851",
   895 => x"80c8ff3f",
   896 => x"81b1e408",
   897 => x"80c01108",
   898 => x"525380ca",
   899 => x"bb3fb008",
   900 => x"81ff0653",
   901 => x"72982794",
   902 => x"38a05180",
   903 => x"c8c63f81",
   904 => x"137081ff",
   905 => x"06515398",
   906 => x"7326ee38",
   907 => x"81b1e408",
   908 => x"80c81108",
   909 => x"525480ca",
   910 => x"8f3fb008",
   911 => x"81ff0653",
   912 => x"72982794",
   913 => x"38a05180",
   914 => x"c89a3f81",
   915 => x"137081ff",
   916 => x"06515398",
   917 => x"7326ee38",
   918 => x"819dd451",
   919 => x"80c89f3f",
   920 => x"81b1e408",
   921 => x"80c41108",
   922 => x"525480c9",
   923 => x"db3fb008",
   924 => x"81ff0653",
   925 => x"72982794",
   926 => x"38a05180",
   927 => x"c7e63f81",
   928 => x"137081ff",
   929 => x"06515398",
   930 => x"7326ee38",
   931 => x"81b1e408",
   932 => x"80cc1108",
   933 => x"525480c9",
   934 => x"af3fb008",
   935 => x"81ff0653",
   936 => x"72982794",
   937 => x"38a05180",
   938 => x"c7ba3f81",
   939 => x"137081ff",
   940 => x"06515398",
   941 => x"7326ee38",
   942 => x"8a5180c7",
   943 => x"a73f81b1",
   944 => x"e408b411",
   945 => x"087081ff",
   946 => x"06819df0",
   947 => x"54525553",
   948 => x"80c7ab3f",
   949 => x"725180c8",
   950 => x"ef3fa051",
   951 => x"80c7853f",
   952 => x"72862694",
   953 => x"38721010",
   954 => x"81a2b005",
   955 => x"54730804",
   956 => x"819e8451",
   957 => x"80c7873f",
   958 => x"81b1e408",
   959 => x"b8110870",
   960 => x"81ff0681",
   961 => x"9e905452",
   962 => x"545480c6",
   963 => x"f13f7352",
   964 => x"885180c7",
   965 => x"8c3f7381",
   966 => x"06537280",
   967 => x"f2387381",
   968 => x"2a708106",
   969 => x"51537280",
   970 => x"ce387382",
   971 => x"2a708106",
   972 => x"515372ae",
   973 => x"3873832a",
   974 => x"81065473",
   975 => x"8f388a51",
   976 => x"80c6a13f",
   977 => x"800bb00c",
   978 => x"853d0d04",
   979 => x"819ea451",
   980 => x"80c6ab3f",
   981 => x"8a5180c6",
   982 => x"8b3f800b",
   983 => x"b00c853d",
   984 => x"0d04819e",
   985 => x"b85180c6",
   986 => x"953f7383",
   987 => x"2a810654",
   988 => x"73802eca",
   989 => x"38d63981",
   990 => x"9ed85180",
   991 => x"c6803f73",
   992 => x"822a7081",
   993 => x"06515372",
   994 => x"802effa9",
   995 => x"38d43981",
   996 => x"9ef05180",
   997 => x"c5e83f73",
   998 => x"812a7081",
   999 => x"06515372",
  1000 => x"802eff86",
  1001 => x"38d13981",
  1002 => x"9f845180",
  1003 => x"c5d03ffe",
  1004 => x"c739819f",
  1005 => x"905180c5",
  1006 => x"c53ffebc",
  1007 => x"39819f9c",
  1008 => x"5180c5ba",
  1009 => x"3ffeb139",
  1010 => x"819fa051",
  1011 => x"80c5af3f",
  1012 => x"fea63981",
  1013 => x"9fac5180",
  1014 => x"c5a43ffe",
  1015 => x"9b39819f",
  1016 => x"b85180c5",
  1017 => x"993ffe90",
  1018 => x"39fe3d0d",
  1019 => x"880a5384",
  1020 => x"0a0b81b1",
  1021 => x"e0088c11",
  1022 => x"08515252",
  1023 => x"80712795",
  1024 => x"38807370",
  1025 => x"8405550c",
  1026 => x"80727084",
  1027 => x"05540cff",
  1028 => x"115170ed",
  1029 => x"38800bb0",
  1030 => x"0c843d0d",
  1031 => x"04fa3d0d",
  1032 => x"880a5784",
  1033 => x"0a568151",
  1034 => x"96ae3fb0",
  1035 => x"0883ffff",
  1036 => x"06547383",
  1037 => x"38905480",
  1038 => x"55747427",
  1039 => x"81c23875",
  1040 => x"0870902c",
  1041 => x"525380c5",
  1042 => x"ff3fb008",
  1043 => x"81ff0652",
  1044 => x"718a2794",
  1045 => x"38a05180",
  1046 => x"c48a3f81",
  1047 => x"127081ff",
  1048 => x"0651528a",
  1049 => x"7226ee38",
  1050 => x"72902b70",
  1051 => x"902c5252",
  1052 => x"80c5d53f",
  1053 => x"b00881ff",
  1054 => x"0652718a",
  1055 => x"279438a0",
  1056 => x"5180c3e0",
  1057 => x"3f811270",
  1058 => x"81ff0653",
  1059 => x"538a7226",
  1060 => x"ee387608",
  1061 => x"70902c52",
  1062 => x"5380c5ac",
  1063 => x"3fb00881",
  1064 => x"ff065271",
  1065 => x"8a279438",
  1066 => x"a05180c3",
  1067 => x"b73f8112",
  1068 => x"7081ff06",
  1069 => x"51528a72",
  1070 => x"26ee3872",
  1071 => x"902b7090",
  1072 => x"2c525280",
  1073 => x"c5823fb0",
  1074 => x"0881ff06",
  1075 => x"52718a27",
  1076 => x"9438a051",
  1077 => x"80c38d3f",
  1078 => x"81127081",
  1079 => x"ff065353",
  1080 => x"8a7226ee",
  1081 => x"388a5180",
  1082 => x"c2fa3f84",
  1083 => x"17841781",
  1084 => x"177083ff",
  1085 => x"ff065854",
  1086 => x"57577375",
  1087 => x"26fec038",
  1088 => x"73b00c88",
  1089 => x"3d0d04fd",
  1090 => x"3d0d81b1",
  1091 => x"e0088c11",
  1092 => x"0870822b",
  1093 => x"83fffc06",
  1094 => x"819fc454",
  1095 => x"51545480",
  1096 => x"c2dc3f72",
  1097 => x"52880a51",
  1098 => x"9af63fb0",
  1099 => x"0854b008",
  1100 => x"fe2eab38",
  1101 => x"b008ff2e",
  1102 => x"96387251",
  1103 => x"80c4893f",
  1104 => x"819fd851",
  1105 => x"80c2b73f",
  1106 => x"73b00c85",
  1107 => x"3d0d0481",
  1108 => x"9fec5180",
  1109 => x"c2a83f73",
  1110 => x"b00c853d",
  1111 => x"0d04819f",
  1112 => x"f45180c2",
  1113 => x"993f73b0",
  1114 => x"0c853d0d",
  1115 => x"04fc3d0d",
  1116 => x"81b1e008",
  1117 => x"8c110870",
  1118 => x"822b83ff",
  1119 => x"fc0681a0",
  1120 => x"80545155",
  1121 => x"5580c1f6",
  1122 => x"3f81b2a4",
  1123 => x"08881108",
  1124 => x"7080c007",
  1125 => x"88130c54",
  1126 => x"55735288",
  1127 => x"0a519d82",
  1128 => x"3fb00881",
  1129 => x"b2a40888",
  1130 => x"110870ff",
  1131 => x"bf068813",
  1132 => x"0c555555",
  1133 => x"b008fe2e",
  1134 => x"80c938b0",
  1135 => x"08fe249c",
  1136 => x"38b008fd",
  1137 => x"2eae3874",
  1138 => x"5180c2fc",
  1139 => x"3f81a094",
  1140 => x"5180c1aa",
  1141 => x"3f74b00c",
  1142 => x"863d0d04",
  1143 => x"b008ff2e",
  1144 => x"098106e3",
  1145 => x"38819fec",
  1146 => x"5180c192",
  1147 => x"3f74b00c",
  1148 => x"863d0d04",
  1149 => x"81a0a851",
  1150 => x"80c1833f",
  1151 => x"74b00c86",
  1152 => x"3d0d0481",
  1153 => x"a0b85180",
  1154 => x"c0f43f74",
  1155 => x"b00c863d",
  1156 => x"0d04fd3d",
  1157 => x"0d815192",
  1158 => x"bf3fb008",
  1159 => x"81ff0654",
  1160 => x"73802ea4",
  1161 => x"38738426",
  1162 => x"903881b1",
  1163 => x"e0087471",
  1164 => x"0c5373b0",
  1165 => x"0c853d0d",
  1166 => x"0481b1e0",
  1167 => x"08538073",
  1168 => x"0c73b00c",
  1169 => x"853d0d04",
  1170 => x"81a0c451",
  1171 => x"80c0af3f",
  1172 => x"81a0d451",
  1173 => x"80c0a73f",
  1174 => x"81b1e008",
  1175 => x"70085253",
  1176 => x"80c1e53f",
  1177 => x"81a0e451",
  1178 => x"80c0933f",
  1179 => x"81b1e008",
  1180 => x"84110853",
  1181 => x"53a05180",
  1182 => x"c0a73f81",
  1183 => x"a0f851bf",
  1184 => x"fd3f81b1",
  1185 => x"e0088811",
  1186 => x"085353a0",
  1187 => x"5180c091",
  1188 => x"3f81a18c",
  1189 => x"51bfe73f",
  1190 => x"81b1e008",
  1191 => x"8c110852",
  1192 => x"5380c1a4",
  1193 => x"3f8a51bf",
  1194 => x"bb3f73b0",
  1195 => x"0c853d0d",
  1196 => x"04f63d0d",
  1197 => x"880a5681",
  1198 => x"51919d3f",
  1199 => x"b0088b3d",
  1200 => x"23825191",
  1201 => x"933fb008",
  1202 => x"028405a6",
  1203 => x"05238351",
  1204 => x"91863fb0",
  1205 => x"088c3d23",
  1206 => x"845190fc",
  1207 => x"3fb00889",
  1208 => x"3d238551",
  1209 => x"90f23fb0",
  1210 => x"08028405",
  1211 => x"9e052386",
  1212 => x"5190e53f",
  1213 => x"b0088a3d",
  1214 => x"23800b81",
  1215 => x"b1e0088c",
  1216 => x"11085153",
  1217 => x"55747227",
  1218 => x"b8387154",
  1219 => x"8c3d7510",
  1220 => x"05f81122",
  1221 => x"70902bf0",
  1222 => x"13227084",
  1223 => x"80802972",
  1224 => x"902c057a",
  1225 => x"0c525558",
  1226 => x"81167081",
  1227 => x"ff065254",
  1228 => x"5274822e",
  1229 => x"94387184",
  1230 => x"17ff1656",
  1231 => x"575573cc",
  1232 => x"38800bb0",
  1233 => x"0c8c3d0d",
  1234 => x"04800b84",
  1235 => x"17ff1656",
  1236 => x"575573ff",
  1237 => x"b738ea39",
  1238 => x"fe3d0d81",
  1239 => x"518ff93f",
  1240 => x"b00881ff",
  1241 => x"0681b1dc",
  1242 => x"08718812",
  1243 => x"0c53b00c",
  1244 => x"843d0d04",
  1245 => x"803d0d81",
  1246 => x"51918f3f",
  1247 => x"b00883ff",
  1248 => x"ff0651ea",
  1249 => x"c83fb008",
  1250 => x"83ffff06",
  1251 => x"b00c823d",
  1252 => x"0d04803d",
  1253 => x"0d81518f",
  1254 => x"bf3fb008",
  1255 => x"81ff0651",
  1256 => x"a0b93f80",
  1257 => x"0bb00c82",
  1258 => x"3d0d0480",
  1259 => x"3d0d81b2",
  1260 => x"a80851f8",
  1261 => x"bb9586a1",
  1262 => x"710c810b",
  1263 => x"b00c823d",
  1264 => x"0d04fc3d",
  1265 => x"0d81518f",
  1266 => x"8f3fb008",
  1267 => x"81ff0654",
  1268 => x"82518f84",
  1269 => x"3fb00881",
  1270 => x"ff0681b2",
  1271 => x"9c088411",
  1272 => x"0870fe8f",
  1273 => x"0a067798",
  1274 => x"2b075154",
  1275 => x"56537280",
  1276 => x"2e863871",
  1277 => x"810a0752",
  1278 => x"7184160c",
  1279 => x"71b00c86",
  1280 => x"3d0d04fd",
  1281 => x"3d0d81b2",
  1282 => x"9c088411",
  1283 => x"08555381",
  1284 => x"518ec53f",
  1285 => x"b00881ff",
  1286 => x"0674dfff",
  1287 => x"ff065452",
  1288 => x"71802e87",
  1289 => x"3873a080",
  1290 => x"80075382",
  1291 => x"518ea93f",
  1292 => x"b00881ff",
  1293 => x"0673efff",
  1294 => x"0a065552",
  1295 => x"71802e87",
  1296 => x"38729080",
  1297 => x"0a075483",
  1298 => x"518e8d3f",
  1299 => x"b00881ff",
  1300 => x"0674f7ff",
  1301 => x"0a065452",
  1302 => x"71802e87",
  1303 => x"38738880",
  1304 => x"0a075384",
  1305 => x"518df13f",
  1306 => x"b00881ff",
  1307 => x"0673fbff",
  1308 => x"0a065552",
  1309 => x"71802e87",
  1310 => x"38728480",
  1311 => x"0a075485",
  1312 => x"518dd53f",
  1313 => x"b00881ff",
  1314 => x"0674fdff",
  1315 => x"0a065452",
  1316 => x"71802e87",
  1317 => x"38738280",
  1318 => x"0a075381",
  1319 => x"b29c0873",
  1320 => x"84120c54",
  1321 => x"72b00c85",
  1322 => x"3d0d04fc",
  1323 => x"3d0d81b2",
  1324 => x"9c087008",
  1325 => x"81a19c53",
  1326 => x"5555bbc2",
  1327 => x"3f739e2a",
  1328 => x"81065271",
  1329 => x"802eb638",
  1330 => x"81a1ac51",
  1331 => x"bbb03f81",
  1332 => x"518d853f",
  1333 => x"b00881ff",
  1334 => x"0681b29c",
  1335 => x"08841108",
  1336 => x"70fd0a06",
  1337 => x"56565652",
  1338 => x"71802e86",
  1339 => x"3873820a",
  1340 => x"07537284",
  1341 => x"160c72b0",
  1342 => x"0c863d0d",
  1343 => x"0481a1b4",
  1344 => x"51bafb3f",
  1345 => x"c339fd3d",
  1346 => x"0d81c1f4",
  1347 => x"0852f881",
  1348 => x"c08e800b",
  1349 => x"81b29c08",
  1350 => x"55537180",
  1351 => x"2e80f738",
  1352 => x"7281ff06",
  1353 => x"84150c81",
  1354 => x"b1d83370",
  1355 => x"81ff0651",
  1356 => x"5271802e",
  1357 => x"80c23872",
  1358 => x"9f2a7310",
  1359 => x"075381c1",
  1360 => x"f8337081",
  1361 => x"ff065152",
  1362 => x"71802ed4",
  1363 => x"38800b81",
  1364 => x"c1f83490",
  1365 => x"883f81b1",
  1366 => x"e8335473",
  1367 => x"80e23881",
  1368 => x"b29c0873",
  1369 => x"81ff0684",
  1370 => x"120c81b1",
  1371 => x"d8337081",
  1372 => x"ff065153",
  1373 => x"5471c038",
  1374 => x"72812a73",
  1375 => x"9f2b0753",
  1376 => x"ffbc3972",
  1377 => x"812a739f",
  1378 => x"2b075380",
  1379 => x"fd51bd81",
  1380 => x"3f81b29c",
  1381 => x"08547281",
  1382 => x"ff068415",
  1383 => x"0c81b1d8",
  1384 => x"337081ff",
  1385 => x"06535471",
  1386 => x"802ed838",
  1387 => x"729f2a73",
  1388 => x"10075380",
  1389 => x"fd51bcd9",
  1390 => x"3f81b29c",
  1391 => x"0854d739",
  1392 => x"800bb00c",
  1393 => x"853d0d04",
  1394 => x"f73d0d85",
  1395 => x"3d549653",
  1396 => x"81a1bc52",
  1397 => x"735180c0",
  1398 => x"bd3fa3b8",
  1399 => x"3f81518a",
  1400 => x"f73f8052",
  1401 => x"8051a289",
  1402 => x"3f735380",
  1403 => x"5281a6bc",
  1404 => x"51b4f43f",
  1405 => x"80528151",
  1406 => x"a1f73f73",
  1407 => x"53825281",
  1408 => x"a6bc51b4",
  1409 => x"e23f8052",
  1410 => x"8251a1e5",
  1411 => x"3f735381",
  1412 => x"5281a6bc",
  1413 => x"51b4d03f",
  1414 => x"80528451",
  1415 => x"a1d33f73",
  1416 => x"53845281",
  1417 => x"a6bc51b4",
  1418 => x"be3f8052",
  1419 => x"8551a1c1",
  1420 => x"3f735390",
  1421 => x"5281a6bc",
  1422 => x"51b4ac3f",
  1423 => x"80528651",
  1424 => x"a1af3f73",
  1425 => x"53835281",
  1426 => x"a6bc51b4",
  1427 => x"9a3f8b3d",
  1428 => x"0d04fef4",
  1429 => x"3f800bb0",
  1430 => x"0c04fc3d",
  1431 => x"0d818dec",
  1432 => x"54805584",
  1433 => x"527451a1",
  1434 => x"883f8053",
  1435 => x"73708105",
  1436 => x"553351a2",
  1437 => x"823f8113",
  1438 => x"7081ff06",
  1439 => x"515380dc",
  1440 => x"7327e938",
  1441 => x"81157081",
  1442 => x"ff065653",
  1443 => x"877527d3",
  1444 => x"38800bb0",
  1445 => x"0c863d0d",
  1446 => x"04fd3d0d",
  1447 => x"81b1d833",
  1448 => x"7081ff06",
  1449 => x"5454729f",
  1450 => x"26ab3881",
  1451 => x"b1d83370",
  1452 => x"81ff0681",
  1453 => x"b1dc0852",
  1454 => x"88120c54",
  1455 => x"80e452ad",
  1456 => x"99518df9",
  1457 => x"3f81b1d8",
  1458 => x"33810553",
  1459 => x"7281b1d8",
  1460 => x"34853d0d",
  1461 => x"0480e452",
  1462 => x"adee518d",
  1463 => x"e03f81b1",
  1464 => x"d8338105",
  1465 => x"537281b1",
  1466 => x"d834853d",
  1467 => x"0d04fd3d",
  1468 => x"0d81b1d8",
  1469 => x"337081ff",
  1470 => x"06545472",
  1471 => x"9f26b738",
  1472 => x"81b1d833",
  1473 => x"7081ff06",
  1474 => x"81b1dc08",
  1475 => x"5688160c",
  1476 => x"5381b1d8",
  1477 => x"33810554",
  1478 => x"7381b1d8",
  1479 => x"3481b1d8",
  1480 => x"33bf0654",
  1481 => x"7381b1d8",
  1482 => x"3480e452",
  1483 => x"adee518d",
  1484 => x"8c3f853d",
  1485 => x"0d0481b1",
  1486 => x"d8337081",
  1487 => x"ff06bf71",
  1488 => x"3181b1dc",
  1489 => x"08528812",
  1490 => x"0c555381",
  1491 => x"b1d83381",
  1492 => x"05547381",
  1493 => x"b1d83481",
  1494 => x"b1d833bf",
  1495 => x"06547381",
  1496 => x"b1d83480",
  1497 => x"e452adee",
  1498 => x"518cd23f",
  1499 => x"853d0d04",
  1500 => x"810b81b1",
  1501 => x"e83404fe",
  1502 => x"3d0d81b2",
  1503 => x"a0089811",
  1504 => x"0870842a",
  1505 => x"70810651",
  1506 => x"53535370",
  1507 => x"802e8d38",
  1508 => x"71ef0698",
  1509 => x"140c810b",
  1510 => x"81c1f834",
  1511 => x"843d0d04",
  1512 => x"fc3d0d81",
  1513 => x"b29c0870",
  1514 => x"08810a06",
  1515 => x"81c1f40c",
  1516 => x"53b9813f",
  1517 => x"b9a43f8d",
  1518 => x"c13f81b2",
  1519 => x"a0089811",
  1520 => x"08880798",
  1521 => x"120c5481",
  1522 => x"c1f40880",
  1523 => x"e4ce5553",
  1524 => x"72843888",
  1525 => x"80547381",
  1526 => x"d5f40c72",
  1527 => x"802e82e4",
  1528 => x"38819acc",
  1529 => x"51b5973f",
  1530 => x"8c51b4f8",
  1531 => x"3f81a1bc",
  1532 => x"51b58b3f",
  1533 => x"81c1f408",
  1534 => x"802e81b7",
  1535 => x"3881a1d4",
  1536 => x"51b4fb3f",
  1537 => x"81c1f408",
  1538 => x"802e8295",
  1539 => x"3881b29c",
  1540 => x"08841108",
  1541 => x"55558053",
  1542 => x"73fe8f0a",
  1543 => x"0673982b",
  1544 => x"07708417",
  1545 => x"0c811470",
  1546 => x"81ff0651",
  1547 => x"54548f73",
  1548 => x"27e63883",
  1549 => x"52aef051",
  1550 => x"8b833ff8",
  1551 => x"81c08e80",
  1552 => x"0b81b29c",
  1553 => x"08565481",
  1554 => x"c1f40880",
  1555 => x"2e81a838",
  1556 => x"7381ff06",
  1557 => x"84160c81",
  1558 => x"b1d83370",
  1559 => x"81ff0651",
  1560 => x"5372802e",
  1561 => x"80c23873",
  1562 => x"9f2a7410",
  1563 => x"075481c1",
  1564 => x"f8337081",
  1565 => x"ff065153",
  1566 => x"72802ed4",
  1567 => x"38800b81",
  1568 => x"c1f83489",
  1569 => x"d83f81b1",
  1570 => x"e8335574",
  1571 => x"81c23881",
  1572 => x"b29c0874",
  1573 => x"81ff0684",
  1574 => x"120c81b1",
  1575 => x"d8337081",
  1576 => x"ff065154",
  1577 => x"5572c038",
  1578 => x"73812a74",
  1579 => x"9f2b0754",
  1580 => x"ffbc3981",
  1581 => x"a1e051b3",
  1582 => x"c53f81a2",
  1583 => x"8451b3be",
  1584 => x"3fb451b5",
  1585 => x"833f81a2",
  1586 => x"9451b3b2",
  1587 => x"3f81a29c",
  1588 => x"51b3ab3f",
  1589 => x"81a2a851",
  1590 => x"b3a43f81",
  1591 => x"c1f408fe",
  1592 => x"ac38be39",
  1593 => x"73812a74",
  1594 => x"9f2b0754",
  1595 => x"80fd51b6",
  1596 => x"a03f81b2",
  1597 => x"9c085573",
  1598 => x"81ff0684",
  1599 => x"160c81b1",
  1600 => x"d8337081",
  1601 => x"ff065653",
  1602 => x"74802ed8",
  1603 => x"38739f2a",
  1604 => x"74100754",
  1605 => x"80fd51b5",
  1606 => x"f83f81b2",
  1607 => x"9c0855d7",
  1608 => x"39b6d852",
  1609 => x"acda5189",
  1610 => x"943f87e8",
  1611 => x"52ad9951",
  1612 => x"898b3fd5",
  1613 => x"e63f81b2",
  1614 => x"9c088411",
  1615 => x"08555580",
  1616 => x"53fdd539",
  1617 => x"b7d23f99",
  1618 => x"b03f9cc8",
  1619 => x"3ffd9239",
  1620 => x"b9b73f80",
  1621 => x"0b81d590",
  1622 => x"34800b81",
  1623 => x"d58c3480",
  1624 => x"0b81d594",
  1625 => x"0c04fc3d",
  1626 => x"0d765281",
  1627 => x"d58c3370",
  1628 => x"10101071",
  1629 => x"100581c1",
  1630 => x"fc055254",
  1631 => x"bea63f77",
  1632 => x"5281d58c",
  1633 => x"33709029",
  1634 => x"71317010",
  1635 => x"1081c4bc",
  1636 => x"05535555",
  1637 => x"be8e3f81",
  1638 => x"d58c3370",
  1639 => x"101081d3",
  1640 => x"bc057a71",
  1641 => x"0c548105",
  1642 => x"537281d5",
  1643 => x"8c34863d",
  1644 => x"0d04803d",
  1645 => x"0d81a2dc",
  1646 => x"51b1c33f",
  1647 => x"823d0d04",
  1648 => x"fe3d0d81",
  1649 => x"d5940853",
  1650 => x"72853884",
  1651 => x"3d0d0472",
  1652 => x"2db00853",
  1653 => x"800b81d5",
  1654 => x"940cb008",
  1655 => x"8c3881a2",
  1656 => x"dc51b19a",
  1657 => x"3f843d0d",
  1658 => x"0481a5f0",
  1659 => x"51b18f3f",
  1660 => x"7283ffff",
  1661 => x"26aa3881",
  1662 => x"ff732796",
  1663 => x"38725290",
  1664 => x"51b19e3f",
  1665 => x"8a51b0dc",
  1666 => x"3f81a2dc",
  1667 => x"51b0ef3f",
  1668 => x"d4397252",
  1669 => x"8851b189",
  1670 => x"3f8a51b0",
  1671 => x"c73fea39",
  1672 => x"7252a051",
  1673 => x"b0fb3f8a",
  1674 => x"51b0b93f",
  1675 => x"dc39fa3d",
  1676 => x"0d02a305",
  1677 => x"3356758d",
  1678 => x"2e80f438",
  1679 => x"75883270",
  1680 => x"307780ff",
  1681 => x"32703072",
  1682 => x"80257180",
  1683 => x"25075451",
  1684 => x"56585574",
  1685 => x"95389f76",
  1686 => x"278c3881",
  1687 => x"d5903355",
  1688 => x"80ce7527",
  1689 => x"ae38883d",
  1690 => x"0d0481d5",
  1691 => x"90335675",
  1692 => x"802ef338",
  1693 => x"8851afec",
  1694 => x"3fa051af",
  1695 => x"e73f8851",
  1696 => x"afe23f81",
  1697 => x"d59033ff",
  1698 => x"05577681",
  1699 => x"d5903488",
  1700 => x"3d0d0475",
  1701 => x"51afcd3f",
  1702 => x"81d59033",
  1703 => x"81115557",
  1704 => x"7381d590",
  1705 => x"347581d4",
  1706 => x"bc183488",
  1707 => x"3d0d048a",
  1708 => x"51afb13f",
  1709 => x"81d59033",
  1710 => x"81115654",
  1711 => x"7481d590",
  1712 => x"34800b81",
  1713 => x"d4bc1534",
  1714 => x"8056800b",
  1715 => x"81d4bc17",
  1716 => x"33565474",
  1717 => x"a02e8338",
  1718 => x"81547480",
  1719 => x"2e903873",
  1720 => x"802e8b38",
  1721 => x"81167081",
  1722 => x"ff065757",
  1723 => x"dd397580",
  1724 => x"2ebf3880",
  1725 => x"0b81d58c",
  1726 => x"33555574",
  1727 => x"7427ab38",
  1728 => x"73577410",
  1729 => x"10107510",
  1730 => x"05765481",
  1731 => x"d4bc5381",
  1732 => x"c1fc0551",
  1733 => x"bcda3fb0",
  1734 => x"08802ea6",
  1735 => x"38811570",
  1736 => x"81ff0656",
  1737 => x"54767526",
  1738 => x"d93881a2",
  1739 => x"e051aece",
  1740 => x"3f81a2dc",
  1741 => x"51aec73f",
  1742 => x"800b81d5",
  1743 => x"9034883d",
  1744 => x"0d047410",
  1745 => x"1081d3bc",
  1746 => x"05700881",
  1747 => x"d5940c56",
  1748 => x"800b81d5",
  1749 => x"9034e739",
  1750 => x"f73d0d02",
  1751 => x"af053359",
  1752 => x"800b81d4",
  1753 => x"bc3381d4",
  1754 => x"bc595556",
  1755 => x"73a02e09",
  1756 => x"81069638",
  1757 => x"81167081",
  1758 => x"ff0681d4",
  1759 => x"bc117033",
  1760 => x"53595754",
  1761 => x"73a02eec",
  1762 => x"38805877",
  1763 => x"792780ea",
  1764 => x"38807733",
  1765 => x"56547474",
  1766 => x"2e833881",
  1767 => x"5474a02e",
  1768 => x"9a387380",
  1769 => x"c53874a0",
  1770 => x"2e913881",
  1771 => x"187081ff",
  1772 => x"06595578",
  1773 => x"7826da38",
  1774 => x"80c03981",
  1775 => x"167081ff",
  1776 => x"0681d4bc",
  1777 => x"11703357",
  1778 => x"52575773",
  1779 => x"a02e0981",
  1780 => x"06d93881",
  1781 => x"167081ff",
  1782 => x"0681d4bc",
  1783 => x"11703357",
  1784 => x"52575773",
  1785 => x"a02ed438",
  1786 => x"c2398116",
  1787 => x"7081ff06",
  1788 => x"81d4bc11",
  1789 => x"595755ff",
  1790 => x"98398a53",
  1791 => x"8b3dfc05",
  1792 => x"527651bf",
  1793 => x"b03f8b3d",
  1794 => x"0d04f73d",
  1795 => x"0d02af05",
  1796 => x"3359800b",
  1797 => x"81d4bc33",
  1798 => x"81d4bc59",
  1799 => x"555673a0",
  1800 => x"2e098106",
  1801 => x"96388116",
  1802 => x"7081ff06",
  1803 => x"81d4bc11",
  1804 => x"70335359",
  1805 => x"575473a0",
  1806 => x"2eec3880",
  1807 => x"58777927",
  1808 => x"80ea3880",
  1809 => x"77335654",
  1810 => x"74742e83",
  1811 => x"38815474",
  1812 => x"a02e9a38",
  1813 => x"7380c538",
  1814 => x"74a02e91",
  1815 => x"38811870",
  1816 => x"81ff0659",
  1817 => x"55787826",
  1818 => x"da3880c0",
  1819 => x"39811670",
  1820 => x"81ff0681",
  1821 => x"d4bc1170",
  1822 => x"33575257",
  1823 => x"5773a02e",
  1824 => x"098106d9",
  1825 => x"38811670",
  1826 => x"81ff0681",
  1827 => x"d4bc1170",
  1828 => x"33575257",
  1829 => x"5773a02e",
  1830 => x"d438c239",
  1831 => x"81167081",
  1832 => x"ff0681d4",
  1833 => x"bc115957",
  1834 => x"55ff9839",
  1835 => x"90538b3d",
  1836 => x"fc055276",
  1837 => x"5180c19a",
  1838 => x"3f8b3d0d",
  1839 => x"04fc3d0d",
  1840 => x"8a51aba0",
  1841 => x"3f81a2f4",
  1842 => x"51abb33f",
  1843 => x"800b81d5",
  1844 => x"8c335353",
  1845 => x"72722780",
  1846 => x"f5387210",
  1847 => x"10107310",
  1848 => x"0581c1fc",
  1849 => x"05705254",
  1850 => x"ab943f72",
  1851 => x"842b7074",
  1852 => x"31822b81",
  1853 => x"c4bc1133",
  1854 => x"51535571",
  1855 => x"802eb738",
  1856 => x"7351b88d",
  1857 => x"3fb00881",
  1858 => x"ff065271",
  1859 => x"89269338",
  1860 => x"a051aad0",
  1861 => x"3f811270",
  1862 => x"81ff0653",
  1863 => x"54897227",
  1864 => x"ef3881a3",
  1865 => x"8c51aad6",
  1866 => x"3f747331",
  1867 => x"822b81c4",
  1868 => x"bc0551aa",
  1869 => x"c93f8a51",
  1870 => x"aaaa3f81",
  1871 => x"137081ff",
  1872 => x"0681d58c",
  1873 => x"33545455",
  1874 => x"717326ff",
  1875 => x"8d388a51",
  1876 => x"aa923f81",
  1877 => x"d58c33b0",
  1878 => x"0c863d0d",
  1879 => x"04fe3d0d",
  1880 => x"81d5ec22",
  1881 => x"ff055170",
  1882 => x"81d5ec23",
  1883 => x"7083ffff",
  1884 => x"06517080",
  1885 => x"c43881d5",
  1886 => x"f0335170",
  1887 => x"81ff2eb9",
  1888 => x"38701010",
  1889 => x"1081d59c",
  1890 => x"05527133",
  1891 => x"81d5f034",
  1892 => x"fe723481",
  1893 => x"d5f03370",
  1894 => x"10101081",
  1895 => x"d59c0552",
  1896 => x"53821122",
  1897 => x"81d5ec23",
  1898 => x"84120853",
  1899 => x"722d81d5",
  1900 => x"ec225170",
  1901 => x"802effbe",
  1902 => x"38843d0d",
  1903 => x"04f93d0d",
  1904 => x"02aa0522",
  1905 => x"56805574",
  1906 => x"10101081",
  1907 => x"d59c0570",
  1908 => x"33525270",
  1909 => x"81fe2e99",
  1910 => x"38811570",
  1911 => x"81ff0656",
  1912 => x"52748a2e",
  1913 => x"098106df",
  1914 => x"38810bb0",
  1915 => x"0c893d0d",
  1916 => x"0481d5f0",
  1917 => x"337081ff",
  1918 => x"0681d5ec",
  1919 => x"22535458",
  1920 => x"7281ff2e",
  1921 => x"b0387283",
  1922 => x"2b547076",
  1923 => x"2780de38",
  1924 => x"75713170",
  1925 => x"83ffff06",
  1926 => x"7481d59c",
  1927 => x"17337083",
  1928 => x"2b81d59e",
  1929 => x"11225658",
  1930 => x"56525757",
  1931 => x"7281ff2e",
  1932 => x"098106d6",
  1933 => x"38727234",
  1934 => x"75821323",
  1935 => x"7984130c",
  1936 => x"7781ff06",
  1937 => x"5473732e",
  1938 => x"96387610",
  1939 => x"101081d5",
  1940 => x"9c055374",
  1941 => x"73348051",
  1942 => x"70b00c89",
  1943 => x"3d0d0474",
  1944 => x"81d5f034",
  1945 => x"7581d5ec",
  1946 => x"238051ec",
  1947 => x"39707631",
  1948 => x"517081d5",
  1949 => x"9e1523ff",
  1950 => x"bc39ff3d",
  1951 => x"0d8a5271",
  1952 => x"10101081",
  1953 => x"d5940551",
  1954 => x"fe7134ff",
  1955 => x"127081ff",
  1956 => x"06535171",
  1957 => x"ea38ff0b",
  1958 => x"81d5f034",
  1959 => x"833d0d04",
  1960 => x"f53d0d7d",
  1961 => x"598a5481",
  1962 => x"028405ba",
  1963 => x"0522575c",
  1964 => x"80e45380",
  1965 => x"52abb93f",
  1966 => x"b008722e",
  1967 => x"09810683",
  1968 => x"38815272",
  1969 => x"802eb138",
  1970 => x"71802e91",
  1971 => x"3880e451",
  1972 => x"aabf3fff",
  1973 => x"137081ff",
  1974 => x"065452d7",
  1975 => x"3972802e",
  1976 => x"9738ab9f",
  1977 => x"3fb00881",
  1978 => x"ff065271",
  1979 => x"952e829a",
  1980 => x"387180c3",
  1981 => x"2e81ec38",
  1982 => x"ff147081",
  1983 => x"ff065553",
  1984 => x"73ffad38",
  1985 => x"75802e81",
  1986 => x"cc388a7c",
  1987 => x"095c5a81",
  1988 => x"51ab923f",
  1989 => x"7b51ab8d",
  1990 => x"3f7a51ab",
  1991 => x"883f8070",
  1992 => x"55578180",
  1993 => x"55ff1570",
  1994 => x"81ff0656",
  1995 => x"529a5375",
  1996 => x"802e9138",
  1997 => x"78708105",
  1998 => x"5a33ff17",
  1999 => x"7083ffff",
  2000 => x"06585353",
  2001 => x"7251aadd",
  2002 => x"3f77802e",
  2003 => x"81a93872",
  2004 => x"882b7432",
  2005 => x"53875472",
  2006 => x"902b5280",
  2007 => x"72248188",
  2008 => x"38721083",
  2009 => x"fffe0653",
  2010 => x"ff145473",
  2011 => x"8025e838",
  2012 => x"7283ffff",
  2013 => x"065474ff",
  2014 => x"ac387780",
  2015 => x"2e818338",
  2016 => x"73882a51",
  2017 => x"aa9f3f73",
  2018 => x"81ff0651",
  2019 => x"aa973fa9",
  2020 => x"df3fb008",
  2021 => x"fa38a9eb",
  2022 => x"3fb00881",
  2023 => x"ff065271",
  2024 => x"862e80eb",
  2025 => x"3871982e",
  2026 => x"80f038ff",
  2027 => x"1a7081ff",
  2028 => x"065b5479",
  2029 => x"fed938fe",
  2030 => x"5271b00c",
  2031 => x"8d3d0d04",
  2032 => x"a9ae3fb0",
  2033 => x"08fa38a9",
  2034 => x"ba3fb008",
  2035 => x"81ff0652",
  2036 => x"71862ee5",
  2037 => x"388451a9",
  2038 => x"cc3fa994",
  2039 => x"3fb008e0",
  2040 => x"38e53981",
  2041 => x"58fe9d39",
  2042 => x"7210a0a1",
  2043 => x"327083ff",
  2044 => x"ff065452",
  2045 => x"fef23972",
  2046 => x"177081ff",
  2047 => x"065852fe",
  2048 => x"f5397651",
  2049 => x"a99f3fff",
  2050 => x"86398058",
  2051 => x"fdf63981",
  2052 => x"1c7081ff",
  2053 => x"065d55fd",
  2054 => x"eb39ff0b",
  2055 => x"b00c8d3d",
  2056 => x"0d04f63d",
  2057 => x"0d7c7e5b",
  2058 => x"5980c357",
  2059 => x"8a55815b",
  2060 => x"805880e4",
  2061 => x"53805477",
  2062 => x"7a2482aa",
  2063 => x"387651a8",
  2064 => x"e43f8052",
  2065 => x"a8aa3fb0",
  2066 => x"08722e09",
  2067 => x"81068338",
  2068 => x"81527280",
  2069 => x"2e81e638",
  2070 => x"71802e91",
  2071 => x"3880e451",
  2072 => x"a7af3fff",
  2073 => x"137081ff",
  2074 => x"065452d6",
  2075 => x"3972802e",
  2076 => x"81cb38a8",
  2077 => x"8e3fb008",
  2078 => x"81ff0652",
  2079 => x"71842e82",
  2080 => x"81387184",
  2081 => x"2481ca38",
  2082 => x"71812e09",
  2083 => x"810681ad",
  2084 => x"388657a7",
  2085 => x"ee3fb008",
  2086 => x"81ff0653",
  2087 => x"7a732e83",
  2088 => x"389557a7",
  2089 => x"de3fb008",
  2090 => x"097081ff",
  2091 => x"0657527a",
  2092 => x"762e8338",
  2093 => x"95578053",
  2094 => x"a7c93f78",
  2095 => x"1356b008",
  2096 => x"76348113",
  2097 => x"7081ff06",
  2098 => x"70982b58",
  2099 => x"54527580",
  2100 => x"25e63880",
  2101 => x"56781670",
  2102 => x"3370882b",
  2103 => x"76325253",
  2104 => x"53875472",
  2105 => x"902b5280",
  2106 => x"72248187",
  2107 => x"38721083",
  2108 => x"fffe0653",
  2109 => x"ff145473",
  2110 => x"8025e838",
  2111 => x"7283ffff",
  2112 => x"06811770",
  2113 => x"81ff0670",
  2114 => x"982b5658",
  2115 => x"53547280",
  2116 => x"25c338a6",
  2117 => x"ee3fb008",
  2118 => x"81ff0674",
  2119 => x"882a5753",
  2120 => x"72762e83",
  2121 => x"389557a6",
  2122 => x"da3fb008",
  2123 => x"81ff0674",
  2124 => x"81ff0653",
  2125 => x"5675722e",
  2126 => x"80d43895",
  2127 => x"57ff1570",
  2128 => x"81ff0656",
  2129 => x"5274fdea",
  2130 => x"38fe0bb0",
  2131 => x"0c8c3d0d",
  2132 => x"0471982e",
  2133 => x"098106e5",
  2134 => x"388651a6",
  2135 => x"c83fff0b",
  2136 => x"b00c8c3d",
  2137 => x"0d049851",
  2138 => x"a6bb3ffd",
  2139 => x"0bb00c8c",
  2140 => x"3d0d0472",
  2141 => x"10a0a132",
  2142 => x"7083ffff",
  2143 => x"065452fe",
  2144 => x"f3398651",
  2145 => x"a69f3f77",
  2146 => x"b00c8c3d",
  2147 => x"0d047686",
  2148 => x"2e098106",
  2149 => x"ffa73877",
  2150 => x"84808029",
  2151 => x"82800a05",
  2152 => x"70902c81",
  2153 => x"801b811e",
  2154 => x"7081ff06",
  2155 => x"5f575b59",
  2156 => x"5374fcfe",
  2157 => x"38ff9239",
  2158 => x"fe3d0d02",
  2159 => x"93053302",
  2160 => x"84059705",
  2161 => x"33545271",
  2162 => x"812e9238",
  2163 => x"7180d52e",
  2164 => x"bb3881a3",
  2165 => x"9051a1a6",
  2166 => x"3f843d0d",
  2167 => x"0481a39c",
  2168 => x"51a19b3f",
  2169 => x"72912e81",
  2170 => x"d9387291",
  2171 => x"24b53872",
  2172 => x"8c2e81e4",
  2173 => x"38728c24",
  2174 => x"80dc3872",
  2175 => x"862e81b7",
  2176 => x"3881a3a8",
  2177 => x"51a0f73f",
  2178 => x"843d0d04",
  2179 => x"81a3b851",
  2180 => x"a0ec3f72",
  2181 => x"8726ea38",
  2182 => x"72101081",
  2183 => x"a69c0552",
  2184 => x"71080472",
  2185 => x"a82e81a5",
  2186 => x"3872a824",
  2187 => x"9438729a",
  2188 => x"2e098106",
  2189 => x"cc3881a3",
  2190 => x"c451a0c2",
  2191 => x"3f843d0d",
  2192 => x"047280e1",
  2193 => x"2e098106",
  2194 => x"ffb73881",
  2195 => x"a3e051a0",
  2196 => x"ad3f843d",
  2197 => x"0d04728f",
  2198 => x"2e098106",
  2199 => x"ffa33881",
  2200 => x"a3f051a0",
  2201 => x"993f843d",
  2202 => x"0d0481a4",
  2203 => x"8c51a08e",
  2204 => x"3f843d0d",
  2205 => x"0481a1bc",
  2206 => x"51a0833f",
  2207 => x"843d0d04",
  2208 => x"81a4a451",
  2209 => x"9ff83f84",
  2210 => x"3d0d0481",
  2211 => x"a4b8519f",
  2212 => x"ed3f843d",
  2213 => x"0d0481a4",
  2214 => x"c8519fe2",
  2215 => x"3f843d0d",
  2216 => x"0481a4e0",
  2217 => x"519fd73f",
  2218 => x"843d0d04",
  2219 => x"81a4f451",
  2220 => x"9fcc3f84",
  2221 => x"3d0d0481",
  2222 => x"a584519f",
  2223 => x"c13f843d",
  2224 => x"0d0481a5",
  2225 => x"94519fb6",
  2226 => x"3f843d0d",
  2227 => x"0481a5a8",
  2228 => x"519fab3f",
  2229 => x"843d0d04",
  2230 => x"81a5c851",
  2231 => x"9fa03f84",
  2232 => x"3d0d04f7",
  2233 => x"3d0d02b3",
  2234 => x"05337c70",
  2235 => x"08c08080",
  2236 => x"0659545a",
  2237 => x"80567583",
  2238 => x"2b7707bf",
  2239 => x"e0800770",
  2240 => x"70840552",
  2241 => x"0871088c",
  2242 => x"2abffe80",
  2243 => x"06790771",
  2244 => x"982a728c",
  2245 => x"2a9fff06",
  2246 => x"73852a70",
  2247 => x"8f06759f",
  2248 => x"06565158",
  2249 => x"5d585255",
  2250 => x"58748d38",
  2251 => x"8116568f",
  2252 => x"7627c338",
  2253 => x"8b3d0d04",
  2254 => x"81a5d851",
  2255 => x"9ec03f75",
  2256 => x"51a0853f",
  2257 => x"8452b008",
  2258 => x"51d0943f",
  2259 => x"81a5e451",
  2260 => x"9eac3f74",
  2261 => x"5288519e",
  2262 => x"c83f8452",
  2263 => x"b00851cf",
  2264 => x"fe3f81a5",
  2265 => x"ec519e96",
  2266 => x"3f785290",
  2267 => x"519eb23f",
  2268 => x"8652b008",
  2269 => x"51cfe83f",
  2270 => x"81a5f451",
  2271 => x"9e803f72",
  2272 => x"519fc53f",
  2273 => x"8452b008",
  2274 => x"51cfd43f",
  2275 => x"81a5fc51",
  2276 => x"9dec3f73",
  2277 => x"519fb13f",
  2278 => x"8452b008",
  2279 => x"51cfc03f",
  2280 => x"81a68451",
  2281 => x"9dd83f77",
  2282 => x"52a0519d",
  2283 => x"f43f8a52",
  2284 => x"b00851cf",
  2285 => x"aa3f7992",
  2286 => x"388a519d",
  2287 => x"a73f8116",
  2288 => x"568f7627",
  2289 => x"feb038fe",
  2290 => x"eb397881",
  2291 => x"ff065274",
  2292 => x"51fbe53f",
  2293 => x"8a519d8c",
  2294 => x"3fe439f8",
  2295 => x"3d0d02ab",
  2296 => x"05335980",
  2297 => x"5675852b",
  2298 => x"e09011e0",
  2299 => x"80120870",
  2300 => x"982a718c",
  2301 => x"2a9fff06",
  2302 => x"72852a70",
  2303 => x"8f06749f",
  2304 => x"06555158",
  2305 => x"5b535659",
  2306 => x"5574802e",
  2307 => x"81a13875",
  2308 => x"bf2681a9",
  2309 => x"3881a68c",
  2310 => x"519ce33f",
  2311 => x"75519ea8",
  2312 => x"3f8652b0",
  2313 => x"0851ceb7",
  2314 => x"3f81a5e4",
  2315 => x"519ccf3f",
  2316 => x"74528851",
  2317 => x"9ceb3f84",
  2318 => x"52b00851",
  2319 => x"cea13f81",
  2320 => x"a5ec519c",
  2321 => x"b93f7652",
  2322 => x"90519cd5",
  2323 => x"3f8652b0",
  2324 => x"0851ce8b",
  2325 => x"3f81a5f4",
  2326 => x"519ca33f",
  2327 => x"72519de8",
  2328 => x"3f8452b0",
  2329 => x"0851cdf7",
  2330 => x"3f81a5fc",
  2331 => x"519c8f3f",
  2332 => x"73519dd4",
  2333 => x"3f8452b0",
  2334 => x"0851cde3",
  2335 => x"3f81a684",
  2336 => x"519bfb3f",
  2337 => x"7708c080",
  2338 => x"800652a0",
  2339 => x"519c923f",
  2340 => x"8a52b008",
  2341 => x"51cdc83f",
  2342 => x"7881ac38",
  2343 => x"8a519bc4",
  2344 => x"3f805374",
  2345 => x"812e81d9",
  2346 => x"3876862e",
  2347 => x"81b53881",
  2348 => x"165680ff",
  2349 => x"7627fead",
  2350 => x"388a3d0d",
  2351 => x"0481a694",
  2352 => x"519bbb3f",
  2353 => x"c016519c",
  2354 => x"ff3f8652",
  2355 => x"b00851cd",
  2356 => x"8e3f81a5",
  2357 => x"e4519ba6",
  2358 => x"3f745288",
  2359 => x"519bc23f",
  2360 => x"8452b008",
  2361 => x"51ccf83f",
  2362 => x"81a5ec51",
  2363 => x"9b903f76",
  2364 => x"5290519b",
  2365 => x"ac3f8652",
  2366 => x"b00851cc",
  2367 => x"e23f81a5",
  2368 => x"f4519afa",
  2369 => x"3f72519c",
  2370 => x"bf3f8452",
  2371 => x"b00851cc",
  2372 => x"ce3f81a5",
  2373 => x"fc519ae6",
  2374 => x"3f73519c",
  2375 => x"ab3f8452",
  2376 => x"b00851cc",
  2377 => x"ba3f81a6",
  2378 => x"84519ad2",
  2379 => x"3f7708c0",
  2380 => x"80800652",
  2381 => x"a0519ae9",
  2382 => x"3f8a52b0",
  2383 => x"0851cc9f",
  2384 => x"3f78802e",
  2385 => x"fed63876",
  2386 => x"81ff0652",
  2387 => x"7451f8e8",
  2388 => x"3f8a519a",
  2389 => x"8f3f8053",
  2390 => x"74812e09",
  2391 => x"8106fec9",
  2392 => x"389f3972",
  2393 => x"81065776",
  2394 => x"802efec3",
  2395 => x"38785277",
  2396 => x"51faf03f",
  2397 => x"81165680",
  2398 => x"ff7627fc",
  2399 => x"e838feb9",
  2400 => x"39745376",
  2401 => x"862e0981",
  2402 => x"06fea438",
  2403 => x"d639803d",
  2404 => x"0d81b294",
  2405 => x"08519971",
  2406 => x"0c81800b",
  2407 => x"84120c81",
  2408 => x"b2900851",
  2409 => x"99710c81",
  2410 => x"800b8412",
  2411 => x"0c823d0d",
  2412 => x"04fe3d0d",
  2413 => x"74028405",
  2414 => x"97053302",
  2415 => x"88059b05",
  2416 => x"3388130c",
  2417 => x"8c120c53",
  2418 => x"8c130870",
  2419 => x"812a8106",
  2420 => x"515271f4",
  2421 => x"388c1308",
  2422 => x"7081ff06",
  2423 => x"b00c5184",
  2424 => x"3d0d0480",
  2425 => x"3d0d728c",
  2426 => x"11087087",
  2427 => x"2a813281",
  2428 => x"06b00c51",
  2429 => x"51823d0d",
  2430 => x"04fe3d0d",
  2431 => x"ff903f81",
  2432 => x"ec538190",
  2433 => x"5281b294",
  2434 => x"0851ffa5",
  2435 => x"3f9d5390",
  2436 => x"5281b294",
  2437 => x"0851ff99",
  2438 => x"3f80c553",
  2439 => x"80d05281",
  2440 => x"b2940851",
  2441 => x"ff8b3f81",
  2442 => x"ec538190",
  2443 => x"5281b294",
  2444 => x"0851fefd",
  2445 => x"3fa15390",
  2446 => x"5281b294",
  2447 => x"0851fef1",
  2448 => x"3f895380",
  2449 => x"d05281b2",
  2450 => x"940851fe",
  2451 => x"e43f81ec",
  2452 => x"53819052",
  2453 => x"81b29408",
  2454 => x"51fed63f",
  2455 => x"b3539052",
  2456 => x"81b29408",
  2457 => x"51feca3f",
  2458 => x"885380d0",
  2459 => x"5281b294",
  2460 => x"0851febd",
  2461 => x"3f81ec53",
  2462 => x"81905281",
  2463 => x"b2940851",
  2464 => x"feaf3fb4",
  2465 => x"53905281",
  2466 => x"b2940851",
  2467 => x"fea33f96",
  2468 => x"5380d052",
  2469 => x"81b29408",
  2470 => x"51fe963f",
  2471 => x"81ec5381",
  2472 => x"905281b2",
  2473 => x"940851fe",
  2474 => x"883fb653",
  2475 => x"905281b2",
  2476 => x"940851fd",
  2477 => x"fc3f80e0",
  2478 => x"5380d052",
  2479 => x"81b29408",
  2480 => x"51fdee3f",
  2481 => x"81ec5381",
  2482 => x"905281b2",
  2483 => x"940851fd",
  2484 => x"e03f80c9",
  2485 => x"53905281",
  2486 => x"b2940851",
  2487 => x"fdd33f81",
  2488 => x"c05380d0",
  2489 => x"5281b294",
  2490 => x"0851fdc5",
  2491 => x"3f843d0d",
  2492 => x"04fd3d0d",
  2493 => x"02970533",
  2494 => x"0284059b",
  2495 => x"05337181",
  2496 => x"b00781bf",
  2497 => x"06535454",
  2498 => x"f8808098",
  2499 => x"8071710c",
  2500 => x"73842a90",
  2501 => x"07710c73",
  2502 => x"8f06710c",
  2503 => x"527281b1",
  2504 => x"f0347381",
  2505 => x"b1f43485",
  2506 => x"3d0d04fd",
  2507 => x"3d0d0297",
  2508 => x"053381b1",
  2509 => x"f4335473",
  2510 => x"05870602",
  2511 => x"84059a05",
  2512 => x"2281b1f0",
  2513 => x"33547305",
  2514 => x"7081ff06",
  2515 => x"7281b007",
  2516 => x"54515454",
  2517 => x"f8808098",
  2518 => x"8071710c",
  2519 => x"73842a90",
  2520 => x"07710c73",
  2521 => x"8f06710c",
  2522 => x"527281b1",
  2523 => x"f0347381",
  2524 => x"b1f43485",
  2525 => x"3d0d04ff",
  2526 => x"3d0d028f",
  2527 => x"0533f880",
  2528 => x"8098840c",
  2529 => x"81b1f033",
  2530 => x"81055170",
  2531 => x"81b1f034",
  2532 => x"833d0d04",
  2533 => x"ff3d0d80",
  2534 => x"c00bf880",
  2535 => x"8098800c",
  2536 => x"81a10bf8",
  2537 => x"80809880",
  2538 => x"0c81c00b",
  2539 => x"f8808098",
  2540 => x"800c81a4",
  2541 => x"0bf88080",
  2542 => x"98800c81",
  2543 => x"a60bf880",
  2544 => x"8098800c",
  2545 => x"81a20bf8",
  2546 => x"80809880",
  2547 => x"0caf0bf8",
  2548 => x"80809880",
  2549 => x"0ca50bf8",
  2550 => x"80809880",
  2551 => x"0c81810b",
  2552 => x"f8808098",
  2553 => x"800c9d0b",
  2554 => x"f8808098",
  2555 => x"800c81fa",
  2556 => x"0bf88080",
  2557 => x"98800c80",
  2558 => x"0bf88080",
  2559 => x"98800c80",
  2560 => x"527181b0",
  2561 => x"0781bf06",
  2562 => x"f8808098",
  2563 => x"800c900b",
  2564 => x"f8808098",
  2565 => x"800c800b",
  2566 => x"f8808098",
  2567 => x"800c8051",
  2568 => x"800bf880",
  2569 => x"8098840c",
  2570 => x"81117081",
  2571 => x"ff065151",
  2572 => x"80e57127",
  2573 => x"eb388112",
  2574 => x"7081ff06",
  2575 => x"53518772",
  2576 => x"27ffbe38",
  2577 => x"81b00bf8",
  2578 => x"80809880",
  2579 => x"0c900bf8",
  2580 => x"80809880",
  2581 => x"0c800bf8",
  2582 => x"80809880",
  2583 => x"0c800b81",
  2584 => x"b1f03480",
  2585 => x"0b81b1f4",
  2586 => x"3481af0b",
  2587 => x"f8808098",
  2588 => x"800c833d",
  2589 => x"0d04ed3d",
  2590 => x"0d650284",
  2591 => x"0580db05",
  2592 => x"33028805",
  2593 => x"80df0533",
  2594 => x"5f5a5680",
  2595 => x"7981067a",
  2596 => x"812a8106",
  2597 => x"7b832b81",
  2598 => x"80067c82",
  2599 => x"2a810657",
  2600 => x"5e435f5c",
  2601 => x"81ff4272",
  2602 => x"7c2e0981",
  2603 => x"0683387b",
  2604 => x"42881608",
  2605 => x"5574802e",
  2606 => x"839f3885",
  2607 => x"16335aff",
  2608 => x"537c7a26",
  2609 => x"8e388416",
  2610 => x"3354737d",
  2611 => x"2685387c",
  2612 => x"74315374",
  2613 => x"13703354",
  2614 => x"577281ff",
  2615 => x"06831733",
  2616 => x"70982b81",
  2617 => x"ff0a119b",
  2618 => x"2a810551",
  2619 => x"5a404081",
  2620 => x"53748338",
  2621 => x"74537281",
  2622 => x"ff064380",
  2623 => x"7a81ff06",
  2624 => x"4557ff54",
  2625 => x"7c64268b",
  2626 => x"38841633",
  2627 => x"537c7327",
  2628 => x"83ce3873",
  2629 => x"7481ff06",
  2630 => x"5553805a",
  2631 => x"797324ab",
  2632 => x"38747a2e",
  2633 => x"09810682",
  2634 => x"bb387e98",
  2635 => x"2b81ff0a",
  2636 => x"119b2a82",
  2637 => x"18337171",
  2638 => x"29117081",
  2639 => x"ff067871",
  2640 => x"298c1c08",
  2641 => x"0552435d",
  2642 => x"5758447f",
  2643 => x"63057081",
  2644 => x"ff067063",
  2645 => x"2b7081ff",
  2646 => x"067b622b",
  2647 => x"7081ff06",
  2648 => x"7e832a81",
  2649 => x"065c5557",
  2650 => x"5256455f",
  2651 => x"75802e8f",
  2652 => x"3881b1f0",
  2653 => x"33640559",
  2654 => x"7880e624",
  2655 => x"8dc6387f",
  2656 => x"78296430",
  2657 => x"5e577b7e",
  2658 => x"2c982b70",
  2659 => x"982c5540",
  2660 => x"73772580",
  2661 => x"fc38ff1f",
  2662 => x"7c81065a",
  2663 => x"537b732e",
  2664 => x"83843860",
  2665 => x"85da3861",
  2666 => x"84a5387d",
  2667 => x"802e81fe",
  2668 => x"38791470",
  2669 => x"33705254",
  2670 => x"56805578",
  2671 => x"752e8538",
  2672 => x"72842a56",
  2673 => x"75832a81",
  2674 => x"06407f80",
  2675 => x"2e843881",
  2676 => x"c0557582",
  2677 => x"2a810640",
  2678 => x"7f802e85",
  2679 => x"3874b007",
  2680 => x"5575812a",
  2681 => x"8106407f",
  2682 => x"802e8538",
  2683 => x"748c0755",
  2684 => x"75810653",
  2685 => x"72802e85",
  2686 => x"38748307",
  2687 => x"557451fa",
  2688 => x"f63f7714",
  2689 => x"982b7098",
  2690 => x"2c555576",
  2691 => x"7424ffa1",
  2692 => x"3862802e",
  2693 => x"9638617f",
  2694 => x"ff055654",
  2695 => x"7b752e81",
  2696 => x"e3387351",
  2697 => x"fad13f60",
  2698 => x"81bd387c",
  2699 => x"528151f9",
  2700 => x"fa3f811c",
  2701 => x"7081ff06",
  2702 => x"5d547e7c",
  2703 => x"26fec738",
  2704 => x"63527e30",
  2705 => x"70982b70",
  2706 => x"982c535c",
  2707 => x"5cf9dc3f",
  2708 => x"635372b0",
  2709 => x"0c953d0d",
  2710 => x"04821633",
  2711 => x"8517335b",
  2712 => x"53fcf639",
  2713 => x"73802eaf",
  2714 => x"38ff1470",
  2715 => x"81ff0655",
  2716 => x"537381ff",
  2717 => x"2ea13874",
  2718 => x"70810556",
  2719 => x"33770570",
  2720 => x"83ffff06",
  2721 => x"ff167081",
  2722 => x"ff065755",
  2723 => x"585a7381",
  2724 => x"ff2e0981",
  2725 => x"06e1387e",
  2726 => x"982b81ff",
  2727 => x"0a119b2a",
  2728 => x"70792919",
  2729 => x"8c190805",
  2730 => x"5c4055fd",
  2731 => x"9e397914",
  2732 => x"70335259",
  2733 => x"f9c13f77",
  2734 => x"14982b70",
  2735 => x"982c5553",
  2736 => x"737725fe",
  2737 => x"cc387914",
  2738 => x"70335259",
  2739 => x"f9a93f77",
  2740 => x"14982b70",
  2741 => x"982c5553",
  2742 => x"767424d2",
  2743 => x"38feb239",
  2744 => x"7c733154",
  2745 => x"fcad3973",
  2746 => x"51f98c3f",
  2747 => x"7c528151",
  2748 => x"f8b93f81",
  2749 => x"1c7081ff",
  2750 => x"065d547e",
  2751 => x"7c26fd86",
  2752 => x"38febd39",
  2753 => x"617b3270",
  2754 => x"81ff0655",
  2755 => x"567d802e",
  2756 => x"fe90387a",
  2757 => x"812a7432",
  2758 => x"705254f8",
  2759 => x"da3f6080",
  2760 => x"2efe8838",
  2761 => x"c2396087",
  2762 => x"8f386185",
  2763 => x"d3387d80",
  2764 => x"2e80e638",
  2765 => x"79147033",
  2766 => x"7c077052",
  2767 => x"54568055",
  2768 => x"78752e85",
  2769 => x"3872842a",
  2770 => x"5675832a",
  2771 => x"81065372",
  2772 => x"802e8438",
  2773 => x"81c05575",
  2774 => x"822a8106",
  2775 => x"5372802e",
  2776 => x"853874b0",
  2777 => x"07557581",
  2778 => x"2a810653",
  2779 => x"72802e85",
  2780 => x"38748c07",
  2781 => x"55758106",
  2782 => x"407f802e",
  2783 => x"85387483",
  2784 => x"07557451",
  2785 => x"f7f13f77",
  2786 => x"14982b70",
  2787 => x"982c5553",
  2788 => x"767424ff",
  2789 => x"9f38fcf9",
  2790 => x"39791470",
  2791 => x"337c0752",
  2792 => x"55f7d43f",
  2793 => x"7714982b",
  2794 => x"70982c55",
  2795 => x"59737725",
  2796 => x"fcdf3879",
  2797 => x"1470337c",
  2798 => x"075255f7",
  2799 => x"ba3f7714",
  2800 => x"982b7098",
  2801 => x"2c555976",
  2802 => x"7424ce38",
  2803 => x"fcc3397d",
  2804 => x"802e80ea",
  2805 => x"38791470",
  2806 => x"33705854",
  2807 => x"55805578",
  2808 => x"752e8538",
  2809 => x"72842a56",
  2810 => x"75832a81",
  2811 => x"06537280",
  2812 => x"2e843881",
  2813 => x"c0557582",
  2814 => x"2a810653",
  2815 => x"72802e85",
  2816 => x"3874b007",
  2817 => x"5575812a",
  2818 => x"81065372",
  2819 => x"802e8538",
  2820 => x"748c0755",
  2821 => x"75810640",
  2822 => x"7f802e85",
  2823 => x"38748307",
  2824 => x"55740970",
  2825 => x"81ff0652",
  2826 => x"53f6cc3f",
  2827 => x"7714982b",
  2828 => x"70982c55",
  2829 => x"56767424",
  2830 => x"ff9b38fb",
  2831 => x"d4397914",
  2832 => x"70337009",
  2833 => x"7081ff06",
  2834 => x"54585440",
  2835 => x"f6a93f77",
  2836 => x"14982b70",
  2837 => x"982c5559",
  2838 => x"737725fb",
  2839 => x"b4387914",
  2840 => x"70337009",
  2841 => x"7081ff06",
  2842 => x"54585440",
  2843 => x"f6893f77",
  2844 => x"14982b70",
  2845 => x"982c5559",
  2846 => x"767424c2",
  2847 => x"38fb9239",
  2848 => x"61802e81",
  2849 => x"c8387d80",
  2850 => x"2e80f138",
  2851 => x"79147033",
  2852 => x"70585455",
  2853 => x"80557875",
  2854 => x"2e853872",
  2855 => x"842a5675",
  2856 => x"832a8106",
  2857 => x"407f802e",
  2858 => x"843881c0",
  2859 => x"5575822a",
  2860 => x"8106407f",
  2861 => x"802e8538",
  2862 => x"74b00755",
  2863 => x"75812a81",
  2864 => x"06407f80",
  2865 => x"2e853874",
  2866 => x"8c075575",
  2867 => x"81065372",
  2868 => x"802e8538",
  2869 => x"74830755",
  2870 => x"74097081",
  2871 => x"ff067053",
  2872 => x"4156f593",
  2873 => x"3f7f51f5",
  2874 => x"8e3f7714",
  2875 => x"982b7098",
  2876 => x"2c555376",
  2877 => x"7424ff94",
  2878 => x"38fa9639",
  2879 => x"79147033",
  2880 => x"70097081",
  2881 => x"ff067055",
  2882 => x"59554155",
  2883 => x"f4e93f75",
  2884 => x"51f4e43f",
  2885 => x"7714982b",
  2886 => x"70982c55",
  2887 => x"59737725",
  2888 => x"f9ef3879",
  2889 => x"14703370",
  2890 => x"097081ff",
  2891 => x"06705559",
  2892 => x"554155f4",
  2893 => x"c23f7551",
  2894 => x"f4bd3f77",
  2895 => x"14982b70",
  2896 => x"982c5559",
  2897 => x"767424ff",
  2898 => x"b338f9c5",
  2899 => x"397d802e",
  2900 => x"80ee3879",
  2901 => x"14703370",
  2902 => x"58545580",
  2903 => x"5578752e",
  2904 => x"85387284",
  2905 => x"2a567583",
  2906 => x"2a810653",
  2907 => x"72802e84",
  2908 => x"3881c055",
  2909 => x"75822a81",
  2910 => x"06537280",
  2911 => x"2e853874",
  2912 => x"b0075575",
  2913 => x"812a8106",
  2914 => x"5372802e",
  2915 => x"8538748c",
  2916 => x"07557581",
  2917 => x"06407f80",
  2918 => x"2e853874",
  2919 => x"83075574",
  2920 => x"81ff0670",
  2921 => x"5256f3cf",
  2922 => x"3f7551f3",
  2923 => x"ca3f7714",
  2924 => x"982b7098",
  2925 => x"2c555376",
  2926 => x"7424ff97",
  2927 => x"38f8d239",
  2928 => x"79147033",
  2929 => x"70535740",
  2930 => x"f3ad3f75",
  2931 => x"51f3a83f",
  2932 => x"7714982b",
  2933 => x"70982c55",
  2934 => x"59737725",
  2935 => x"f8b33879",
  2936 => x"14703370",
  2937 => x"535740f3",
  2938 => x"8e3f7551",
  2939 => x"f3893f77",
  2940 => x"14982b70",
  2941 => x"982c5559",
  2942 => x"767424c4",
  2943 => x"38f89239",
  2944 => x"7d802e80",
  2945 => x"ec387914",
  2946 => x"70337c07",
  2947 => x"70525456",
  2948 => x"80557875",
  2949 => x"2e853872",
  2950 => x"842a5675",
  2951 => x"832a8106",
  2952 => x"5372802e",
  2953 => x"843881c0",
  2954 => x"5575822a",
  2955 => x"81065372",
  2956 => x"802e8538",
  2957 => x"74b00755",
  2958 => x"75812a81",
  2959 => x"06537280",
  2960 => x"2e853874",
  2961 => x"8c075575",
  2962 => x"8106407f",
  2963 => x"802e8538",
  2964 => x"74830755",
  2965 => x"74097081",
  2966 => x"ff065253",
  2967 => x"f2993f77",
  2968 => x"14982b70",
  2969 => x"982c5556",
  2970 => x"767424ff",
  2971 => x"9938f7a1",
  2972 => x"39791470",
  2973 => x"337c0770",
  2974 => x"097081ff",
  2975 => x"06545541",
  2976 => x"56f1f43f",
  2977 => x"7714982b",
  2978 => x"70982c55",
  2979 => x"59737725",
  2980 => x"f6ff3879",
  2981 => x"1470337c",
  2982 => x"07700970",
  2983 => x"81ff0654",
  2984 => x"554156f1",
  2985 => x"d23f7714",
  2986 => x"982b7098",
  2987 => x"2c555976",
  2988 => x"7424ffbd",
  2989 => x"38f6da39",
  2990 => x"61802e80",
  2991 => x"f9387d80",
  2992 => x"2e81e838",
  2993 => x"79147033",
  2994 => x"7c077052",
  2995 => x"54568055",
  2996 => x"78752e85",
  2997 => x"3872842a",
  2998 => x"5675832a",
  2999 => x"81065372",
  3000 => x"802e8438",
  3001 => x"81c05575",
  3002 => x"822a8106",
  3003 => x"5372802e",
  3004 => x"853874b0",
  3005 => x"07557581",
  3006 => x"2a810653",
  3007 => x"72802e85",
  3008 => x"38748c07",
  3009 => x"55758106",
  3010 => x"407f802e",
  3011 => x"85387483",
  3012 => x"07557409",
  3013 => x"7081ff06",
  3014 => x"70535456",
  3015 => x"f0d93f72",
  3016 => x"51f0d43f",
  3017 => x"7714982b",
  3018 => x"70982c55",
  3019 => x"40767424",
  3020 => x"ff9238f5",
  3021 => x"dc397d80",
  3022 => x"2e81c538",
  3023 => x"79147033",
  3024 => x"7c077052",
  3025 => x"54568055",
  3026 => x"78752e85",
  3027 => x"3872842a",
  3028 => x"5675832a",
  3029 => x"81065372",
  3030 => x"802e8438",
  3031 => x"81c05575",
  3032 => x"822a8106",
  3033 => x"5372802e",
  3034 => x"853874b0",
  3035 => x"07557581",
  3036 => x"2a810653",
  3037 => x"72802e85",
  3038 => x"38748c07",
  3039 => x"55758106",
  3040 => x"407f802e",
  3041 => x"85387483",
  3042 => x"07557481",
  3043 => x"ff067052",
  3044 => x"53efe43f",
  3045 => x"7251efdf",
  3046 => x"3f771498",
  3047 => x"2b70982c",
  3048 => x"55567674",
  3049 => x"24ff9538",
  3050 => x"f4e73979",
  3051 => x"1470337c",
  3052 => x"07700970",
  3053 => x"81ff0670",
  3054 => x"55564256",
  3055 => x"59efb83f",
  3056 => x"7251efb3",
  3057 => x"3f771498",
  3058 => x"2b70982c",
  3059 => x"55597377",
  3060 => x"25f4be38",
  3061 => x"79147033",
  3062 => x"7c077009",
  3063 => x"7081ff06",
  3064 => x"70555642",
  3065 => x"5659ef8f",
  3066 => x"3f7251ef",
  3067 => x"8a3f7714",
  3068 => x"982b7098",
  3069 => x"2c555976",
  3070 => x"7424ffaf",
  3071 => x"38f49239",
  3072 => x"79147033",
  3073 => x"7c077053",
  3074 => x"5455eeeb",
  3075 => x"3f7251ee",
  3076 => x"e63f7714",
  3077 => x"982b7098",
  3078 => x"2c555973",
  3079 => x"7725f3f1",
  3080 => x"38791470",
  3081 => x"337c0770",
  3082 => x"535455ee",
  3083 => x"ca3f7251",
  3084 => x"eec53f77",
  3085 => x"14982b70",
  3086 => x"982c5559",
  3087 => x"767424c0",
  3088 => x"38f3ce39",
  3089 => x"81b1f433",
  3090 => x"7f055680",
  3091 => x"527581ff",
  3092 => x"0651ed9d",
  3093 => x"3f80537c",
  3094 => x"a02ef3f6",
  3095 => x"387f7829",
  3096 => x"64305e57",
  3097 => x"f2a039f8",
  3098 => x"3d0d7a7d",
  3099 => x"028805af",
  3100 => x"05335a55",
  3101 => x"59807470",
  3102 => x"81055633",
  3103 => x"75585657",
  3104 => x"74772e09",
  3105 => x"81068838",
  3106 => x"76b00c8a",
  3107 => x"3d0d0474",
  3108 => x"53775278",
  3109 => x"51efdf3f",
  3110 => x"b00881ff",
  3111 => x"06770570",
  3112 => x"83ffff06",
  3113 => x"77708105",
  3114 => x"59335258",
  3115 => x"5574802e",
  3116 => x"d7387453",
  3117 => x"77527851",
  3118 => x"efbc3fb0",
  3119 => x"0881ff06",
  3120 => x"77057083",
  3121 => x"ffff0677",
  3122 => x"70810559",
  3123 => x"33525855",
  3124 => x"74ffbc38",
  3125 => x"ffb239cd",
  3126 => x"c73f04fb",
  3127 => x"3d0d7779",
  3128 => x"55558056",
  3129 => x"757524ab",
  3130 => x"38807424",
  3131 => x"9d388053",
  3132 => x"73527451",
  3133 => x"80e13fb0",
  3134 => x"08547580",
  3135 => x"2e8538b0",
  3136 => x"08305473",
  3137 => x"b00c873d",
  3138 => x"0d047330",
  3139 => x"76813257",
  3140 => x"54dc3974",
  3141 => x"30558156",
  3142 => x"738025d2",
  3143 => x"38ec39fa",
  3144 => x"3d0d787a",
  3145 => x"57558057",
  3146 => x"767524a4",
  3147 => x"38759f2c",
  3148 => x"54815375",
  3149 => x"74327431",
  3150 => x"5274519b",
  3151 => x"3fb00854",
  3152 => x"76802e85",
  3153 => x"38b00830",
  3154 => x"5473b00c",
  3155 => x"883d0d04",
  3156 => x"74305581",
  3157 => x"57d739fc",
  3158 => x"3d0d7678",
  3159 => x"53548153",
  3160 => x"80747326",
  3161 => x"52557280",
  3162 => x"2e983870",
  3163 => x"802ea938",
  3164 => x"807224a4",
  3165 => x"38711073",
  3166 => x"10757226",
  3167 => x"53545272",
  3168 => x"ea387351",
  3169 => x"78833874",
  3170 => x"5170b00c",
  3171 => x"863d0d04",
  3172 => x"72812a72",
  3173 => x"812a5353",
  3174 => x"72802ee6",
  3175 => x"38717426",
  3176 => x"ef387372",
  3177 => x"31757407",
  3178 => x"74812a74",
  3179 => x"812a5555",
  3180 => x"5654e539",
  3181 => x"10101010",
  3182 => x"10101010",
  3183 => x"10101010",
  3184 => x"10101010",
  3185 => x"10101010",
  3186 => x"10101010",
  3187 => x"10101010",
  3188 => x"10101053",
  3189 => x"51047381",
  3190 => x"ff067383",
  3191 => x"06098105",
  3192 => x"83051010",
  3193 => x"102b0772",
  3194 => x"fc060c51",
  3195 => x"51043c04",
  3196 => x"72728072",
  3197 => x"8106ff05",
  3198 => x"09720605",
  3199 => x"71105272",
  3200 => x"0a100a53",
  3201 => x"72ed3851",
  3202 => x"51535104",
  3203 => x"b008b408",
  3204 => x"b8087575",
  3205 => x"80e29f2d",
  3206 => x"5050b008",
  3207 => x"56b80cb4",
  3208 => x"0cb00c51",
  3209 => x"04b008b4",
  3210 => x"08b80875",
  3211 => x"7580e1db",
  3212 => x"2d5050b0",
  3213 => x"0856b80c",
  3214 => x"b40cb00c",
  3215 => x"5104b008",
  3216 => x"b408b808",
  3217 => x"aef72db8",
  3218 => x"0cb40cb0",
  3219 => x"0c04ff3d",
  3220 => x"0d028f05",
  3221 => x"3381b2ac",
  3222 => x"0852710c",
  3223 => x"800bb00c",
  3224 => x"833d0d04",
  3225 => x"ff3d0d02",
  3226 => x"8f053351",
  3227 => x"81d5f408",
  3228 => x"52712db0",
  3229 => x"0881ff06",
  3230 => x"b00c833d",
  3231 => x"0d04fe3d",
  3232 => x"0d747033",
  3233 => x"53537180",
  3234 => x"2e933881",
  3235 => x"13725281",
  3236 => x"d5f40853",
  3237 => x"53712d72",
  3238 => x"335271ef",
  3239 => x"38843d0d",
  3240 => x"04f43d0d",
  3241 => x"7f028405",
  3242 => x"bb053355",
  3243 => x"57880b8c",
  3244 => x"3d5b5989",
  3245 => x"5381afc4",
  3246 => x"52795186",
  3247 => x"d93f7379",
  3248 => x"2e80ff38",
  3249 => x"78567390",
  3250 => x"2e80ec38",
  3251 => x"02a70558",
  3252 => x"768f0654",
  3253 => x"73892680",
  3254 => x"c2387518",
  3255 => x"b0155555",
  3256 => x"73753476",
  3257 => x"842aff17",
  3258 => x"7081ff06",
  3259 => x"58555775",
  3260 => x"df38781a",
  3261 => x"55757534",
  3262 => x"79703355",
  3263 => x"5573802e",
  3264 => x"93388115",
  3265 => x"745281d5",
  3266 => x"f4085755",
  3267 => x"752d7433",
  3268 => x"5473ef38",
  3269 => x"78b00c8e",
  3270 => x"3d0d0475",
  3271 => x"18b71555",
  3272 => x"55737534",
  3273 => x"76842aff",
  3274 => x"177081ff",
  3275 => x"06585557",
  3276 => x"75ff9d38",
  3277 => x"ffbc3984",
  3278 => x"70575902",
  3279 => x"a70558ff",
  3280 => x"8f398270",
  3281 => x"5759f439",
  3282 => x"f13d0d61",
  3283 => x"8d3d705b",
  3284 => x"5c5a807a",
  3285 => x"5657767a",
  3286 => x"24818538",
  3287 => x"7817548a",
  3288 => x"52745184",
  3289 => x"ff3fb008",
  3290 => x"b0055372",
  3291 => x"74348117",
  3292 => x"578a5274",
  3293 => x"5184c83f",
  3294 => x"b00855b0",
  3295 => x"08de38b0",
  3296 => x"08779f2a",
  3297 => x"1870812c",
  3298 => x"5a565680",
  3299 => x"78259e38",
  3300 => x"7817ff05",
  3301 => x"55751970",
  3302 => x"33555374",
  3303 => x"33733473",
  3304 => x"75348116",
  3305 => x"ff165656",
  3306 => x"777624e9",
  3307 => x"38761958",
  3308 => x"80783480",
  3309 => x"7a241770",
  3310 => x"81ff067c",
  3311 => x"70335657",
  3312 => x"55567280",
  3313 => x"2e933881",
  3314 => x"15735281",
  3315 => x"d5f40858",
  3316 => x"55762d74",
  3317 => x"335372ef",
  3318 => x"3873b00c",
  3319 => x"913d0d04",
  3320 => x"ad7b3402",
  3321 => x"ad057a30",
  3322 => x"71195656",
  3323 => x"598a5274",
  3324 => x"5183f13f",
  3325 => x"b008b005",
  3326 => x"53727434",
  3327 => x"8117578a",
  3328 => x"52745183",
  3329 => x"ba3fb008",
  3330 => x"55b008fe",
  3331 => x"cf38feef",
  3332 => x"39fd3d0d",
  3333 => x"81b2a008",
  3334 => x"76b2e429",
  3335 => x"94120c54",
  3336 => x"850b9815",
  3337 => x"0c981408",
  3338 => x"70810651",
  3339 => x"5372f638",
  3340 => x"853d0d04",
  3341 => x"803d0d81",
  3342 => x"b2a00851",
  3343 => x"870b8412",
  3344 => x"0cff0ba4",
  3345 => x"120ca70b",
  3346 => x"a8120cb2",
  3347 => x"e40b9412",
  3348 => x"0c870b98",
  3349 => x"120c823d",
  3350 => x"0d04803d",
  3351 => x"0d81b2a4",
  3352 => x"0851b80b",
  3353 => x"8c120c83",
  3354 => x"0b88120c",
  3355 => x"823d0d04",
  3356 => x"803d0d81",
  3357 => x"b2a40884",
  3358 => x"11088106",
  3359 => x"b00c5182",
  3360 => x"3d0d04ff",
  3361 => x"3d0d81b2",
  3362 => x"a4085284",
  3363 => x"12087081",
  3364 => x"06515170",
  3365 => x"802ef438",
  3366 => x"71087081",
  3367 => x"ff06b00c",
  3368 => x"51833d0d",
  3369 => x"04fe3d0d",
  3370 => x"02930533",
  3371 => x"81b2a408",
  3372 => x"53538412",
  3373 => x"0870892a",
  3374 => x"70810651",
  3375 => x"515170f2",
  3376 => x"3872720c",
  3377 => x"843d0d04",
  3378 => x"fe3d0d02",
  3379 => x"93053353",
  3380 => x"728a2e9c",
  3381 => x"3881b2a4",
  3382 => x"08528412",
  3383 => x"0870892a",
  3384 => x"70810651",
  3385 => x"515170f2",
  3386 => x"3872720c",
  3387 => x"843d0d04",
  3388 => x"81b2a408",
  3389 => x"52841208",
  3390 => x"70892a70",
  3391 => x"81065151",
  3392 => x"5170f238",
  3393 => x"8d720c84",
  3394 => x"12087089",
  3395 => x"2a708106",
  3396 => x"51515170",
  3397 => x"c538d239",
  3398 => x"803d0d81",
  3399 => x"b2980851",
  3400 => x"800b8412",
  3401 => x"0c83fe80",
  3402 => x"0b88120c",
  3403 => x"800b81d5",
  3404 => x"f834800b",
  3405 => x"81d5fc34",
  3406 => x"823d0d04",
  3407 => x"fa3d0d02",
  3408 => x"a3053381",
  3409 => x"b2980881",
  3410 => x"d5f83370",
  3411 => x"81ff0670",
  3412 => x"10101181",
  3413 => x"d5fc3370",
  3414 => x"81ff0672",
  3415 => x"90291170",
  3416 => x"882b7807",
  3417 => x"770c535b",
  3418 => x"5b555559",
  3419 => x"5454738a",
  3420 => x"2e983874",
  3421 => x"80cf2e92",
  3422 => x"38738c2e",
  3423 => x"a4388116",
  3424 => x"537281d5",
  3425 => x"fc34883d",
  3426 => x"0d0471a3",
  3427 => x"26a33881",
  3428 => x"17527181",
  3429 => x"d5f83480",
  3430 => x"0b81d5fc",
  3431 => x"34883d0d",
  3432 => x"04805271",
  3433 => x"882b730c",
  3434 => x"81125297",
  3435 => x"907226f3",
  3436 => x"38800b81",
  3437 => x"d5f83480",
  3438 => x"0b81d5fc",
  3439 => x"34df39bc",
  3440 => x"0802bc0c",
  3441 => x"fd3d0d80",
  3442 => x"53bc088c",
  3443 => x"050852bc",
  3444 => x"08880508",
  3445 => x"51f7803f",
  3446 => x"b00870b0",
  3447 => x"0c54853d",
  3448 => x"0dbc0c04",
  3449 => x"bc0802bc",
  3450 => x"0cfd3d0d",
  3451 => x"8153bc08",
  3452 => x"8c050852",
  3453 => x"bc088805",
  3454 => x"0851f6db",
  3455 => x"3fb00870",
  3456 => x"b00c5485",
  3457 => x"3d0dbc0c",
  3458 => x"04803d0d",
  3459 => x"86518496",
  3460 => x"3f8151a1",
  3461 => x"d33ffc3d",
  3462 => x"0d767079",
  3463 => x"7b555555",
  3464 => x"558f7227",
  3465 => x"8c387275",
  3466 => x"07830651",
  3467 => x"70802ea7",
  3468 => x"38ff1252",
  3469 => x"71ff2e98",
  3470 => x"38727081",
  3471 => x"05543374",
  3472 => x"70810556",
  3473 => x"34ff1252",
  3474 => x"71ff2e09",
  3475 => x"8106ea38",
  3476 => x"74b00c86",
  3477 => x"3d0d0474",
  3478 => x"51727084",
  3479 => x"05540871",
  3480 => x"70840553",
  3481 => x"0c727084",
  3482 => x"05540871",
  3483 => x"70840553",
  3484 => x"0c727084",
  3485 => x"05540871",
  3486 => x"70840553",
  3487 => x"0c727084",
  3488 => x"05540871",
  3489 => x"70840553",
  3490 => x"0cf01252",
  3491 => x"718f26c9",
  3492 => x"38837227",
  3493 => x"95387270",
  3494 => x"84055408",
  3495 => x"71708405",
  3496 => x"530cfc12",
  3497 => x"52718326",
  3498 => x"ed387054",
  3499 => x"ff8339fd",
  3500 => x"3d0d7553",
  3501 => x"84d81308",
  3502 => x"802e8a38",
  3503 => x"805372b0",
  3504 => x"0c853d0d",
  3505 => x"04818052",
  3506 => x"72518d9b",
  3507 => x"3fb00884",
  3508 => x"d8140cff",
  3509 => x"53b00880",
  3510 => x"2ee438b0",
  3511 => x"08549f53",
  3512 => x"80747084",
  3513 => x"05560cff",
  3514 => x"13538073",
  3515 => x"24ce3880",
  3516 => x"74708405",
  3517 => x"560cff13",
  3518 => x"53728025",
  3519 => x"e338ffbc",
  3520 => x"39fd3d0d",
  3521 => x"75775553",
  3522 => x"9f74278d",
  3523 => x"3896730c",
  3524 => x"ff5271b0",
  3525 => x"0c853d0d",
  3526 => x"0484d813",
  3527 => x"08527180",
  3528 => x"2e933873",
  3529 => x"10101270",
  3530 => x"0879720c",
  3531 => x"515271b0",
  3532 => x"0c853d0d",
  3533 => x"047251fe",
  3534 => x"f63fff52",
  3535 => x"b008d338",
  3536 => x"84d81308",
  3537 => x"74101011",
  3538 => x"70087a72",
  3539 => x"0c515152",
  3540 => x"dd39f93d",
  3541 => x"0d797b58",
  3542 => x"56769f26",
  3543 => x"80e83884",
  3544 => x"d8160854",
  3545 => x"73802eaa",
  3546 => x"38761010",
  3547 => x"14700855",
  3548 => x"5573802e",
  3549 => x"ba388058",
  3550 => x"73812e8f",
  3551 => x"3873ff2e",
  3552 => x"a3388075",
  3553 => x"0c765173",
  3554 => x"2d805877",
  3555 => x"b00c893d",
  3556 => x"0d047551",
  3557 => x"fe993fff",
  3558 => x"58b008ef",
  3559 => x"3884d816",
  3560 => x"0854c639",
  3561 => x"96760c81",
  3562 => x"0bb00c89",
  3563 => x"3d0d0475",
  3564 => x"5181ed3f",
  3565 => x"7653b008",
  3566 => x"52755181",
  3567 => x"ad3fb008",
  3568 => x"b00c893d",
  3569 => x"0d049676",
  3570 => x"0cff0bb0",
  3571 => x"0c893d0d",
  3572 => x"04fc3d0d",
  3573 => x"76785653",
  3574 => x"ff54749f",
  3575 => x"26b13884",
  3576 => x"d8130852",
  3577 => x"71802eae",
  3578 => x"38741010",
  3579 => x"12700853",
  3580 => x"53815471",
  3581 => x"802e9838",
  3582 => x"825471ff",
  3583 => x"2e913883",
  3584 => x"5471812e",
  3585 => x"8a388073",
  3586 => x"0c745171",
  3587 => x"2d805473",
  3588 => x"b00c863d",
  3589 => x"0d047251",
  3590 => x"fd953fb0",
  3591 => x"08f13884",
  3592 => x"d8130852",
  3593 => x"c439ff3d",
  3594 => x"0d735281",
  3595 => x"b2b00851",
  3596 => x"fea03f83",
  3597 => x"3d0d04fe",
  3598 => x"3d0d7553",
  3599 => x"745281b2",
  3600 => x"b00851fd",
  3601 => x"bc3f843d",
  3602 => x"0d04803d",
  3603 => x"0d81b2b0",
  3604 => x"0851fcdb",
  3605 => x"3f823d0d",
  3606 => x"04ff3d0d",
  3607 => x"735281b2",
  3608 => x"b00851fe",
  3609 => x"ec3f833d",
  3610 => x"0d04fc3d",
  3611 => x"0d800b81",
  3612 => x"d6840c78",
  3613 => x"5277519c",
  3614 => x"aa3fb008",
  3615 => x"54b008ff",
  3616 => x"2e883873",
  3617 => x"b00c863d",
  3618 => x"0d0481d6",
  3619 => x"84085574",
  3620 => x"802ef038",
  3621 => x"7675710c",
  3622 => x"5373b00c",
  3623 => x"863d0d04",
  3624 => x"9bfc3f04",
  3625 => x"fc3d0d76",
  3626 => x"70797073",
  3627 => x"07830654",
  3628 => x"54545570",
  3629 => x"80c33871",
  3630 => x"70087009",
  3631 => x"70f7fbfd",
  3632 => x"ff130670",
  3633 => x"f8848281",
  3634 => x"80065151",
  3635 => x"53535470",
  3636 => x"a6388414",
  3637 => x"72747084",
  3638 => x"05560c70",
  3639 => x"08700970",
  3640 => x"f7fbfdff",
  3641 => x"130670f8",
  3642 => x"84828180",
  3643 => x"06515153",
  3644 => x"53547080",
  3645 => x"2edc3873",
  3646 => x"52717081",
  3647 => x"05533351",
  3648 => x"70737081",
  3649 => x"05553470",
  3650 => x"f03874b0",
  3651 => x"0c863d0d",
  3652 => x"04fd3d0d",
  3653 => x"75707183",
  3654 => x"06535552",
  3655 => x"70b83871",
  3656 => x"70087009",
  3657 => x"f7fbfdff",
  3658 => x"120670f8",
  3659 => x"84828180",
  3660 => x"06515152",
  3661 => x"53709d38",
  3662 => x"84137008",
  3663 => x"7009f7fb",
  3664 => x"fdff1206",
  3665 => x"70f88482",
  3666 => x"81800651",
  3667 => x"51525370",
  3668 => x"802ee538",
  3669 => x"72527133",
  3670 => x"5170802e",
  3671 => x"8a388112",
  3672 => x"70335252",
  3673 => x"70f83871",
  3674 => x"7431b00c",
  3675 => x"853d0d04",
  3676 => x"fa3d0d78",
  3677 => x"7a7c7054",
  3678 => x"55555272",
  3679 => x"802e80d9",
  3680 => x"38717407",
  3681 => x"83065170",
  3682 => x"802e80d4",
  3683 => x"38ff1353",
  3684 => x"72ff2eb1",
  3685 => x"38713374",
  3686 => x"33565174",
  3687 => x"712e0981",
  3688 => x"06a93872",
  3689 => x"802e8187",
  3690 => x"387081ff",
  3691 => x"06517080",
  3692 => x"2e80fc38",
  3693 => x"81128115",
  3694 => x"ff155555",
  3695 => x"5272ff2e",
  3696 => x"098106d1",
  3697 => x"38713374",
  3698 => x"33565170",
  3699 => x"81ff0675",
  3700 => x"81ff0671",
  3701 => x"71315152",
  3702 => x"5270b00c",
  3703 => x"883d0d04",
  3704 => x"71745755",
  3705 => x"83732788",
  3706 => x"38710874",
  3707 => x"082e8838",
  3708 => x"74765552",
  3709 => x"ff9739fc",
  3710 => x"13537280",
  3711 => x"2eb13874",
  3712 => x"087009f7",
  3713 => x"fbfdff12",
  3714 => x"0670f884",
  3715 => x"82818006",
  3716 => x"51515170",
  3717 => x"9a388415",
  3718 => x"84175755",
  3719 => x"837327d0",
  3720 => x"38740876",
  3721 => x"082ed038",
  3722 => x"74765552",
  3723 => x"fedf3980",
  3724 => x"0bb00c88",
  3725 => x"3d0d04f3",
  3726 => x"3d0d6062",
  3727 => x"64725a5a",
  3728 => x"5e5e805c",
  3729 => x"76708105",
  3730 => x"583381af",
  3731 => x"d1113370",
  3732 => x"832a7081",
  3733 => x"06515555",
  3734 => x"5672e938",
  3735 => x"75ad2e82",
  3736 => x"883875ab",
  3737 => x"2e828438",
  3738 => x"77307079",
  3739 => x"07802579",
  3740 => x"90327030",
  3741 => x"70720780",
  3742 => x"25730753",
  3743 => x"57575153",
  3744 => x"72802e87",
  3745 => x"3875b02e",
  3746 => x"81eb3877",
  3747 => x"8a388858",
  3748 => x"75b02e83",
  3749 => x"388a5881",
  3750 => x"0a5a7b84",
  3751 => x"38fe0a5a",
  3752 => x"77527951",
  3753 => x"f6be3fb0",
  3754 => x"0878537a",
  3755 => x"525bf68f",
  3756 => x"3fb0085a",
  3757 => x"807081af",
  3758 => x"d1183370",
  3759 => x"822a7081",
  3760 => x"06515656",
  3761 => x"5a557280",
  3762 => x"2e80c138",
  3763 => x"d0165675",
  3764 => x"782580d7",
  3765 => x"38807924",
  3766 => x"757b2607",
  3767 => x"53729338",
  3768 => x"747a2e80",
  3769 => x"eb387a76",
  3770 => x"2580ed38",
  3771 => x"72802e80",
  3772 => x"e738ff77",
  3773 => x"70810559",
  3774 => x"33575981",
  3775 => x"afd11633",
  3776 => x"70822a70",
  3777 => x"81065154",
  3778 => x"5472c138",
  3779 => x"73830653",
  3780 => x"72802e97",
  3781 => x"38738106",
  3782 => x"c9175553",
  3783 => x"728538ff",
  3784 => x"a9165473",
  3785 => x"56777624",
  3786 => x"ffab3880",
  3787 => x"792480f0",
  3788 => x"387b802e",
  3789 => x"84387430",
  3790 => x"557c802e",
  3791 => x"8c38ff17",
  3792 => x"53788338",
  3793 => x"7d53727d",
  3794 => x"0c74b00c",
  3795 => x"8f3d0d04",
  3796 => x"8153757b",
  3797 => x"24ff9538",
  3798 => x"81757929",
  3799 => x"17787081",
  3800 => x"055a3358",
  3801 => x"5659ff93",
  3802 => x"39815c76",
  3803 => x"70810558",
  3804 => x"3356fdf4",
  3805 => x"39807733",
  3806 => x"54547280",
  3807 => x"f82eb238",
  3808 => x"7280d832",
  3809 => x"70307080",
  3810 => x"25760751",
  3811 => x"51537280",
  3812 => x"2efdf838",
  3813 => x"81173382",
  3814 => x"18585690",
  3815 => x"58fdf839",
  3816 => x"810a557b",
  3817 => x"8438fe0a",
  3818 => x"557f53a2",
  3819 => x"730cff89",
  3820 => x"398154cc",
  3821 => x"39fd3d0d",
  3822 => x"77547653",
  3823 => x"755281b2",
  3824 => x"b00851fc",
  3825 => x"f23f853d",
  3826 => x"0d04f33d",
  3827 => x"0d606264",
  3828 => x"725a5a5d",
  3829 => x"5d805e76",
  3830 => x"70810558",
  3831 => x"3381afd1",
  3832 => x"11337083",
  3833 => x"2a708106",
  3834 => x"51555556",
  3835 => x"72e93875",
  3836 => x"ad2e81ff",
  3837 => x"3875ab2e",
  3838 => x"81fb3877",
  3839 => x"30707907",
  3840 => x"80257990",
  3841 => x"32703070",
  3842 => x"72078025",
  3843 => x"73075357",
  3844 => x"57515372",
  3845 => x"802e8738",
  3846 => x"75b02e81",
  3847 => x"e238778a",
  3848 => x"38885875",
  3849 => x"b02e8338",
  3850 => x"8a587752",
  3851 => x"ff51f38f",
  3852 => x"3fb00878",
  3853 => x"535aff51",
  3854 => x"f3aa3fb0",
  3855 => x"085b8070",
  3856 => x"5a5581af",
  3857 => x"d1163370",
  3858 => x"822a7081",
  3859 => x"06515454",
  3860 => x"72802e80",
  3861 => x"c138d016",
  3862 => x"56757825",
  3863 => x"80d73880",
  3864 => x"7924757b",
  3865 => x"26075372",
  3866 => x"9338747a",
  3867 => x"2e80eb38",
  3868 => x"7a762580",
  3869 => x"ed387280",
  3870 => x"2e80e738",
  3871 => x"ff777081",
  3872 => x"05593357",
  3873 => x"5981afd1",
  3874 => x"16337082",
  3875 => x"2a708106",
  3876 => x"51545472",
  3877 => x"c1387383",
  3878 => x"06537280",
  3879 => x"2e973873",
  3880 => x"8106c917",
  3881 => x"55537285",
  3882 => x"38ffa916",
  3883 => x"54735677",
  3884 => x"7624ffab",
  3885 => x"38807924",
  3886 => x"8189387d",
  3887 => x"802e8438",
  3888 => x"7430557b",
  3889 => x"802e8c38",
  3890 => x"ff175378",
  3891 => x"83387c53",
  3892 => x"727c0c74",
  3893 => x"b00c8f3d",
  3894 => x"0d048153",
  3895 => x"757b24ff",
  3896 => x"95388175",
  3897 => x"79291778",
  3898 => x"7081055a",
  3899 => x"33585659",
  3900 => x"ff933981",
  3901 => x"5e767081",
  3902 => x"05583356",
  3903 => x"fdfd3980",
  3904 => x"77335454",
  3905 => x"7280f82e",
  3906 => x"80c33872",
  3907 => x"80d83270",
  3908 => x"30708025",
  3909 => x"76075151",
  3910 => x"5372802e",
  3911 => x"fe803881",
  3912 => x"17338218",
  3913 => x"58569070",
  3914 => x"5358ff51",
  3915 => x"f1913fb0",
  3916 => x"0878535a",
  3917 => x"ff51f1ac",
  3918 => x"3fb0085b",
  3919 => x"80705a55",
  3920 => x"fe8039ff",
  3921 => x"605455a2",
  3922 => x"730cfef7",
  3923 => x"398154ff",
  3924 => x"ba39fd3d",
  3925 => x"0d775476",
  3926 => x"53755281",
  3927 => x"b2b00851",
  3928 => x"fce83f85",
  3929 => x"3d0d04f3",
  3930 => x"3d0d7f61",
  3931 => x"8b1170f8",
  3932 => x"065c5555",
  3933 => x"5e729626",
  3934 => x"83389059",
  3935 => x"80792474",
  3936 => x"7a260753",
  3937 => x"80547274",
  3938 => x"2e098106",
  3939 => x"80cb387d",
  3940 => x"518bca3f",
  3941 => x"7883f726",
  3942 => x"80c63878",
  3943 => x"832a7010",
  3944 => x"101081b9",
  3945 => x"ec058c11",
  3946 => x"0859595a",
  3947 => x"76782e83",
  3948 => x"b0388417",
  3949 => x"08fc0656",
  3950 => x"8c170888",
  3951 => x"1808718c",
  3952 => x"120c8812",
  3953 => x"0c587517",
  3954 => x"84110881",
  3955 => x"0784120c",
  3956 => x"537d518b",
  3957 => x"893f8817",
  3958 => x"5473b00c",
  3959 => x"8f3d0d04",
  3960 => x"78892a79",
  3961 => x"832a5b53",
  3962 => x"72802ebf",
  3963 => x"3878862a",
  3964 => x"b8055a84",
  3965 => x"7327b438",
  3966 => x"80db135a",
  3967 => x"947327ab",
  3968 => x"38788c2a",
  3969 => x"80ee055a",
  3970 => x"80d47327",
  3971 => x"9e38788f",
  3972 => x"2a80f705",
  3973 => x"5a82d473",
  3974 => x"27913878",
  3975 => x"922a80fc",
  3976 => x"055a8ad4",
  3977 => x"73278438",
  3978 => x"80fe5a79",
  3979 => x"10101081",
  3980 => x"b9ec058c",
  3981 => x"11085855",
  3982 => x"76752ea3",
  3983 => x"38841708",
  3984 => x"fc06707a",
  3985 => x"31555673",
  3986 => x"8f2488d5",
  3987 => x"38738025",
  3988 => x"fee6388c",
  3989 => x"17085776",
  3990 => x"752e0981",
  3991 => x"06df3881",
  3992 => x"1a5a81b9",
  3993 => x"fc085776",
  3994 => x"81b9f42e",
  3995 => x"82c03884",
  3996 => x"1708fc06",
  3997 => x"707a3155",
  3998 => x"56738f24",
  3999 => x"81f93881",
  4000 => x"b9f40b81",
  4001 => x"ba800c81",
  4002 => x"b9f40b81",
  4003 => x"b9fc0c73",
  4004 => x"8025feb2",
  4005 => x"3883ff76",
  4006 => x"2783df38",
  4007 => x"75892a76",
  4008 => x"832a5553",
  4009 => x"72802ebf",
  4010 => x"3875862a",
  4011 => x"b8055484",
  4012 => x"7327b438",
  4013 => x"80db1354",
  4014 => x"947327ab",
  4015 => x"38758c2a",
  4016 => x"80ee0554",
  4017 => x"80d47327",
  4018 => x"9e38758f",
  4019 => x"2a80f705",
  4020 => x"5482d473",
  4021 => x"27913875",
  4022 => x"922a80fc",
  4023 => x"05548ad4",
  4024 => x"73278438",
  4025 => x"80fe5473",
  4026 => x"10101081",
  4027 => x"b9ec0588",
  4028 => x"11085658",
  4029 => x"74782e86",
  4030 => x"cf388415",
  4031 => x"08fc0653",
  4032 => x"7573278d",
  4033 => x"38881508",
  4034 => x"5574782e",
  4035 => x"098106ea",
  4036 => x"388c1508",
  4037 => x"81b9ec0b",
  4038 => x"84050871",
  4039 => x"8c1a0c76",
  4040 => x"881a0c78",
  4041 => x"88130c78",
  4042 => x"8c180c5d",
  4043 => x"58795380",
  4044 => x"7a2483e6",
  4045 => x"3872822c",
  4046 => x"81712b5c",
  4047 => x"537a7c26",
  4048 => x"8198387b",
  4049 => x"7b065372",
  4050 => x"82f13879",
  4051 => x"fc068405",
  4052 => x"5a7a1070",
  4053 => x"7d06545b",
  4054 => x"7282e038",
  4055 => x"841a5af1",
  4056 => x"3988178c",
  4057 => x"11085858",
  4058 => x"76782e09",
  4059 => x"8106fcc2",
  4060 => x"38821a5a",
  4061 => x"fdec3978",
  4062 => x"17798107",
  4063 => x"84190c70",
  4064 => x"81ba800c",
  4065 => x"7081b9fc",
  4066 => x"0c81b9f4",
  4067 => x"0b8c120c",
  4068 => x"8c110888",
  4069 => x"120c7481",
  4070 => x"0784120c",
  4071 => x"74117571",
  4072 => x"0c51537d",
  4073 => x"5187b73f",
  4074 => x"881754fc",
  4075 => x"ac3981b9",
  4076 => x"ec0b8405",
  4077 => x"087a545c",
  4078 => x"798025fe",
  4079 => x"f83882da",
  4080 => x"397a097c",
  4081 => x"067081b9",
  4082 => x"ec0b8405",
  4083 => x"0c5c7a10",
  4084 => x"5b7a7c26",
  4085 => x"85387a85",
  4086 => x"b83881b9",
  4087 => x"ec0b8805",
  4088 => x"08708412",
  4089 => x"08fc0670",
  4090 => x"7c317c72",
  4091 => x"268f7225",
  4092 => x"0757575c",
  4093 => x"5d557280",
  4094 => x"2e80db38",
  4095 => x"797a1681",
  4096 => x"b9e4081b",
  4097 => x"90115a55",
  4098 => x"575b81b9",
  4099 => x"e008ff2e",
  4100 => x"8838a08f",
  4101 => x"13e08006",
  4102 => x"5776527d",
  4103 => x"5186c03f",
  4104 => x"b00854b0",
  4105 => x"08ff2e90",
  4106 => x"38b00876",
  4107 => x"27829938",
  4108 => x"7481b9ec",
  4109 => x"2e829138",
  4110 => x"81b9ec0b",
  4111 => x"88050855",
  4112 => x"841508fc",
  4113 => x"06707a31",
  4114 => x"7a72268f",
  4115 => x"72250752",
  4116 => x"55537283",
  4117 => x"e6387479",
  4118 => x"81078417",
  4119 => x"0c791670",
  4120 => x"81b9ec0b",
  4121 => x"88050c75",
  4122 => x"81078412",
  4123 => x"0c547e52",
  4124 => x"5785eb3f",
  4125 => x"881754fa",
  4126 => x"e0397583",
  4127 => x"2a705454",
  4128 => x"80742481",
  4129 => x"9b387282",
  4130 => x"2c81712b",
  4131 => x"81b9f008",
  4132 => x"077081b9",
  4133 => x"ec0b8405",
  4134 => x"0c751010",
  4135 => x"1081b9ec",
  4136 => x"05881108",
  4137 => x"585a5d53",
  4138 => x"778c180c",
  4139 => x"7488180c",
  4140 => x"7688190c",
  4141 => x"768c160c",
  4142 => x"fcf33979",
  4143 => x"7a101010",
  4144 => x"81b9ec05",
  4145 => x"7057595d",
  4146 => x"8c150857",
  4147 => x"76752ea3",
  4148 => x"38841708",
  4149 => x"fc06707a",
  4150 => x"31555673",
  4151 => x"8f2483ca",
  4152 => x"38738025",
  4153 => x"8481388c",
  4154 => x"17085776",
  4155 => x"752e0981",
  4156 => x"06df3888",
  4157 => x"15811b70",
  4158 => x"8306555b",
  4159 => x"5572c938",
  4160 => x"7c830653",
  4161 => x"72802efd",
  4162 => x"b838ff1d",
  4163 => x"f819595d",
  4164 => x"88180878",
  4165 => x"2eea38fd",
  4166 => x"b539831a",
  4167 => x"53fc9639",
  4168 => x"83147082",
  4169 => x"2c81712b",
  4170 => x"81b9f008",
  4171 => x"077081b9",
  4172 => x"ec0b8405",
  4173 => x"0c761010",
  4174 => x"1081b9ec",
  4175 => x"05881108",
  4176 => x"595b5e51",
  4177 => x"53fee139",
  4178 => x"81b9b008",
  4179 => x"1758b008",
  4180 => x"762e818d",
  4181 => x"3881b9e0",
  4182 => x"08ff2e83",
  4183 => x"ec387376",
  4184 => x"311881b9",
  4185 => x"b00c7387",
  4186 => x"06705753",
  4187 => x"72802e88",
  4188 => x"38887331",
  4189 => x"70155556",
  4190 => x"76149fff",
  4191 => x"06a08071",
  4192 => x"31177054",
  4193 => x"7f535753",
  4194 => x"83d53fb0",
  4195 => x"0853b008",
  4196 => x"ff2e81a0",
  4197 => x"3881b9b0",
  4198 => x"08167081",
  4199 => x"b9b00c74",
  4200 => x"7581b9ec",
  4201 => x"0b88050c",
  4202 => x"74763118",
  4203 => x"70810751",
  4204 => x"5556587b",
  4205 => x"81b9ec2e",
  4206 => x"839c3879",
  4207 => x"8f2682cb",
  4208 => x"38810b84",
  4209 => x"150c8415",
  4210 => x"08fc0670",
  4211 => x"7a317a72",
  4212 => x"268f7225",
  4213 => x"07525553",
  4214 => x"72802efc",
  4215 => x"f93880db",
  4216 => x"39b0089f",
  4217 => x"ff065372",
  4218 => x"feeb3877",
  4219 => x"81b9b00c",
  4220 => x"81b9ec0b",
  4221 => x"8805087b",
  4222 => x"18810784",
  4223 => x"120c5581",
  4224 => x"b9dc0878",
  4225 => x"27863877",
  4226 => x"81b9dc0c",
  4227 => x"81b9d808",
  4228 => x"7827fcac",
  4229 => x"387781b9",
  4230 => x"d80c8415",
  4231 => x"08fc0670",
  4232 => x"7a317a72",
  4233 => x"268f7225",
  4234 => x"07525553",
  4235 => x"72802efc",
  4236 => x"a5388839",
  4237 => x"80745456",
  4238 => x"fedb397d",
  4239 => x"51829f3f",
  4240 => x"800bb00c",
  4241 => x"8f3d0d04",
  4242 => x"73538074",
  4243 => x"24a93872",
  4244 => x"822c8171",
  4245 => x"2b81b9f0",
  4246 => x"08077081",
  4247 => x"b9ec0b84",
  4248 => x"050c5d53",
  4249 => x"778c180c",
  4250 => x"7488180c",
  4251 => x"7688190c",
  4252 => x"768c160c",
  4253 => x"f9b73983",
  4254 => x"1470822c",
  4255 => x"81712b81",
  4256 => x"b9f00807",
  4257 => x"7081b9ec",
  4258 => x"0b84050c",
  4259 => x"5e5153d4",
  4260 => x"397b7b06",
  4261 => x"5372fca3",
  4262 => x"38841a7b",
  4263 => x"105c5af1",
  4264 => x"39ff1a81",
  4265 => x"11515af7",
  4266 => x"b9397817",
  4267 => x"79810784",
  4268 => x"190c8c18",
  4269 => x"08881908",
  4270 => x"718c120c",
  4271 => x"88120c59",
  4272 => x"7081ba80",
  4273 => x"0c7081b9",
  4274 => x"fc0c81b9",
  4275 => x"f40b8c12",
  4276 => x"0c8c1108",
  4277 => x"88120c74",
  4278 => x"81078412",
  4279 => x"0c741175",
  4280 => x"710c5153",
  4281 => x"f9bd3975",
  4282 => x"17841108",
  4283 => x"81078412",
  4284 => x"0c538c17",
  4285 => x"08881808",
  4286 => x"718c120c",
  4287 => x"88120c58",
  4288 => x"7d5180da",
  4289 => x"3f881754",
  4290 => x"f5cf3972",
  4291 => x"84150cf4",
  4292 => x"1af80670",
  4293 => x"841e0881",
  4294 => x"0607841e",
  4295 => x"0c701d54",
  4296 => x"5b850b84",
  4297 => x"140c850b",
  4298 => x"88140c8f",
  4299 => x"7b27fdcf",
  4300 => x"38881c52",
  4301 => x"7d518290",
  4302 => x"3f81b9ec",
  4303 => x"0b880508",
  4304 => x"81b9b008",
  4305 => x"5955fdb7",
  4306 => x"397781b9",
  4307 => x"b00c7381",
  4308 => x"b9e00cfc",
  4309 => x"91397284",
  4310 => x"150cfda3",
  4311 => x"390404fd",
  4312 => x"3d0d800b",
  4313 => x"81d6840c",
  4314 => x"765186cb",
  4315 => x"3fb00853",
  4316 => x"b008ff2e",
  4317 => x"883872b0",
  4318 => x"0c853d0d",
  4319 => x"0481d684",
  4320 => x"08547380",
  4321 => x"2ef03875",
  4322 => x"74710c52",
  4323 => x"72b00c85",
  4324 => x"3d0d04fb",
  4325 => x"3d0d7770",
  4326 => x"5256c23f",
  4327 => x"81b9ec0b",
  4328 => x"88050884",
  4329 => x"1108fc06",
  4330 => x"707b319f",
  4331 => x"ef05e080",
  4332 => x"06e08005",
  4333 => x"565653a0",
  4334 => x"80742494",
  4335 => x"38805275",
  4336 => x"51ff9c3f",
  4337 => x"81b9f408",
  4338 => x"155372b0",
  4339 => x"082e8f38",
  4340 => x"7551ff8a",
  4341 => x"3f805372",
  4342 => x"b00c873d",
  4343 => x"0d047330",
  4344 => x"527551fe",
  4345 => x"fa3fb008",
  4346 => x"ff2ea838",
  4347 => x"81b9ec0b",
  4348 => x"88050875",
  4349 => x"75318107",
  4350 => x"84120c53",
  4351 => x"81b9b008",
  4352 => x"743181b9",
  4353 => x"b00c7551",
  4354 => x"fed43f81",
  4355 => x"0bb00c87",
  4356 => x"3d0d0480",
  4357 => x"527551fe",
  4358 => x"c63f81b9",
  4359 => x"ec0b8805",
  4360 => x"08b00871",
  4361 => x"3156538f",
  4362 => x"7525ffa4",
  4363 => x"38b00881",
  4364 => x"b9e00831",
  4365 => x"81b9b00c",
  4366 => x"74810784",
  4367 => x"140c7551",
  4368 => x"fe9c3f80",
  4369 => x"53ff9039",
  4370 => x"f63d0d7c",
  4371 => x"7e545b72",
  4372 => x"802e8283",
  4373 => x"387a51fe",
  4374 => x"843ff813",
  4375 => x"84110870",
  4376 => x"fe067013",
  4377 => x"841108fc",
  4378 => x"065d5859",
  4379 => x"545881b9",
  4380 => x"f408752e",
  4381 => x"82de3878",
  4382 => x"84160c80",
  4383 => x"73810654",
  4384 => x"5a727a2e",
  4385 => x"81d53878",
  4386 => x"15841108",
  4387 => x"81065153",
  4388 => x"72a03878",
  4389 => x"17577981",
  4390 => x"e6388815",
  4391 => x"08537281",
  4392 => x"b9f42e82",
  4393 => x"f9388c15",
  4394 => x"08708c15",
  4395 => x"0c738812",
  4396 => x"0c567681",
  4397 => x"0784190c",
  4398 => x"76187771",
  4399 => x"0c537981",
  4400 => x"913883ff",
  4401 => x"772781c8",
  4402 => x"3876892a",
  4403 => x"77832a56",
  4404 => x"5372802e",
  4405 => x"bf387686",
  4406 => x"2ab80555",
  4407 => x"847327b4",
  4408 => x"3880db13",
  4409 => x"55947327",
  4410 => x"ab38768c",
  4411 => x"2a80ee05",
  4412 => x"5580d473",
  4413 => x"279e3876",
  4414 => x"8f2a80f7",
  4415 => x"055582d4",
  4416 => x"73279138",
  4417 => x"76922a80",
  4418 => x"fc05558a",
  4419 => x"d4732784",
  4420 => x"3880fe55",
  4421 => x"74101010",
  4422 => x"81b9ec05",
  4423 => x"88110855",
  4424 => x"5673762e",
  4425 => x"82b33884",
  4426 => x"1408fc06",
  4427 => x"53767327",
  4428 => x"8d388814",
  4429 => x"08547376",
  4430 => x"2e098106",
  4431 => x"ea388c14",
  4432 => x"08708c1a",
  4433 => x"0c74881a",
  4434 => x"0c788812",
  4435 => x"0c56778c",
  4436 => x"150c7a51",
  4437 => x"fc883f8c",
  4438 => x"3d0d0477",
  4439 => x"08787131",
  4440 => x"59770588",
  4441 => x"19085457",
  4442 => x"7281b9f4",
  4443 => x"2e80e038",
  4444 => x"8c180870",
  4445 => x"8c150c73",
  4446 => x"88120c56",
  4447 => x"fe893988",
  4448 => x"15088c16",
  4449 => x"08708c13",
  4450 => x"0c578817",
  4451 => x"0cfea339",
  4452 => x"76832a70",
  4453 => x"54558075",
  4454 => x"24819838",
  4455 => x"72822c81",
  4456 => x"712b81b9",
  4457 => x"f0080781",
  4458 => x"b9ec0b84",
  4459 => x"050c5374",
  4460 => x"10101081",
  4461 => x"b9ec0588",
  4462 => x"11085556",
  4463 => x"758c190c",
  4464 => x"7388190c",
  4465 => x"7788170c",
  4466 => x"778c150c",
  4467 => x"ff843981",
  4468 => x"5afdb439",
  4469 => x"78177381",
  4470 => x"06545772",
  4471 => x"98387708",
  4472 => x"78713159",
  4473 => x"77058c19",
  4474 => x"08881a08",
  4475 => x"718c120c",
  4476 => x"88120c57",
  4477 => x"57768107",
  4478 => x"84190c77",
  4479 => x"81b9ec0b",
  4480 => x"88050c81",
  4481 => x"b9e80877",
  4482 => x"26fec738",
  4483 => x"81b9e408",
  4484 => x"527a51fa",
  4485 => x"fe3f7a51",
  4486 => x"fac43ffe",
  4487 => x"ba398178",
  4488 => x"8c150c78",
  4489 => x"88150c73",
  4490 => x"8c1a0c73",
  4491 => x"881a0c5a",
  4492 => x"fd803983",
  4493 => x"1570822c",
  4494 => x"81712b81",
  4495 => x"b9f00807",
  4496 => x"81b9ec0b",
  4497 => x"84050c51",
  4498 => x"53741010",
  4499 => x"1081b9ec",
  4500 => x"05881108",
  4501 => x"5556fee4",
  4502 => x"39745380",
  4503 => x"7524a738",
  4504 => x"72822c81",
  4505 => x"712b81b9",
  4506 => x"f0080781",
  4507 => x"b9ec0b84",
  4508 => x"050c5375",
  4509 => x"8c190c73",
  4510 => x"88190c77",
  4511 => x"88170c77",
  4512 => x"8c150cfd",
  4513 => x"cd398315",
  4514 => x"70822c81",
  4515 => x"712b81b9",
  4516 => x"f0080781",
  4517 => x"b9ec0b84",
  4518 => x"050c5153",
  4519 => x"d639810b",
  4520 => x"b00c0480",
  4521 => x"3d0d7281",
  4522 => x"2e893880",
  4523 => x"0bb00c82",
  4524 => x"3d0d0473",
  4525 => x"51b23ffe",
  4526 => x"3d0d81d6",
  4527 => x"80085170",
  4528 => x"8a3881d6",
  4529 => x"887081d6",
  4530 => x"800c5170",
  4531 => x"75125252",
  4532 => x"ff537087",
  4533 => x"fb808026",
  4534 => x"88387081",
  4535 => x"d6800c71",
  4536 => x"5372b00c",
  4537 => x"843d0d04",
  4538 => x"00ff3900",
  4539 => x"00000000",
  4540 => x"00000000",
  4541 => x"00000000",
  4542 => x"00000000",
  4543 => x"00cac5ca",
  4544 => x"c5c0c0c0",
  4545 => x"c0c0c0c0",
  4546 => x"c0c0c0cf",
  4547 => x"cfcfcf00",
  4548 => x"00000f0f",
  4549 => x"0f0f8f8f",
  4550 => x"cfcfcfcf",
  4551 => x"cfcf4f0f",
  4552 => x"0f0f0000",
  4553 => x"cfcfcfcf",
  4554 => x"0f0f0f0f",
  4555 => x"0f0f0f0f",
  4556 => x"0f0ffefe",
  4557 => x"fefc0000",
  4558 => x"cfcfcfcf",
  4559 => x"cfcfcfcf",
  4560 => x"cfcfcfcf",
  4561 => x"cfffff7e",
  4562 => x"7e000000",
  4563 => x"00000000",
  4564 => x"00000000",
  4565 => x"00000000",
  4566 => x"00003f3f",
  4567 => x"3f3f0101",
  4568 => x"01010101",
  4569 => x"01010101",
  4570 => x"3f3f3f3f",
  4571 => x"0000383c",
  4572 => x"3e3e3f3f",
  4573 => x"3f3b3b39",
  4574 => x"39383838",
  4575 => x"38383800",
  4576 => x"003f3f3f",
  4577 => x"3f383838",
  4578 => x"38383838",
  4579 => x"38383c3f",
  4580 => x"3f1f0f00",
  4581 => x"003f3f3f",
  4582 => x"3f030303",
  4583 => x"03030303",
  4584 => x"03033f3f",
  4585 => x"3f3e0000",
  4586 => x"00000000",
  4587 => x"00000000",
  4588 => x"00000000",
  4589 => x"00000000",
  4590 => x"00000000",
  4591 => x"00000000",
  4592 => x"00000000",
  4593 => x"00000000",
  4594 => x"00000000",
  4595 => x"00000000",
  4596 => x"00000000",
  4597 => x"00000000",
  4598 => x"00000000",
  4599 => x"00000000",
  4600 => x"00000000",
  4601 => x"00000000",
  4602 => x"00000000",
  4603 => x"00000000",
  4604 => x"00000000",
  4605 => x"00000000",
  4606 => x"00000000",
  4607 => x"00000000",
  4608 => x"00000000",
  4609 => x"00000000",
  4610 => x"8080c0c0",
  4611 => x"e0e06000",
  4612 => x"00000000",
  4613 => x"00000000",
  4614 => x"00000000",
  4615 => x"00000000",
  4616 => x"00000000",
  4617 => x"00000000",
  4618 => x"00000000",
  4619 => x"00000000",
  4620 => x"00000000",
  4621 => x"00000000",
  4622 => x"00000000",
  4623 => x"00000000",
  4624 => x"00000000",
  4625 => x"00000000",
  4626 => x"00000000",
  4627 => x"00000000",
  4628 => x"00000000",
  4629 => x"00000000",
  4630 => x"00000000",
  4631 => x"00000000",
  4632 => x"806098ee",
  4633 => x"77bbddec",
  4634 => x"ee6e0200",
  4635 => x"00000000",
  4636 => x"00e08080",
  4637 => x"e00000e0",
  4638 => x"a0a00000",
  4639 => x"e0000000",
  4640 => x"00e0c000",
  4641 => x"c0e00000",
  4642 => x"e08080e0",
  4643 => x"0000c020",
  4644 => x"20c00000",
  4645 => x"e0000000",
  4646 => x"20e02000",
  4647 => x"0020a060",
  4648 => x"20000000",
  4649 => x"00000000",
  4650 => x"00000000",
  4651 => x"00000000",
  4652 => x"00000000",
  4653 => x"00000000",
  4654 => x"00000000",
  4655 => x"00030007",
  4656 => x"00070701",
  4657 => x"00000000",
  4658 => x"00000000",
  4659 => x"00000300",
  4660 => x"c0030000",
  4661 => x"034242c0",
  4662 => x"00c34242",
  4663 => x"0000c380",
  4664 => x"01c00340",
  4665 => x"c04300c0",
  4666 => x"43408001",
  4667 => x"c20201c0",
  4668 => x"00c38202",
  4669 => x"80c00300",
  4670 => x"00c04342",
  4671 => x"8202c040",
  4672 => x"40800000",
  4673 => x"c0404000",
  4674 => x"80404000",
  4675 => x"00c04040",
  4676 => x"8000c040",
  4677 => x"4000c080",
  4678 => x"00c00000",
  4679 => x"00000000",
  4680 => x"00000000",
  4681 => x"00000000",
  4682 => x"00000000",
  4683 => x"00ff0000",
  4684 => x"0000c645",
  4685 => x"44800785",
  4686 => x"45408007",
  4687 => x"80424700",
  4688 => x"80474000",
  4689 => x"07c14344",
  4690 => x"00c38404",
  4691 => x"c30007c1",
  4692 => x"42418700",
  4693 => x"80404784",
  4694 => x"04c34047",
  4695 => x"8101c640",
  4696 => x"40070505",
  4697 => x"00040502",
  4698 => x"00000704",
  4699 => x"04030007",
  4700 => x"05050007",
  4701 => x"00020700",
  4702 => x"00000000",
  4703 => x"00000000",
  4704 => x"00000000",
  4705 => x"00000000",
  4706 => x"0000ff00",
  4707 => x"00000007",
  4708 => x"01030500",
  4709 => x"03040403",
  4710 => x"00040502",
  4711 => x"00040502",
  4712 => x"00000705",
  4713 => x"05000700",
  4714 => x"02070000",
  4715 => x"07040403",
  4716 => x"00030404",
  4717 => x"03000701",
  4718 => x"03050007",
  4719 => x"01010000",
  4720 => x"00000000",
  4721 => x"00000000",
  4722 => x"00000000",
  4723 => x"00000000",
  4724 => x"00000000",
  4725 => x"71756974",
  4726 => x"00000000",
  4727 => x"68656c70",
  4728 => x"00000000",
  4729 => x"73686f77",
  4730 => x"2042504d",
  4731 => x"20726567",
  4732 => x"69737465",
  4733 => x"72730000",
  4734 => x"62706d00",
  4735 => x"73686f77",
  4736 => x"2f736574",
  4737 => x"20646562",
  4738 => x"75672072",
  4739 => x"65676973",
  4740 => x"74657273",
  4741 => x"203c7365",
  4742 => x"74206d6f",
  4743 => x"64653e00",
  4744 => x"64656275",
  4745 => x"67000000",
  4746 => x"73797374",
  4747 => x"656d2072",
  4748 => x"65736574",
  4749 => x"00000000",
  4750 => x"72657365",
  4751 => x"74000000",
  4752 => x"73686f77",
  4753 => x"20646562",
  4754 => x"75672062",
  4755 => x"75666665",
  4756 => x"72203c6c",
  4757 => x"656e6774",
  4758 => x"683e0000",
  4759 => x"646f776e",
  4760 => x"6c6f6164",
  4761 => x"20646562",
  4762 => x"75672062",
  4763 => x"75666665",
  4764 => x"72202878",
  4765 => x"6d6f6465",
  4766 => x"6d290000",
  4767 => x"62726561",
  4768 => x"64000000",
  4769 => x"75706c6f",
  4770 => x"61642064",
  4771 => x"65627567",
  4772 => x"20627566",
  4773 => x"66657220",
  4774 => x"28786d6f",
  4775 => x"64656d29",
  4776 => x"00000000",
  4777 => x"62777269",
  4778 => x"74650000",
  4779 => x"636c6561",
  4780 => x"72206465",
  4781 => x"62756720",
  4782 => x"62756666",
  4783 => x"65720000",
  4784 => x"62636c65",
  4785 => x"61720000",
  4786 => x"73657475",
  4787 => x"70206368",
  4788 => x"616e6e65",
  4789 => x"6c207465",
  4790 => x"7374203c",
  4791 => x"70302e2e",
  4792 => x"353e0000",
  4793 => x"63687465",
  4794 => x"73740000",
  4795 => x"74657374",
  4796 => x"67656e65",
  4797 => x"7261746f",
  4798 => x"72203c73",
  4799 => x"63616c65",
  4800 => x"723e203c",
  4801 => x"72657374",
  4802 => x"6172743e",
  4803 => x"00000000",
  4804 => x"74657374",
  4805 => x"67656e00",
  4806 => x"3c6d7574",
  4807 => x"655f6e3e",
  4808 => x"203c7273",
  4809 => x"745f6e3e",
  4810 => x"203c6270",
  4811 => x"625f6e3e",
  4812 => x"203c6f73",
  4813 => x"72313e20",
  4814 => x"3c6f7372",
  4815 => x"323e0000",
  4816 => x"64616363",
  4817 => x"6f6e6600",
  4818 => x"636c6b20",
  4819 => x"3c73656c",
  4820 => x"6563743e",
  4821 => x"2030203d",
  4822 => x"20696e74",
  4823 => x"2c203120",
  4824 => x"3d206578",
  4825 => x"74000000",
  4826 => x"636c6b00",
  4827 => x"73686f77",
  4828 => x"20737973",
  4829 => x"74656d20",
  4830 => x"696e666f",
  4831 => x"203c7665",
  4832 => x"72626f73",
  4833 => x"653e0000",
  4834 => x"73797369",
  4835 => x"6e666f00",
  4836 => x"72756e6e",
  4837 => x"696e6720",
  4838 => x"6c696768",
  4839 => x"74000000",
  4840 => x"72756e00",
  4841 => x"72756e20",
  4842 => x"64697370",
  4843 => x"6c617920",
  4844 => x"74657374",
  4845 => x"2066756e",
  4846 => x"6374696f",
  4847 => x"6e000000",
  4848 => x"64697370",
  4849 => x"6c617900",
  4850 => x"73657420",
  4851 => x"6261636b",
  4852 => x"6c696768",
  4853 => x"74203c30",
  4854 => x"2e2e3331",
  4855 => x"3e000000",
  4856 => x"6261636b",
  4857 => x"00000000",
  4858 => x"73686f77",
  4859 => x"206c6f67",
  4860 => x"6f206f6e",
  4861 => x"20676c63",
  4862 => x"64000000",
  4863 => x"6c6f676f",
  4864 => x"00000000",
  4865 => x"63686563",
  4866 => x"6b204932",
  4867 => x"43206164",
  4868 => x"64726573",
  4869 => x"73000000",
  4870 => x"69326300",
  4871 => x"72656164",
  4872 => x"20454550",
  4873 => x"524f4d20",
  4874 => x"3c627573",
  4875 => x"3e203c69",
  4876 => x"32635f61",
  4877 => x"6464723e",
  4878 => x"203c6c65",
  4879 => x"6e677468",
  4880 => x"3e000000",
  4881 => x"65657072",
  4882 => x"6f6d0000",
  4883 => x"41444320",
  4884 => x"72656769",
  4885 => x"73746572",
  4886 => x"20747261",
  4887 => x"6e736665",
  4888 => x"72203c76",
  4889 => x"616c7565",
  4890 => x"3e000000",
  4891 => x"61747261",
  4892 => x"6e730000",
  4893 => x"696e6974",
  4894 => x"20414443",
  4895 => x"20726567",
  4896 => x"69737465",
  4897 => x"72730000",
  4898 => x"61696e69",
  4899 => x"74000000",
  4900 => x"616c6961",
  4901 => x"7320666f",
  4902 => x"72207800",
  4903 => x"6d656d00",
  4904 => x"77726974",
  4905 => x"6520776f",
  4906 => x"7264203c",
  4907 => x"61646472",
  4908 => x"3e203c6c",
  4909 => x"656e6774",
  4910 => x"683e203c",
  4911 => x"76616c75",
  4912 => x"65287329",
  4913 => x"3e000000",
  4914 => x"776d656d",
  4915 => x"00000000",
  4916 => x"6558616d",
  4917 => x"696e6520",
  4918 => x"6d656d6f",
  4919 => x"72790000",
  4920 => x"636c6561",
  4921 => x"72207363",
  4922 => x"7265656e",
  4923 => x"00000000",
  4924 => x"636c6561",
  4925 => x"72000000",
  4926 => x"0a307800",
  4927 => x"69326320",
  4928 => x"464d430a",
  4929 => x"00000000",
  4930 => x"61646472",
  4931 => x"6573733a",
  4932 => x"20307800",
  4933 => x"2020202d",
  4934 => x"2d3e2020",
  4935 => x"2041434b",
  4936 => x"0a000000",
  4937 => x"72656164",
  4938 => x"20646174",
  4939 => x"61202800",
  4940 => x"20627974",
  4941 => x"65732920",
  4942 => x"66726f6d",
  4943 => x"20493243",
  4944 => x"2d616464",
  4945 => x"72657373",
  4946 => x"20307800",
  4947 => x"0a0a0000",
  4948 => x"6e6f6163",
  4949 => x"6b200000",
  4950 => x"6368726f",
  4951 => x"6e74656c",
  4952 => x"20726567",
  4953 => x"20307800",
  4954 => x"3a203078",
  4955 => x"00000000",
  4956 => x"206e6163",
  4957 => x"6b000000",
  4958 => x"6572726f",
  4959 => x"7220286e",
  4960 => x"61636b29",
  4961 => x"0a000000",
  4962 => x"6265616d",
  4963 => x"20706f73",
  4964 => x"6974696f",
  4965 => x"6e206d6f",
  4966 => x"6e69746f",
  4967 => x"72207265",
  4968 => x"67697374",
  4969 => x"65727300",
  4970 => x"0a202020",
  4971 => x"20202020",
  4972 => x"20202020",
  4973 => x"20202020",
  4974 => x"20202020",
  4975 => x"20202020",
  4976 => x"20636861",
  4977 => x"6e6e656c",
  4978 => x"20302020",
  4979 => x"20636861",
  4980 => x"6e6e656c",
  4981 => x"20312020",
  4982 => x"20636861",
  4983 => x"6e6e656c",
  4984 => x"20322020",
  4985 => x"20636861",
  4986 => x"6e6e656c",
  4987 => x"20330000",
  4988 => x"0a202020",
  4989 => x"20202020",
  4990 => x"20202020",
  4991 => x"20202020",
  4992 => x"20202020",
  4993 => x"20202020",
  4994 => x"202d2d2d",
  4995 => x"2d20686f",
  4996 => x"72697a6f",
  4997 => x"6e74616c",
  4998 => x"202d2d2d",
  4999 => x"2d2d2020",
  5000 => x"202d2d2d",
  5001 => x"2d2d2d20",
  5002 => x"76657274",
  5003 => x"6963616c",
  5004 => x"202d2d2d",
  5005 => x"2d2d0000",
  5006 => x"0a736361",
  5007 => x"6c657220",
  5008 => x"76616c75",
  5009 => x"65732020",
  5010 => x"20202020",
  5011 => x"20202020",
  5012 => x"20000000",
  5013 => x"0a6e6f69",
  5014 => x"73652063",
  5015 => x"6f6d7065",
  5016 => x"6e736174",
  5017 => x"696f6e20",
  5018 => x"20202020",
  5019 => x"20000000",
  5020 => x"0a6d6561",
  5021 => x"73757265",
  5022 => x"6d656e74",
  5023 => x"20202020",
  5024 => x"20202020",
  5025 => x"20202020",
  5026 => x"20000000",
  5027 => x"0a73756d",
  5028 => x"20636861",
  5029 => x"6e6e656c",
  5030 => x"2020203a",
  5031 => x"20000000",
  5032 => x"0a706f73",
  5033 => x"6974696f",
  5034 => x"6e20636f",
  5035 => x"6d707574",
  5036 => x"6174696f",
  5037 => x"6e000000",
  5038 => x"0a202073",
  5039 => x"63616c65",
  5040 => x"72207661",
  5041 => x"6c756573",
  5042 => x"20202020",
  5043 => x"20202020",
  5044 => x"20000000",
  5045 => x"0a20206f",
  5046 => x"66667365",
  5047 => x"74202020",
  5048 => x"20202020",
  5049 => x"20202020",
  5050 => x"20202020",
  5051 => x"20000000",
  5052 => x"0a6f7574",
  5053 => x"70757420",
  5054 => x"73656c65",
  5055 => x"6374203a",
  5056 => x"20000000",
  5057 => x"6368616e",
  5058 => x"6e656c20",
  5059 => x"30000000",
  5060 => x"0a63616c",
  5061 => x"63207374",
  5062 => x"61746520",
  5063 => x"2020203a",
  5064 => x"20307800",
  5065 => x"0a202064",
  5066 => x"69766964",
  5067 => x"656e6420",
  5068 => x"63757474",
  5069 => x"65640000",
  5070 => x"0a20206e",
  5071 => x"6f697365",
  5072 => x"20636f6d",
  5073 => x"70656e73",
  5074 => x"6174696f",
  5075 => x"6e20746f",
  5076 => x"20626967",
  5077 => x"00000000",
  5078 => x"0a20206e",
  5079 => x"6f697365",
  5080 => x"2076616c",
  5081 => x"75652063",
  5082 => x"75747465",
  5083 => x"64000000",
  5084 => x"0a202073",
  5085 => x"756d2076",
  5086 => x"616c7565",
  5087 => x"20637574",
  5088 => x"74656400",
  5089 => x"76657274",
  5090 => x"6963616c",
  5091 => x"00000000",
  5092 => x"686f7269",
  5093 => x"7a6f6e74",
  5094 => x"616c0000",
  5095 => x"73756d00",
  5096 => x"6368616e",
  5097 => x"6e656c20",
  5098 => x"33000000",
  5099 => x"6368616e",
  5100 => x"6e656c20",
  5101 => x"32000000",
  5102 => x"6368616e",
  5103 => x"6e656c20",
  5104 => x"31000000",
  5105 => x"786d6f64",
  5106 => x"656d2074",
  5107 => x"72616e73",
  5108 => x"6d69742e",
  5109 => x"2e2e0a00",
  5110 => x"20627974",
  5111 => x"65732074",
  5112 => x"72616e73",
  5113 => x"6d697474",
  5114 => x"65640a00",
  5115 => x"63616e63",
  5116 => x"656c0a00",
  5117 => x"72657472",
  5118 => x"79206f75",
  5119 => x"740a0000",
  5120 => x"786d6f64",
  5121 => x"656d2072",
  5122 => x"65636569",
  5123 => x"76652e2e",
  5124 => x"2e0a0000",
  5125 => x"20627974",
  5126 => x"65732072",
  5127 => x"65636569",
  5128 => x"7665640a",
  5129 => x"00000000",
  5130 => x"72782062",
  5131 => x"75666665",
  5132 => x"72206675",
  5133 => x"6c6c0a00",
  5134 => x"74696d65",
  5135 => x"206f7574",
  5136 => x"0a000000",
  5137 => x"64656275",
  5138 => x"67207265",
  5139 => x"67697374",
  5140 => x"65727300",
  5141 => x"0a6d6f64",
  5142 => x"65202020",
  5143 => x"20202020",
  5144 => x"203a2000",
  5145 => x"0a616464",
  5146 => x"72657373",
  5147 => x"20302020",
  5148 => x"203a2030",
  5149 => x"78000000",
  5150 => x"0a616464",
  5151 => x"72657373",
  5152 => x"20312020",
  5153 => x"203a2030",
  5154 => x"78000000",
  5155 => x"0a627566",
  5156 => x"66657220",
  5157 => x"73697a65",
  5158 => x"203a2000",
  5159 => x"65787465",
  5160 => x"726e616c",
  5161 => x"20636c6f",
  5162 => x"636b2000",
  5163 => x"61637469",
  5164 => x"76650a00",
  5165 => x"4e4f5420",
  5166 => x"00000000",
  5167 => x"6265616d",
  5168 => x"20706f73",
  5169 => x"6974696f",
  5170 => x"6e206d6f",
  5171 => x"6e69746f",
  5172 => x"72000000",
  5173 => x"20286f6e",
  5174 => x"2073696d",
  5175 => x"290a0000",
  5176 => x"0a636f6d",
  5177 => x"70696c65",
  5178 => x"643a204a",
  5179 => x"756c2020",
  5180 => x"31203230",
  5181 => x"31312020",
  5182 => x"30393a30",
  5183 => x"353a3030",
  5184 => x"00000000",
  5185 => x"0a737973",
  5186 => x"74656d20",
  5187 => x"636c6f63",
  5188 => x"6b3a2000",
  5189 => x"204d487a",
  5190 => x"0a000000",
  5191 => x"44454255",
  5192 => x"47204d4f",
  5193 => x"44450000",
  5194 => x"204f4e0a",
  5195 => x"00000000",
  5196 => x"00000ef0",
  5197 => x"00000fde",
  5198 => x"00000fd3",
  5199 => x"00000fc8",
  5200 => x"00000fbd",
  5201 => x"00000fb2",
  5202 => x"00000fa7",
  5203 => x"0187fc09",
  5204 => x"026f0000",
  5205 => x"0003fff6",
  5206 => x"00060000",
  5207 => x"3e200000",
  5208 => x"636f6d6d",
  5209 => x"616e6420",
  5210 => x"6e6f7420",
  5211 => x"666f756e",
  5212 => x"642e0a00",
  5213 => x"73757070",
  5214 => x"6f727465",
  5215 => x"6420636f",
  5216 => x"6d6d616e",
  5217 => x"64733a0a",
  5218 => x"0a000000",
  5219 => x"202d2000",
  5220 => x"76656e64",
  5221 => x"6f723f20",
  5222 => x"20000000",
  5223 => x"67616973",
  5224 => x"6c657220",
  5225 => x"20000000",
  5226 => x"756e6b6e",
  5227 => x"6f776e20",
  5228 => x"64657669",
  5229 => x"63650000",
  5230 => x"485a4452",
  5231 => x"20202020",
  5232 => x"20000000",
  5233 => x"47656e65",
  5234 => x"72616c20",
  5235 => x"50757270",
  5236 => x"6f736520",
  5237 => x"492f4f20",
  5238 => x"706f7274",
  5239 => x"00000000",
  5240 => x"56474120",
  5241 => x"636f6e74",
  5242 => x"726f6c6c",
  5243 => x"65720000",
  5244 => x"4475616c",
  5245 => x"2d706f72",
  5246 => x"74204148",
  5247 => x"42205352",
  5248 => x"414d206d",
  5249 => x"6f64756c",
  5250 => x"65000000",
  5251 => x"64656275",
  5252 => x"67206275",
  5253 => x"66666572",
  5254 => x"20636f6e",
  5255 => x"74726f6c",
  5256 => x"00000000",
  5257 => x"74726967",
  5258 => x"67657220",
  5259 => x"67656e65",
  5260 => x"7261746f",
  5261 => x"72000000",
  5262 => x"64656275",
  5263 => x"6720636f",
  5264 => x"6e736f6c",
  5265 => x"65000000",
  5266 => x"44434d20",
  5267 => x"70686173",
  5268 => x"65207368",
  5269 => x"69667420",
  5270 => x"636f6e74",
  5271 => x"726f6c00",
  5272 => x"5a505520",
  5273 => x"4d656d6f",
  5274 => x"72792077",
  5275 => x"72617070",
  5276 => x"65720000",
  5277 => x"5a505520",
  5278 => x"41484220",
  5279 => x"57726170",
  5280 => x"70657200",
  5281 => x"4148422f",
  5282 => x"41504220",
  5283 => x"42726964",
  5284 => x"67650000",
  5285 => x"4d6f6475",
  5286 => x"6c617220",
  5287 => x"54696d65",
  5288 => x"7220556e",
  5289 => x"69740000",
  5290 => x"414d4241",
  5291 => x"20577261",
  5292 => x"70706572",
  5293 => x"20666f72",
  5294 => x"204f4320",
  5295 => x"4932432d",
  5296 => x"6d617374",
  5297 => x"65720000",
  5298 => x"47656e65",
  5299 => x"72696320",
  5300 => x"55415254",
  5301 => x"00000000",
  5302 => x"20206170",
  5303 => x"62736c76",
  5304 => x"00000000",
  5305 => x"76656e64",
  5306 => x"20307800",
  5307 => x"64657620",
  5308 => x"30780000",
  5309 => x"76657220",
  5310 => x"00000000",
  5311 => x"69727120",
  5312 => x"00000000",
  5313 => x"61646472",
  5314 => x"20307800",
  5315 => x"6168626d",
  5316 => x"73740000",
  5317 => x"61686273",
  5318 => x"6c760000",
  5319 => x"00002201",
  5320 => x"000022ac",
  5321 => x"000022a1",
  5322 => x"00002296",
  5323 => x"0000228b",
  5324 => x"00002280",
  5325 => x"00002275",
  5326 => x"0000226a",
  5327 => x"04580808",
  5328 => x"20ff0000",
  5329 => x"0000534c",
  5330 => x"0000542c",
  5331 => x"02010305",
  5332 => x"05070501",
  5333 => x"03030505",
  5334 => x"02030104",
  5335 => x"05050505",
  5336 => x"05050505",
  5337 => x"05050101",
  5338 => x"04050404",
  5339 => x"07050505",
  5340 => x"05050505",
  5341 => x"05030405",
  5342 => x"05050505",
  5343 => x"05050505",
  5344 => x"05050505",
  5345 => x"05050503",
  5346 => x"04030505",
  5347 => x"02050504",
  5348 => x"05050405",
  5349 => x"04010204",
  5350 => x"02050404",
  5351 => x"05050404",
  5352 => x"04040507",
  5353 => x"05040404",
  5354 => x"02040500",
  5355 => x"04050200",
  5356 => x"04080303",
  5357 => x"04090003",
  5358 => x"06000000",
  5359 => x"00020204",
  5360 => x"04040400",
  5361 => x"04060003",
  5362 => x"05000000",
  5363 => x"00000404",
  5364 => x"05050204",
  5365 => x"05060305",
  5366 => x"04030705",
  5367 => x"04050303",
  5368 => x"02040502",
  5369 => x"03020405",
  5370 => x"06060604",
  5371 => x"05050505",
  5372 => x"05050504",
  5373 => x"04040404",
  5374 => x"03030303",
  5375 => x"05050505",
  5376 => x"05050505",
  5377 => x"05040404",
  5378 => x"04050404",
  5379 => x"04040404",
  5380 => x"04040503",
  5381 => x"04040404",
  5382 => x"02020303",
  5383 => x"04040404",
  5384 => x"04040405",
  5385 => x"04040404",
  5386 => x"04030303",
  5387 => x"00005f07",
  5388 => x"0007741c",
  5389 => x"771c172e",
  5390 => x"6a3e2b3a",
  5391 => x"06493608",
  5392 => x"36493036",
  5393 => x"49597648",
  5394 => x"073c4281",
  5395 => x"81423c0a",
  5396 => x"041f040a",
  5397 => x"08083e08",
  5398 => x"08806008",
  5399 => x"080840c0",
  5400 => x"300c033e",
  5401 => x"4141413e",
  5402 => x"44427f40",
  5403 => x"40466151",
  5404 => x"49462241",
  5405 => x"49493618",
  5406 => x"14127f10",
  5407 => x"27454545",
  5408 => x"393e4949",
  5409 => x"49300101",
  5410 => x"710d0336",
  5411 => x"49494936",
  5412 => x"06494929",
  5413 => x"1e36d008",
  5414 => x"14224114",
  5415 => x"14141414",
  5416 => x"41221408",
  5417 => x"02510906",
  5418 => x"3c4299a5",
  5419 => x"bd421c7c",
  5420 => x"1211127c",
  5421 => x"7f494949",
  5422 => x"363e4141",
  5423 => x"41227f41",
  5424 => x"41413e7f",
  5425 => x"49494941",
  5426 => x"7f090909",
  5427 => x"013e4149",
  5428 => x"497a7f08",
  5429 => x"08087f41",
  5430 => x"7f414041",
  5431 => x"413f7f08",
  5432 => x"1422417f",
  5433 => x"40404040",
  5434 => x"7f060c06",
  5435 => x"7f7f0608",
  5436 => x"307f3e41",
  5437 => x"41413e7f",
  5438 => x"09090906",
  5439 => x"3e4161c1",
  5440 => x"be7f0919",
  5441 => x"29462649",
  5442 => x"49493201",
  5443 => x"017f0101",
  5444 => x"3f404040",
  5445 => x"3f073840",
  5446 => x"38071f60",
  5447 => x"1f601f63",
  5448 => x"14081463",
  5449 => x"01067806",
  5450 => x"01615149",
  5451 => x"45437f41",
  5452 => x"41030c30",
  5453 => x"c041417f",
  5454 => x"04020102",
  5455 => x"04808080",
  5456 => x"80800102",
  5457 => x"20545454",
  5458 => x"787f4444",
  5459 => x"44383844",
  5460 => x"44443844",
  5461 => x"44447f38",
  5462 => x"54545458",
  5463 => x"087e0901",
  5464 => x"18a4a4a4",
  5465 => x"787f0404",
  5466 => x"787d807d",
  5467 => x"7f102844",
  5468 => x"3f407c04",
  5469 => x"7804787c",
  5470 => x"04047838",
  5471 => x"444438fc",
  5472 => x"24242418",
  5473 => x"18242424",
  5474 => x"fc7c0804",
  5475 => x"04485454",
  5476 => x"24043f44",
  5477 => x"403c4040",
  5478 => x"7c1c2040",
  5479 => x"201c1c60",
  5480 => x"601c6060",
  5481 => x"1c442810",
  5482 => x"28449ca0",
  5483 => x"601c6454",
  5484 => x"544c187e",
  5485 => x"8181ffff",
  5486 => x"81817e18",
  5487 => x"18040810",
  5488 => x"0c143e55",
  5489 => x"55ff8181",
  5490 => x"81ff8060",
  5491 => x"80608060",
  5492 => x"60600060",
  5493 => x"60006060",
  5494 => x"047f0414",
  5495 => x"7f140201",
  5496 => x"01024629",
  5497 => x"1608344a",
  5498 => x"31483000",
  5499 => x"18243e41",
  5500 => x"227f4941",
  5501 => x"03040403",
  5502 => x"03040304",
  5503 => x"04030403",
  5504 => x"183c3c18",
  5505 => x"08080808",
  5506 => x"03010203",
  5507 => x"020e020e",
  5508 => x"060e0048",
  5509 => x"30384438",
  5510 => x"54483844",
  5511 => x"fe44487e",
  5512 => x"49014438",
  5513 => x"28384403",
  5514 => x"147c1403",
  5515 => x"e7e74e55",
  5516 => x"55390101",
  5517 => x"0001011c",
  5518 => x"2a555522",
  5519 => x"1c1d151e",
  5520 => x"18240018",
  5521 => x"24080808",
  5522 => x"18080808",
  5523 => x"3c42bd95",
  5524 => x"a9423c01",
  5525 => x"01010101",
  5526 => x"06090906",
  5527 => x"44445f44",
  5528 => x"44191512",
  5529 => x"15150a02",
  5530 => x"01fc2020",
  5531 => x"1c0e7f01",
  5532 => x"7f011818",
  5533 => x"00804002",
  5534 => x"1f060909",
  5535 => x"06241800",
  5536 => x"2418824f",
  5537 => x"304c62f1",
  5538 => x"824f300c",
  5539 => x"d2b1955f",
  5540 => x"304c62f1",
  5541 => x"30484520",
  5542 => x"60392e38",
  5543 => x"6060382e",
  5544 => x"3960701d",
  5545 => x"131d7072",
  5546 => x"1d121e71",
  5547 => x"701d121d",
  5548 => x"70603b25",
  5549 => x"3b607e11",
  5550 => x"7f49411e",
  5551 => x"2161927c",
  5552 => x"5556447c",
  5553 => x"5655447c",
  5554 => x"5655467d",
  5555 => x"54544545",
  5556 => x"7e44447e",
  5557 => x"45467d46",
  5558 => x"457c4508",
  5559 => x"7f49413e",
  5560 => x"7e091222",
  5561 => x"7d384546",
  5562 => x"44383844",
  5563 => x"46453838",
  5564 => x"46454638",
  5565 => x"3a454546",
  5566 => x"39384544",
  5567 => x"45382214",
  5568 => x"081422bc",
  5569 => x"625a463d",
  5570 => x"3c41423c",
  5571 => x"3c42413c",
  5572 => x"3c42413e",
  5573 => x"3d40403d",
  5574 => x"0608f209",
  5575 => x"067f2222",
  5576 => x"1cfe0989",
  5577 => x"76205556",
  5578 => x"78205655",
  5579 => x"78225555",
  5580 => x"7a235556",
  5581 => x"7b205554",
  5582 => x"79275557",
  5583 => x"78205438",
  5584 => x"54483844",
  5585 => x"c4385556",
  5586 => x"58385655",
  5587 => x"583a5555",
  5588 => x"5a395454",
  5589 => x"59017a7a",
  5590 => x"01027902",
  5591 => x"02780260",
  5592 => x"91927c7b",
  5593 => x"090a7338",
  5594 => x"45463838",
  5595 => x"4645383a",
  5596 => x"45453a3b",
  5597 => x"45463b39",
  5598 => x"44443908",
  5599 => x"082a0808",
  5600 => x"b8644c3a",
  5601 => x"3c41427c",
  5602 => x"3c42417c",
  5603 => x"3a41417a",
  5604 => x"3d40407d",
  5605 => x"986219ff",
  5606 => x"423c9a60",
  5607 => x"1a000000",
  5608 => x"30622020",
  5609 => x"20202020",
  5610 => x"20202020",
  5611 => x"20202020",
  5612 => x"20202020",
  5613 => x"20202020",
  5614 => x"20202020",
  5615 => x"20202020",
  5616 => x"20200000",
  5617 => x"20202020",
  5618 => x"20202020",
  5619 => x"00000000",
  5620 => x"00202020",
  5621 => x"20202020",
  5622 => x"20202828",
  5623 => x"28282820",
  5624 => x"20202020",
  5625 => x"20202020",
  5626 => x"20202020",
  5627 => x"20202020",
  5628 => x"20881010",
  5629 => x"10101010",
  5630 => x"10101010",
  5631 => x"10101010",
  5632 => x"10040404",
  5633 => x"04040404",
  5634 => x"04040410",
  5635 => x"10101010",
  5636 => x"10104141",
  5637 => x"41414141",
  5638 => x"01010101",
  5639 => x"01010101",
  5640 => x"01010101",
  5641 => x"01010101",
  5642 => x"01010101",
  5643 => x"10101010",
  5644 => x"10104242",
  5645 => x"42424242",
  5646 => x"02020202",
  5647 => x"02020202",
  5648 => x"02020202",
  5649 => x"02020202",
  5650 => x"02020202",
  5651 => x"10101010",
  5652 => x"20000000",
  5653 => x"00000000",
  5654 => x"00000000",
  5655 => x"00000000",
  5656 => x"00000000",
  5657 => x"00000000",
  5658 => x"00000000",
  5659 => x"00000000",
  5660 => x"00000000",
  5661 => x"00000000",
  5662 => x"00000000",
  5663 => x"00000000",
  5664 => x"00000000",
  5665 => x"00000000",
  5666 => x"00000000",
  5667 => x"00000000",
  5668 => x"00000000",
  5669 => x"00000000",
  5670 => x"00000000",
  5671 => x"00000000",
  5672 => x"00000000",
  5673 => x"00000000",
  5674 => x"00000000",
  5675 => x"00000000",
  5676 => x"00000000",
  5677 => x"00000000",
  5678 => x"00000000",
  5679 => x"00000000",
  5680 => x"00000000",
  5681 => x"00000000",
  5682 => x"00000000",
  5683 => x"00000000",
  5684 => x"00000000",
  5685 => x"43000000",
  5686 => x"00000000",
  5687 => x"80000c00",
  5688 => x"80000b00",
  5689 => x"80000800",
  5690 => x"00000000",
  5691 => x"ff000000",
  5692 => x"00000000",
  5693 => x"00000000",
  5694 => x"00ffffff",
  5695 => x"ff00ffff",
  5696 => x"ffff00ff",
  5697 => x"ffffff00",
  5698 => x"00000000",
  5699 => x"00000000",
  5700 => x"80000a00",
  5701 => x"80000700",
  5702 => x"80000600",
  5703 => x"80000400",
  5704 => x"80000200",
  5705 => x"80000100",
  5706 => x"80000004",
  5707 => x"80000000",
  5708 => x"00005934",
  5709 => x"00000000",
  5710 => x"00005b9c",
  5711 => x"00005bf8",
  5712 => x"00005c54",
  5713 => x"00000000",
  5714 => x"00000000",
  5715 => x"00000000",
  5716 => x"00000000",
  5717 => x"00000000",
  5718 => x"00000000",
  5719 => x"00000000",
  5720 => x"00000000",
  5721 => x"00000000",
  5722 => x"000058d4",
  5723 => x"00000000",
  5724 => x"00000000",
  5725 => x"00000000",
  5726 => x"00000000",
  5727 => x"00000000",
  5728 => x"00000000",
  5729 => x"00000000",
  5730 => x"00000000",
  5731 => x"00000000",
  5732 => x"00000000",
  5733 => x"00000000",
  5734 => x"00000000",
  5735 => x"00000000",
  5736 => x"00000000",
  5737 => x"00000000",
  5738 => x"00000000",
  5739 => x"00000000",
  5740 => x"00000000",
  5741 => x"00000000",
  5742 => x"00000000",
  5743 => x"00000000",
  5744 => x"00000000",
  5745 => x"00000000",
  5746 => x"00000000",
  5747 => x"00000000",
  5748 => x"00000000",
  5749 => x"00000000",
  5750 => x"00000000",
  5751 => x"00000001",
  5752 => x"330eabcd",
  5753 => x"1234e66d",
  5754 => x"deec0005",
  5755 => x"000b0000",
  5756 => x"00000000",
  5757 => x"00000000",
  5758 => x"00000000",
  5759 => x"00000000",
  5760 => x"00000000",
  5761 => x"00000000",
  5762 => x"00000000",
  5763 => x"00000000",
  5764 => x"00000000",
  5765 => x"00000000",
  5766 => x"00000000",
  5767 => x"00000000",
  5768 => x"00000000",
  5769 => x"00000000",
  5770 => x"00000000",
  5771 => x"00000000",
  5772 => x"00000000",
  5773 => x"00000000",
  5774 => x"00000000",
  5775 => x"00000000",
  5776 => x"00000000",
  5777 => x"00000000",
  5778 => x"00000000",
  5779 => x"00000000",
  5780 => x"00000000",
  5781 => x"00000000",
  5782 => x"00000000",
  5783 => x"00000000",
  5784 => x"00000000",
  5785 => x"00000000",
  5786 => x"00000000",
  5787 => x"00000000",
  5788 => x"00000000",
  5789 => x"00000000",
  5790 => x"00000000",
  5791 => x"00000000",
  5792 => x"00000000",
  5793 => x"00000000",
  5794 => x"00000000",
  5795 => x"00000000",
  5796 => x"00000000",
  5797 => x"00000000",
  5798 => x"00000000",
  5799 => x"00000000",
  5800 => x"00000000",
  5801 => x"00000000",
  5802 => x"00000000",
  5803 => x"00000000",
  5804 => x"00000000",
  5805 => x"00000000",
  5806 => x"00000000",
  5807 => x"00000000",
  5808 => x"00000000",
  5809 => x"00000000",
  5810 => x"00000000",
  5811 => x"00000000",
  5812 => x"00000000",
  5813 => x"00000000",
  5814 => x"00000000",
  5815 => x"00000000",
  5816 => x"00000000",
  5817 => x"00000000",
  5818 => x"00000000",
  5819 => x"00000000",
  5820 => x"00000000",
  5821 => x"00000000",
  5822 => x"00000000",
  5823 => x"00000000",
  5824 => x"00000000",
  5825 => x"00000000",
  5826 => x"00000000",
  5827 => x"00000000",
  5828 => x"00000000",
  5829 => x"00000000",
  5830 => x"00000000",
  5831 => x"00000000",
  5832 => x"00000000",
  5833 => x"00000000",
  5834 => x"00000000",
  5835 => x"00000000",
  5836 => x"00000000",
  5837 => x"00000000",
  5838 => x"00000000",
  5839 => x"00000000",
  5840 => x"00000000",
  5841 => x"00000000",
  5842 => x"00000000",
  5843 => x"00000000",
  5844 => x"00000000",
  5845 => x"00000000",
  5846 => x"00000000",
  5847 => x"00000000",
  5848 => x"00000000",
  5849 => x"00000000",
  5850 => x"00000000",
  5851 => x"00000000",
  5852 => x"00000000",
  5853 => x"00000000",
  5854 => x"00000000",
  5855 => x"00000000",
  5856 => x"00000000",
  5857 => x"00000000",
  5858 => x"00000000",
  5859 => x"00000000",
  5860 => x"00000000",
  5861 => x"00000000",
  5862 => x"00000000",
  5863 => x"00000000",
  5864 => x"00000000",
  5865 => x"00000000",
  5866 => x"00000000",
  5867 => x"00000000",
  5868 => x"00000000",
  5869 => x"00000000",
  5870 => x"00000000",
  5871 => x"00000000",
  5872 => x"00000000",
  5873 => x"00000000",
  5874 => x"00000000",
  5875 => x"00000000",
  5876 => x"00000000",
  5877 => x"00000000",
  5878 => x"00000000",
  5879 => x"00000000",
  5880 => x"00000000",
  5881 => x"00000000",
  5882 => x"00000000",
  5883 => x"00000000",
  5884 => x"00000000",
  5885 => x"00000000",
  5886 => x"00000000",
  5887 => x"00000000",
  5888 => x"00000000",
  5889 => x"00000000",
  5890 => x"00000000",
  5891 => x"00000000",
  5892 => x"00000000",
  5893 => x"00000000",
  5894 => x"00000000",
  5895 => x"00000000",
  5896 => x"00000000",
  5897 => x"00000000",
  5898 => x"00000000",
  5899 => x"00000000",
  5900 => x"00000000",
  5901 => x"00000000",
  5902 => x"00000000",
  5903 => x"00000000",
  5904 => x"00000000",
  5905 => x"00000000",
  5906 => x"00000000",
  5907 => x"00000000",
  5908 => x"00000000",
  5909 => x"00000000",
  5910 => x"00000000",
  5911 => x"00000000",
  5912 => x"00000000",
  5913 => x"00000000",
  5914 => x"00000000",
  5915 => x"00000000",
  5916 => x"00000000",
  5917 => x"00000000",
  5918 => x"00000000",
  5919 => x"00000000",
  5920 => x"00000000",
  5921 => x"00000000",
  5922 => x"00000000",
  5923 => x"00000000",
  5924 => x"00000000",
  5925 => x"00000000",
  5926 => x"00000000",
  5927 => x"00000000",
  5928 => x"00000000",
  5929 => x"00000000",
  5930 => x"00000000",
  5931 => x"00000000",
  5932 => x"00000000",
  5933 => x"00000000",
  5934 => x"00000000",
  5935 => x"00000000",
  5936 => x"00000000",
  5937 => x"00000000",
  5938 => x"00000000",
  5939 => x"00000000",
  5940 => x"00000000",
  5941 => x"00000000",
  5942 => x"00000000",
  5943 => x"00000000",
  5944 => x"ffffffff",
  5945 => x"00000000",
  5946 => x"00020000",
  5947 => x"00000000",
  5948 => x"00000000",
  5949 => x"00005cec",
  5950 => x"00005cec",
  5951 => x"00005cf4",
  5952 => x"00005cf4",
  5953 => x"00005cfc",
  5954 => x"00005cfc",
  5955 => x"00005d04",
  5956 => x"00005d04",
  5957 => x"00005d0c",
  5958 => x"00005d0c",
  5959 => x"00005d14",
  5960 => x"00005d14",
  5961 => x"00005d1c",
  5962 => x"00005d1c",
  5963 => x"00005d24",
  5964 => x"00005d24",
  5965 => x"00005d2c",
  5966 => x"00005d2c",
  5967 => x"00005d34",
  5968 => x"00005d34",
  5969 => x"00005d3c",
  5970 => x"00005d3c",
  5971 => x"00005d44",
  5972 => x"00005d44",
  5973 => x"00005d4c",
  5974 => x"00005d4c",
  5975 => x"00005d54",
  5976 => x"00005d54",
  5977 => x"00005d5c",
  5978 => x"00005d5c",
  5979 => x"00005d64",
  5980 => x"00005d64",
  5981 => x"00005d6c",
  5982 => x"00005d6c",
  5983 => x"00005d74",
  5984 => x"00005d74",
  5985 => x"00005d7c",
  5986 => x"00005d7c",
  5987 => x"00005d84",
  5988 => x"00005d84",
  5989 => x"00005d8c",
  5990 => x"00005d8c",
  5991 => x"00005d94",
  5992 => x"00005d94",
  5993 => x"00005d9c",
  5994 => x"00005d9c",
  5995 => x"00005da4",
  5996 => x"00005da4",
  5997 => x"00005dac",
  5998 => x"00005dac",
  5999 => x"00005db4",
  6000 => x"00005db4",
  6001 => x"00005dbc",
  6002 => x"00005dbc",
  6003 => x"00005dc4",
  6004 => x"00005dc4",
  6005 => x"00005dcc",
  6006 => x"00005dcc",
  6007 => x"00005dd4",
  6008 => x"00005dd4",
  6009 => x"00005ddc",
  6010 => x"00005ddc",
  6011 => x"00005de4",
  6012 => x"00005de4",
  6013 => x"00005dec",
  6014 => x"00005dec",
  6015 => x"00005df4",
  6016 => x"00005df4",
  6017 => x"00005dfc",
  6018 => x"00005dfc",
  6019 => x"00005e04",
  6020 => x"00005e04",
  6021 => x"00005e0c",
  6022 => x"00005e0c",
  6023 => x"00005e14",
  6024 => x"00005e14",
  6025 => x"00005e1c",
  6026 => x"00005e1c",
  6027 => x"00005e24",
  6028 => x"00005e24",
  6029 => x"00005e2c",
  6030 => x"00005e2c",
  6031 => x"00005e34",
  6032 => x"00005e34",
  6033 => x"00005e3c",
  6034 => x"00005e3c",
  6035 => x"00005e44",
  6036 => x"00005e44",
  6037 => x"00005e4c",
  6038 => x"00005e4c",
  6039 => x"00005e54",
  6040 => x"00005e54",
  6041 => x"00005e5c",
  6042 => x"00005e5c",
  6043 => x"00005e64",
  6044 => x"00005e64",
  6045 => x"00005e6c",
  6046 => x"00005e6c",
  6047 => x"00005e74",
  6048 => x"00005e74",
  6049 => x"00005e7c",
  6050 => x"00005e7c",
  6051 => x"00005e84",
  6052 => x"00005e84",
  6053 => x"00005e8c",
  6054 => x"00005e8c",
  6055 => x"00005e94",
  6056 => x"00005e94",
  6057 => x"00005e9c",
  6058 => x"00005e9c",
  6059 => x"00005ea4",
  6060 => x"00005ea4",
  6061 => x"00005eac",
  6062 => x"00005eac",
  6063 => x"00005eb4",
  6064 => x"00005eb4",
  6065 => x"00005ebc",
  6066 => x"00005ebc",
  6067 => x"00005ec4",
  6068 => x"00005ec4",
  6069 => x"00005ecc",
  6070 => x"00005ecc",
  6071 => x"00005ed4",
  6072 => x"00005ed4",
  6073 => x"00005edc",
  6074 => x"00005edc",
  6075 => x"00005ee4",
  6076 => x"00005ee4",
  6077 => x"00005eec",
  6078 => x"00005eec",
  6079 => x"00005ef4",
  6080 => x"00005ef4",
  6081 => x"00005efc",
  6082 => x"00005efc",
  6083 => x"00005f04",
  6084 => x"00005f04",
  6085 => x"00005f0c",
  6086 => x"00005f0c",
  6087 => x"00005f14",
  6088 => x"00005f14",
  6089 => x"00005f1c",
  6090 => x"00005f1c",
  6091 => x"00005f24",
  6092 => x"00005f24",
  6093 => x"00005f2c",
  6094 => x"00005f2c",
  6095 => x"00005f34",
  6096 => x"00005f34",
  6097 => x"00005f3c",
  6098 => x"00005f3c",
  6099 => x"00005f44",
  6100 => x"00005f44",
  6101 => x"00005f4c",
  6102 => x"00005f4c",
  6103 => x"00005f54",
  6104 => x"00005f54",
  6105 => x"00005f5c",
  6106 => x"00005f5c",
  6107 => x"00005f64",
  6108 => x"00005f64",
  6109 => x"00005f6c",
  6110 => x"00005f6c",
  6111 => x"00005f74",
  6112 => x"00005f74",
  6113 => x"00005f7c",
  6114 => x"00005f7c",
  6115 => x"00005f84",
  6116 => x"00005f84",
  6117 => x"00005f8c",
  6118 => x"00005f8c",
  6119 => x"00005f94",
  6120 => x"00005f94",
  6121 => x"00005f9c",
  6122 => x"00005f9c",
  6123 => x"00005fa4",
  6124 => x"00005fa4",
  6125 => x"00005fac",
  6126 => x"00005fac",
  6127 => x"00005fb4",
  6128 => x"00005fb4",
  6129 => x"00005fbc",
  6130 => x"00005fbc",
  6131 => x"00005fc4",
  6132 => x"00005fc4",
  6133 => x"00005fcc",
  6134 => x"00005fcc",
  6135 => x"00005fd4",
  6136 => x"00005fd4",
  6137 => x"00005fdc",
  6138 => x"00005fdc",
  6139 => x"00005fe4",
  6140 => x"00005fe4",
  6141 => x"00005fec",
  6142 => x"00005fec",
  6143 => x"00005ff4",
  6144 => x"00005ff4",
  6145 => x"00005ffc",
  6146 => x"00005ffc",
  6147 => x"00006004",
  6148 => x"00006004",
  6149 => x"0000600c",
  6150 => x"0000600c",
  6151 => x"00006014",
  6152 => x"00006014",
  6153 => x"0000601c",
  6154 => x"0000601c",
  6155 => x"00006024",
  6156 => x"00006024",
  6157 => x"0000602c",
  6158 => x"0000602c",
  6159 => x"00006034",
  6160 => x"00006034",
  6161 => x"0000603c",
  6162 => x"0000603c",
  6163 => x"00006044",
  6164 => x"00006044",
  6165 => x"0000604c",
  6166 => x"0000604c",
  6167 => x"00006054",
  6168 => x"00006054",
  6169 => x"0000605c",
  6170 => x"0000605c",
  6171 => x"00006064",
  6172 => x"00006064",
  6173 => x"0000606c",
  6174 => x"0000606c",
  6175 => x"00006074",
  6176 => x"00006074",
  6177 => x"0000607c",
  6178 => x"0000607c",
  6179 => x"00006084",
  6180 => x"00006084",
  6181 => x"0000608c",
  6182 => x"0000608c",
  6183 => x"00006094",
  6184 => x"00006094",
  6185 => x"0000609c",
  6186 => x"0000609c",
  6187 => x"000060a4",
  6188 => x"000060a4",
  6189 => x"000060ac",
  6190 => x"000060ac",
  6191 => x"000060b4",
  6192 => x"000060b4",
  6193 => x"000060bc",
  6194 => x"000060bc",
  6195 => x"000060c4",
  6196 => x"000060c4",
  6197 => x"000060cc",
  6198 => x"000060cc",
  6199 => x"000060d4",
  6200 => x"000060d4",
  6201 => x"000060dc",
  6202 => x"000060dc",
  6203 => x"000060e4",
  6204 => x"000060e4",
	--others => x"aaaaaaaa" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
