-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0bba",
     1 => x"c5040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"aa040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0bbc",
    73 => x"de040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0bbcc1",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80fb",
   162 => x"f0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"bcc40400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0bbd",
   169 => x"92040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0bbc",
   177 => x"fa040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80fc800c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053351",
   258 => x"bade3f71",
   259 => x"b00c833d",
   260 => x"0d04fd3d",
   261 => x"0d818be4",
   262 => x"0852f881",
   263 => x"c08e800b",
   264 => x"80fc8c08",
   265 => x"55537180",
   266 => x"2e80f738",
   267 => x"7281ff06",
   268 => x"84150c80",
   269 => x"fbe03370",
   270 => x"81ff0651",
   271 => x"5271802e",
   272 => x"80c23872",
   273 => x"9f2a7310",
   274 => x"0753818b",
   275 => x"e8337081",
   276 => x"ff065152",
   277 => x"71802ed4",
   278 => x"38800b81",
   279 => x"8be83493",
   280 => x"ee3f80fb",
   281 => x"dc335473",
   282 => x"80e23880",
   283 => x"fc8c0873",
   284 => x"81ff0684",
   285 => x"120c80fb",
   286 => x"e0337081",
   287 => x"ff065153",
   288 => x"5471c038",
   289 => x"72812a73",
   290 => x"9f2b0753",
   291 => x"ffbc3972",
   292 => x"812a739f",
   293 => x"2b075380",
   294 => x"fd51b8b5",
   295 => x"3f80fc8c",
   296 => x"08547281",
   297 => x"ff068415",
   298 => x"0c80fbe0",
   299 => x"337081ff",
   300 => x"06535471",
   301 => x"802ed838",
   302 => x"729f2a73",
   303 => x"10075380",
   304 => x"fd51b88d",
   305 => x"3f80fc8c",
   306 => x"0854d739",
   307 => x"800bb00c",
   308 => x"853d0d04",
   309 => x"fb3d0d8a",
   310 => x"51b3f53f",
   311 => x"8ad73fac",
   312 => x"87530b0b",
   313 => x"80e5ec52",
   314 => x"0b0b80e5",
   315 => x"fc518ad8",
   316 => x"3fac9e53",
   317 => x"0b0b80e6",
   318 => x"84520b0b",
   319 => x"80e6a051",
   320 => x"8ac63fb4",
   321 => x"af530b0b",
   322 => x"80e6a852",
   323 => x"0b0b80f2",
   324 => x"84518ab4",
   325 => x"3fb69753",
   326 => x"0b0b80e6",
   327 => x"c0520b0b",
   328 => x"80e6b851",
   329 => x"8aa23fb8",
   330 => x"b8530b0b",
   331 => x"80e6cc52",
   332 => x"0b0b80e6",
   333 => x"ec518a90",
   334 => x"3fb9a353",
   335 => x"0b0b80e6",
   336 => x"f4520b0b",
   337 => x"80e79851",
   338 => x"89fe3fb9",
   339 => x"dc530b0b",
   340 => x"80e7a052",
   341 => x"0b0b80e7",
   342 => x"bc5189ec",
   343 => x"3fba9253",
   344 => x"0b0b80e7",
   345 => x"c4520b0b",
   346 => x"80e7e851",
   347 => x"89da3fb8",
   348 => x"f8530b0b",
   349 => x"80e7f052",
   350 => x"0b0b80e8",
   351 => x"885189c8",
   352 => x"3fb99153",
   353 => x"0b0b80e8",
   354 => x"90520b0b",
   355 => x"80e8ac51",
   356 => x"89b63fb7",
   357 => x"8d530b0b",
   358 => x"80e8b452",
   359 => x"0b0b80e8",
   360 => x"cc5189a4",
   361 => x"3fb7e353",
   362 => x"0b0b80e8",
   363 => x"d4520b0b",
   364 => x"80e8f051",
   365 => x"89923f91",
   366 => x"a2530b0b",
   367 => x"80e8f852",
   368 => x"0b0b80e9",
   369 => x"8c518980",
   370 => x"3f90e253",
   371 => x"0b0b80e9",
   372 => x"94520b0b",
   373 => x"80e9bc51",
   374 => x"88ee3fb3",
   375 => x"90530b0b",
   376 => x"80e9c452",
   377 => x"0b0b80e9",
   378 => x"d85188dc",
   379 => x"3f889253",
   380 => x"0b0b80e9",
   381 => x"e0520b0b",
   382 => x"80e9f051",
   383 => x"88ca3fa6",
   384 => x"c0530b0b",
   385 => x"80e9f452",
   386 => x"0b0b80ea",
   387 => x"885188b8",
   388 => x"3fa9c853",
   389 => x"0b0b80ea",
   390 => x"8c520b0b",
   391 => x"80eab451",
   392 => x"88a63fb4",
   393 => x"83530b0b",
   394 => x"80eabc52",
   395 => x"0b0b80ea",
   396 => x"cc518894",
   397 => x"3f929c53",
   398 => x"0b0b80ea",
   399 => x"d0520b0b",
   400 => x"80eae851",
   401 => x"88823faa",
   402 => x"82530b0b",
   403 => x"80eaf052",
   404 => x"0b0b80ea",
   405 => x"fc5187f0",
   406 => x"3fabb153",
   407 => x"0b0b80eb",
   408 => x"80520b0b",
   409 => x"80eba851",
   410 => x"87de3faa",
   411 => x"82530b0b",
   412 => x"80ebb052",
   413 => x"0b0b80eb",
   414 => x"d05187cc",
   415 => x"3fabf753",
   416 => x"0b0b80eb",
   417 => x"d4520b0b",
   418 => x"80ebe451",
   419 => x"87ba3f90",
   420 => x"ae530b0b",
   421 => x"80f5fc52",
   422 => x"0b0b80e5",
   423 => x"e45187a8",
   424 => x"3f8e8c3f",
   425 => x"87ff3f81",
   426 => x"0b81a3d8",
   427 => x"34818be8",
   428 => x"337081ff",
   429 => x"06555573",
   430 => x"81ea38b4",
   431 => x"f63fb008",
   432 => x"81d33887",
   433 => x"ee3f80fc",
   434 => x"8c087008",
   435 => x"70842a81",
   436 => x"06515556",
   437 => x"73802e80",
   438 => x"f238f881",
   439 => x"c08e8055",
   440 => x"818be408",
   441 => x"802e8183",
   442 => x"387481ff",
   443 => x"0684170c",
   444 => x"80fbe033",
   445 => x"7081ff06",
   446 => x"51547380",
   447 => x"2e80c138",
   448 => x"749f2a75",
   449 => x"10075581",
   450 => x"8be83370",
   451 => x"81ff0651",
   452 => x"5473802e",
   453 => x"d438800b",
   454 => x"818be834",
   455 => x"8eb13f80",
   456 => x"fbdc3356",
   457 => x"75a53880",
   458 => x"fc8c0875",
   459 => x"81ff0684",
   460 => x"120c80fb",
   461 => x"e0337081",
   462 => x"ff065155",
   463 => x"5673c138",
   464 => x"74812a75",
   465 => x"9f2b0755",
   466 => x"ffbd3981",
   467 => x"a3d83355",
   468 => x"74feda38",
   469 => x"873d0d04",
   470 => x"74812a75",
   471 => x"9f2b0755",
   472 => x"80fd51b2",
   473 => x"ec3f80fc",
   474 => x"8c085674",
   475 => x"81ff0684",
   476 => x"170c80fb",
   477 => x"e0337081",
   478 => x"ff065754",
   479 => x"75802ed8",
   480 => x"38749f2a",
   481 => x"75100755",
   482 => x"80fd51b2",
   483 => x"c43f80fc",
   484 => x"8c0856d7",
   485 => x"39b3af3f",
   486 => x"b00881ff",
   487 => x"06518781",
   488 => x"3ffea039",
   489 => x"800b818b",
   490 => x"e8348da3",
   491 => x"3fb3843f",
   492 => x"b008802e",
   493 => x"fe8d38dd",
   494 => x"39803d0d",
   495 => x"0b0b80eb",
   496 => x"ec51aea6",
   497 => x"3f8c51ae",
   498 => x"873f0b0b",
   499 => x"80ebf051",
   500 => x"ae983f81",
   501 => x"8be40880",
   502 => x"2e8e380b",
   503 => x"0b80ec88",
   504 => x"51ae873f",
   505 => x"823d0d04",
   506 => x"0b0b80ec",
   507 => x"9451adfa",
   508 => x"3f810a51",
   509 => x"adf43f0b",
   510 => x"0b80eca8",
   511 => x"51adeb3f",
   512 => x"0b0b80ec",
   513 => x"d051ade2",
   514 => x"3f80e451",
   515 => x"afa63f0b",
   516 => x"0b80ece4",
   517 => x"51add33f",
   518 => x"0b0b80ec",
   519 => x"ec51adca",
   520 => x"3f0b0b80",
   521 => x"ecf851ad",
   522 => x"c13f823d",
   523 => x"0d04ff89",
   524 => x"3f8afc3f",
   525 => x"800bb00c",
   526 => x"04fe3d0d",
   527 => x"80fc9008",
   528 => x"98110870",
   529 => x"842a7081",
   530 => x"06515353",
   531 => x"5370802e",
   532 => x"8d3871ef",
   533 => x"0698140c",
   534 => x"810b818b",
   535 => x"e834843d",
   536 => x"0d04f93d",
   537 => x"0d815189",
   538 => x"943fb008",
   539 => x"55825189",
   540 => x"8c3f74b0",
   541 => x"08075399",
   542 => x"cc57fce2",
   543 => x"97f68058",
   544 => x"72802e90",
   545 => x"38747554",
   546 => x"57805480",
   547 => x"770774b0",
   548 => x"08075957",
   549 => x"76517752",
   550 => x"9bfa3f72",
   551 => x"b00c893d",
   552 => x"0d04fb3d",
   553 => x"0d815187",
   554 => x"a23fb008",
   555 => x"56815382",
   556 => x"528051a5",
   557 => x"a83f80fb",
   558 => x"ec085589",
   559 => x"750c80fc",
   560 => x"8c088411",
   561 => x"0870810a",
   562 => x"0784130c",
   563 => x"55557551",
   564 => x"afd93f80",
   565 => x"fc8c0884",
   566 => x"110870fe",
   567 => x"0a068413",
   568 => x"0c555581",
   569 => x"53825280",
   570 => x"51a4f23f",
   571 => x"80fbec08",
   572 => x"5589750c",
   573 => x"80fc8c08",
   574 => x"84110870",
   575 => x"810a0784",
   576 => x"130c5555",
   577 => x"7551afa3",
   578 => x"3f80fc8c",
   579 => x"08841108",
   580 => x"70fe0a06",
   581 => x"84130c55",
   582 => x"55ff9239",
   583 => x"fe3d0d81",
   584 => x"5186a83f",
   585 => x"80fc8c08",
   586 => x"84110870",
   587 => x"810a0784",
   588 => x"130c5353",
   589 => x"b00851ae",
   590 => x"f23f80fc",
   591 => x"8c088411",
   592 => x"0870fe0a",
   593 => x"06708414",
   594 => x"0cb00c53",
   595 => x"53843d0d",
   596 => x"04fc3d0d",
   597 => x"80fc8c08",
   598 => x"7008810a",
   599 => x"06818be4",
   600 => x"0c54af91",
   601 => x"3fafb53f",
   602 => x"8ac53f93",
   603 => x"8c3f80fc",
   604 => x"90089811",
   605 => x"08708807",
   606 => x"98130c55",
   607 => x"55818be4",
   608 => x"0880d538",
   609 => x"88800b81",
   610 => x"a4b40cfc",
   611 => x"ac3f818b",
   612 => x"e408802e",
   613 => x"80d33881",
   614 => x"53825280",
   615 => x"51a3be3f",
   616 => x"80fbec08",
   617 => x"5589750c",
   618 => x"80fc8c08",
   619 => x"84110870",
   620 => x"810a0784",
   621 => x"130c5555",
   622 => x"8051adef",
   623 => x"3f80fc8c",
   624 => x"08841108",
   625 => x"70fe0a06",
   626 => x"84130c55",
   627 => x"5580fbec",
   628 => x"08558075",
   629 => x"0cb0ab3f",
   630 => x"bdba0b81",
   631 => x"a4b40cfb",
   632 => x"d83f818b",
   633 => x"e408ffaf",
   634 => x"3880c2e8",
   635 => x"0b81a4b4",
   636 => x"0cf5e13f",
   637 => x"81538252",
   638 => x"8051a2e1",
   639 => x"3f80fbec",
   640 => x"08558975",
   641 => x"0c80fc8c",
   642 => x"08841108",
   643 => x"70810a07",
   644 => x"84130c55",
   645 => x"558051ad",
   646 => x"923f80fc",
   647 => x"8c088411",
   648 => x"0870fe0a",
   649 => x"0684130c",
   650 => x"555580fb",
   651 => x"ec085580",
   652 => x"750cafce",
   653 => x"3f800b81",
   654 => x"a3d03480",
   655 => x"0b81a3cc",
   656 => x"34800b81",
   657 => x"a3d40c04",
   658 => x"fc3d0d81",
   659 => x"a3cc3353",
   660 => x"72a72680",
   661 => x"c5387652",
   662 => x"72101010",
   663 => x"73100581",
   664 => x"8bec0551",
   665 => x"b4b73f77",
   666 => x"5281a3cc",
   667 => x"33709029",
   668 => x"71317010",
   669 => x"10818efc",
   670 => x"05535654",
   671 => x"b49f3f81",
   672 => x"a3cc3370",
   673 => x"101081a1",
   674 => x"dc057a71",
   675 => x"0c548105",
   676 => x"537281a3",
   677 => x"cc34863d",
   678 => x"0d0480ed",
   679 => x"8051a8ca",
   680 => x"3f863d0d",
   681 => x"04803d0d",
   682 => x"80ed9c51",
   683 => x"a8bc3f82",
   684 => x"3d0d04fe",
   685 => x"3d0d81a3",
   686 => x"d4085372",
   687 => x"8538843d",
   688 => x"0d04722d",
   689 => x"b0085380",
   690 => x"0b81a3d4",
   691 => x"0cb0088c",
   692 => x"3880ed9c",
   693 => x"51a8933f",
   694 => x"843d0d04",
   695 => x"80f8cc51",
   696 => x"a8883f72",
   697 => x"83ffff26",
   698 => x"aa3881ff",
   699 => x"73279638",
   700 => x"72529051",
   701 => x"a8973f8a",
   702 => x"51a7d53f",
   703 => x"80ed9c51",
   704 => x"a7e83fd4",
   705 => x"39725288",
   706 => x"51a8823f",
   707 => x"8a51a7c0",
   708 => x"3fea3972",
   709 => x"52a051a7",
   710 => x"f43f8a51",
   711 => x"a7b23fdc",
   712 => x"39fa3d0d",
   713 => x"02a30533",
   714 => x"56758d2e",
   715 => x"80f43875",
   716 => x"88327030",
   717 => x"7780ff32",
   718 => x"70307280",
   719 => x"25718025",
   720 => x"07545156",
   721 => x"58557495",
   722 => x"389f7627",
   723 => x"8c3881a3",
   724 => x"d0335580",
   725 => x"ce7527ae",
   726 => x"38883d0d",
   727 => x"0481a3d0",
   728 => x"33567580",
   729 => x"2ef33888",
   730 => x"51a6e53f",
   731 => x"a051a6e0",
   732 => x"3f8851a6",
   733 => x"db3f81a3",
   734 => x"d033ff05",
   735 => x"577681a3",
   736 => x"d034883d",
   737 => x"0d047551",
   738 => x"a6c63f81",
   739 => x"a3d03381",
   740 => x"11555773",
   741 => x"81a3d034",
   742 => x"7581a2fc",
   743 => x"1834883d",
   744 => x"0d048a51",
   745 => x"a6aa3f81",
   746 => x"a3d03381",
   747 => x"11565474",
   748 => x"81a3d034",
   749 => x"800b81a2",
   750 => x"fc153480",
   751 => x"56800b81",
   752 => x"a2fc1733",
   753 => x"565474a0",
   754 => x"2e833881",
   755 => x"5474802e",
   756 => x"90387380",
   757 => x"2e8b3881",
   758 => x"167081ff",
   759 => x"065757dd",
   760 => x"3975802e",
   761 => x"bf38800b",
   762 => x"81a3cc33",
   763 => x"55557474",
   764 => x"27ab3873",
   765 => x"57741010",
   766 => x"10751005",
   767 => x"765481a2",
   768 => x"fc53818b",
   769 => x"ec0551b2",
   770 => x"e03fb008",
   771 => x"802ea638",
   772 => x"81157081",
   773 => x"ff065654",
   774 => x"767526d9",
   775 => x"3880eda0",
   776 => x"51a5c73f",
   777 => x"80ed9c51",
   778 => x"a5c03f80",
   779 => x"0b81a3d0",
   780 => x"34883d0d",
   781 => x"04741010",
   782 => x"81a1dc05",
   783 => x"700881a3",
   784 => x"d40c5680",
   785 => x"0b81a3d0",
   786 => x"34e739f7",
   787 => x"3d0d02af",
   788 => x"05335980",
   789 => x"0b81a2fc",
   790 => x"3381a2fc",
   791 => x"59555673",
   792 => x"a02e0981",
   793 => x"06963881",
   794 => x"167081ff",
   795 => x"0681a2fc",
   796 => x"11703353",
   797 => x"59575473",
   798 => x"a02eec38",
   799 => x"80587779",
   800 => x"2780ea38",
   801 => x"80773356",
   802 => x"5474742e",
   803 => x"83388154",
   804 => x"74a02e9a",
   805 => x"387380c5",
   806 => x"3874a02e",
   807 => x"91388118",
   808 => x"7081ff06",
   809 => x"59557878",
   810 => x"26da3880",
   811 => x"c0398116",
   812 => x"7081ff06",
   813 => x"81a2fc11",
   814 => x"70335752",
   815 => x"575773a0",
   816 => x"2e098106",
   817 => x"d9388116",
   818 => x"7081ff06",
   819 => x"81a2fc11",
   820 => x"70335752",
   821 => x"575773a0",
   822 => x"2ed438c2",
   823 => x"39811670",
   824 => x"81ff0681",
   825 => x"a2fc1159",
   826 => x"5755ff98",
   827 => x"3980538b",
   828 => x"3dfc0552",
   829 => x"7651b5b6",
   830 => x"3f8b3d0d",
   831 => x"04f73d0d",
   832 => x"02af0533",
   833 => x"59800b81",
   834 => x"a2fc3381",
   835 => x"a2fc5955",
   836 => x"5673a02e",
   837 => x"09810696",
   838 => x"38811670",
   839 => x"81ff0681",
   840 => x"a2fc1170",
   841 => x"33535957",
   842 => x"5473a02e",
   843 => x"ec388058",
   844 => x"77792780",
   845 => x"ea388077",
   846 => x"33565474",
   847 => x"742e8338",
   848 => x"815474a0",
   849 => x"2e9a3873",
   850 => x"80c53874",
   851 => x"a02e9138",
   852 => x"81187081",
   853 => x"ff065955",
   854 => x"787826da",
   855 => x"3880c039",
   856 => x"81167081",
   857 => x"ff0681a2",
   858 => x"fc117033",
   859 => x"57525757",
   860 => x"73a02e09",
   861 => x"8106d938",
   862 => x"81167081",
   863 => x"ff0681a2",
   864 => x"fc117033",
   865 => x"57525757",
   866 => x"73a02ed4",
   867 => x"38c23981",
   868 => x"167081ff",
   869 => x"0681a2fc",
   870 => x"11595755",
   871 => x"ff983990",
   872 => x"538b3dfc",
   873 => x"05527651",
   874 => x"b7a13f8b",
   875 => x"3d0d04fc",
   876 => x"3d0d8a51",
   877 => x"a29a3f80",
   878 => x"edb451a2",
   879 => x"ad3f800b",
   880 => x"81a3cc33",
   881 => x"53537272",
   882 => x"2780f538",
   883 => x"72101010",
   884 => x"73100581",
   885 => x"8bec0570",
   886 => x"5254a28e",
   887 => x"3f72842b",
   888 => x"70743182",
   889 => x"2b818efc",
   890 => x"11335153",
   891 => x"5571802e",
   892 => x"b7387351",
   893 => x"ae943fb0",
   894 => x"0881ff06",
   895 => x"52718926",
   896 => x"9338a051",
   897 => x"a1ca3f81",
   898 => x"127081ff",
   899 => x"06535489",
   900 => x"7227ef38",
   901 => x"80edcc51",
   902 => x"a1d03f74",
   903 => x"7331822b",
   904 => x"818efc05",
   905 => x"51a1c33f",
   906 => x"8a51a1a4",
   907 => x"3f811370",
   908 => x"81ff0681",
   909 => x"a3cc3354",
   910 => x"54557173",
   911 => x"26ff8d38",
   912 => x"8a51a18c",
   913 => x"3f81a3cc",
   914 => x"33b00c86",
   915 => x"3d0d04fe",
   916 => x"3d0d81a4",
   917 => x"ac22ff05",
   918 => x"517081a4",
   919 => x"ac237083",
   920 => x"ffff0651",
   921 => x"7080c438",
   922 => x"81a4b033",
   923 => x"517081ff",
   924 => x"2eb93870",
   925 => x"10101081",
   926 => x"a3dc0552",
   927 => x"713381a4",
   928 => x"b034fe72",
   929 => x"3481a4b0",
   930 => x"33701010",
   931 => x"1081a3dc",
   932 => x"05525382",
   933 => x"112281a4",
   934 => x"ac238412",
   935 => x"0853722d",
   936 => x"81a4ac22",
   937 => x"5170802e",
   938 => x"ffbe3884",
   939 => x"3d0d04ff",
   940 => x"3d0d8a52",
   941 => x"71101010",
   942 => x"81a3d405",
   943 => x"51fe7134",
   944 => x"ff127081",
   945 => x"ff065351",
   946 => x"71ea38ff",
   947 => x"0b81a4b0",
   948 => x"34833d0d",
   949 => x"04fe3d0d",
   950 => x"02930533",
   951 => x"02840597",
   952 => x"05335452",
   953 => x"71842e80",
   954 => x"d1387184",
   955 => x"24913871",
   956 => x"812eac38",
   957 => x"80edd051",
   958 => x"9ff03f84",
   959 => x"3d0d0471",
   960 => x"80d52e09",
   961 => x"8106ed38",
   962 => x"80eddc51",
   963 => x"9fdc3f72",
   964 => x"8c26b338",
   965 => x"72101080",
   966 => x"f2d00552",
   967 => x"71080480",
   968 => x"ede8519f",
   969 => x"c53ffa13",
   970 => x"527180db",
   971 => x"26983871",
   972 => x"101080f3",
   973 => x"84055271",
   974 => x"080480ed",
   975 => x"f4519faa",
   976 => x"3f728f2e",
   977 => x"8c3880ee",
   978 => x"80519f9e",
   979 => x"3f843d0d",
   980 => x"0480ee90",
   981 => x"519f933f",
   982 => x"843d0d04",
   983 => x"80eea851",
   984 => x"9f883f84",
   985 => x"3d0d0480",
   986 => x"eeb8519e",
   987 => x"fd3f843d",
   988 => x"0d0480ee",
   989 => x"d0519ef2",
   990 => x"3f843d0d",
   991 => x"0480eee0",
   992 => x"519ee73f",
   993 => x"843d0d04",
   994 => x"80ef8051",
   995 => x"9edc3f84",
   996 => x"3d0d0480",
   997 => x"ef9c519e",
   998 => x"d13f843d",
   999 => x"0d0480ef",
  1000 => x"b8519ec6",
  1001 => x"3f843d0d",
  1002 => x"0480efcc",
  1003 => x"519ebb3f",
  1004 => x"843d0d04",
  1005 => x"80efe851",
  1006 => x"9eb03f84",
  1007 => x"3d0d0480",
  1008 => x"eff8519e",
  1009 => x"a53f843d",
  1010 => x"0d0480f0",
  1011 => x"88519e9a",
  1012 => x"3f843d0d",
  1013 => x"0480f0a8",
  1014 => x"519e8f3f",
  1015 => x"843d0d04",
  1016 => x"80f0bc51",
  1017 => x"9e843f84",
  1018 => x"3d0d0480",
  1019 => x"f0d8519d",
  1020 => x"f93f843d",
  1021 => x"0d0480f0",
  1022 => x"f0519dee",
  1023 => x"3f843d0d",
  1024 => x"0480f184",
  1025 => x"519de33f",
  1026 => x"843d0d04",
  1027 => x"80f19451",
  1028 => x"9dd83f84",
  1029 => x"3d0d0480",
  1030 => x"f1a8519d",
  1031 => x"cd3f843d",
  1032 => x"0d0480f1",
  1033 => x"b8519dc2",
  1034 => x"3f843d0d",
  1035 => x"0480f1d0",
  1036 => x"519db73f",
  1037 => x"843d0d04",
  1038 => x"80f1e451",
  1039 => x"9dac3f84",
  1040 => x"3d0d0480",
  1041 => x"f1f4519d",
  1042 => x"a13f843d",
  1043 => x"0d04f73d",
  1044 => x"0d02b305",
  1045 => x"337c7008",
  1046 => x"c0808006",
  1047 => x"59545a80",
  1048 => x"5675832b",
  1049 => x"7707bfe0",
  1050 => x"80077070",
  1051 => x"84055208",
  1052 => x"71088c2a",
  1053 => x"bffe8006",
  1054 => x"79077198",
  1055 => x"2a728c2a",
  1056 => x"9fff0673",
  1057 => x"852a708f",
  1058 => x"06759f06",
  1059 => x"5651585d",
  1060 => x"58525558",
  1061 => x"748d3881",
  1062 => x"16568f76",
  1063 => x"27c3388b",
  1064 => x"3d0d0480",
  1065 => x"f28c519c",
  1066 => x"c13f7551",
  1067 => x"9e863f84",
  1068 => x"52b00851",
  1069 => x"9fc73f80",
  1070 => x"f298519c",
  1071 => x"ad3f7452",
  1072 => x"88519cc9",
  1073 => x"3f8452b0",
  1074 => x"08519fb1",
  1075 => x"3f80f2a0",
  1076 => x"519c973f",
  1077 => x"78529051",
  1078 => x"9cb33f86",
  1079 => x"52b00851",
  1080 => x"9f9b3f80",
  1081 => x"f2a8519c",
  1082 => x"813f7251",
  1083 => x"9dc63f84",
  1084 => x"52b00851",
  1085 => x"9f873f80",
  1086 => x"f2b0519b",
  1087 => x"ed3f7351",
  1088 => x"9db23f84",
  1089 => x"52b00851",
  1090 => x"9ef33f80",
  1091 => x"f2b8519b",
  1092 => x"d93f7752",
  1093 => x"a0519bf5",
  1094 => x"3f8a52b0",
  1095 => x"08519edd",
  1096 => x"3f799238",
  1097 => x"8a519ba8",
  1098 => x"3f811656",
  1099 => x"8f7627fe",
  1100 => x"b038feeb",
  1101 => x"397881ff",
  1102 => x"06527451",
  1103 => x"fb973f8a",
  1104 => x"519b8d3f",
  1105 => x"e439f83d",
  1106 => x"0d02ab05",
  1107 => x"33598056",
  1108 => x"75852be0",
  1109 => x"9011e080",
  1110 => x"12087098",
  1111 => x"2a718c2a",
  1112 => x"9fff0672",
  1113 => x"852a708f",
  1114 => x"06749f06",
  1115 => x"5551585b",
  1116 => x"53565955",
  1117 => x"74802e81",
  1118 => x"a13875bf",
  1119 => x"2681a938",
  1120 => x"80f2c051",
  1121 => x"9ae43f75",
  1122 => x"519ca93f",
  1123 => x"8652b008",
  1124 => x"519dea3f",
  1125 => x"80f29851",
  1126 => x"9ad03f74",
  1127 => x"5288519a",
  1128 => x"ec3f8452",
  1129 => x"b008519d",
  1130 => x"d43f80f2",
  1131 => x"a0519aba",
  1132 => x"3f765290",
  1133 => x"519ad63f",
  1134 => x"8652b008",
  1135 => x"519dbe3f",
  1136 => x"80f2a851",
  1137 => x"9aa43f72",
  1138 => x"519be93f",
  1139 => x"8452b008",
  1140 => x"519daa3f",
  1141 => x"80f2b051",
  1142 => x"9a903f73",
  1143 => x"519bd53f",
  1144 => x"8452b008",
  1145 => x"519d963f",
  1146 => x"80f2b851",
  1147 => x"99fc3f77",
  1148 => x"08c08080",
  1149 => x"0652a051",
  1150 => x"9a933f8a",
  1151 => x"52b00851",
  1152 => x"9cfb3f78",
  1153 => x"81ac388a",
  1154 => x"5199c53f",
  1155 => x"80537481",
  1156 => x"2e81d938",
  1157 => x"76862e81",
  1158 => x"b5388116",
  1159 => x"5680ff76",
  1160 => x"27fead38",
  1161 => x"8a3d0d04",
  1162 => x"80f2c851",
  1163 => x"99bc3fc0",
  1164 => x"16519b80",
  1165 => x"3f8652b0",
  1166 => x"08519cc1",
  1167 => x"3f80f298",
  1168 => x"5199a73f",
  1169 => x"74528851",
  1170 => x"99c33f84",
  1171 => x"52b00851",
  1172 => x"9cab3f80",
  1173 => x"f2a05199",
  1174 => x"913f7652",
  1175 => x"905199ad",
  1176 => x"3f8652b0",
  1177 => x"08519c95",
  1178 => x"3f80f2a8",
  1179 => x"5198fb3f",
  1180 => x"72519ac0",
  1181 => x"3f8452b0",
  1182 => x"08519c81",
  1183 => x"3f80f2b0",
  1184 => x"5198e73f",
  1185 => x"73519aac",
  1186 => x"3f8452b0",
  1187 => x"08519bed",
  1188 => x"3f80f2b8",
  1189 => x"5198d33f",
  1190 => x"7708c080",
  1191 => x"800652a0",
  1192 => x"5198ea3f",
  1193 => x"8a52b008",
  1194 => x"519bd23f",
  1195 => x"78802efe",
  1196 => x"d6387681",
  1197 => x"ff065274",
  1198 => x"51f89a3f",
  1199 => x"8a519890",
  1200 => x"3f805374",
  1201 => x"812e0981",
  1202 => x"06fec938",
  1203 => x"9f397281",
  1204 => x"06577680",
  1205 => x"2efec338",
  1206 => x"78527751",
  1207 => x"faf03f81",
  1208 => x"165680ff",
  1209 => x"7627fce8",
  1210 => x"38feb939",
  1211 => x"74537686",
  1212 => x"2e098106",
  1213 => x"fea438d6",
  1214 => x"39803d0d",
  1215 => x"80fc8808",
  1216 => x"51b1710c",
  1217 => x"81800b84",
  1218 => x"120c823d",
  1219 => x"0d04fe3d",
  1220 => x"0d740284",
  1221 => x"05970533",
  1222 => x"0288059b",
  1223 => x"05338813",
  1224 => x"0c8c120c",
  1225 => x"538c1308",
  1226 => x"70812a81",
  1227 => x"06515271",
  1228 => x"f4388c13",
  1229 => x"087081ff",
  1230 => x"06b00c51",
  1231 => x"843d0d04",
  1232 => x"fb3d0d80",
  1233 => x"0b80f5f4",
  1234 => x"5256979e",
  1235 => x"3f755574",
  1236 => x"105381d0",
  1237 => x"5280fc88",
  1238 => x"0851ffb2",
  1239 => x"3fb00887",
  1240 => x"2a708106",
  1241 => x"51547380",
  1242 => x"2e993881",
  1243 => x"157081ff",
  1244 => x"0670982b",
  1245 => x"52565473",
  1246 => x"8025d438",
  1247 => x"75b00c87",
  1248 => x"3d0d0480",
  1249 => x"f6805196",
  1250 => x"e13f7452",
  1251 => x"885196fd",
  1252 => x"3f80f68c",
  1253 => x"5196d33f",
  1254 => x"81167083",
  1255 => x"ffff0681",
  1256 => x"177081ff",
  1257 => x"0670982b",
  1258 => x"52585257",
  1259 => x"54738025",
  1260 => x"ff9d38c8",
  1261 => x"39f33d0d",
  1262 => x"7f028405",
  1263 => x"80c30533",
  1264 => x"02880580",
  1265 => x"c6052280",
  1266 => x"f69c545b",
  1267 => x"5558969a",
  1268 => x"3f785197",
  1269 => x"df3f80f6",
  1270 => x"a851968e",
  1271 => x"3f735288",
  1272 => x"5196aa3f",
  1273 => x"80ebec51",
  1274 => x"96803f80",
  1275 => x"57767927",
  1276 => x"81913873",
  1277 => x"108e3d5c",
  1278 => x"5a795381",
  1279 => x"90527751",
  1280 => x"fe8c3f76",
  1281 => x"882a5390",
  1282 => x"527751fe",
  1283 => x"813f7681",
  1284 => x"ff065390",
  1285 => x"527751fd",
  1286 => x"f53f811a",
  1287 => x"53819052",
  1288 => x"7751fdea",
  1289 => x"3f805380",
  1290 => x"e0527751",
  1291 => x"fde03fb0",
  1292 => x"08872a81",
  1293 => x"0654738a",
  1294 => x"38881808",
  1295 => x"7081ff06",
  1296 => x"5d567b81",
  1297 => x"ff0680f8",
  1298 => x"cc525695",
  1299 => x"9d3f7552",
  1300 => x"885195b9",
  1301 => x"3f80edfc",
  1302 => x"51958f3f",
  1303 => x"e0165480",
  1304 => x"df7427b6",
  1305 => x"38768706",
  1306 => x"701c5755",
  1307 => x"a0763474",
  1308 => x"872eb938",
  1309 => x"81177083",
  1310 => x"ffff0658",
  1311 => x"55787726",
  1312 => x"fef73880",
  1313 => x"e00b8c19",
  1314 => x"0c8c1808",
  1315 => x"70812a81",
  1316 => x"06585a76",
  1317 => x"f4388f3d",
  1318 => x"0d047687",
  1319 => x"06701c55",
  1320 => x"55757434",
  1321 => x"74872e09",
  1322 => x"8106c938",
  1323 => x"7a5194ba",
  1324 => x"3f8a5194",
  1325 => x"9b3f8117",
  1326 => x"7083ffff",
  1327 => x"06585578",
  1328 => x"7726feb5",
  1329 => x"38ffbc39",
  1330 => x"fb3d0d81",
  1331 => x"51eefc3f",
  1332 => x"8251f0a9",
  1333 => x"3fb00881",
  1334 => x"ff065683",
  1335 => x"51eeec3f",
  1336 => x"b00883ff",
  1337 => x"ff0680fc",
  1338 => x"88085654",
  1339 => x"73843881",
  1340 => x"80547353",
  1341 => x"75527451",
  1342 => x"fdbb3f73",
  1343 => x"b00c873d",
  1344 => x"0d04fb3d",
  1345 => x"0d8151ef",
  1346 => x"f43fb008",
  1347 => x"538251ef",
  1348 => x"ec3fb008",
  1349 => x"56b00883",
  1350 => x"38905672",
  1351 => x"fc065575",
  1352 => x"812e80f1",
  1353 => x"38805473",
  1354 => x"7627aa38",
  1355 => x"73830653",
  1356 => x"72802eae",
  1357 => x"3880f8cc",
  1358 => x"5193af3f",
  1359 => x"74708405",
  1360 => x"560852a0",
  1361 => x"5193c63f",
  1362 => x"a0519384",
  1363 => x"3f811454",
  1364 => x"757426d8",
  1365 => x"388a5192",
  1366 => x"f73f800b",
  1367 => x"b00c873d",
  1368 => x"0d0480f6",
  1369 => x"c4519382",
  1370 => x"3f7452a0",
  1371 => x"51939e3f",
  1372 => x"80f88c51",
  1373 => x"92f43f80",
  1374 => x"f8cc5192",
  1375 => x"ed3f7470",
  1376 => x"84055608",
  1377 => x"52a05193",
  1378 => x"843fa051",
  1379 => x"92c23f81",
  1380 => x"1454ffbc",
  1381 => x"3980f8cc",
  1382 => x"5192cf3f",
  1383 => x"740852a0",
  1384 => x"5192ea3f",
  1385 => x"8a5192a8",
  1386 => x"3f800bb0",
  1387 => x"0c873d0d",
  1388 => x"04fc3d0d",
  1389 => x"8151eec5",
  1390 => x"3fb00852",
  1391 => x"8251ed8b",
  1392 => x"3fb00881",
  1393 => x"ff067256",
  1394 => x"53835472",
  1395 => x"802ea138",
  1396 => x"7351eea9",
  1397 => x"3f811470",
  1398 => x"81ff06ff",
  1399 => x"157081ff",
  1400 => x"06b00879",
  1401 => x"7084055b",
  1402 => x"0c565255",
  1403 => x"5272e138",
  1404 => x"72b00c86",
  1405 => x"3d0d0480",
  1406 => x"3d0d8c51",
  1407 => x"91d23f80",
  1408 => x"0bb00c82",
  1409 => x"3d0d0480",
  1410 => x"3d0d80fc",
  1411 => x"980851f8",
  1412 => x"bb9586a1",
  1413 => x"710c810b",
  1414 => x"b00c823d",
  1415 => x"0d04803d",
  1416 => x"0d8151ec",
  1417 => x"a63fb008",
  1418 => x"81ff0651",
  1419 => x"f6983f80",
  1420 => x"0bb00c82",
  1421 => x"3d0d04ff",
  1422 => x"3d0d80fb",
  1423 => x"e408a011",
  1424 => x"087080ff",
  1425 => x"0a06a013",
  1426 => x"0c5252bb",
  1427 => x"c880800b",
  1428 => x"a0130c83",
  1429 => x"3d0d04ff",
  1430 => x"3d0d028f",
  1431 => x"05337098",
  1432 => x"2b80fbe4",
  1433 => x"0852b012",
  1434 => x"0c51833d",
  1435 => x"0d04ff3d",
  1436 => x"0d80fbe4",
  1437 => x"0852a412",
  1438 => x"0870892a",
  1439 => x"70810651",
  1440 => x"51517080",
  1441 => x"2ef038b4",
  1442 => x"12087090",
  1443 => x"2ab00c51",
  1444 => x"833d0d04",
  1445 => x"f83d0d7a",
  1446 => x"7c5755ff",
  1447 => x"9a3f80fc",
  1448 => x"8c088411",
  1449 => x"08828080",
  1450 => x"0784120c",
  1451 => x"841108fd",
  1452 => x"ffff0684",
  1453 => x"120c8411",
  1454 => x"08818080",
  1455 => x"0784120c",
  1456 => x"841108fe",
  1457 => x"ffff0684",
  1458 => x"120c5390",
  1459 => x"0b893d34",
  1460 => x"94028405",
  1461 => x"9d053480",
  1462 => x"0284059e",
  1463 => x"053480e1",
  1464 => x"0284059f",
  1465 => x"0534883d",
  1466 => x"80fbe408",
  1467 => x"5457a413",
  1468 => x"0870882a",
  1469 => x"81065152",
  1470 => x"71802ef2",
  1471 => x"388751fe",
  1472 => x"d63f800b",
  1473 => x"80f6cf33",
  1474 => x"53537272",
  1475 => x"27993871",
  1476 => x"54761370",
  1477 => x"335252fe",
  1478 => x"be3f8113",
  1479 => x"7081ff06",
  1480 => x"54527373",
  1481 => x"26eb38fe",
  1482 => x"c53f800b",
  1483 => x"80f6cf33",
  1484 => x"53537272",
  1485 => x"27933871",
  1486 => x"54feb33f",
  1487 => x"81137081",
  1488 => x"ff065452",
  1489 => x"737326f1",
  1490 => x"3874882a",
  1491 => x"5473893d",
  1492 => x"34740284",
  1493 => x"059d0534",
  1494 => x"74882b76",
  1495 => x"982a0752",
  1496 => x"71028405",
  1497 => x"9e053474",
  1498 => x"902b7690",
  1499 => x"2a075473",
  1500 => x"0284059f",
  1501 => x"05347498",
  1502 => x"2b76882a",
  1503 => x"0753728a",
  1504 => x"3d347502",
  1505 => x"8405a105",
  1506 => x"3480fbe4",
  1507 => x"0853a413",
  1508 => x"0870882a",
  1509 => x"81065652",
  1510 => x"74802ef2",
  1511 => x"388251fd",
  1512 => x"b63f800b",
  1513 => x"80f6ca33",
  1514 => x"53537272",
  1515 => x"27993871",
  1516 => x"54761370",
  1517 => x"335256fd",
  1518 => x"9e3f8113",
  1519 => x"7081ff06",
  1520 => x"54557373",
  1521 => x"26eb38fd",
  1522 => x"a53f800b",
  1523 => x"80f6ca33",
  1524 => x"53537272",
  1525 => x"27933871",
  1526 => x"54fd933f",
  1527 => x"81137081",
  1528 => x"ff065452",
  1529 => x"737326f1",
  1530 => x"388a0b89",
  1531 => x"3d34ff8c",
  1532 => x"0284059d",
  1533 => x"053480fb",
  1534 => x"e40853a4",
  1535 => x"13087088",
  1536 => x"2a810655",
  1537 => x"5673802e",
  1538 => x"f2388851",
  1539 => x"fcc93f80",
  1540 => x"0b80f6d0",
  1541 => x"33535372",
  1542 => x"72279938",
  1543 => x"71547613",
  1544 => x"70335255",
  1545 => x"fcb13f81",
  1546 => x"137081ff",
  1547 => x"06545273",
  1548 => x"7326eb38",
  1549 => x"fcb83f80",
  1550 => x"0b80f6d0",
  1551 => x"33535372",
  1552 => x"72279338",
  1553 => x"7154fca6",
  1554 => x"3f811370",
  1555 => x"81ff0654",
  1556 => x"56737326",
  1557 => x"f1388a0b",
  1558 => x"893d34ff",
  1559 => x"8c028405",
  1560 => x"9d053480",
  1561 => x"fbe40853",
  1562 => x"a4130870",
  1563 => x"882a8106",
  1564 => x"55557380",
  1565 => x"2ef23889",
  1566 => x"51fbdc3f",
  1567 => x"800b80f6",
  1568 => x"d1335353",
  1569 => x"72722799",
  1570 => x"38715476",
  1571 => x"13703352",
  1572 => x"52fbc43f",
  1573 => x"81137081",
  1574 => x"ff065456",
  1575 => x"737326eb",
  1576 => x"38fbcb3f",
  1577 => x"800b80f6",
  1578 => x"d1335353",
  1579 => x"72722793",
  1580 => x"387154fb",
  1581 => x"b93f8113",
  1582 => x"7081ff06",
  1583 => x"54577373",
  1584 => x"26f13880",
  1585 => x"fc8c0884",
  1586 => x"110880c0",
  1587 => x"80078412",
  1588 => x"0c841108",
  1589 => x"ffbfff06",
  1590 => x"84120c54",
  1591 => x"800bb00c",
  1592 => x"8a3d0d04",
  1593 => x"f83d0d02",
  1594 => x"ab053389",
  1595 => x"3d80fbe4",
  1596 => x"08565856",
  1597 => x"a4140870",
  1598 => x"882a8106",
  1599 => x"51537280",
  1600 => x"2ef23875",
  1601 => x"81800751",
  1602 => x"facd3f80",
  1603 => x"0b80f6c8",
  1604 => x"17335454",
  1605 => x"73732795",
  1606 => x"38725580",
  1607 => x"51fab83f",
  1608 => x"81147081",
  1609 => x"ff065553",
  1610 => x"747426ef",
  1611 => x"38fabf3f",
  1612 => x"800b80f6",
  1613 => x"c8173370",
  1614 => x"81ff0655",
  1615 => x"57547373",
  1616 => x"279a3872",
  1617 => x"55761453",
  1618 => x"faa43fb0",
  1619 => x"08733481",
  1620 => x"147081ff",
  1621 => x"06555374",
  1622 => x"7426ea38",
  1623 => x"7581ff06",
  1624 => x"80f8cc52",
  1625 => x"558b833f",
  1626 => x"80547375",
  1627 => x"27993873",
  1628 => x"17703353",
  1629 => x"5388518b",
  1630 => x"943f8114",
  1631 => x"7081ff06",
  1632 => x"55567474",
  1633 => x"26e9388a",
  1634 => x"518ac53f",
  1635 => x"8a3d0d04",
  1636 => x"fe3d0d80",
  1637 => x"fc8c0884",
  1638 => x"11087081",
  1639 => x"80800784",
  1640 => x"130c5484",
  1641 => x"110870fe",
  1642 => x"ffff0684",
  1643 => x"130c5452",
  1644 => x"f9853f80",
  1645 => x"f6d4518a",
  1646 => x"b13f8751",
  1647 => x"fea63f80",
  1648 => x"f6e4518a",
  1649 => x"a53f8251",
  1650 => x"fe9a3f80",
  1651 => x"f6f4518a",
  1652 => x"993f8551",
  1653 => x"fe8e3f80",
  1654 => x"f784518a",
  1655 => x"8d3f8651",
  1656 => x"fe823f80",
  1657 => x"f794518a",
  1658 => x"813f8851",
  1659 => x"fdf63f80",
  1660 => x"f7a45189",
  1661 => x"f53f8951",
  1662 => x"fdea3f80",
  1663 => x"0bb00c84",
  1664 => x"3d0d04fe",
  1665 => x"3d0d80fc",
  1666 => x"8c088411",
  1667 => x"08820a07",
  1668 => x"84120c70",
  1669 => x"0870902a",
  1670 => x"84130870",
  1671 => x"fd0a0684",
  1672 => x"150c5481",
  1673 => x"ffff06b0",
  1674 => x"0c535384",
  1675 => x"3d0d04ff",
  1676 => x"3d0d80fb",
  1677 => x"ec087008",
  1678 => x"7081ff06",
  1679 => x"51515271",
  1680 => x"89268c38",
  1681 => x"71101080",
  1682 => x"f8f40552",
  1683 => x"71080480",
  1684 => x"f7b45189",
  1685 => x"953f8a51",
  1686 => x"88f63f80",
  1687 => x"0bb00c83",
  1688 => x"3d0d0480",
  1689 => x"e7e85189",
  1690 => x"813f8a51",
  1691 => x"88e23f80",
  1692 => x"0bb00c83",
  1693 => x"3d0d0480",
  1694 => x"f7bc5188",
  1695 => x"ed3f8a51",
  1696 => x"88ce3f80",
  1697 => x"0bb00c83",
  1698 => x"3d0d0480",
  1699 => x"f7c45188",
  1700 => x"d93f8a51",
  1701 => x"88ba3f80",
  1702 => x"0bb00c83",
  1703 => x"3d0d0480",
  1704 => x"f7d05188",
  1705 => x"c53f8a51",
  1706 => x"88a63f80",
  1707 => x"0bb00c83",
  1708 => x"3d0d0480",
  1709 => x"f7d85188",
  1710 => x"b13f8a51",
  1711 => x"88923f80",
  1712 => x"0bb00c83",
  1713 => x"3d0d0480",
  1714 => x"f7e05188",
  1715 => x"9d3f8a51",
  1716 => x"87fe3f80",
  1717 => x"0bb00c83",
  1718 => x"3d0d0480",
  1719 => x"f7e85188",
  1720 => x"893f8a51",
  1721 => x"87ea3f80",
  1722 => x"0bb00c83",
  1723 => x"3d0d0480",
  1724 => x"f7f05187",
  1725 => x"f53f8a51",
  1726 => x"87d63f80",
  1727 => x"0bb00c83",
  1728 => x"3d0d0480",
  1729 => x"f7f85187",
  1730 => x"e13f8a51",
  1731 => x"87c23f80",
  1732 => x"0bb00c83",
  1733 => x"3d0d04fe",
  1734 => x"3d0d80fb",
  1735 => x"ec088411",
  1736 => x"0880f880",
  1737 => x"53545287",
  1738 => x"c13f7282",
  1739 => x"2a810651",
  1740 => x"89823f80",
  1741 => x"f8905187",
  1742 => x"b13f7281",
  1743 => x"2a810651",
  1744 => x"88f23f80",
  1745 => x"f8a45187",
  1746 => x"a13f7281",
  1747 => x"065188e4",
  1748 => x"3f8a5186",
  1749 => x"fb3f72b0",
  1750 => x"0c843d0d",
  1751 => x"04fe3d0d",
  1752 => x"02930533",
  1753 => x"02840597",
  1754 => x"053380fb",
  1755 => x"ec085553",
  1756 => x"5180730c",
  1757 => x"7688140c",
  1758 => x"70832b72",
  1759 => x"078c140c",
  1760 => x"72085170",
  1761 => x"fb3870b0",
  1762 => x"0c843d0d",
  1763 => x"04fe3d0d",
  1764 => x"80f8b851",
  1765 => x"86d43f80",
  1766 => x"fbec08a0",
  1767 => x"11085353",
  1768 => x"a05186e9",
  1769 => x"3f80fbec",
  1770 => x"08a41108",
  1771 => x"5353a051",
  1772 => x"86db3f80",
  1773 => x"f8d05186",
  1774 => x"b13f80fb",
  1775 => x"ec08a811",
  1776 => x"085353a0",
  1777 => x"5186c63f",
  1778 => x"80fbec08",
  1779 => x"ac110853",
  1780 => x"53a05186",
  1781 => x"b83f8a51",
  1782 => x"85f63f80",
  1783 => x"0bb00c84",
  1784 => x"3d0d04fc",
  1785 => x"3d0d80fb",
  1786 => x"ec089c11",
  1787 => x"087081ff",
  1788 => x"0680f8e8",
  1789 => x"54575353",
  1790 => x"85f03f74",
  1791 => x"5187b53f",
  1792 => x"8a5185cc",
  1793 => x"3f800bff",
  1794 => x"16555372",
  1795 => x"7425a238",
  1796 => x"72101080",
  1797 => x"fbe80805",
  1798 => x"70085252",
  1799 => x"87963f8a",
  1800 => x"5185ad3f",
  1801 => x"81137081",
  1802 => x"ff065452",
  1803 => x"737324e0",
  1804 => x"3874b00c",
  1805 => x"863d0d04",
  1806 => x"fd3d0d81",
  1807 => x"51e08c3f",
  1808 => x"b00881ff",
  1809 => x"06528251",
  1810 => x"e1b33fb0",
  1811 => x"0881ff06",
  1812 => x"538351e1",
  1813 => x"a83f80fb",
  1814 => x"ec085480",
  1815 => x"740cb008",
  1816 => x"88150c71",
  1817 => x"832b7307",
  1818 => x"8c150c73",
  1819 => x"085271fb",
  1820 => x"3871b00c",
  1821 => x"853d0d04",
  1822 => x"ff3d0d81",
  1823 => x"51dfcc3f",
  1824 => x"80fbec08",
  1825 => x"b0089012",
  1826 => x"0c528272",
  1827 => x"0c833d0d",
  1828 => x"04803d0d",
  1829 => x"80fbec08",
  1830 => x"5180710c",
  1831 => x"70b00c82",
  1832 => x"3d0d04fd",
  1833 => x"3d0d800b",
  1834 => x"80fbec08",
  1835 => x"54548073",
  1836 => x"0cfecac0",
  1837 => x"90860b88",
  1838 => x"140c7383",
  1839 => x"2b82078c",
  1840 => x"140c7208",
  1841 => x"5271fb38",
  1842 => x"81147081",
  1843 => x"ff065551",
  1844 => x"a27427da",
  1845 => x"3871b00c",
  1846 => x"853d0d04",
  1847 => x"fd3d0d80",
  1848 => x"0b80fbec",
  1849 => x"08545480",
  1850 => x"730c880a",
  1851 => x"0b88140c",
  1852 => x"73832b81",
  1853 => x"078c140c",
  1854 => x"72085271",
  1855 => x"fb388114",
  1856 => x"7081ff06",
  1857 => x"5551a274",
  1858 => x"27dd3871",
  1859 => x"b00c853d",
  1860 => x"0d04fe3d",
  1861 => x"0d8151de",
  1862 => x"b23f80fb",
  1863 => x"ec085380",
  1864 => x"730c810b",
  1865 => x"88140cb0",
  1866 => x"08832b8f",
  1867 => x"f8067082",
  1868 => x"078c150c",
  1869 => x"52720852",
  1870 => x"71fb3889",
  1871 => x"730c71b0",
  1872 => x"0c843d0d",
  1873 => x"04d88a3f",
  1874 => x"04fb3d0d",
  1875 => x"77795555",
  1876 => x"80567575",
  1877 => x"24ab3880",
  1878 => x"74249d38",
  1879 => x"80537352",
  1880 => x"745180e1",
  1881 => x"3fb00854",
  1882 => x"75802e85",
  1883 => x"38b00830",
  1884 => x"5473b00c",
  1885 => x"873d0d04",
  1886 => x"73307681",
  1887 => x"325754dc",
  1888 => x"39743055",
  1889 => x"81567380",
  1890 => x"25d238ec",
  1891 => x"39fa3d0d",
  1892 => x"787a5755",
  1893 => x"80577675",
  1894 => x"24a43875",
  1895 => x"9f2c5481",
  1896 => x"53757432",
  1897 => x"74315274",
  1898 => x"519b3fb0",
  1899 => x"08547680",
  1900 => x"2e8538b0",
  1901 => x"08305473",
  1902 => x"b00c883d",
  1903 => x"0d047430",
  1904 => x"558157d7",
  1905 => x"39fc3d0d",
  1906 => x"76785354",
  1907 => x"81538074",
  1908 => x"73265255",
  1909 => x"72802e98",
  1910 => x"3870802e",
  1911 => x"a9388072",
  1912 => x"24a43871",
  1913 => x"10731075",
  1914 => x"72265354",
  1915 => x"5272ea38",
  1916 => x"73517883",
  1917 => x"38745170",
  1918 => x"b00c863d",
  1919 => x"0d047281",
  1920 => x"2a72812a",
  1921 => x"53537280",
  1922 => x"2ee63871",
  1923 => x"7426ef38",
  1924 => x"73723175",
  1925 => x"74077481",
  1926 => x"2a74812a",
  1927 => x"55555654",
  1928 => x"e5391010",
  1929 => x"10101010",
  1930 => x"10101010",
  1931 => x"10101010",
  1932 => x"10101010",
  1933 => x"10101010",
  1934 => x"10101010",
  1935 => x"10101010",
  1936 => x"10535104",
  1937 => x"7381ff06",
  1938 => x"73830609",
  1939 => x"81058305",
  1940 => x"1010102b",
  1941 => x"0772fc06",
  1942 => x"0c515104",
  1943 => x"3c047272",
  1944 => x"80728106",
  1945 => x"ff050972",
  1946 => x"06057110",
  1947 => x"52720a10",
  1948 => x"0a5372ed",
  1949 => x"38515153",
  1950 => x"5104b008",
  1951 => x"b408b808",
  1952 => x"7575bb8d",
  1953 => x"2d5050b0",
  1954 => x"0856b80c",
  1955 => x"b40cb00c",
  1956 => x"5104b008",
  1957 => x"b408b808",
  1958 => x"7575bac9",
  1959 => x"2d5050b0",
  1960 => x"0856b80c",
  1961 => x"b40cb00c",
  1962 => x"5104b008",
  1963 => x"b408b808",
  1964 => x"90b92db8",
  1965 => x"0cb40cb0",
  1966 => x"0c04ff3d",
  1967 => x"0d028f05",
  1968 => x"3380fc9c",
  1969 => x"0852710c",
  1970 => x"800bb00c",
  1971 => x"833d0d04",
  1972 => x"ff3d0d02",
  1973 => x"8f053351",
  1974 => x"81a4b408",
  1975 => x"52712db0",
  1976 => x"0881ff06",
  1977 => x"b00c833d",
  1978 => x"0d04fe3d",
  1979 => x"0d747033",
  1980 => x"53537180",
  1981 => x"2e933881",
  1982 => x"13725281",
  1983 => x"a4b40853",
  1984 => x"53712d72",
  1985 => x"335271ef",
  1986 => x"38843d0d",
  1987 => x"04f43d0d",
  1988 => x"7f028405",
  1989 => x"bb053355",
  1990 => x"57880b8c",
  1991 => x"3d5b5989",
  1992 => x"5380f9c0",
  1993 => x"52795185",
  1994 => x"e63f7379",
  1995 => x"2e80ff38",
  1996 => x"78567390",
  1997 => x"2e80ec38",
  1998 => x"02a70558",
  1999 => x"768f0654",
  2000 => x"73892680",
  2001 => x"c2387518",
  2002 => x"b0155555",
  2003 => x"73753476",
  2004 => x"842aff17",
  2005 => x"7081ff06",
  2006 => x"58555775",
  2007 => x"df38781a",
  2008 => x"55757534",
  2009 => x"79703355",
  2010 => x"5573802e",
  2011 => x"93388115",
  2012 => x"745281a4",
  2013 => x"b4085755",
  2014 => x"752d7433",
  2015 => x"5473ef38",
  2016 => x"78b00c8e",
  2017 => x"3d0d0475",
  2018 => x"18b71555",
  2019 => x"55737534",
  2020 => x"76842aff",
  2021 => x"177081ff",
  2022 => x"06585557",
  2023 => x"75ff9d38",
  2024 => x"ffbc3984",
  2025 => x"70575902",
  2026 => x"a70558ff",
  2027 => x"8f398270",
  2028 => x"5759f439",
  2029 => x"f13d0d61",
  2030 => x"8d3d705b",
  2031 => x"5c5a807a",
  2032 => x"5657767a",
  2033 => x"24818538",
  2034 => x"7817548a",
  2035 => x"52745184",
  2036 => x"8c3fb008",
  2037 => x"b0055372",
  2038 => x"74348117",
  2039 => x"578a5274",
  2040 => x"5183d53f",
  2041 => x"b00855b0",
  2042 => x"08de38b0",
  2043 => x"08779f2a",
  2044 => x"1870812c",
  2045 => x"5a565680",
  2046 => x"78259e38",
  2047 => x"7817ff05",
  2048 => x"55751970",
  2049 => x"33555374",
  2050 => x"33733473",
  2051 => x"75348116",
  2052 => x"ff165656",
  2053 => x"777624e9",
  2054 => x"38761958",
  2055 => x"80783480",
  2056 => x"7a241770",
  2057 => x"81ff067c",
  2058 => x"70335657",
  2059 => x"55567280",
  2060 => x"2e933881",
  2061 => x"15735281",
  2062 => x"a4b40858",
  2063 => x"55762d74",
  2064 => x"335372ef",
  2065 => x"3873b00c",
  2066 => x"913d0d04",
  2067 => x"ad7b3402",
  2068 => x"ad057a30",
  2069 => x"71195656",
  2070 => x"598a5274",
  2071 => x"5182fe3f",
  2072 => x"b008b005",
  2073 => x"53727434",
  2074 => x"8117578a",
  2075 => x"52745182",
  2076 => x"c73fb008",
  2077 => x"55b008fe",
  2078 => x"cf38feef",
  2079 => x"39fd3d0d",
  2080 => x"02970533",
  2081 => x"0284059b",
  2082 => x"05335553",
  2083 => x"72742797",
  2084 => x"38a05181",
  2085 => x"a4b40852",
  2086 => x"712d8113",
  2087 => x"7081ff06",
  2088 => x"54527373",
  2089 => x"26eb3885",
  2090 => x"3d0d04ff",
  2091 => x"3d0d80fc",
  2092 => x"90087410",
  2093 => x"1570822b",
  2094 => x"94130c52",
  2095 => x"52850b98",
  2096 => x"130c9812",
  2097 => x"08708106",
  2098 => x"515170f6",
  2099 => x"38833d0d",
  2100 => x"04fd3d0d",
  2101 => x"80fc9008",
  2102 => x"7680e1d4",
  2103 => x"2994120c",
  2104 => x"54850b98",
  2105 => x"150c9814",
  2106 => x"08708106",
  2107 => x"515372f6",
  2108 => x"38853d0d",
  2109 => x"04803d0d",
  2110 => x"80fc9008",
  2111 => x"51870b84",
  2112 => x"120cff0b",
  2113 => x"a4120ca7",
  2114 => x"0ba8120c",
  2115 => x"80e1d40b",
  2116 => x"94120c87",
  2117 => x"0b98120c",
  2118 => x"823d0d04",
  2119 => x"803d0d80",
  2120 => x"fc940851",
  2121 => x"80ec0b8c",
  2122 => x"120c830b",
  2123 => x"88120c82",
  2124 => x"3d0d0480",
  2125 => x"3d0d80fc",
  2126 => x"94088411",
  2127 => x"088106b0",
  2128 => x"0c51823d",
  2129 => x"0d04ff3d",
  2130 => x"0d80fc94",
  2131 => x"08528412",
  2132 => x"08708106",
  2133 => x"51517080",
  2134 => x"2ef43871",
  2135 => x"087081ff",
  2136 => x"06b00c51",
  2137 => x"833d0d04",
  2138 => x"fe3d0d02",
  2139 => x"93053353",
  2140 => x"728a2e9c",
  2141 => x"3880fc94",
  2142 => x"08528412",
  2143 => x"0870892a",
  2144 => x"70810651",
  2145 => x"515170f2",
  2146 => x"3872720c",
  2147 => x"843d0d04",
  2148 => x"80fc9408",
  2149 => x"52841208",
  2150 => x"70892a70",
  2151 => x"81065151",
  2152 => x"5170f238",
  2153 => x"8d720c84",
  2154 => x"12087089",
  2155 => x"2a708106",
  2156 => x"51515170",
  2157 => x"c538d239",
  2158 => x"bc0802bc",
  2159 => x"0cfd3d0d",
  2160 => x"8053bc08",
  2161 => x"8c050852",
  2162 => x"bc088805",
  2163 => x"0851f7f5",
  2164 => x"3fb00870",
  2165 => x"b00c5485",
  2166 => x"3d0dbc0c",
  2167 => x"04bc0802",
  2168 => x"bc0cfd3d",
  2169 => x"0d8153bc",
  2170 => x"088c0508",
  2171 => x"52bc0888",
  2172 => x"050851f7",
  2173 => x"d03fb008",
  2174 => x"70b00c54",
  2175 => x"853d0dbc",
  2176 => x"0c04803d",
  2177 => x"0d865184",
  2178 => x"963f8151",
  2179 => x"a1d33ffc",
  2180 => x"3d0d7670",
  2181 => x"797b5555",
  2182 => x"55558f72",
  2183 => x"278c3872",
  2184 => x"75078306",
  2185 => x"5170802e",
  2186 => x"a738ff12",
  2187 => x"5271ff2e",
  2188 => x"98387270",
  2189 => x"81055433",
  2190 => x"74708105",
  2191 => x"5634ff12",
  2192 => x"5271ff2e",
  2193 => x"098106ea",
  2194 => x"3874b00c",
  2195 => x"863d0d04",
  2196 => x"74517270",
  2197 => x"84055408",
  2198 => x"71708405",
  2199 => x"530c7270",
  2200 => x"84055408",
  2201 => x"71708405",
  2202 => x"530c7270",
  2203 => x"84055408",
  2204 => x"71708405",
  2205 => x"530c7270",
  2206 => x"84055408",
  2207 => x"71708405",
  2208 => x"530cf012",
  2209 => x"52718f26",
  2210 => x"c9388372",
  2211 => x"27953872",
  2212 => x"70840554",
  2213 => x"08717084",
  2214 => x"05530cfc",
  2215 => x"12527183",
  2216 => x"26ed3870",
  2217 => x"54ff8339",
  2218 => x"fd3d0d75",
  2219 => x"5384d813",
  2220 => x"08802e8a",
  2221 => x"38805372",
  2222 => x"b00c853d",
  2223 => x"0d048180",
  2224 => x"5272518d",
  2225 => x"9b3fb008",
  2226 => x"84d8140c",
  2227 => x"ff53b008",
  2228 => x"802ee438",
  2229 => x"b008549f",
  2230 => x"53807470",
  2231 => x"8405560c",
  2232 => x"ff135380",
  2233 => x"7324ce38",
  2234 => x"80747084",
  2235 => x"05560cff",
  2236 => x"13537280",
  2237 => x"25e338ff",
  2238 => x"bc39fd3d",
  2239 => x"0d757755",
  2240 => x"539f7427",
  2241 => x"8d389673",
  2242 => x"0cff5271",
  2243 => x"b00c853d",
  2244 => x"0d0484d8",
  2245 => x"13085271",
  2246 => x"802e9338",
  2247 => x"73101012",
  2248 => x"70087972",
  2249 => x"0c515271",
  2250 => x"b00c853d",
  2251 => x"0d047251",
  2252 => x"fef63fff",
  2253 => x"52b008d3",
  2254 => x"3884d813",
  2255 => x"08741010",
  2256 => x"1170087a",
  2257 => x"720c5151",
  2258 => x"52dd39f9",
  2259 => x"3d0d797b",
  2260 => x"5856769f",
  2261 => x"2680e838",
  2262 => x"84d81608",
  2263 => x"5473802e",
  2264 => x"aa387610",
  2265 => x"10147008",
  2266 => x"55557380",
  2267 => x"2eba3880",
  2268 => x"5873812e",
  2269 => x"8f3873ff",
  2270 => x"2ea33880",
  2271 => x"750c7651",
  2272 => x"732d8058",
  2273 => x"77b00c89",
  2274 => x"3d0d0475",
  2275 => x"51fe993f",
  2276 => x"ff58b008",
  2277 => x"ef3884d8",
  2278 => x"160854c6",
  2279 => x"3996760c",
  2280 => x"810bb00c",
  2281 => x"893d0d04",
  2282 => x"755181ed",
  2283 => x"3f7653b0",
  2284 => x"08527551",
  2285 => x"81ad3fb0",
  2286 => x"08b00c89",
  2287 => x"3d0d0496",
  2288 => x"760cff0b",
  2289 => x"b00c893d",
  2290 => x"0d04fc3d",
  2291 => x"0d767856",
  2292 => x"53ff5474",
  2293 => x"9f26b138",
  2294 => x"84d81308",
  2295 => x"5271802e",
  2296 => x"ae387410",
  2297 => x"10127008",
  2298 => x"53538154",
  2299 => x"71802e98",
  2300 => x"38825471",
  2301 => x"ff2e9138",
  2302 => x"83547181",
  2303 => x"2e8a3880",
  2304 => x"730c7451",
  2305 => x"712d8054",
  2306 => x"73b00c86",
  2307 => x"3d0d0472",
  2308 => x"51fd953f",
  2309 => x"b008f138",
  2310 => x"84d81308",
  2311 => x"52c439ff",
  2312 => x"3d0d7352",
  2313 => x"80fca008",
  2314 => x"51fea03f",
  2315 => x"833d0d04",
  2316 => x"fe3d0d75",
  2317 => x"53745280",
  2318 => x"fca00851",
  2319 => x"fdbc3f84",
  2320 => x"3d0d0480",
  2321 => x"3d0d80fc",
  2322 => x"a00851fc",
  2323 => x"db3f823d",
  2324 => x"0d04ff3d",
  2325 => x"0d735280",
  2326 => x"fca00851",
  2327 => x"feec3f83",
  2328 => x"3d0d04fc",
  2329 => x"3d0d800b",
  2330 => x"81a4bc0c",
  2331 => x"78527751",
  2332 => x"9caa3fb0",
  2333 => x"0854b008",
  2334 => x"ff2e8838",
  2335 => x"73b00c86",
  2336 => x"3d0d0481",
  2337 => x"a4bc0855",
  2338 => x"74802ef0",
  2339 => x"38767571",
  2340 => x"0c5373b0",
  2341 => x"0c863d0d",
  2342 => x"049bfc3f",
  2343 => x"04fc3d0d",
  2344 => x"76707970",
  2345 => x"73078306",
  2346 => x"54545455",
  2347 => x"7080c338",
  2348 => x"71700870",
  2349 => x"0970f7fb",
  2350 => x"fdff1306",
  2351 => x"70f88482",
  2352 => x"81800651",
  2353 => x"51535354",
  2354 => x"70a63884",
  2355 => x"14727470",
  2356 => x"8405560c",
  2357 => x"70087009",
  2358 => x"70f7fbfd",
  2359 => x"ff130670",
  2360 => x"f8848281",
  2361 => x"80065151",
  2362 => x"53535470",
  2363 => x"802edc38",
  2364 => x"73527170",
  2365 => x"81055333",
  2366 => x"51707370",
  2367 => x"81055534",
  2368 => x"70f03874",
  2369 => x"b00c863d",
  2370 => x"0d04fd3d",
  2371 => x"0d757071",
  2372 => x"83065355",
  2373 => x"5270b838",
  2374 => x"71700870",
  2375 => x"09f7fbfd",
  2376 => x"ff120670",
  2377 => x"f8848281",
  2378 => x"80065151",
  2379 => x"5253709d",
  2380 => x"38841370",
  2381 => x"087009f7",
  2382 => x"fbfdff12",
  2383 => x"0670f884",
  2384 => x"82818006",
  2385 => x"51515253",
  2386 => x"70802ee5",
  2387 => x"38725271",
  2388 => x"33517080",
  2389 => x"2e8a3881",
  2390 => x"12703352",
  2391 => x"5270f838",
  2392 => x"717431b0",
  2393 => x"0c853d0d",
  2394 => x"04fa3d0d",
  2395 => x"787a7c70",
  2396 => x"54555552",
  2397 => x"72802e80",
  2398 => x"d9387174",
  2399 => x"07830651",
  2400 => x"70802e80",
  2401 => x"d438ff13",
  2402 => x"5372ff2e",
  2403 => x"b1387133",
  2404 => x"74335651",
  2405 => x"74712e09",
  2406 => x"8106a938",
  2407 => x"72802e81",
  2408 => x"87387081",
  2409 => x"ff065170",
  2410 => x"802e80fc",
  2411 => x"38811281",
  2412 => x"15ff1555",
  2413 => x"555272ff",
  2414 => x"2e098106",
  2415 => x"d1387133",
  2416 => x"74335651",
  2417 => x"7081ff06",
  2418 => x"7581ff06",
  2419 => x"71713151",
  2420 => x"525270b0",
  2421 => x"0c883d0d",
  2422 => x"04717457",
  2423 => x"55837327",
  2424 => x"88387108",
  2425 => x"74082e88",
  2426 => x"38747655",
  2427 => x"52ff9739",
  2428 => x"fc135372",
  2429 => x"802eb138",
  2430 => x"74087009",
  2431 => x"f7fbfdff",
  2432 => x"120670f8",
  2433 => x"84828180",
  2434 => x"06515151",
  2435 => x"709a3884",
  2436 => x"15841757",
  2437 => x"55837327",
  2438 => x"d0387408",
  2439 => x"76082ed0",
  2440 => x"38747655",
  2441 => x"52fedf39",
  2442 => x"800bb00c",
  2443 => x"883d0d04",
  2444 => x"f33d0d60",
  2445 => x"6264725a",
  2446 => x"5a5e5e80",
  2447 => x"5c767081",
  2448 => x"05583380",
  2449 => x"f9d51133",
  2450 => x"70832a70",
  2451 => x"81065155",
  2452 => x"555672e9",
  2453 => x"3875ad2e",
  2454 => x"82883875",
  2455 => x"ab2e8284",
  2456 => x"38773070",
  2457 => x"79078025",
  2458 => x"79903270",
  2459 => x"30707207",
  2460 => x"80257307",
  2461 => x"53575751",
  2462 => x"5372802e",
  2463 => x"873875b0",
  2464 => x"2e81eb38",
  2465 => x"778a3888",
  2466 => x"5875b02e",
  2467 => x"83388a58",
  2468 => x"810a5a7b",
  2469 => x"8438fe0a",
  2470 => x"5a775279",
  2471 => x"51f6be3f",
  2472 => x"b0087853",
  2473 => x"7a525bf6",
  2474 => x"8f3fb008",
  2475 => x"5a807080",
  2476 => x"f9d51833",
  2477 => x"70822a70",
  2478 => x"81065156",
  2479 => x"565a5572",
  2480 => x"802e80c1",
  2481 => x"38d01656",
  2482 => x"75782580",
  2483 => x"d7388079",
  2484 => x"24757b26",
  2485 => x"07537293",
  2486 => x"38747a2e",
  2487 => x"80eb387a",
  2488 => x"762580ed",
  2489 => x"3872802e",
  2490 => x"80e738ff",
  2491 => x"77708105",
  2492 => x"59335759",
  2493 => x"80f9d516",
  2494 => x"3370822a",
  2495 => x"70810651",
  2496 => x"545472c1",
  2497 => x"38738306",
  2498 => x"5372802e",
  2499 => x"97387381",
  2500 => x"06c91755",
  2501 => x"53728538",
  2502 => x"ffa91654",
  2503 => x"73567776",
  2504 => x"24ffab38",
  2505 => x"80792480",
  2506 => x"f0387b80",
  2507 => x"2e843874",
  2508 => x"30557c80",
  2509 => x"2e8c38ff",
  2510 => x"17537883",
  2511 => x"387d5372",
  2512 => x"7d0c74b0",
  2513 => x"0c8f3d0d",
  2514 => x"04815375",
  2515 => x"7b24ff95",
  2516 => x"38817579",
  2517 => x"29177870",
  2518 => x"81055a33",
  2519 => x"585659ff",
  2520 => x"9339815c",
  2521 => x"76708105",
  2522 => x"583356fd",
  2523 => x"f4398077",
  2524 => x"33545472",
  2525 => x"80f82eb2",
  2526 => x"387280d8",
  2527 => x"32703070",
  2528 => x"80257607",
  2529 => x"51515372",
  2530 => x"802efdf8",
  2531 => x"38811733",
  2532 => x"82185856",
  2533 => x"9058fdf8",
  2534 => x"39810a55",
  2535 => x"7b8438fe",
  2536 => x"0a557f53",
  2537 => x"a2730cff",
  2538 => x"89398154",
  2539 => x"cc39fd3d",
  2540 => x"0d775476",
  2541 => x"53755280",
  2542 => x"fca00851",
  2543 => x"fcf23f85",
  2544 => x"3d0d04f3",
  2545 => x"3d0d6062",
  2546 => x"64725a5a",
  2547 => x"5d5d805e",
  2548 => x"76708105",
  2549 => x"583380f9",
  2550 => x"d5113370",
  2551 => x"832a7081",
  2552 => x"06515555",
  2553 => x"5672e938",
  2554 => x"75ad2e81",
  2555 => x"ff3875ab",
  2556 => x"2e81fb38",
  2557 => x"77307079",
  2558 => x"07802579",
  2559 => x"90327030",
  2560 => x"70720780",
  2561 => x"25730753",
  2562 => x"57575153",
  2563 => x"72802e87",
  2564 => x"3875b02e",
  2565 => x"81e23877",
  2566 => x"8a388858",
  2567 => x"75b02e83",
  2568 => x"388a5877",
  2569 => x"52ff51f3",
  2570 => x"8f3fb008",
  2571 => x"78535aff",
  2572 => x"51f3aa3f",
  2573 => x"b0085b80",
  2574 => x"705a5580",
  2575 => x"f9d51633",
  2576 => x"70822a70",
  2577 => x"81065154",
  2578 => x"5472802e",
  2579 => x"80c138d0",
  2580 => x"16567578",
  2581 => x"2580d738",
  2582 => x"80792475",
  2583 => x"7b260753",
  2584 => x"72933874",
  2585 => x"7a2e80eb",
  2586 => x"387a7625",
  2587 => x"80ed3872",
  2588 => x"802e80e7",
  2589 => x"38ff7770",
  2590 => x"81055933",
  2591 => x"575980f9",
  2592 => x"d5163370",
  2593 => x"822a7081",
  2594 => x"06515454",
  2595 => x"72c13873",
  2596 => x"83065372",
  2597 => x"802e9738",
  2598 => x"738106c9",
  2599 => x"17555372",
  2600 => x"8538ffa9",
  2601 => x"16547356",
  2602 => x"777624ff",
  2603 => x"ab388079",
  2604 => x"24818938",
  2605 => x"7d802e84",
  2606 => x"38743055",
  2607 => x"7b802e8c",
  2608 => x"38ff1753",
  2609 => x"7883387c",
  2610 => x"53727c0c",
  2611 => x"74b00c8f",
  2612 => x"3d0d0481",
  2613 => x"53757b24",
  2614 => x"ff953881",
  2615 => x"75792917",
  2616 => x"78708105",
  2617 => x"5a335856",
  2618 => x"59ff9339",
  2619 => x"815e7670",
  2620 => x"81055833",
  2621 => x"56fdfd39",
  2622 => x"80773354",
  2623 => x"547280f8",
  2624 => x"2e80c338",
  2625 => x"7280d832",
  2626 => x"70307080",
  2627 => x"25760751",
  2628 => x"51537280",
  2629 => x"2efe8038",
  2630 => x"81173382",
  2631 => x"18585690",
  2632 => x"705358ff",
  2633 => x"51f1913f",
  2634 => x"b0087853",
  2635 => x"5aff51f1",
  2636 => x"ac3fb008",
  2637 => x"5b80705a",
  2638 => x"55fe8039",
  2639 => x"ff605455",
  2640 => x"a2730cfe",
  2641 => x"f7398154",
  2642 => x"ffba39fd",
  2643 => x"3d0d7754",
  2644 => x"76537552",
  2645 => x"80fca008",
  2646 => x"51fce83f",
  2647 => x"853d0d04",
  2648 => x"f33d0d7f",
  2649 => x"618b1170",
  2650 => x"f8065c55",
  2651 => x"555e7296",
  2652 => x"26833890",
  2653 => x"59807924",
  2654 => x"747a2607",
  2655 => x"53805472",
  2656 => x"742e0981",
  2657 => x"0680cb38",
  2658 => x"7d518bca",
  2659 => x"3f7883f7",
  2660 => x"2680c638",
  2661 => x"78832a70",
  2662 => x"10101081",
  2663 => x"83dc058c",
  2664 => x"11085959",
  2665 => x"5a76782e",
  2666 => x"83b03884",
  2667 => x"1708fc06",
  2668 => x"568c1708",
  2669 => x"88180871",
  2670 => x"8c120c88",
  2671 => x"120c5875",
  2672 => x"17841108",
  2673 => x"81078412",
  2674 => x"0c537d51",
  2675 => x"8b893f88",
  2676 => x"175473b0",
  2677 => x"0c8f3d0d",
  2678 => x"0478892a",
  2679 => x"79832a5b",
  2680 => x"5372802e",
  2681 => x"bf387886",
  2682 => x"2ab8055a",
  2683 => x"847327b4",
  2684 => x"3880db13",
  2685 => x"5a947327",
  2686 => x"ab38788c",
  2687 => x"2a80ee05",
  2688 => x"5a80d473",
  2689 => x"279e3878",
  2690 => x"8f2a80f7",
  2691 => x"055a82d4",
  2692 => x"73279138",
  2693 => x"78922a80",
  2694 => x"fc055a8a",
  2695 => x"d4732784",
  2696 => x"3880fe5a",
  2697 => x"79101010",
  2698 => x"8183dc05",
  2699 => x"8c110858",
  2700 => x"5576752e",
  2701 => x"a3388417",
  2702 => x"08fc0670",
  2703 => x"7a315556",
  2704 => x"738f2488",
  2705 => x"d5387380",
  2706 => x"25fee638",
  2707 => x"8c170857",
  2708 => x"76752e09",
  2709 => x"8106df38",
  2710 => x"811a5a81",
  2711 => x"83ec0857",
  2712 => x"768183e4",
  2713 => x"2e82c038",
  2714 => x"841708fc",
  2715 => x"06707a31",
  2716 => x"5556738f",
  2717 => x"2481f938",
  2718 => x"8183e40b",
  2719 => x"8183f00c",
  2720 => x"8183e40b",
  2721 => x"8183ec0c",
  2722 => x"738025fe",
  2723 => x"b23883ff",
  2724 => x"762783df",
  2725 => x"3875892a",
  2726 => x"76832a55",
  2727 => x"5372802e",
  2728 => x"bf387586",
  2729 => x"2ab80554",
  2730 => x"847327b4",
  2731 => x"3880db13",
  2732 => x"54947327",
  2733 => x"ab38758c",
  2734 => x"2a80ee05",
  2735 => x"5480d473",
  2736 => x"279e3875",
  2737 => x"8f2a80f7",
  2738 => x"055482d4",
  2739 => x"73279138",
  2740 => x"75922a80",
  2741 => x"fc05548a",
  2742 => x"d4732784",
  2743 => x"3880fe54",
  2744 => x"73101010",
  2745 => x"8183dc05",
  2746 => x"88110856",
  2747 => x"5874782e",
  2748 => x"86cf3884",
  2749 => x"1508fc06",
  2750 => x"53757327",
  2751 => x"8d388815",
  2752 => x"08557478",
  2753 => x"2e098106",
  2754 => x"ea388c15",
  2755 => x"088183dc",
  2756 => x"0b840508",
  2757 => x"718c1a0c",
  2758 => x"76881a0c",
  2759 => x"7888130c",
  2760 => x"788c180c",
  2761 => x"5d587953",
  2762 => x"807a2483",
  2763 => x"e6387282",
  2764 => x"2c81712b",
  2765 => x"5c537a7c",
  2766 => x"26819838",
  2767 => x"7b7b0653",
  2768 => x"7282f138",
  2769 => x"79fc0684",
  2770 => x"055a7a10",
  2771 => x"707d0654",
  2772 => x"5b7282e0",
  2773 => x"38841a5a",
  2774 => x"f1398817",
  2775 => x"8c110858",
  2776 => x"5876782e",
  2777 => x"098106fc",
  2778 => x"c238821a",
  2779 => x"5afdec39",
  2780 => x"78177981",
  2781 => x"0784190c",
  2782 => x"708183f0",
  2783 => x"0c708183",
  2784 => x"ec0c8183",
  2785 => x"e40b8c12",
  2786 => x"0c8c1108",
  2787 => x"88120c74",
  2788 => x"81078412",
  2789 => x"0c741175",
  2790 => x"710c5153",
  2791 => x"7d5187b7",
  2792 => x"3f881754",
  2793 => x"fcac3981",
  2794 => x"83dc0b84",
  2795 => x"05087a54",
  2796 => x"5c798025",
  2797 => x"fef83882",
  2798 => x"da397a09",
  2799 => x"7c067081",
  2800 => x"83dc0b84",
  2801 => x"050c5c7a",
  2802 => x"105b7a7c",
  2803 => x"2685387a",
  2804 => x"85b83881",
  2805 => x"83dc0b88",
  2806 => x"05087084",
  2807 => x"1208fc06",
  2808 => x"707c317c",
  2809 => x"72268f72",
  2810 => x"25075757",
  2811 => x"5c5d5572",
  2812 => x"802e80db",
  2813 => x"38797a16",
  2814 => x"8183d408",
  2815 => x"1b90115a",
  2816 => x"55575b81",
  2817 => x"83d008ff",
  2818 => x"2e8838a0",
  2819 => x"8f13e080",
  2820 => x"06577652",
  2821 => x"7d5186c0",
  2822 => x"3fb00854",
  2823 => x"b008ff2e",
  2824 => x"9038b008",
  2825 => x"76278299",
  2826 => x"38748183",
  2827 => x"dc2e8291",
  2828 => x"388183dc",
  2829 => x"0b880508",
  2830 => x"55841508",
  2831 => x"fc06707a",
  2832 => x"317a7226",
  2833 => x"8f722507",
  2834 => x"52555372",
  2835 => x"83e63874",
  2836 => x"79810784",
  2837 => x"170c7916",
  2838 => x"708183dc",
  2839 => x"0b88050c",
  2840 => x"75810784",
  2841 => x"120c547e",
  2842 => x"525785eb",
  2843 => x"3f881754",
  2844 => x"fae03975",
  2845 => x"832a7054",
  2846 => x"54807424",
  2847 => x"819b3872",
  2848 => x"822c8171",
  2849 => x"2b8183e0",
  2850 => x"08077081",
  2851 => x"83dc0b84",
  2852 => x"050c7510",
  2853 => x"10108183",
  2854 => x"dc058811",
  2855 => x"08585a5d",
  2856 => x"53778c18",
  2857 => x"0c748818",
  2858 => x"0c768819",
  2859 => x"0c768c16",
  2860 => x"0cfcf339",
  2861 => x"797a1010",
  2862 => x"108183dc",
  2863 => x"05705759",
  2864 => x"5d8c1508",
  2865 => x"5776752e",
  2866 => x"a3388417",
  2867 => x"08fc0670",
  2868 => x"7a315556",
  2869 => x"738f2483",
  2870 => x"ca387380",
  2871 => x"25848138",
  2872 => x"8c170857",
  2873 => x"76752e09",
  2874 => x"8106df38",
  2875 => x"8815811b",
  2876 => x"70830655",
  2877 => x"5b5572c9",
  2878 => x"387c8306",
  2879 => x"5372802e",
  2880 => x"fdb838ff",
  2881 => x"1df81959",
  2882 => x"5d881808",
  2883 => x"782eea38",
  2884 => x"fdb53983",
  2885 => x"1a53fc96",
  2886 => x"39831470",
  2887 => x"822c8171",
  2888 => x"2b8183e0",
  2889 => x"08077081",
  2890 => x"83dc0b84",
  2891 => x"050c7610",
  2892 => x"10108183",
  2893 => x"dc058811",
  2894 => x"08595b5e",
  2895 => x"5153fee1",
  2896 => x"398183a0",
  2897 => x"081758b0",
  2898 => x"08762e81",
  2899 => x"8d388183",
  2900 => x"d008ff2e",
  2901 => x"83ec3873",
  2902 => x"76311881",
  2903 => x"83a00c73",
  2904 => x"87067057",
  2905 => x"5372802e",
  2906 => x"88388873",
  2907 => x"31701555",
  2908 => x"5676149f",
  2909 => x"ff06a080",
  2910 => x"71311770",
  2911 => x"547f5357",
  2912 => x"5383d53f",
  2913 => x"b00853b0",
  2914 => x"08ff2e81",
  2915 => x"a0388183",
  2916 => x"a0081670",
  2917 => x"8183a00c",
  2918 => x"74758183",
  2919 => x"dc0b8805",
  2920 => x"0c747631",
  2921 => x"18708107",
  2922 => x"51555658",
  2923 => x"7b8183dc",
  2924 => x"2e839c38",
  2925 => x"798f2682",
  2926 => x"cb38810b",
  2927 => x"84150c84",
  2928 => x"1508fc06",
  2929 => x"707a317a",
  2930 => x"72268f72",
  2931 => x"25075255",
  2932 => x"5372802e",
  2933 => x"fcf93880",
  2934 => x"db39b008",
  2935 => x"9fff0653",
  2936 => x"72feeb38",
  2937 => x"778183a0",
  2938 => x"0c8183dc",
  2939 => x"0b880508",
  2940 => x"7b188107",
  2941 => x"84120c55",
  2942 => x"8183cc08",
  2943 => x"78278638",
  2944 => x"778183cc",
  2945 => x"0c8183c8",
  2946 => x"087827fc",
  2947 => x"ac387781",
  2948 => x"83c80c84",
  2949 => x"1508fc06",
  2950 => x"707a317a",
  2951 => x"72268f72",
  2952 => x"25075255",
  2953 => x"5372802e",
  2954 => x"fca53888",
  2955 => x"39807454",
  2956 => x"56fedb39",
  2957 => x"7d51829f",
  2958 => x"3f800bb0",
  2959 => x"0c8f3d0d",
  2960 => x"04735380",
  2961 => x"7424a938",
  2962 => x"72822c81",
  2963 => x"712b8183",
  2964 => x"e0080770",
  2965 => x"8183dc0b",
  2966 => x"84050c5d",
  2967 => x"53778c18",
  2968 => x"0c748818",
  2969 => x"0c768819",
  2970 => x"0c768c16",
  2971 => x"0cf9b739",
  2972 => x"83147082",
  2973 => x"2c81712b",
  2974 => x"8183e008",
  2975 => x"07708183",
  2976 => x"dc0b8405",
  2977 => x"0c5e5153",
  2978 => x"d4397b7b",
  2979 => x"065372fc",
  2980 => x"a338841a",
  2981 => x"7b105c5a",
  2982 => x"f139ff1a",
  2983 => x"8111515a",
  2984 => x"f7b93978",
  2985 => x"17798107",
  2986 => x"84190c8c",
  2987 => x"18088819",
  2988 => x"08718c12",
  2989 => x"0c88120c",
  2990 => x"59708183",
  2991 => x"f00c7081",
  2992 => x"83ec0c81",
  2993 => x"83e40b8c",
  2994 => x"120c8c11",
  2995 => x"0888120c",
  2996 => x"74810784",
  2997 => x"120c7411",
  2998 => x"75710c51",
  2999 => x"53f9bd39",
  3000 => x"75178411",
  3001 => x"08810784",
  3002 => x"120c538c",
  3003 => x"17088818",
  3004 => x"08718c12",
  3005 => x"0c88120c",
  3006 => x"587d5180",
  3007 => x"da3f8817",
  3008 => x"54f5cf39",
  3009 => x"7284150c",
  3010 => x"f41af806",
  3011 => x"70841e08",
  3012 => x"81060784",
  3013 => x"1e0c701d",
  3014 => x"545b850b",
  3015 => x"84140c85",
  3016 => x"0b88140c",
  3017 => x"8f7b27fd",
  3018 => x"cf38881c",
  3019 => x"527d5182",
  3020 => x"903f8183",
  3021 => x"dc0b8805",
  3022 => x"088183a0",
  3023 => x"085955fd",
  3024 => x"b7397781",
  3025 => x"83a00c73",
  3026 => x"8183d00c",
  3027 => x"fc913972",
  3028 => x"84150cfd",
  3029 => x"a3390404",
  3030 => x"fd3d0d80",
  3031 => x"0b81a4bc",
  3032 => x"0c765186",
  3033 => x"cb3fb008",
  3034 => x"53b008ff",
  3035 => x"2e883872",
  3036 => x"b00c853d",
  3037 => x"0d0481a4",
  3038 => x"bc085473",
  3039 => x"802ef038",
  3040 => x"7574710c",
  3041 => x"5272b00c",
  3042 => x"853d0d04",
  3043 => x"fb3d0d77",
  3044 => x"705256c2",
  3045 => x"3f8183dc",
  3046 => x"0b880508",
  3047 => x"841108fc",
  3048 => x"06707b31",
  3049 => x"9fef05e0",
  3050 => x"8006e080",
  3051 => x"05565653",
  3052 => x"a0807424",
  3053 => x"94388052",
  3054 => x"7551ff9c",
  3055 => x"3f8183e4",
  3056 => x"08155372",
  3057 => x"b0082e8f",
  3058 => x"387551ff",
  3059 => x"8a3f8053",
  3060 => x"72b00c87",
  3061 => x"3d0d0473",
  3062 => x"30527551",
  3063 => x"fefa3fb0",
  3064 => x"08ff2ea8",
  3065 => x"388183dc",
  3066 => x"0b880508",
  3067 => x"75753181",
  3068 => x"0784120c",
  3069 => x"538183a0",
  3070 => x"08743181",
  3071 => x"83a00c75",
  3072 => x"51fed43f",
  3073 => x"810bb00c",
  3074 => x"873d0d04",
  3075 => x"80527551",
  3076 => x"fec63f81",
  3077 => x"83dc0b88",
  3078 => x"0508b008",
  3079 => x"71315653",
  3080 => x"8f7525ff",
  3081 => x"a438b008",
  3082 => x"8183d008",
  3083 => x"318183a0",
  3084 => x"0c748107",
  3085 => x"84140c75",
  3086 => x"51fe9c3f",
  3087 => x"8053ff90",
  3088 => x"39f63d0d",
  3089 => x"7c7e545b",
  3090 => x"72802e82",
  3091 => x"83387a51",
  3092 => x"fe843ff8",
  3093 => x"13841108",
  3094 => x"70fe0670",
  3095 => x"13841108",
  3096 => x"fc065d58",
  3097 => x"59545881",
  3098 => x"83e40875",
  3099 => x"2e82de38",
  3100 => x"7884160c",
  3101 => x"80738106",
  3102 => x"545a727a",
  3103 => x"2e81d538",
  3104 => x"78158411",
  3105 => x"08810651",
  3106 => x"5372a038",
  3107 => x"78175779",
  3108 => x"81e63888",
  3109 => x"15085372",
  3110 => x"8183e42e",
  3111 => x"82f9388c",
  3112 => x"1508708c",
  3113 => x"150c7388",
  3114 => x"120c5676",
  3115 => x"81078419",
  3116 => x"0c761877",
  3117 => x"710c5379",
  3118 => x"81913883",
  3119 => x"ff772781",
  3120 => x"c8387689",
  3121 => x"2a77832a",
  3122 => x"56537280",
  3123 => x"2ebf3876",
  3124 => x"862ab805",
  3125 => x"55847327",
  3126 => x"b43880db",
  3127 => x"13559473",
  3128 => x"27ab3876",
  3129 => x"8c2a80ee",
  3130 => x"055580d4",
  3131 => x"73279e38",
  3132 => x"768f2a80",
  3133 => x"f7055582",
  3134 => x"d4732791",
  3135 => x"3876922a",
  3136 => x"80fc0555",
  3137 => x"8ad47327",
  3138 => x"843880fe",
  3139 => x"55741010",
  3140 => x"108183dc",
  3141 => x"05881108",
  3142 => x"55567376",
  3143 => x"2e82b338",
  3144 => x"841408fc",
  3145 => x"06537673",
  3146 => x"278d3888",
  3147 => x"14085473",
  3148 => x"762e0981",
  3149 => x"06ea388c",
  3150 => x"1408708c",
  3151 => x"1a0c7488",
  3152 => x"1a0c7888",
  3153 => x"120c5677",
  3154 => x"8c150c7a",
  3155 => x"51fc883f",
  3156 => x"8c3d0d04",
  3157 => x"77087871",
  3158 => x"31597705",
  3159 => x"88190854",
  3160 => x"57728183",
  3161 => x"e42e80e0",
  3162 => x"388c1808",
  3163 => x"708c150c",
  3164 => x"7388120c",
  3165 => x"56fe8939",
  3166 => x"8815088c",
  3167 => x"1608708c",
  3168 => x"130c5788",
  3169 => x"170cfea3",
  3170 => x"3976832a",
  3171 => x"70545580",
  3172 => x"75248198",
  3173 => x"3872822c",
  3174 => x"81712b81",
  3175 => x"83e00807",
  3176 => x"8183dc0b",
  3177 => x"84050c53",
  3178 => x"74101010",
  3179 => x"8183dc05",
  3180 => x"88110855",
  3181 => x"56758c19",
  3182 => x"0c738819",
  3183 => x"0c778817",
  3184 => x"0c778c15",
  3185 => x"0cff8439",
  3186 => x"815afdb4",
  3187 => x"39781773",
  3188 => x"81065457",
  3189 => x"72983877",
  3190 => x"08787131",
  3191 => x"5977058c",
  3192 => x"1908881a",
  3193 => x"08718c12",
  3194 => x"0c88120c",
  3195 => x"57577681",
  3196 => x"0784190c",
  3197 => x"778183dc",
  3198 => x"0b88050c",
  3199 => x"8183d808",
  3200 => x"7726fec7",
  3201 => x"388183d4",
  3202 => x"08527a51",
  3203 => x"fafe3f7a",
  3204 => x"51fac43f",
  3205 => x"feba3981",
  3206 => x"788c150c",
  3207 => x"7888150c",
  3208 => x"738c1a0c",
  3209 => x"73881a0c",
  3210 => x"5afd8039",
  3211 => x"83157082",
  3212 => x"2c81712b",
  3213 => x"8183e008",
  3214 => x"078183dc",
  3215 => x"0b84050c",
  3216 => x"51537410",
  3217 => x"10108183",
  3218 => x"dc058811",
  3219 => x"085556fe",
  3220 => x"e4397453",
  3221 => x"807524a7",
  3222 => x"3872822c",
  3223 => x"81712b81",
  3224 => x"83e00807",
  3225 => x"8183dc0b",
  3226 => x"84050c53",
  3227 => x"758c190c",
  3228 => x"7388190c",
  3229 => x"7788170c",
  3230 => x"778c150c",
  3231 => x"fdcd3983",
  3232 => x"1570822c",
  3233 => x"81712b81",
  3234 => x"83e00807",
  3235 => x"8183dc0b",
  3236 => x"84050c51",
  3237 => x"53d63981",
  3238 => x"0bb00c04",
  3239 => x"803d0d72",
  3240 => x"812e8938",
  3241 => x"800bb00c",
  3242 => x"823d0d04",
  3243 => x"7351b23f",
  3244 => x"fe3d0d81",
  3245 => x"a4b80851",
  3246 => x"708a3881",
  3247 => x"a4c07081",
  3248 => x"a4b80c51",
  3249 => x"70751252",
  3250 => x"52ff5370",
  3251 => x"87fb8080",
  3252 => x"26883870",
  3253 => x"81a4b80c",
  3254 => x"715372b0",
  3255 => x"0c843d0d",
  3256 => x"0400ff39",
  3257 => x"68656c70",
  3258 => x"00000000",
  3259 => x"73797374",
  3260 => x"656d2072",
  3261 => x"65736574",
  3262 => x"00000000",
  3263 => x"72657365",
  3264 => x"74000000",
  3265 => x"73686f77",
  3266 => x"20737973",
  3267 => x"74656d20",
  3268 => x"696e666f",
  3269 => x"203c7665",
  3270 => x"72626f73",
  3271 => x"653e0000",
  3272 => x"73797369",
  3273 => x"6e666f00",
  3274 => x"72656e61",
  3275 => x"20636f6e",
  3276 => x"74726f6c",
  3277 => x"6c657220",
  3278 => x"73746174",
  3279 => x"75730000",
  3280 => x"72656e61",
  3281 => x"20737461",
  3282 => x"74757300",
  3283 => x"3c636861",
  3284 => x"6e6e656c",
  3285 => x"3e203c68",
  3286 => x"6967683e",
  3287 => x"203c6c6f",
  3288 => x"775f636f",
  3289 => x"6e666967",
  3290 => x"3e000000",
  3291 => x"636f6e66",
  3292 => x"69670000",
  3293 => x"646f2063",
  3294 => x"6f6d706c",
  3295 => x"65746520",
  3296 => x"64656d6f",
  3297 => x"20636f6e",
  3298 => x"66696720",
  3299 => x"666f7220",
  3300 => x"52454e41",
  3301 => x"00000000",
  3302 => x"64656d6f",
  3303 => x"00000000",
  3304 => x"73657420",
  3305 => x"52454e41",
  3306 => x"20746f20",
  3307 => x"706f7765",
  3308 => x"7220646f",
  3309 => x"776e206d",
  3310 => x"6f646500",
  3311 => x"706f6666",
  3312 => x"00000000",
  3313 => x"73657420",
  3314 => x"72656e61",
  3315 => x"20636861",
  3316 => x"6e6e656c",
  3317 => x"20302074",
  3318 => x"6f20666f",
  3319 => x"6c6c6f77",
  3320 => x"6572206d",
  3321 => x"6f646500",
  3322 => x"666f6c6c",
  3323 => x"6f770000",
  3324 => x"3c74696d",
  3325 => x"653e2061",
  3326 => x"63746976",
  3327 => x"61746520",
  3328 => x"52454e41",
  3329 => x"00000000",
  3330 => x"61637175",
  3331 => x"69726500",
  3332 => x"73657420",
  3333 => x"52454e41",
  3334 => x"20636f6e",
  3335 => x"74726f6c",
  3336 => x"6c657220",
  3337 => x"746f2049",
  3338 => x"444c4500",
  3339 => x"73746f70",
  3340 => x"00000000",
  3341 => x"7072696e",
  3342 => x"74207472",
  3343 => x"69676765",
  3344 => x"72206368",
  3345 => x"61696e73",
  3346 => x"00000000",
  3347 => x"63686169",
  3348 => x"6e730000",
  3349 => x"7072696e",
  3350 => x"74207361",
  3351 => x"6d706c65",
  3352 => x"64205245",
  3353 => x"4e412074",
  3354 => x"6f6b656e",
  3355 => x"73000000",
  3356 => x"746f6b65",
  3357 => x"6e000000",
  3358 => x"74726f75",
  3359 => x"626c6573",
  3360 => x"65617263",
  3361 => x"68205245",
  3362 => x"4e410000",
  3363 => x"74726f75",
  3364 => x"626c6500",
  3365 => x"696e6974",
  3366 => x"616c697a",
  3367 => x"65204444",
  3368 => x"53206368",
  3369 => x"6970203c",
  3370 => x"66726571",
  3371 => x"2074756e",
  3372 => x"696e6720",
  3373 => x"776f7264",
  3374 => x"3e000000",
  3375 => x"64647369",
  3376 => x"6e697400",
  3377 => x"72656164",
  3378 => x"20646473",
  3379 => x"20726567",
  3380 => x"69737465",
  3381 => x"72730000",
  3382 => x"64647369",
  3383 => x"6e666f00",
  3384 => x"72756e6e",
  3385 => x"696e6720",
  3386 => x"6c696768",
  3387 => x"74000000",
  3388 => x"72756e00",
  3389 => x"63686563",
  3390 => x"6b204932",
  3391 => x"43206164",
  3392 => x"64726573",
  3393 => x"73000000",
  3394 => x"69326300",
  3395 => x"72656164",
  3396 => x"20454550",
  3397 => x"524f4d20",
  3398 => x"3c627573",
  3399 => x"3e203c69",
  3400 => x"32635f61",
  3401 => x"6464723e",
  3402 => x"203c6c65",
  3403 => x"6e677468",
  3404 => x"3e000000",
  3405 => x"65657072",
  3406 => x"6f6d0000",
  3407 => x"72656164",
  3408 => x"20616463",
  3409 => x"2076616c",
  3410 => x"75650000",
  3411 => x"61646300",
  3412 => x"67656e65",
  3413 => x"72617465",
  3414 => x"20746573",
  3415 => x"7420696d",
  3416 => x"70756c73",
  3417 => x"65000000",
  3418 => x"74657374",
  3419 => x"67656e00",
  3420 => x"616c6961",
  3421 => x"7320666f",
  3422 => x"72207800",
  3423 => x"6d656d00",
  3424 => x"77726974",
  3425 => x"6520776f",
  3426 => x"7264203c",
  3427 => x"61646472",
  3428 => x"3e203c6c",
  3429 => x"656e6774",
  3430 => x"683e203c",
  3431 => x"76616c75",
  3432 => x"65287329",
  3433 => x"3e000000",
  3434 => x"776d656d",
  3435 => x"00000000",
  3436 => x"6558616d",
  3437 => x"696e6520",
  3438 => x"6d656d6f",
  3439 => x"7279203c",
  3440 => x"61646472",
  3441 => x"3e203c6c",
  3442 => x"656e6774",
  3443 => x"683e0000",
  3444 => x"78000000",
  3445 => x"636c6561",
  3446 => x"72207363",
  3447 => x"7265656e",
  3448 => x"00000000",
  3449 => x"636c6561",
  3450 => x"72000000",
  3451 => x"0a0a0000",
  3452 => x"72656e61",
  3453 => x"3320636f",
  3454 => x"6e74726f",
  3455 => x"6c6c6572",
  3456 => x"20626f61",
  3457 => x"72640000",
  3458 => x"20286f6e",
  3459 => x"2073696d",
  3460 => x"290a0000",
  3461 => x"0a485720",
  3462 => x"73796e74",
  3463 => x"68657369",
  3464 => x"7a65643a",
  3465 => x"20000000",
  3466 => x"0a535720",
  3467 => x"636f6d70",
  3468 => x"696c6564",
  3469 => x"2020203a",
  3470 => x"20446563",
  3471 => x"20323120",
  3472 => x"32303131",
  3473 => x"20203135",
  3474 => x"3a30303a",
  3475 => x"35390000",
  3476 => x"0a737973",
  3477 => x"74656d20",
  3478 => x"636c6f63",
  3479 => x"6b20203a",
  3480 => x"20000000",
  3481 => x"204d487a",
  3482 => x"0a000000",
  3483 => x"44454255",
  3484 => x"47204d4f",
  3485 => x"44450000",
  3486 => x"204f4e0a",
  3487 => x"00000000",
  3488 => x"4552524f",
  3489 => x"523a2074",
  3490 => x"6f6f206d",
  3491 => x"75636820",
  3492 => x"636f6d6d",
  3493 => x"616e6473",
  3494 => x"2e0a0000",
  3495 => x"3e200000",
  3496 => x"636f6d6d",
  3497 => x"616e6420",
  3498 => x"6e6f7420",
  3499 => x"666f756e",
  3500 => x"642e0a00",
  3501 => x"73757070",
  3502 => x"6f727465",
  3503 => x"6420636f",
  3504 => x"6d6d616e",
  3505 => x"64733a0a",
  3506 => x"0a000000",
  3507 => x"202d2000",
  3508 => x"76656e64",
  3509 => x"6f723f20",
  3510 => x"20000000",
  3511 => x"485a4452",
  3512 => x"20202020",
  3513 => x"20000000",
  3514 => x"67616973",
  3515 => x"6c657220",
  3516 => x"20000000",
  3517 => x"45534120",
  3518 => x"20202020",
  3519 => x"20000000",
  3520 => x"756e6b6e",
  3521 => x"6f776e20",
  3522 => x"64657669",
  3523 => x"63650000",
  3524 => x"4c656f6e",
  3525 => x"32204d65",
  3526 => x"6d6f7279",
  3527 => x"20436f6e",
  3528 => x"74726f6c",
  3529 => x"6c657200",
  3530 => x"56474120",
  3531 => x"636f6e74",
  3532 => x"726f6c6c",
  3533 => x"65720000",
  3534 => x"53504920",
  3535 => x"4d656d6f",
  3536 => x"72792043",
  3537 => x"6f6e7472",
  3538 => x"6f6c6c65",
  3539 => x"72000000",
  3540 => x"53504920",
  3541 => x"436f6e74",
  3542 => x"726f6c6c",
  3543 => x"65720000",
  3544 => x"414d4241",
  3545 => x"20577261",
  3546 => x"70706572",
  3547 => x"20666f72",
  3548 => x"204f4320",
  3549 => x"4932432d",
  3550 => x"6d617374",
  3551 => x"65720000",
  3552 => x"47522031",
  3553 => x"302f3130",
  3554 => x"30204d62",
  3555 => x"69742045",
  3556 => x"74686572",
  3557 => x"6e657420",
  3558 => x"4d414300",
  3559 => x"47656e65",
  3560 => x"72616c20",
  3561 => x"50757270",
  3562 => x"6f736520",
  3563 => x"492f4f20",
  3564 => x"706f7274",
  3565 => x"00000000",
  3566 => x"4d6f6475",
  3567 => x"6c617220",
  3568 => x"54696d65",
  3569 => x"7220556e",
  3570 => x"69740000",
  3571 => x"4475616c",
  3572 => x"2d706f72",
  3573 => x"74204148",
  3574 => x"42205352",
  3575 => x"414d206d",
  3576 => x"6f64756c",
  3577 => x"65000000",
  3578 => x"47656e65",
  3579 => x"72696320",
  3580 => x"55415254",
  3581 => x"00000000",
  3582 => x"4148422f",
  3583 => x"41504220",
  3584 => x"42726964",
  3585 => x"67650000",
  3586 => x"64696666",
  3587 => x"6572656e",
  3588 => x"7469616c",
  3589 => x"20637572",
  3590 => x"72656e74",
  3591 => x"206d6f6e",
  3592 => x"69746f72",
  3593 => x"00000000",
  3594 => x"64656275",
  3595 => x"67207472",
  3596 => x"61636572",
  3597 => x"206d656d",
  3598 => x"6f727900",
  3599 => x"4541444f",
  3600 => x"47533130",
  3601 => x"32206469",
  3602 => x"73706c61",
  3603 => x"79206472",
  3604 => x"69766572",
  3605 => x"00000000",
  3606 => x"64656275",
  3607 => x"67206275",
  3608 => x"66666572",
  3609 => x"20636f6e",
  3610 => x"74726f6c",
  3611 => x"00000000",
  3612 => x"52454e41",
  3613 => x"3320636f",
  3614 => x"6e74726f",
  3615 => x"6c6c6572",
  3616 => x"00000000",
  3617 => x"53465020",
  3618 => x"636f6e74",
  3619 => x"726f6c6c",
  3620 => x"65720000",
  3621 => x"5a505520",
  3622 => x"4d656d6f",
  3623 => x"72792077",
  3624 => x"72617070",
  3625 => x"65720000",
  3626 => x"5a505520",
  3627 => x"41484220",
  3628 => x"57726170",
  3629 => x"70657200",
  3630 => x"6265616d",
  3631 => x"20706f73",
  3632 => x"6974696f",
  3633 => x"6e206d6f",
  3634 => x"6e69746f",
  3635 => x"72000000",
  3636 => x"74726967",
  3637 => x"67657220",
  3638 => x"67656e65",
  3639 => x"7261746f",
  3640 => x"72000000",
  3641 => x"64656275",
  3642 => x"6720636f",
  3643 => x"6e736f6c",
  3644 => x"65000000",
  3645 => x"44434d20",
  3646 => x"70686173",
  3647 => x"65207368",
  3648 => x"69667420",
  3649 => x"636f6e74",
  3650 => x"726f6c00",
  3651 => x"20206170",
  3652 => x"62736c76",
  3653 => x"00000000",
  3654 => x"76656e64",
  3655 => x"20307800",
  3656 => x"64657620",
  3657 => x"30780000",
  3658 => x"76657220",
  3659 => x"00000000",
  3660 => x"69727120",
  3661 => x"00000000",
  3662 => x"61646472",
  3663 => x"20307800",
  3664 => x"6168626d",
  3665 => x"73740000",
  3666 => x"61686273",
  3667 => x"6c760000",
  3668 => x"00000f46",
  3669 => x"00001017",
  3670 => x"0000100c",
  3671 => x"00001043",
  3672 => x"00001038",
  3673 => x"0000102d",
  3674 => x"00001022",
  3675 => x"00000feb",
  3676 => x"00000fe0",
  3677 => x"00000fd5",
  3678 => x"00000fca",
  3679 => x"00001001",
  3680 => x"00000ff6",
  3681 => x"00000fbf",
  3682 => x"00000f46",
  3683 => x"00000f46",
  3684 => x"00000f46",
  3685 => x"00000f46",
  3686 => x"00000f46",
  3687 => x"00000fb4",
  3688 => x"00000f46",
  3689 => x"00000f46",
  3690 => x"00000fa9",
  3691 => x"00000f46",
  3692 => x"00000f9e",
  3693 => x"00000f46",
  3694 => x"00000f46",
  3695 => x"00000f46",
  3696 => x"00000f46",
  3697 => x"00000f46",
  3698 => x"00000f46",
  3699 => x"00000f46",
  3700 => x"00000f46",
  3701 => x"00000f93",
  3702 => x"00000f46",
  3703 => x"00000f46",
  3704 => x"00000f88",
  3705 => x"00000f46",
  3706 => x"00000f46",
  3707 => x"00000f46",
  3708 => x"00000f46",
  3709 => x"00000f46",
  3710 => x"00000f46",
  3711 => x"00000f46",
  3712 => x"00000f46",
  3713 => x"00000f46",
  3714 => x"00000f46",
  3715 => x"00000f7d",
  3716 => x"00000f46",
  3717 => x"00000f46",
  3718 => x"00000f46",
  3719 => x"00000f46",
  3720 => x"00000f72",
  3721 => x"00000f46",
  3722 => x"00000f46",
  3723 => x"00000f46",
  3724 => x"00000f46",
  3725 => x"00000f46",
  3726 => x"00000f46",
  3727 => x"00000f46",
  3728 => x"00000f46",
  3729 => x"00000f46",
  3730 => x"00000f46",
  3731 => x"00000f46",
  3732 => x"00000f46",
  3733 => x"00000f46",
  3734 => x"00000f46",
  3735 => x"00000f46",
  3736 => x"00000f46",
  3737 => x"00000f46",
  3738 => x"00000f46",
  3739 => x"00000f46",
  3740 => x"00000f46",
  3741 => x"00000f46",
  3742 => x"00000f46",
  3743 => x"00000f46",
  3744 => x"00000f67",
  3745 => x"00000f46",
  3746 => x"00000f46",
  3747 => x"00000f46",
  3748 => x"00000f46",
  3749 => x"00000f46",
  3750 => x"00000f46",
  3751 => x"00000f46",
  3752 => x"00000f46",
  3753 => x"00000f46",
  3754 => x"00000f46",
  3755 => x"00000f46",
  3756 => x"00000f46",
  3757 => x"00000f46",
  3758 => x"00000f46",
  3759 => x"00000f46",
  3760 => x"00000f46",
  3761 => x"00000f46",
  3762 => x"00000f46",
  3763 => x"00000f46",
  3764 => x"00000f46",
  3765 => x"00000f46",
  3766 => x"00000f46",
  3767 => x"00000f46",
  3768 => x"00000f46",
  3769 => x"00000f46",
  3770 => x"00000f46",
  3771 => x"00000f46",
  3772 => x"00000f5c",
  3773 => x"69326320",
  3774 => x"464d430a",
  3775 => x"00000000",
  3776 => x"61646472",
  3777 => x"6573733a",
  3778 => x"20307800",
  3779 => x"2020202d",
  3780 => x"2d3e2020",
  3781 => x"2041434b",
  3782 => x"0a000000",
  3783 => x"72656164",
  3784 => x"20646174",
  3785 => x"61202800",
  3786 => x"20627974",
  3787 => x"65732920",
  3788 => x"66726f6d",
  3789 => x"20493243",
  3790 => x"2d616464",
  3791 => x"72657373",
  3792 => x"20307800",
  3793 => x"0a307800",
  3794 => x"02020606",
  3795 => x"06040304",
  3796 => x"02020102",
  3797 => x"636f6e74",
  3798 => x"726f6c20",
  3799 => x"2020203a",
  3800 => x"20000000",
  3801 => x"66726571",
  3802 => x"75656e63",
  3803 => x"7920203a",
  3804 => x"20000000",
  3805 => x"75706461",
  3806 => x"74652063",
  3807 => x"6c6b203a",
  3808 => x"20000000",
  3809 => x"72616d70",
  3810 => x"20726174",
  3811 => x"6520203a",
  3812 => x"20000000",
  3813 => x"49206d75",
  3814 => x"6c742072",
  3815 => x"6567203a",
  3816 => x"20000000",
  3817 => x"51206d75",
  3818 => x"6c742072",
  3819 => x"6567203a",
  3820 => x"20000000",
  3821 => x"554e4b4e",
  3822 => x"4f574e00",
  3823 => x"69646c65",
  3824 => x"00000000",
  3825 => x"636f6e66",
  3826 => x"69677572",
  3827 => x"65000000",
  3828 => x"64657465",
  3829 => x"63740000",
  3830 => x"61717569",
  3831 => x"72650000",
  3832 => x"616e616c",
  3833 => x"797a6500",
  3834 => x"64657369",
  3835 => x"72650000",
  3836 => x"72656164",
  3837 => x"6f757400",
  3838 => x"72656164",
  3839 => x"6c616700",
  3840 => x"66617374",
  3841 => x"20747269",
  3842 => x"67676572",
  3843 => x"203a2000",
  3844 => x"0a736c6f",
  3845 => x"77207472",
  3846 => x"69676765",
  3847 => x"72203a20",
  3848 => x"00000000",
  3849 => x"0a6f7665",
  3850 => x"72666c6f",
  3851 => x"77202020",
  3852 => x"20203a20",
  3853 => x"00000000",
  3854 => x"66617374",
  3855 => x"20747269",
  3856 => x"67676572",
  3857 => x"20636861",
  3858 => x"696e3a20",
  3859 => x"30780000",
  3860 => x"0a736c6f",
  3861 => x"77207472",
  3862 => x"69676765",
  3863 => x"72206368",
  3864 => x"61696e3a",
  3865 => x"20307800",
  3866 => x"746f6b65",
  3867 => x"6e733a20",
  3868 => x"00000000",
  3869 => x"00001a77",
  3870 => x"00001a8b",
  3871 => x"00001a4f",
  3872 => x"00001a9f",
  3873 => x"00001ab3",
  3874 => x"00001ac7",
  3875 => x"00001adb",
  3876 => x"00001aef",
  3877 => x"00001b03",
  3878 => x"00001a63",
  3879 => x"30622020",
  3880 => x"20202020",
  3881 => x"20202020",
  3882 => x"20202020",
  3883 => x"20202020",
  3884 => x"20202020",
  3885 => x"20202020",
  3886 => x"20202020",
  3887 => x"20200000",
  3888 => x"20202020",
  3889 => x"20202020",
  3890 => x"00000000",
  3891 => x"79657300",
  3892 => x"6e6f0000",
  3893 => x"00202020",
  3894 => x"20202020",
  3895 => x"20202828",
  3896 => x"28282820",
  3897 => x"20202020",
  3898 => x"20202020",
  3899 => x"20202020",
  3900 => x"20202020",
  3901 => x"20881010",
  3902 => x"10101010",
  3903 => x"10101010",
  3904 => x"10101010",
  3905 => x"10040404",
  3906 => x"04040404",
  3907 => x"04040410",
  3908 => x"10101010",
  3909 => x"10104141",
  3910 => x"41414141",
  3911 => x"01010101",
  3912 => x"01010101",
  3913 => x"01010101",
  3914 => x"01010101",
  3915 => x"01010101",
  3916 => x"10101010",
  3917 => x"10104242",
  3918 => x"42424242",
  3919 => x"02020202",
  3920 => x"02020202",
  3921 => x"02020202",
  3922 => x"02020202",
  3923 => x"02020202",
  3924 => x"10101010",
  3925 => x"20000000",
  3926 => x"00000000",
  3927 => x"00000000",
  3928 => x"00000000",
  3929 => x"00000000",
  3930 => x"00000000",
  3931 => x"00000000",
  3932 => x"00000000",
  3933 => x"00000000",
  3934 => x"00000000",
  3935 => x"00000000",
  3936 => x"00000000",
  3937 => x"00000000",
  3938 => x"00000000",
  3939 => x"00000000",
  3940 => x"00000000",
  3941 => x"00000000",
  3942 => x"00000000",
  3943 => x"00000000",
  3944 => x"00000000",
  3945 => x"00000000",
  3946 => x"00000000",
  3947 => x"00000000",
  3948 => x"00000000",
  3949 => x"00000000",
  3950 => x"00000000",
  3951 => x"00000000",
  3952 => x"00000000",
  3953 => x"00000000",
  3954 => x"00000000",
  3955 => x"00000000",
  3956 => x"00000000",
  3957 => x"00000000",
  3958 => x"43000000",
  3959 => x"00000000",
  3960 => x"00000000",
  3961 => x"80000b00",
  3962 => x"10000000",
  3963 => x"80000d00",
  3964 => x"00ffffff",
  3965 => x"ff00ffff",
  3966 => x"ffff00ff",
  3967 => x"ffffff00",
  3968 => x"00000000",
  3969 => x"00000000",
  3970 => x"80000a00",
  3971 => x"80000400",
  3972 => x"80000200",
  3973 => x"80000100",
  3974 => x"80000004",
  3975 => x"80000000",
  3976 => x"00003e24",
  3977 => x"00000000",
  3978 => x"0000408c",
  3979 => x"000040e8",
  3980 => x"00004144",
  3981 => x"00000000",
  3982 => x"00000000",
  3983 => x"00000000",
  3984 => x"00000000",
  3985 => x"00000000",
  3986 => x"00000000",
  3987 => x"00000000",
  3988 => x"00000000",
  3989 => x"00000000",
  3990 => x"00003dd8",
  3991 => x"00000000",
  3992 => x"00000000",
  3993 => x"00000000",
  3994 => x"00000000",
  3995 => x"00000000",
  3996 => x"00000000",
  3997 => x"00000000",
  3998 => x"00000000",
  3999 => x"00000000",
  4000 => x"00000000",
  4001 => x"00000000",
  4002 => x"00000000",
  4003 => x"00000000",
  4004 => x"00000000",
  4005 => x"00000000",
  4006 => x"00000000",
  4007 => x"00000000",
  4008 => x"00000000",
  4009 => x"00000000",
  4010 => x"00000000",
  4011 => x"00000000",
  4012 => x"00000000",
  4013 => x"00000000",
  4014 => x"00000000",
  4015 => x"00000000",
  4016 => x"00000000",
  4017 => x"00000000",
  4018 => x"00000000",
  4019 => x"00000001",
  4020 => x"330eabcd",
  4021 => x"1234e66d",
  4022 => x"deec0005",
  4023 => x"000b0000",
  4024 => x"00000000",
  4025 => x"00000000",
  4026 => x"00000000",
  4027 => x"00000000",
  4028 => x"00000000",
  4029 => x"00000000",
  4030 => x"00000000",
  4031 => x"00000000",
  4032 => x"00000000",
  4033 => x"00000000",
  4034 => x"00000000",
  4035 => x"00000000",
  4036 => x"00000000",
  4037 => x"00000000",
  4038 => x"00000000",
  4039 => x"00000000",
  4040 => x"00000000",
  4041 => x"00000000",
  4042 => x"00000000",
  4043 => x"00000000",
  4044 => x"00000000",
  4045 => x"00000000",
  4046 => x"00000000",
  4047 => x"00000000",
  4048 => x"00000000",
  4049 => x"00000000",
  4050 => x"00000000",
  4051 => x"00000000",
  4052 => x"00000000",
  4053 => x"00000000",
  4054 => x"00000000",
  4055 => x"00000000",
  4056 => x"00000000",
  4057 => x"00000000",
  4058 => x"00000000",
  4059 => x"00000000",
  4060 => x"00000000",
  4061 => x"00000000",
  4062 => x"00000000",
  4063 => x"00000000",
  4064 => x"00000000",
  4065 => x"00000000",
  4066 => x"00000000",
  4067 => x"00000000",
  4068 => x"00000000",
  4069 => x"00000000",
  4070 => x"00000000",
  4071 => x"00000000",
  4072 => x"00000000",
  4073 => x"00000000",
  4074 => x"00000000",
  4075 => x"00000000",
  4076 => x"00000000",
  4077 => x"00000000",
  4078 => x"00000000",
  4079 => x"00000000",
  4080 => x"00000000",
  4081 => x"00000000",
  4082 => x"00000000",
  4083 => x"00000000",
  4084 => x"00000000",
  4085 => x"00000000",
  4086 => x"00000000",
  4087 => x"00000000",
  4088 => x"00000000",
  4089 => x"00000000",
  4090 => x"00000000",
  4091 => x"00000000",
  4092 => x"00000000",
  4093 => x"00000000",
  4094 => x"00000000",
  4095 => x"00000000",
  4096 => x"00000000",
  4097 => x"00000000",
  4098 => x"00000000",
  4099 => x"00000000",
  4100 => x"00000000",
  4101 => x"00000000",
  4102 => x"00000000",
  4103 => x"00000000",
  4104 => x"00000000",
  4105 => x"00000000",
  4106 => x"00000000",
  4107 => x"00000000",
  4108 => x"00000000",
  4109 => x"00000000",
  4110 => x"00000000",
  4111 => x"00000000",
  4112 => x"00000000",
  4113 => x"00000000",
  4114 => x"00000000",
  4115 => x"00000000",
  4116 => x"00000000",
  4117 => x"00000000",
  4118 => x"00000000",
  4119 => x"00000000",
  4120 => x"00000000",
  4121 => x"00000000",
  4122 => x"00000000",
  4123 => x"00000000",
  4124 => x"00000000",
  4125 => x"00000000",
  4126 => x"00000000",
  4127 => x"00000000",
  4128 => x"00000000",
  4129 => x"00000000",
  4130 => x"00000000",
  4131 => x"00000000",
  4132 => x"00000000",
  4133 => x"00000000",
  4134 => x"00000000",
  4135 => x"00000000",
  4136 => x"00000000",
  4137 => x"00000000",
  4138 => x"00000000",
  4139 => x"00000000",
  4140 => x"00000000",
  4141 => x"00000000",
  4142 => x"00000000",
  4143 => x"00000000",
  4144 => x"00000000",
  4145 => x"00000000",
  4146 => x"00000000",
  4147 => x"00000000",
  4148 => x"00000000",
  4149 => x"00000000",
  4150 => x"00000000",
  4151 => x"00000000",
  4152 => x"00000000",
  4153 => x"00000000",
  4154 => x"00000000",
  4155 => x"00000000",
  4156 => x"00000000",
  4157 => x"00000000",
  4158 => x"00000000",
  4159 => x"00000000",
  4160 => x"00000000",
  4161 => x"00000000",
  4162 => x"00000000",
  4163 => x"00000000",
  4164 => x"00000000",
  4165 => x"00000000",
  4166 => x"00000000",
  4167 => x"00000000",
  4168 => x"00000000",
  4169 => x"00000000",
  4170 => x"00000000",
  4171 => x"00000000",
  4172 => x"00000000",
  4173 => x"00000000",
  4174 => x"00000000",
  4175 => x"00000000",
  4176 => x"00000000",
  4177 => x"00000000",
  4178 => x"00000000",
  4179 => x"00000000",
  4180 => x"00000000",
  4181 => x"00000000",
  4182 => x"00000000",
  4183 => x"00000000",
  4184 => x"00000000",
  4185 => x"00000000",
  4186 => x"00000000",
  4187 => x"00000000",
  4188 => x"00000000",
  4189 => x"00000000",
  4190 => x"00000000",
  4191 => x"00000000",
  4192 => x"00000000",
  4193 => x"00000000",
  4194 => x"00000000",
  4195 => x"00000000",
  4196 => x"00000000",
  4197 => x"00000000",
  4198 => x"00000000",
  4199 => x"00000000",
  4200 => x"00000000",
  4201 => x"00000000",
  4202 => x"00000000",
  4203 => x"00000000",
  4204 => x"00000000",
  4205 => x"00000000",
  4206 => x"00000000",
  4207 => x"00000000",
  4208 => x"00000000",
  4209 => x"00000000",
  4210 => x"00000000",
  4211 => x"00000000",
  4212 => x"ffffffff",
  4213 => x"00000000",
  4214 => x"00020000",
  4215 => x"00000000",
  4216 => x"00000000",
  4217 => x"000041dc",
  4218 => x"000041dc",
  4219 => x"000041e4",
  4220 => x"000041e4",
  4221 => x"000041ec",
  4222 => x"000041ec",
  4223 => x"000041f4",
  4224 => x"000041f4",
  4225 => x"000041fc",
  4226 => x"000041fc",
  4227 => x"00004204",
  4228 => x"00004204",
  4229 => x"0000420c",
  4230 => x"0000420c",
  4231 => x"00004214",
  4232 => x"00004214",
  4233 => x"0000421c",
  4234 => x"0000421c",
  4235 => x"00004224",
  4236 => x"00004224",
  4237 => x"0000422c",
  4238 => x"0000422c",
  4239 => x"00004234",
  4240 => x"00004234",
  4241 => x"0000423c",
  4242 => x"0000423c",
  4243 => x"00004244",
  4244 => x"00004244",
  4245 => x"0000424c",
  4246 => x"0000424c",
  4247 => x"00004254",
  4248 => x"00004254",
  4249 => x"0000425c",
  4250 => x"0000425c",
  4251 => x"00004264",
  4252 => x"00004264",
  4253 => x"0000426c",
  4254 => x"0000426c",
  4255 => x"00004274",
  4256 => x"00004274",
  4257 => x"0000427c",
  4258 => x"0000427c",
  4259 => x"00004284",
  4260 => x"00004284",
  4261 => x"0000428c",
  4262 => x"0000428c",
  4263 => x"00004294",
  4264 => x"00004294",
  4265 => x"0000429c",
  4266 => x"0000429c",
  4267 => x"000042a4",
  4268 => x"000042a4",
  4269 => x"000042ac",
  4270 => x"000042ac",
  4271 => x"000042b4",
  4272 => x"000042b4",
  4273 => x"000042bc",
  4274 => x"000042bc",
  4275 => x"000042c4",
  4276 => x"000042c4",
  4277 => x"000042cc",
  4278 => x"000042cc",
  4279 => x"000042d4",
  4280 => x"000042d4",
  4281 => x"000042dc",
  4282 => x"000042dc",
  4283 => x"000042e4",
  4284 => x"000042e4",
  4285 => x"000042ec",
  4286 => x"000042ec",
  4287 => x"000042f4",
  4288 => x"000042f4",
  4289 => x"000042fc",
  4290 => x"000042fc",
  4291 => x"00004304",
  4292 => x"00004304",
  4293 => x"0000430c",
  4294 => x"0000430c",
  4295 => x"00004314",
  4296 => x"00004314",
  4297 => x"0000431c",
  4298 => x"0000431c",
  4299 => x"00004324",
  4300 => x"00004324",
  4301 => x"0000432c",
  4302 => x"0000432c",
  4303 => x"00004334",
  4304 => x"00004334",
  4305 => x"0000433c",
  4306 => x"0000433c",
  4307 => x"00004344",
  4308 => x"00004344",
  4309 => x"0000434c",
  4310 => x"0000434c",
  4311 => x"00004354",
  4312 => x"00004354",
  4313 => x"0000435c",
  4314 => x"0000435c",
  4315 => x"00004364",
  4316 => x"00004364",
  4317 => x"0000436c",
  4318 => x"0000436c",
  4319 => x"00004374",
  4320 => x"00004374",
  4321 => x"0000437c",
  4322 => x"0000437c",
  4323 => x"00004384",
  4324 => x"00004384",
  4325 => x"0000438c",
  4326 => x"0000438c",
  4327 => x"00004394",
  4328 => x"00004394",
  4329 => x"0000439c",
  4330 => x"0000439c",
  4331 => x"000043a4",
  4332 => x"000043a4",
  4333 => x"000043ac",
  4334 => x"000043ac",
  4335 => x"000043b4",
  4336 => x"000043b4",
  4337 => x"000043bc",
  4338 => x"000043bc",
  4339 => x"000043c4",
  4340 => x"000043c4",
  4341 => x"000043cc",
  4342 => x"000043cc",
  4343 => x"000043d4",
  4344 => x"000043d4",
  4345 => x"000043dc",
  4346 => x"000043dc",
  4347 => x"000043e4",
  4348 => x"000043e4",
  4349 => x"000043ec",
  4350 => x"000043ec",
  4351 => x"000043f4",
  4352 => x"000043f4",
  4353 => x"000043fc",
  4354 => x"000043fc",
  4355 => x"00004404",
  4356 => x"00004404",
  4357 => x"0000440c",
  4358 => x"0000440c",
  4359 => x"00004414",
  4360 => x"00004414",
  4361 => x"0000441c",
  4362 => x"0000441c",
  4363 => x"00004424",
  4364 => x"00004424",
  4365 => x"0000442c",
  4366 => x"0000442c",
  4367 => x"00004434",
  4368 => x"00004434",
  4369 => x"0000443c",
  4370 => x"0000443c",
  4371 => x"00004444",
  4372 => x"00004444",
  4373 => x"0000444c",
  4374 => x"0000444c",
  4375 => x"00004454",
  4376 => x"00004454",
  4377 => x"0000445c",
  4378 => x"0000445c",
  4379 => x"00004464",
  4380 => x"00004464",
  4381 => x"0000446c",
  4382 => x"0000446c",
  4383 => x"00004474",
  4384 => x"00004474",
  4385 => x"0000447c",
  4386 => x"0000447c",
  4387 => x"00004484",
  4388 => x"00004484",
  4389 => x"0000448c",
  4390 => x"0000448c",
  4391 => x"00004494",
  4392 => x"00004494",
  4393 => x"0000449c",
  4394 => x"0000449c",
  4395 => x"000044a4",
  4396 => x"000044a4",
  4397 => x"000044ac",
  4398 => x"000044ac",
  4399 => x"000044b4",
  4400 => x"000044b4",
  4401 => x"000044bc",
  4402 => x"000044bc",
  4403 => x"000044c4",
  4404 => x"000044c4",
  4405 => x"000044cc",
  4406 => x"000044cc",
  4407 => x"000044d4",
  4408 => x"000044d4",
  4409 => x"000044dc",
  4410 => x"000044dc",
  4411 => x"000044e4",
  4412 => x"000044e4",
  4413 => x"000044ec",
  4414 => x"000044ec",
  4415 => x"000044f4",
  4416 => x"000044f4",
  4417 => x"000044fc",
  4418 => x"000044fc",
  4419 => x"00004504",
  4420 => x"00004504",
  4421 => x"0000450c",
  4422 => x"0000450c",
  4423 => x"00004514",
  4424 => x"00004514",
  4425 => x"0000451c",
  4426 => x"0000451c",
  4427 => x"00004524",
  4428 => x"00004524",
  4429 => x"0000452c",
  4430 => x"0000452c",
  4431 => x"00004534",
  4432 => x"00004534",
  4433 => x"0000453c",
  4434 => x"0000453c",
  4435 => x"00004544",
  4436 => x"00004544",
  4437 => x"0000454c",
  4438 => x"0000454c",
  4439 => x"00004554",
  4440 => x"00004554",
  4441 => x"0000455c",
  4442 => x"0000455c",
  4443 => x"00004564",
  4444 => x"00004564",
  4445 => x"0000456c",
  4446 => x"0000456c",
  4447 => x"00004574",
  4448 => x"00004574",
  4449 => x"0000457c",
  4450 => x"0000457c",
  4451 => x"00004584",
  4452 => x"00004584",
  4453 => x"0000458c",
  4454 => x"0000458c",
  4455 => x"00004594",
  4456 => x"00004594",
  4457 => x"0000459c",
  4458 => x"0000459c",
  4459 => x"000045a4",
  4460 => x"000045a4",
  4461 => x"000045ac",
  4462 => x"000045ac",
  4463 => x"000045b4",
  4464 => x"000045b4",
  4465 => x"000045bc",
  4466 => x"000045bc",
  4467 => x"000045c4",
  4468 => x"000045c4",
  4469 => x"000045cc",
  4470 => x"000045cc",
  4471 => x"000045d4",
  4472 => x"000045d4",
	--others => x"00dead00" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
