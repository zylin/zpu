-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0ba7a40c",
     3 => x"3a0b0b0b",
     4 => x"a4eb0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0ba5ab2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0ba7",
   162 => x"90738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8a",
   171 => x"c42d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8b",
   179 => x"f62d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0ba7a00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f9e",
   257 => x"cb3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104a7",
   280 => x"a008802e",
   281 => x"a138a7a4",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"b78c0c82",
   286 => x"a0800bb7",
   287 => x"900c8290",
   288 => x"800bb794",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0bb7",
   292 => x"8c0cf880",
   293 => x"8082800b",
   294 => x"b7900cf8",
   295 => x"80808480",
   296 => x"0bb7940c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0bb78c",
   300 => x"0c80c0a8",
   301 => x"80940bb7",
   302 => x"900c0b0b",
   303 => x"0ba6fc0b",
   304 => x"b7940c04",
   305 => x"ff3d0db7",
   306 => x"98335170",
   307 => x"a338a7ac",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"a7ac0c70",
   312 => x"2da7ac08",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0bb79834",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0bb7",
   319 => x"8808802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0bb788",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"fd3d0d8a",
   330 => x"54f88080",
   331 => x"908051f8",
   332 => x"80809084",
   333 => x"528a710c",
   334 => x"90720c90",
   335 => x"710c7108",
   336 => x"5383fd3f",
   337 => x"8c08028c",
   338 => x"0cf93d0d",
   339 => x"800b8c08",
   340 => x"fc050c8c",
   341 => x"08880508",
   342 => x"8025ab38",
   343 => x"8c088805",
   344 => x"08308c08",
   345 => x"88050c80",
   346 => x"0b8c08f4",
   347 => x"050c8c08",
   348 => x"fc050888",
   349 => x"38810b8c",
   350 => x"08f4050c",
   351 => x"8c08f405",
   352 => x"088c08fc",
   353 => x"050c8c08",
   354 => x"8c050880",
   355 => x"25ab388c",
   356 => x"088c0508",
   357 => x"308c088c",
   358 => x"050c800b",
   359 => x"8c08f005",
   360 => x"0c8c08fc",
   361 => x"05088838",
   362 => x"810b8c08",
   363 => x"f0050c8c",
   364 => x"08f00508",
   365 => x"8c08fc05",
   366 => x"0c80538c",
   367 => x"088c0508",
   368 => x"528c0888",
   369 => x"05085181",
   370 => x"a73f8008",
   371 => x"708c08f8",
   372 => x"050c548c",
   373 => x"08fc0508",
   374 => x"802e8c38",
   375 => x"8c08f805",
   376 => x"08308c08",
   377 => x"f8050c8c",
   378 => x"08f80508",
   379 => x"70800c54",
   380 => x"893d0d8c",
   381 => x"0c048c08",
   382 => x"028c0cfb",
   383 => x"3d0d800b",
   384 => x"8c08fc05",
   385 => x"0c8c0888",
   386 => x"05088025",
   387 => x"93388c08",
   388 => x"88050830",
   389 => x"8c088805",
   390 => x"0c810b8c",
   391 => x"08fc050c",
   392 => x"8c088c05",
   393 => x"0880258c",
   394 => x"388c088c",
   395 => x"0508308c",
   396 => x"088c050c",
   397 => x"81538c08",
   398 => x"8c050852",
   399 => x"8c088805",
   400 => x"0851ad3f",
   401 => x"8008708c",
   402 => x"08f8050c",
   403 => x"548c08fc",
   404 => x"0508802e",
   405 => x"8c388c08",
   406 => x"f8050830",
   407 => x"8c08f805",
   408 => x"0c8c08f8",
   409 => x"05087080",
   410 => x"0c54873d",
   411 => x"0d8c0c04",
   412 => x"8c08028c",
   413 => x"0cfd3d0d",
   414 => x"810b8c08",
   415 => x"fc050c80",
   416 => x"0b8c08f8",
   417 => x"050c8c08",
   418 => x"8c05088c",
   419 => x"08880508",
   420 => x"27ac388c",
   421 => x"08fc0508",
   422 => x"802ea338",
   423 => x"800b8c08",
   424 => x"8c050824",
   425 => x"99388c08",
   426 => x"8c050810",
   427 => x"8c088c05",
   428 => x"0c8c08fc",
   429 => x"0508108c",
   430 => x"08fc050c",
   431 => x"c9398c08",
   432 => x"fc050880",
   433 => x"2e80c938",
   434 => x"8c088c05",
   435 => x"088c0888",
   436 => x"050826a1",
   437 => x"388c0888",
   438 => x"05088c08",
   439 => x"8c050831",
   440 => x"8c088805",
   441 => x"0c8c08f8",
   442 => x"05088c08",
   443 => x"fc050807",
   444 => x"8c08f805",
   445 => x"0c8c08fc",
   446 => x"0508812a",
   447 => x"8c08fc05",
   448 => x"0c8c088c",
   449 => x"0508812a",
   450 => x"8c088c05",
   451 => x"0cffaf39",
   452 => x"8c089005",
   453 => x"08802e8f",
   454 => x"388c0888",
   455 => x"0508708c",
   456 => x"08f4050c",
   457 => x"518d398c",
   458 => x"08f80508",
   459 => x"708c08f4",
   460 => x"050c518c",
   461 => x"08f40508",
   462 => x"800c853d",
   463 => x"0d8c0c04",
   464 => x"803d0d86",
   465 => x"5182fd3f",
   466 => x"815196dc",
   467 => x"3ffd3d0d",
   468 => x"755384d8",
   469 => x"1308802e",
   470 => x"8a388053",
   471 => x"72800c85",
   472 => x"3d0d0481",
   473 => x"80527251",
   474 => x"83d23f80",
   475 => x"0884d814",
   476 => x"0cff5380",
   477 => x"08802ee4",
   478 => x"38800854",
   479 => x"9f538074",
   480 => x"70840556",
   481 => x"0cff1353",
   482 => x"807324ce",
   483 => x"38807470",
   484 => x"8405560c",
   485 => x"ff135372",
   486 => x"8025e338",
   487 => x"ffbc39fd",
   488 => x"3d0d7577",
   489 => x"55539f74",
   490 => x"278d3896",
   491 => x"730cff52",
   492 => x"71800c85",
   493 => x"3d0d0484",
   494 => x"d8130852",
   495 => x"71802e93",
   496 => x"38731010",
   497 => x"12700879",
   498 => x"720c5152",
   499 => x"71800c85",
   500 => x"3d0d0472",
   501 => x"51fef63f",
   502 => x"ff528008",
   503 => x"d33884d8",
   504 => x"13087410",
   505 => x"10117008",
   506 => x"7a720c51",
   507 => x"5152dd39",
   508 => x"f93d0d79",
   509 => x"7b585676",
   510 => x"9f2680e8",
   511 => x"3884d816",
   512 => x"08547380",
   513 => x"2eaa3876",
   514 => x"10101470",
   515 => x"08555573",
   516 => x"802eba38",
   517 => x"80587381",
   518 => x"2e8f3873",
   519 => x"ff2ea338",
   520 => x"80750c76",
   521 => x"51732d80",
   522 => x"5877800c",
   523 => x"893d0d04",
   524 => x"7551fe99",
   525 => x"3fff5880",
   526 => x"08ef3884",
   527 => x"d8160854",
   528 => x"c6399676",
   529 => x"0c810b80",
   530 => x"0c893d0d",
   531 => x"04755181",
   532 => x"e73f7653",
   533 => x"80085275",
   534 => x"5181a93f",
   535 => x"8008800c",
   536 => x"893d0d04",
   537 => x"96760cff",
   538 => x"0b800c89",
   539 => x"3d0d04fc",
   540 => x"3d0d7678",
   541 => x"5653ff54",
   542 => x"749f26b1",
   543 => x"3884d813",
   544 => x"08527180",
   545 => x"2eae3874",
   546 => x"10101270",
   547 => x"08535381",
   548 => x"5471802e",
   549 => x"98388254",
   550 => x"71ff2e91",
   551 => x"38835471",
   552 => x"812e8a38",
   553 => x"80730c74",
   554 => x"51712d80",
   555 => x"5473800c",
   556 => x"863d0d04",
   557 => x"7251fd95",
   558 => x"3f8008f1",
   559 => x"3884d813",
   560 => x"0852c439",
   561 => x"ff3d0d73",
   562 => x"52a7b008",
   563 => x"51fea13f",
   564 => x"833d0d04",
   565 => x"fe3d0d75",
   566 => x"537452a7",
   567 => x"b00851fd",
   568 => x"be3f843d",
   569 => x"0d04803d",
   570 => x"0da7b008",
   571 => x"51fcde3f",
   572 => x"823d0d04",
   573 => x"ff3d0d73",
   574 => x"52a7b008",
   575 => x"51fef03f",
   576 => x"833d0d04",
   577 => x"fc3d0d80",
   578 => x"0bb7a40c",
   579 => x"78527751",
   580 => x"92973f80",
   581 => x"08548008",
   582 => x"ff2e8838",
   583 => x"73800c86",
   584 => x"3d0d04b7",
   585 => x"a4085574",
   586 => x"802ef138",
   587 => x"7675710c",
   588 => x"5373800c",
   589 => x"863d0d04",
   590 => x"91ea3f04",
   591 => x"f33d0d7f",
   592 => x"618b1170",
   593 => x"f8065c55",
   594 => x"555e7296",
   595 => x"26833890",
   596 => x"59807924",
   597 => x"747a2607",
   598 => x"53805472",
   599 => x"742e0981",
   600 => x"0680ca38",
   601 => x"7d518b96",
   602 => x"3f7883f7",
   603 => x"2680c538",
   604 => x"78832a70",
   605 => x"101010ae",
   606 => x"ec058c11",
   607 => x"0859595a",
   608 => x"76782e83",
   609 => x"a7388417",
   610 => x"08fc0656",
   611 => x"8c170888",
   612 => x"1808718c",
   613 => x"120c8812",
   614 => x"0c587517",
   615 => x"84110881",
   616 => x"0784120c",
   617 => x"537d518a",
   618 => x"d63f8817",
   619 => x"5473800c",
   620 => x"8f3d0d04",
   621 => x"78892a79",
   622 => x"832a5b53",
   623 => x"72802ebf",
   624 => x"3878862a",
   625 => x"b8055a84",
   626 => x"7327b438",
   627 => x"80db135a",
   628 => x"947327ab",
   629 => x"38788c2a",
   630 => x"80ee055a",
   631 => x"80d47327",
   632 => x"9e38788f",
   633 => x"2a80f705",
   634 => x"5a82d473",
   635 => x"27913878",
   636 => x"922a80fc",
   637 => x"055a8ad4",
   638 => x"73278438",
   639 => x"80fe5a79",
   640 => x"101010ae",
   641 => x"ec058c11",
   642 => x"08585576",
   643 => x"752ea338",
   644 => x"841708fc",
   645 => x"06707a31",
   646 => x"5556738f",
   647 => x"2488aa38",
   648 => x"738025fe",
   649 => x"e7388c17",
   650 => x"08577675",
   651 => x"2e098106",
   652 => x"df38811a",
   653 => x"5aaefc08",
   654 => x"5776aef4",
   655 => x"2e82b738",
   656 => x"841708fc",
   657 => x"06707a31",
   658 => x"5556738f",
   659 => x"2481f338",
   660 => x"aef40baf",
   661 => x"800caef4",
   662 => x"0baefc0c",
   663 => x"738025fe",
   664 => x"b93883ff",
   665 => x"762783d2",
   666 => x"3875892a",
   667 => x"76832a55",
   668 => x"5372802e",
   669 => x"bf387586",
   670 => x"2ab80554",
   671 => x"847327b4",
   672 => x"3880db13",
   673 => x"54947327",
   674 => x"ab38758c",
   675 => x"2a80ee05",
   676 => x"5480d473",
   677 => x"279e3875",
   678 => x"8f2a80f7",
   679 => x"055482d4",
   680 => x"73279138",
   681 => x"75922a80",
   682 => x"fc05548a",
   683 => x"d4732784",
   684 => x"3880fe54",
   685 => x"73101010",
   686 => x"aeec0588",
   687 => x"11085658",
   688 => x"74782e86",
   689 => x"af388415",
   690 => x"08fc0653",
   691 => x"7573278d",
   692 => x"38881508",
   693 => x"5574782e",
   694 => x"098106ea",
   695 => x"388c1508",
   696 => x"aeec0b84",
   697 => x"0508718c",
   698 => x"1a0c7688",
   699 => x"1a0c7888",
   700 => x"130c788c",
   701 => x"180c5d58",
   702 => x"7953807a",
   703 => x"2483d738",
   704 => x"72822c81",
   705 => x"712b5c53",
   706 => x"7a7c2681",
   707 => x"93387b7b",
   708 => x"06537282",
   709 => x"e33879fc",
   710 => x"0684055a",
   711 => x"7a10707d",
   712 => x"06545b72",
   713 => x"82d23884",
   714 => x"1a5af139",
   715 => x"88178c11",
   716 => x"08585876",
   717 => x"782e0981",
   718 => x"06fccb38",
   719 => x"821a5afd",
   720 => x"f4397817",
   721 => x"79810784",
   722 => x"190c70af",
   723 => x"800c70ae",
   724 => x"fc0caef4",
   725 => x"0b8c120c",
   726 => x"8c110888",
   727 => x"120c7481",
   728 => x"0784120c",
   729 => x"74117571",
   730 => x"0c51537d",
   731 => x"5187903f",
   732 => x"881754fc",
   733 => x"b839aeec",
   734 => x"0b840508",
   735 => x"7a545c79",
   736 => x"8025fefc",
   737 => x"3882cf39",
   738 => x"7a097c06",
   739 => x"70aeec0b",
   740 => x"84050c5c",
   741 => x"7a105b7a",
   742 => x"7c268538",
   743 => x"7a859a38",
   744 => x"aeec0b88",
   745 => x"05087084",
   746 => x"1208fc06",
   747 => x"707c317c",
   748 => x"72268f72",
   749 => x"25075757",
   750 => x"5c5d5572",
   751 => x"802e80d7",
   752 => x"38797a16",
   753 => x"aee4081b",
   754 => x"90115a55",
   755 => x"575baee0",
   756 => x"08ff2e88",
   757 => x"38a08f13",
   758 => x"e0800657",
   759 => x"76527d51",
   760 => x"869e3f80",
   761 => x"08548008",
   762 => x"ff2e8f38",
   763 => x"80087627",
   764 => x"828f3874",
   765 => x"aeec2e82",
   766 => x"8838aeec",
   767 => x"0b880508",
   768 => x"55841508",
   769 => x"fc06707a",
   770 => x"317a7226",
   771 => x"8f722507",
   772 => x"52555372",
   773 => x"83d13874",
   774 => x"79810784",
   775 => x"170c7916",
   776 => x"70aeec0b",
   777 => x"88050c75",
   778 => x"81078412",
   779 => x"0c547e52",
   780 => x"5785cc3f",
   781 => x"881754fa",
   782 => x"f4397583",
   783 => x"2a705454",
   784 => x"80742481",
   785 => x"97387282",
   786 => x"2c81712b",
   787 => x"aef00807",
   788 => x"70aeec0b",
   789 => x"84050c75",
   790 => x"101010ae",
   791 => x"ec058811",
   792 => x"08585a5d",
   793 => x"53778c18",
   794 => x"0c748818",
   795 => x"0c768819",
   796 => x"0c768c16",
   797 => x"0cfd8139",
   798 => x"797a1010",
   799 => x"10aeec05",
   800 => x"7057595d",
   801 => x"8c150857",
   802 => x"76752ea3",
   803 => x"38841708",
   804 => x"fc06707a",
   805 => x"31555673",
   806 => x"8f2483b6",
   807 => x"38738025",
   808 => x"83ea388c",
   809 => x"17085776",
   810 => x"752e0981",
   811 => x"06df3888",
   812 => x"15811b70",
   813 => x"8306555b",
   814 => x"5572c938",
   815 => x"7c830653",
   816 => x"72802efd",
   817 => x"c338ff1d",
   818 => x"f819595d",
   819 => x"88180878",
   820 => x"2eea38fd",
   821 => x"bf39831a",
   822 => x"53fca539",
   823 => x"83147082",
   824 => x"2c81712b",
   825 => x"aef00807",
   826 => x"70aeec0b",
   827 => x"84050c76",
   828 => x"101010ae",
   829 => x"ec058811",
   830 => x"08595b5e",
   831 => x"5153fee5",
   832 => x"39aeb008",
   833 => x"17588008",
   834 => x"762e8187",
   835 => x"38aee008",
   836 => x"ff2e83d8",
   837 => x"38737631",
   838 => x"18aeb00c",
   839 => x"73870670",
   840 => x"57537280",
   841 => x"2e883888",
   842 => x"73317015",
   843 => x"55567614",
   844 => x"9fff06a0",
   845 => x"80713117",
   846 => x"70547f53",
   847 => x"575383c0",
   848 => x"3f800853",
   849 => x"8008ff2e",
   850 => x"819638ae",
   851 => x"b0081670",
   852 => x"aeb00c74",
   853 => x"75aeec0b",
   854 => x"88050c74",
   855 => x"76311870",
   856 => x"81075155",
   857 => x"56587bae",
   858 => x"ec2e838b",
   859 => x"38798f26",
   860 => x"82be3881",
   861 => x"0b84150c",
   862 => x"841508fc",
   863 => x"06707a31",
   864 => x"7a72268f",
   865 => x"72250752",
   866 => x"55537280",
   867 => x"2efd8838",
   868 => x"80d53980",
   869 => x"089fff06",
   870 => x"5372fef1",
   871 => x"3877aeb0",
   872 => x"0caeec0b",
   873 => x"8805087b",
   874 => x"18810784",
   875 => x"120c55ae",
   876 => x"dc087827",
   877 => x"853877ae",
   878 => x"dc0caed8",
   879 => x"087827fc",
   880 => x"c03877ae",
   881 => x"d80c8415",
   882 => x"08fc0670",
   883 => x"7a317a72",
   884 => x"268f7225",
   885 => x"07525553",
   886 => x"72802efc",
   887 => x"ba388839",
   888 => x"80745456",
   889 => x"fee5397d",
   890 => x"5182943f",
   891 => x"800b800c",
   892 => x"8f3d0d04",
   893 => x"73538074",
   894 => x"24a73872",
   895 => x"822c8171",
   896 => x"2baef008",
   897 => x"0770aeec",
   898 => x"0b84050c",
   899 => x"5d53778c",
   900 => x"180c7488",
   901 => x"180c7688",
   902 => x"190c768c",
   903 => x"160cf9d8",
   904 => x"39831470",
   905 => x"822c8171",
   906 => x"2baef008",
   907 => x"0770aeec",
   908 => x"0b84050c",
   909 => x"5e5153d6",
   910 => x"397b7b06",
   911 => x"5372fcb8",
   912 => x"38841a7b",
   913 => x"105c5af1",
   914 => x"39ff1a81",
   915 => x"11515af7",
   916 => x"e4397817",
   917 => x"79810784",
   918 => x"190c8c18",
   919 => x"08881908",
   920 => x"718c120c",
   921 => x"88120c59",
   922 => x"70af800c",
   923 => x"70aefc0c",
   924 => x"aef40b8c",
   925 => x"120c8c11",
   926 => x"0888120c",
   927 => x"74810784",
   928 => x"120c7411",
   929 => x"75710c51",
   930 => x"53f9e039",
   931 => x"75178411",
   932 => x"08810784",
   933 => x"120c538c",
   934 => x"17088818",
   935 => x"08718c12",
   936 => x"0c88120c",
   937 => x"587d5180",
   938 => x"d63f8817",
   939 => x"54f5fe39",
   940 => x"7284150c",
   941 => x"f41af806",
   942 => x"70841e08",
   943 => x"81060784",
   944 => x"1e0c701d",
   945 => x"545b850b",
   946 => x"84140c85",
   947 => x"0b88140c",
   948 => x"8f7b27fd",
   949 => x"da38881c",
   950 => x"527d5182",
   951 => x"823faeec",
   952 => x"0b880508",
   953 => x"aeb00859",
   954 => x"55fdc439",
   955 => x"77aeb00c",
   956 => x"73aee00c",
   957 => x"fca63972",
   958 => x"84150cfd",
   959 => x"b2390404",
   960 => x"fd3d0d80",
   961 => x"0bb7a40c",
   962 => x"765186b2",
   963 => x"3f800853",
   964 => x"8008ff2e",
   965 => x"88387280",
   966 => x"0c853d0d",
   967 => x"04b7a408",
   968 => x"5473802e",
   969 => x"f1387574",
   970 => x"710c5272",
   971 => x"800c853d",
   972 => x"0d04fb3d",
   973 => x"0d777052",
   974 => x"56c43fae",
   975 => x"ec0b8805",
   976 => x"08841108",
   977 => x"fc06707b",
   978 => x"319fef05",
   979 => x"e08006e0",
   980 => x"80055656",
   981 => x"53a08074",
   982 => x"24933880",
   983 => x"527551ff",
   984 => x"9f3faef4",
   985 => x"08155372",
   986 => x"80082e8f",
   987 => x"387551ff",
   988 => x"8e3f8053",
   989 => x"72800c87",
   990 => x"3d0d0473",
   991 => x"30527551",
   992 => x"fefe3f80",
   993 => x"08ff2ea5",
   994 => x"38aeec0b",
   995 => x"88050875",
   996 => x"75318107",
   997 => x"84120c53",
   998 => x"aeb00874",
   999 => x"31aeb00c",
  1000 => x"7551fedb",
  1001 => x"3f810b80",
  1002 => x"0c873d0d",
  1003 => x"04805275",
  1004 => x"51fecd3f",
  1005 => x"aeec0b88",
  1006 => x"05088008",
  1007 => x"71315653",
  1008 => x"8f7525ff",
  1009 => x"a8388008",
  1010 => x"aee00831",
  1011 => x"aeb00c74",
  1012 => x"81078414",
  1013 => x"0c7551fe",
  1014 => x"a63f8053",
  1015 => x"ff9639f6",
  1016 => x"3d0d7c7e",
  1017 => x"545b7280",
  1018 => x"2e828038",
  1019 => x"7a51fe8e",
  1020 => x"3ff81384",
  1021 => x"110870fe",
  1022 => x"06701384",
  1023 => x"1108fc06",
  1024 => x"5d585954",
  1025 => x"58aef408",
  1026 => x"752e82d8",
  1027 => x"38788416",
  1028 => x"0c807381",
  1029 => x"06545a72",
  1030 => x"7a2e81d3",
  1031 => x"38781584",
  1032 => x"11088106",
  1033 => x"5153729f",
  1034 => x"38781757",
  1035 => x"7981e338",
  1036 => x"88150853",
  1037 => x"72aef42e",
  1038 => x"82f1388c",
  1039 => x"1508708c",
  1040 => x"150c7388",
  1041 => x"120c5676",
  1042 => x"81078419",
  1043 => x"0c761877",
  1044 => x"710c5379",
  1045 => x"81903883",
  1046 => x"ff772781",
  1047 => x"c6387689",
  1048 => x"2a77832a",
  1049 => x"56537280",
  1050 => x"2ebf3876",
  1051 => x"862ab805",
  1052 => x"55847327",
  1053 => x"b43880db",
  1054 => x"13559473",
  1055 => x"27ab3876",
  1056 => x"8c2a80ee",
  1057 => x"055580d4",
  1058 => x"73279e38",
  1059 => x"768f2a80",
  1060 => x"f7055582",
  1061 => x"d4732791",
  1062 => x"3876922a",
  1063 => x"80fc0555",
  1064 => x"8ad47327",
  1065 => x"843880fe",
  1066 => x"55741010",
  1067 => x"10aeec05",
  1068 => x"88110855",
  1069 => x"5673762e",
  1070 => x"82a93884",
  1071 => x"1408fc06",
  1072 => x"53767327",
  1073 => x"8d388814",
  1074 => x"08547376",
  1075 => x"2e098106",
  1076 => x"ea388c14",
  1077 => x"08708c1a",
  1078 => x"0c74881a",
  1079 => x"0c788812",
  1080 => x"0c56778c",
  1081 => x"150c7a51",
  1082 => x"fc953f8c",
  1083 => x"3d0d0477",
  1084 => x"08787131",
  1085 => x"59770588",
  1086 => x"19085457",
  1087 => x"72aef42e",
  1088 => x"80dd388c",
  1089 => x"1808708c",
  1090 => x"150c7388",
  1091 => x"120c56fe",
  1092 => x"8c398815",
  1093 => x"088c1608",
  1094 => x"708c130c",
  1095 => x"5788170c",
  1096 => x"fea53976",
  1097 => x"832a7054",
  1098 => x"55807524",
  1099 => x"81923872",
  1100 => x"822c8171",
  1101 => x"2baef008",
  1102 => x"07aeec0b",
  1103 => x"84050c53",
  1104 => x"74101010",
  1105 => x"aeec0588",
  1106 => x"11085556",
  1107 => x"758c190c",
  1108 => x"7388190c",
  1109 => x"7788170c",
  1110 => x"778c150c",
  1111 => x"ff883981",
  1112 => x"5afdba39",
  1113 => x"78177381",
  1114 => x"06545772",
  1115 => x"98387708",
  1116 => x"78713159",
  1117 => x"77058c19",
  1118 => x"08881a08",
  1119 => x"718c120c",
  1120 => x"88120c57",
  1121 => x"57768107",
  1122 => x"84190c77",
  1123 => x"aeec0b88",
  1124 => x"050caee8",
  1125 => x"087726fe",
  1126 => x"cd38aee4",
  1127 => x"08527a51",
  1128 => x"fb903f7a",
  1129 => x"51fad83f",
  1130 => x"fec13981",
  1131 => x"788c150c",
  1132 => x"7888150c",
  1133 => x"738c1a0c",
  1134 => x"73881a0c",
  1135 => x"5afd8839",
  1136 => x"83157082",
  1137 => x"2c81712b",
  1138 => x"aef00807",
  1139 => x"aeec0b84",
  1140 => x"050c5153",
  1141 => x"74101010",
  1142 => x"aeec0588",
  1143 => x"11085556",
  1144 => x"feea3974",
  1145 => x"53807524",
  1146 => x"a5387282",
  1147 => x"2c81712b",
  1148 => x"aef00807",
  1149 => x"aeec0b84",
  1150 => x"050c5375",
  1151 => x"8c190c73",
  1152 => x"88190c77",
  1153 => x"88170c77",
  1154 => x"8c150cfd",
  1155 => x"d9398315",
  1156 => x"70822c81",
  1157 => x"712baef0",
  1158 => x"0807aeec",
  1159 => x"0b84050c",
  1160 => x"5153d839",
  1161 => x"810b800c",
  1162 => x"04803d0d",
  1163 => x"72812e89",
  1164 => x"38800b80",
  1165 => x"0c823d0d",
  1166 => x"04735180",
  1167 => x"eb3ffe3d",
  1168 => x"0db79c08",
  1169 => x"51708838",
  1170 => x"b7a870b7",
  1171 => x"9c0c5170",
  1172 => x"75125252",
  1173 => x"ff537087",
  1174 => x"fb808026",
  1175 => x"873870b7",
  1176 => x"9c0c7153",
  1177 => x"72800c84",
  1178 => x"3d0d04fd",
  1179 => x"3d0d800b",
  1180 => x"a7a40854",
  1181 => x"5472812e",
  1182 => x"983873b7",
  1183 => x"a00ce3df",
  1184 => x"3fe2fd3f",
  1185 => x"b6f45281",
  1186 => x"51e5993f",
  1187 => x"8008519e",
  1188 => x"3f72b7a0",
  1189 => x"0ce3c83f",
  1190 => x"e2e63fb6",
  1191 => x"f4528151",
  1192 => x"e5823f80",
  1193 => x"0851873f",
  1194 => x"00ff3900",
  1195 => x"ff39f73d",
  1196 => x"0d7ba7b0",
  1197 => x"0882c811",
  1198 => x"085a545a",
  1199 => x"77802e80",
  1200 => x"d9388188",
  1201 => x"18841908",
  1202 => x"ff058171",
  1203 => x"2b595559",
  1204 => x"80742480",
  1205 => x"e9388074",
  1206 => x"24b53873",
  1207 => x"822b7811",
  1208 => x"88055656",
  1209 => x"81801908",
  1210 => x"77065372",
  1211 => x"802eb538",
  1212 => x"78167008",
  1213 => x"53537951",
  1214 => x"74085372",
  1215 => x"2dff14fc",
  1216 => x"17fc1779",
  1217 => x"812c5a57",
  1218 => x"57547380",
  1219 => x"25d63877",
  1220 => x"085877ff",
  1221 => x"ad38a7b0",
  1222 => x"0853bc13",
  1223 => x"08a53879",
  1224 => x"51ff853f",
  1225 => x"74085372",
  1226 => x"2dff14fc",
  1227 => x"17fc1779",
  1228 => x"812c5a57",
  1229 => x"57547380",
  1230 => x"25ffa938",
  1231 => x"d2398057",
  1232 => x"ff943972",
  1233 => x"51bc1308",
  1234 => x"53722d79",
  1235 => x"51fed93f",
  1236 => x"ff3d0db6",
  1237 => x"fc0bfc05",
  1238 => x"70085252",
  1239 => x"70ff2e91",
  1240 => x"38702dfc",
  1241 => x"12700852",
  1242 => x"5270ff2e",
  1243 => x"098106f1",
  1244 => x"38833d0d",
  1245 => x"0404e2cc",
  1246 => x"3f040000",
  1247 => x"00000040",
  1248 => x"43000000",
  1249 => x"64756d6d",
  1250 => x"792e6578",
  1251 => x"65000000",
  1252 => x"00ffffff",
  1253 => x"ff00ffff",
  1254 => x"ffff00ff",
  1255 => x"ffffff00",
  1256 => x"00000000",
  1257 => x"00000000",
  1258 => x"00000000",
  1259 => x"00001b84",
  1260 => x"000013b4",
  1261 => x"00000000",
  1262 => x"0000161c",
  1263 => x"00001678",
  1264 => x"000016d4",
  1265 => x"00000000",
  1266 => x"00000000",
  1267 => x"00000000",
  1268 => x"00000000",
  1269 => x"00000000",
  1270 => x"00000000",
  1271 => x"00000000",
  1272 => x"00000000",
  1273 => x"00000000",
  1274 => x"00001380",
  1275 => x"00000000",
  1276 => x"00000000",
  1277 => x"00000000",
  1278 => x"00000000",
  1279 => x"00000000",
  1280 => x"00000000",
  1281 => x"00000000",
  1282 => x"00000000",
  1283 => x"00000000",
  1284 => x"00000000",
  1285 => x"00000000",
  1286 => x"00000000",
  1287 => x"00000000",
  1288 => x"00000000",
  1289 => x"00000000",
  1290 => x"00000000",
  1291 => x"00000000",
  1292 => x"00000000",
  1293 => x"00000000",
  1294 => x"00000000",
  1295 => x"00000000",
  1296 => x"00000000",
  1297 => x"00000000",
  1298 => x"00000000",
  1299 => x"00000000",
  1300 => x"00000000",
  1301 => x"00000000",
  1302 => x"00000000",
  1303 => x"00000001",
  1304 => x"330eabcd",
  1305 => x"1234e66d",
  1306 => x"deec0005",
  1307 => x"000b0000",
  1308 => x"00000000",
  1309 => x"00000000",
  1310 => x"00000000",
  1311 => x"00000000",
  1312 => x"00000000",
  1313 => x"00000000",
  1314 => x"00000000",
  1315 => x"00000000",
  1316 => x"00000000",
  1317 => x"00000000",
  1318 => x"00000000",
  1319 => x"00000000",
  1320 => x"00000000",
  1321 => x"00000000",
  1322 => x"00000000",
  1323 => x"00000000",
  1324 => x"00000000",
  1325 => x"00000000",
  1326 => x"00000000",
  1327 => x"00000000",
  1328 => x"00000000",
  1329 => x"00000000",
  1330 => x"00000000",
  1331 => x"00000000",
  1332 => x"00000000",
  1333 => x"00000000",
  1334 => x"00000000",
  1335 => x"00000000",
  1336 => x"00000000",
  1337 => x"00000000",
  1338 => x"00000000",
  1339 => x"00000000",
  1340 => x"00000000",
  1341 => x"00000000",
  1342 => x"00000000",
  1343 => x"00000000",
  1344 => x"00000000",
  1345 => x"00000000",
  1346 => x"00000000",
  1347 => x"00000000",
  1348 => x"00000000",
  1349 => x"00000000",
  1350 => x"00000000",
  1351 => x"00000000",
  1352 => x"00000000",
  1353 => x"00000000",
  1354 => x"00000000",
  1355 => x"00000000",
  1356 => x"00000000",
  1357 => x"00000000",
  1358 => x"00000000",
  1359 => x"00000000",
  1360 => x"00000000",
  1361 => x"00000000",
  1362 => x"00000000",
  1363 => x"00000000",
  1364 => x"00000000",
  1365 => x"00000000",
  1366 => x"00000000",
  1367 => x"00000000",
  1368 => x"00000000",
  1369 => x"00000000",
  1370 => x"00000000",
  1371 => x"00000000",
  1372 => x"00000000",
  1373 => x"00000000",
  1374 => x"00000000",
  1375 => x"00000000",
  1376 => x"00000000",
  1377 => x"00000000",
  1378 => x"00000000",
  1379 => x"00000000",
  1380 => x"00000000",
  1381 => x"00000000",
  1382 => x"00000000",
  1383 => x"00000000",
  1384 => x"00000000",
  1385 => x"00000000",
  1386 => x"00000000",
  1387 => x"00000000",
  1388 => x"00000000",
  1389 => x"00000000",
  1390 => x"00000000",
  1391 => x"00000000",
  1392 => x"00000000",
  1393 => x"00000000",
  1394 => x"00000000",
  1395 => x"00000000",
  1396 => x"00000000",
  1397 => x"00000000",
  1398 => x"00000000",
  1399 => x"00000000",
  1400 => x"00000000",
  1401 => x"00000000",
  1402 => x"00000000",
  1403 => x"00000000",
  1404 => x"00000000",
  1405 => x"00000000",
  1406 => x"00000000",
  1407 => x"00000000",
  1408 => x"00000000",
  1409 => x"00000000",
  1410 => x"00000000",
  1411 => x"00000000",
  1412 => x"00000000",
  1413 => x"00000000",
  1414 => x"00000000",
  1415 => x"00000000",
  1416 => x"00000000",
  1417 => x"00000000",
  1418 => x"00000000",
  1419 => x"00000000",
  1420 => x"00000000",
  1421 => x"00000000",
  1422 => x"00000000",
  1423 => x"00000000",
  1424 => x"00000000",
  1425 => x"00000000",
  1426 => x"00000000",
  1427 => x"00000000",
  1428 => x"00000000",
  1429 => x"00000000",
  1430 => x"00000000",
  1431 => x"00000000",
  1432 => x"00000000",
  1433 => x"00000000",
  1434 => x"00000000",
  1435 => x"00000000",
  1436 => x"00000000",
  1437 => x"00000000",
  1438 => x"00000000",
  1439 => x"00000000",
  1440 => x"00000000",
  1441 => x"00000000",
  1442 => x"00000000",
  1443 => x"00000000",
  1444 => x"00000000",
  1445 => x"00000000",
  1446 => x"00000000",
  1447 => x"00000000",
  1448 => x"00000000",
  1449 => x"00000000",
  1450 => x"00000000",
  1451 => x"00000000",
  1452 => x"00000000",
  1453 => x"00000000",
  1454 => x"00000000",
  1455 => x"00000000",
  1456 => x"00000000",
  1457 => x"00000000",
  1458 => x"00000000",
  1459 => x"00000000",
  1460 => x"00000000",
  1461 => x"00000000",
  1462 => x"00000000",
  1463 => x"00000000",
  1464 => x"00000000",
  1465 => x"00000000",
  1466 => x"00000000",
  1467 => x"00000000",
  1468 => x"00000000",
  1469 => x"00000000",
  1470 => x"00000000",
  1471 => x"00000000",
  1472 => x"00000000",
  1473 => x"00000000",
  1474 => x"00000000",
  1475 => x"00000000",
  1476 => x"00000000",
  1477 => x"00000000",
  1478 => x"00000000",
  1479 => x"00000000",
  1480 => x"00000000",
  1481 => x"00000000",
  1482 => x"00000000",
  1483 => x"00000000",
  1484 => x"00000000",
  1485 => x"00000000",
  1486 => x"00000000",
  1487 => x"00000000",
  1488 => x"00000000",
  1489 => x"00000000",
  1490 => x"00000000",
  1491 => x"00000000",
  1492 => x"00000000",
  1493 => x"00000000",
  1494 => x"00000000",
  1495 => x"00000000",
  1496 => x"ffffffff",
  1497 => x"00000000",
  1498 => x"00020000",
  1499 => x"00000000",
  1500 => x"00000000",
  1501 => x"0000176c",
  1502 => x"0000176c",
  1503 => x"00001774",
  1504 => x"00001774",
  1505 => x"0000177c",
  1506 => x"0000177c",
  1507 => x"00001784",
  1508 => x"00001784",
  1509 => x"0000178c",
  1510 => x"0000178c",
  1511 => x"00001794",
  1512 => x"00001794",
  1513 => x"0000179c",
  1514 => x"0000179c",
  1515 => x"000017a4",
  1516 => x"000017a4",
  1517 => x"000017ac",
  1518 => x"000017ac",
  1519 => x"000017b4",
  1520 => x"000017b4",
  1521 => x"000017bc",
  1522 => x"000017bc",
  1523 => x"000017c4",
  1524 => x"000017c4",
  1525 => x"000017cc",
  1526 => x"000017cc",
  1527 => x"000017d4",
  1528 => x"000017d4",
  1529 => x"000017dc",
  1530 => x"000017dc",
  1531 => x"000017e4",
  1532 => x"000017e4",
  1533 => x"000017ec",
  1534 => x"000017ec",
  1535 => x"000017f4",
  1536 => x"000017f4",
  1537 => x"000017fc",
  1538 => x"000017fc",
  1539 => x"00001804",
  1540 => x"00001804",
  1541 => x"0000180c",
  1542 => x"0000180c",
  1543 => x"00001814",
  1544 => x"00001814",
  1545 => x"0000181c",
  1546 => x"0000181c",
  1547 => x"00001824",
  1548 => x"00001824",
  1549 => x"0000182c",
  1550 => x"0000182c",
  1551 => x"00001834",
  1552 => x"00001834",
  1553 => x"0000183c",
  1554 => x"0000183c",
  1555 => x"00001844",
  1556 => x"00001844",
  1557 => x"0000184c",
  1558 => x"0000184c",
  1559 => x"00001854",
  1560 => x"00001854",
  1561 => x"0000185c",
  1562 => x"0000185c",
  1563 => x"00001864",
  1564 => x"00001864",
  1565 => x"0000186c",
  1566 => x"0000186c",
  1567 => x"00001874",
  1568 => x"00001874",
  1569 => x"0000187c",
  1570 => x"0000187c",
  1571 => x"00001884",
  1572 => x"00001884",
  1573 => x"0000188c",
  1574 => x"0000188c",
  1575 => x"00001894",
  1576 => x"00001894",
  1577 => x"0000189c",
  1578 => x"0000189c",
  1579 => x"000018a4",
  1580 => x"000018a4",
  1581 => x"000018ac",
  1582 => x"000018ac",
  1583 => x"000018b4",
  1584 => x"000018b4",
  1585 => x"000018bc",
  1586 => x"000018bc",
  1587 => x"000018c4",
  1588 => x"000018c4",
  1589 => x"000018cc",
  1590 => x"000018cc",
  1591 => x"000018d4",
  1592 => x"000018d4",
  1593 => x"000018dc",
  1594 => x"000018dc",
  1595 => x"000018e4",
  1596 => x"000018e4",
  1597 => x"000018ec",
  1598 => x"000018ec",
  1599 => x"000018f4",
  1600 => x"000018f4",
  1601 => x"000018fc",
  1602 => x"000018fc",
  1603 => x"00001904",
  1604 => x"00001904",
  1605 => x"0000190c",
  1606 => x"0000190c",
  1607 => x"00001914",
  1608 => x"00001914",
  1609 => x"0000191c",
  1610 => x"0000191c",
  1611 => x"00001924",
  1612 => x"00001924",
  1613 => x"0000192c",
  1614 => x"0000192c",
  1615 => x"00001934",
  1616 => x"00001934",
  1617 => x"0000193c",
  1618 => x"0000193c",
  1619 => x"00001944",
  1620 => x"00001944",
  1621 => x"0000194c",
  1622 => x"0000194c",
  1623 => x"00001954",
  1624 => x"00001954",
  1625 => x"0000195c",
  1626 => x"0000195c",
  1627 => x"00001964",
  1628 => x"00001964",
  1629 => x"0000196c",
  1630 => x"0000196c",
  1631 => x"00001974",
  1632 => x"00001974",
  1633 => x"0000197c",
  1634 => x"0000197c",
  1635 => x"00001984",
  1636 => x"00001984",
  1637 => x"0000198c",
  1638 => x"0000198c",
  1639 => x"00001994",
  1640 => x"00001994",
  1641 => x"0000199c",
  1642 => x"0000199c",
  1643 => x"000019a4",
  1644 => x"000019a4",
  1645 => x"000019ac",
  1646 => x"000019ac",
  1647 => x"000019b4",
  1648 => x"000019b4",
  1649 => x"000019bc",
  1650 => x"000019bc",
  1651 => x"000019c4",
  1652 => x"000019c4",
  1653 => x"000019cc",
  1654 => x"000019cc",
  1655 => x"000019d4",
  1656 => x"000019d4",
  1657 => x"000019dc",
  1658 => x"000019dc",
  1659 => x"000019e4",
  1660 => x"000019e4",
  1661 => x"000019ec",
  1662 => x"000019ec",
  1663 => x"000019f4",
  1664 => x"000019f4",
  1665 => x"000019fc",
  1666 => x"000019fc",
  1667 => x"00001a04",
  1668 => x"00001a04",
  1669 => x"00001a0c",
  1670 => x"00001a0c",
  1671 => x"00001a14",
  1672 => x"00001a14",
  1673 => x"00001a1c",
  1674 => x"00001a1c",
  1675 => x"00001a24",
  1676 => x"00001a24",
  1677 => x"00001a2c",
  1678 => x"00001a2c",
  1679 => x"00001a34",
  1680 => x"00001a34",
  1681 => x"00001a3c",
  1682 => x"00001a3c",
  1683 => x"00001a44",
  1684 => x"00001a44",
  1685 => x"00001a4c",
  1686 => x"00001a4c",
  1687 => x"00001a54",
  1688 => x"00001a54",
  1689 => x"00001a5c",
  1690 => x"00001a5c",
  1691 => x"00001a64",
  1692 => x"00001a64",
  1693 => x"00001a6c",
  1694 => x"00001a6c",
  1695 => x"00001a74",
  1696 => x"00001a74",
  1697 => x"00001a7c",
  1698 => x"00001a7c",
  1699 => x"00001a84",
  1700 => x"00001a84",
  1701 => x"00001a8c",
  1702 => x"00001a8c",
  1703 => x"00001a94",
  1704 => x"00001a94",
  1705 => x"00001a9c",
  1706 => x"00001a9c",
  1707 => x"00001aa4",
  1708 => x"00001aa4",
  1709 => x"00001aac",
  1710 => x"00001aac",
  1711 => x"00001ab4",
  1712 => x"00001ab4",
  1713 => x"00001abc",
  1714 => x"00001abc",
  1715 => x"00001ac4",
  1716 => x"00001ac4",
  1717 => x"00001acc",
  1718 => x"00001acc",
  1719 => x"00001ad4",
  1720 => x"00001ad4",
  1721 => x"00001adc",
  1722 => x"00001adc",
  1723 => x"00001ae4",
  1724 => x"00001ae4",
  1725 => x"00001aec",
  1726 => x"00001aec",
  1727 => x"00001af4",
  1728 => x"00001af4",
  1729 => x"00001afc",
  1730 => x"00001afc",
  1731 => x"00001b04",
  1732 => x"00001b04",
  1733 => x"00001b0c",
  1734 => x"00001b0c",
  1735 => x"00001b14",
  1736 => x"00001b14",
  1737 => x"00001b1c",
  1738 => x"00001b1c",
  1739 => x"00001b24",
  1740 => x"00001b24",
  1741 => x"00001b2c",
  1742 => x"00001b2c",
  1743 => x"00001b34",
  1744 => x"00001b34",
  1745 => x"00001b3c",
  1746 => x"00001b3c",
  1747 => x"00001b44",
  1748 => x"00001b44",
  1749 => x"00001b4c",
  1750 => x"00001b4c",
  1751 => x"00001b54",
  1752 => x"00001b54",
  1753 => x"00001b5c",
  1754 => x"00001b5c",
  1755 => x"00001b64",
  1756 => x"00001b64",
  1757 => x"00001384",
  1758 => x"ffffffff",
  1759 => x"00000000",
  1760 => x"ffffffff",
  1761 => x"00000000",
  1762 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
