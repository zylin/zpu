
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 15;
constant bytes : integer := 24820;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B80E1";
    when 16#00001# => romdata <= X"D7040000";
    when 16#00002# => romdata <= X"00000000";
    when 16#00003# => romdata <= X"00000000";
    when 16#00004# => romdata <= X"00000000";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"0B0B80E4";
    when 16#00009# => romdata <= X"BE040000";
    when 16#0000A# => romdata <= X"00000000";
    when 16#0000B# => romdata <= X"00000000";
    when 16#0000C# => romdata <= X"00000000";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B80E3";
    when 16#00049# => romdata <= X"F0040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B80E3D3";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B81B1";
    when 16#000A2# => romdata <= X"F8738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B80";
    when 16#000A5# => romdata <= X"E3D60400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"0B0B80E4";
    when 16#000A9# => romdata <= X"A5040000";
    when 16#000AA# => romdata <= X"00000000";
    when 16#000AB# => romdata <= X"00000000";
    when 16#000AC# => romdata <= X"00000000";
    when 16#000AD# => romdata <= X"00000000";
    when 16#000AE# => romdata <= X"00000000";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"0B0B80E4";
    when 16#000B1# => romdata <= X"8C040000";
    when 16#000B2# => romdata <= X"00000000";
    when 16#000B3# => romdata <= X"00000000";
    when 16#000B4# => romdata <= X"00000000";
    when 16#000B5# => romdata <= X"00000000";
    when 16#000B6# => romdata <= X"00000000";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"81B2880C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"FF3D0D02";
    when 16#00101# => romdata <= X"8F053370";
    when 16#00102# => romdata <= X"525280E1";
    when 16#00103# => romdata <= X"BB3F7151";
    when 16#00104# => romdata <= X"80E2A93F";
    when 16#00105# => romdata <= X"71B00C83";
    when 16#00106# => romdata <= X"3D0D04FD";
    when 16#00107# => romdata <= X"3D0D8A51";
    when 16#00108# => romdata <= X"80DCC13F";
    when 16#00109# => romdata <= X"AAAD3F97";
    when 16#0010A# => romdata <= X"8A538193";
    when 16#0010B# => romdata <= X"E4528193";
    when 16#0010C# => romdata <= X"F851AAB2";
    when 16#0010D# => romdata <= X"3FA49253";
    when 16#0010E# => romdata <= X"8193FC52";
    when 16#0010F# => romdata <= X"8194A051";
    when 16#00110# => romdata <= X"AAA43FA7";
    when 16#00111# => romdata <= X"AB538194";
    when 16#00112# => romdata <= X"A8528194";
    when 16#00113# => romdata <= X"B851AA96";
    when 16#00114# => romdata <= X"3FA09D53";
    when 16#00115# => romdata <= X"8194C052";
    when 16#00116# => romdata <= X"8195B851";
    when 16#00117# => romdata <= X"AA883FA2";
    when 16#00118# => romdata <= X"87538194";
    when 16#00119# => romdata <= X"DC528194";
    when 16#0011A# => romdata <= X"FC51A9FA";
    when 16#0011B# => romdata <= X"3FA2ED53";
    when 16#0011C# => romdata <= X"81958452";
    when 16#0011D# => romdata <= X"8195A451";
    when 16#0011E# => romdata <= X"A9EC3F9F";
    when 16#0011F# => romdata <= X"E9538195";
    when 16#00120# => romdata <= X"AC528195";
    when 16#00121# => romdata <= X"C051A9DE";
    when 16#00122# => romdata <= X"3FA5B153";
    when 16#00123# => romdata <= X"8195C852";
    when 16#00124# => romdata <= X"8195E451";
    when 16#00125# => romdata <= X"A9D03FA7";
    when 16#00126# => romdata <= X"C2538195";
    when 16#00127# => romdata <= X"EC528196";
    when 16#00128# => romdata <= X"9051A9C2";
    when 16#00129# => romdata <= X"3FA88353";
    when 16#0012A# => romdata <= X"81969852";
    when 16#0012B# => romdata <= X"8196C051";
    when 16#0012C# => romdata <= X"A9B43FA9";
    when 16#0012D# => romdata <= X"AB538196";
    when 16#0012E# => romdata <= X"C8528196";
    when 16#0012F# => romdata <= X"E851A9A6";
    when 16#00130# => romdata <= X"3FA79253";
    when 16#00131# => romdata <= X"8196EC52";
    when 16#00132# => romdata <= X"81978851";
    when 16#00133# => romdata <= X"A9983FAA";
    when 16#00134# => romdata <= X"86538197";
    when 16#00135# => romdata <= X"90528197";
    when 16#00136# => romdata <= X"A051A98A";
    when 16#00137# => romdata <= X"3FACD253";
    when 16#00138# => romdata <= X"8197A452";
    when 16#00139# => romdata <= X"8197C051";
    when 16#0013A# => romdata <= X"A8FC3FA6";
    when 16#0013B# => romdata <= X"D8538197";
    when 16#0013C# => romdata <= X"C8528197";
    when 16#0013D# => romdata <= X"E051A8EE";
    when 16#0013E# => romdata <= X"3FACDA53";
    when 16#0013F# => romdata <= X"8197E852";
    when 16#00140# => romdata <= X"8197FC51";
    when 16#00141# => romdata <= X"A8E03F8D";
    when 16#00142# => romdata <= X"F9538198";
    when 16#00143# => romdata <= X"84528198";
    when 16#00144# => romdata <= X"9851A8D2";
    when 16#00145# => romdata <= X"3F918353";
    when 16#00146# => romdata <= X"81989C52";
    when 16#00147# => romdata <= X"8198C451";
    when 16#00148# => romdata <= X"A8C43FA6";
    when 16#00149# => romdata <= X"F4538198";
    when 16#0014A# => romdata <= X"CC528198";
    when 16#0014B# => romdata <= X"EC51A8B6";
    when 16#0014C# => romdata <= X"3F96A753";
    when 16#0014D# => romdata <= X"8198F452";
    when 16#0014E# => romdata <= X"81998851";
    when 16#0014F# => romdata <= X"A8A83F8B";
    when 16#00150# => romdata <= X"FD538199";
    when 16#00151# => romdata <= X"90528199";
    when 16#00152# => romdata <= X"9C51A89A";
    when 16#00153# => romdata <= X"3F8DA253";
    when 16#00154# => romdata <= X"8199A052";
    when 16#00155# => romdata <= X"8199C851";
    when 16#00156# => romdata <= X"A88C3F8B";
    when 16#00157# => romdata <= X"FD538199";
    when 16#00158# => romdata <= X"D05281A0";
    when 16#00159# => romdata <= X"F451A7FE";
    when 16#0015A# => romdata <= X"3F8DE853";
    when 16#0015B# => romdata <= X"8199E052";
    when 16#0015C# => romdata <= X"8199F051";
    when 16#0015D# => romdata <= X"A7F03F8B";
    when 16#0015E# => romdata <= X"F253819A";
    when 16#0015F# => romdata <= X"84528193";
    when 16#00160# => romdata <= X"D451A7E2";
    when 16#00161# => romdata <= X"3FB9BD53";
    when 16#00162# => romdata <= X"819A8452";
    when 16#00163# => romdata <= X"8193DC51";
    when 16#00164# => romdata <= X"A7D43FAE";
    when 16#00165# => romdata <= X"A83FA89A";
    when 16#00166# => romdata <= X"3F810B81";
    when 16#00167# => romdata <= X"D5983481";
    when 16#00168# => romdata <= X"C1F83370";
    when 16#00169# => romdata <= X"81FF0651";
    when 16#0016A# => romdata <= X"5473B238";
    when 16#0016B# => romdata <= X"80DDC13F";
    when 16#0016C# => romdata <= X"B0089038";
    when 16#0016D# => romdata <= X"A88A3F81";
    when 16#0016E# => romdata <= X"D5983354";
    when 16#0016F# => romdata <= X"73E13885";
    when 16#00170# => romdata <= X"3D0D0480";
    when 16#00171# => romdata <= X"DDBD3FB0";
    when 16#00172# => romdata <= X"0881FF06";
    when 16#00173# => romdata <= X"51A8DF3F";
    when 16#00174# => romdata <= X"A7EE3F81";
    when 16#00175# => romdata <= X"D5983354";
    when 16#00176# => romdata <= X"73C538E3";
    when 16#00177# => romdata <= X"39800B81";
    when 16#00178# => romdata <= X"C1F834AE";
    when 16#00179# => romdata <= X"F83F80DD";
    when 16#0017A# => romdata <= X"873FB008";
    when 16#0017B# => romdata <= X"802EC538";
    when 16#0017C# => romdata <= X"D239800B";
    when 16#0017D# => romdata <= X"81D59834";
    when 16#0017E# => romdata <= X"800BB00C";
    when 16#0017F# => romdata <= X"04FB3D0D";
    when 16#00180# => romdata <= X"8151AC86";
    when 16#00181# => romdata <= X"3FB00853";
    when 16#00182# => romdata <= X"8251ABFE";
    when 16#00183# => romdata <= X"3FB00856";
    when 16#00184# => romdata <= X"B0088338";
    when 16#00185# => romdata <= X"905672FC";
    when 16#00186# => romdata <= X"06547581";
    when 16#00187# => romdata <= X"2E80FB38";
    when 16#00188# => romdata <= X"80557476";
    when 16#00189# => romdata <= X"27AD3874";
    when 16#0018A# => romdata <= X"83065372";
    when 16#0018B# => romdata <= X"802EB238";
    when 16#0018C# => romdata <= X"81A5F051";
    when 16#0018D# => romdata <= X"80D8C73F";
    when 16#0018E# => romdata <= X"73708405";
    when 16#0018F# => romdata <= X"550852A0";
    when 16#00190# => romdata <= X"5180D8DD";
    when 16#00191# => romdata <= X"3FA05180";
    when 16#00192# => romdata <= X"D89A3F81";
    when 16#00193# => romdata <= X"15557575";
    when 16#00194# => romdata <= X"26D5388A";
    when 16#00195# => romdata <= X"5180D88C";
    when 16#00196# => romdata <= X"3F800BB0";
    when 16#00197# => romdata <= X"0C873D0D";
    when 16#00198# => romdata <= X"048199F8";
    when 16#00199# => romdata <= X"5180D896";
    when 16#0019A# => romdata <= X"3F7352A0";
    when 16#0019B# => romdata <= X"5180D8B1";
    when 16#0019C# => romdata <= X"3F81A0E0";
    when 16#0019D# => romdata <= X"5180D886";
    when 16#0019E# => romdata <= X"3F81A5F0";
    when 16#0019F# => romdata <= X"5180D7FE";
    when 16#001A0# => romdata <= X"3F737084";
    when 16#001A1# => romdata <= X"05550852";
    when 16#001A2# => romdata <= X"A05180D8";
    when 16#001A3# => romdata <= X"943FA051";
    when 16#001A4# => romdata <= X"80D7D13F";
    when 16#001A5# => romdata <= X"811555FF";
    when 16#001A6# => romdata <= X"B5397308";
    when 16#001A7# => romdata <= X"B00C873D";
    when 16#001A8# => romdata <= X"0D04FC3D";
    when 16#001A9# => romdata <= X"0D8151AA";
    when 16#001AA# => romdata <= X"E13FB008";
    when 16#001AB# => romdata <= X"528251A9";
    when 16#001AC# => romdata <= X"A73FB008";
    when 16#001AD# => romdata <= X"81FF0672";
    when 16#001AE# => romdata <= X"56538354";
    when 16#001AF# => romdata <= X"72802EA1";
    when 16#001B0# => romdata <= X"387351AA";
    when 16#001B1# => romdata <= X"C53F8114";
    when 16#001B2# => romdata <= X"7081FF06";
    when 16#001B3# => romdata <= X"FF157081";
    when 16#001B4# => romdata <= X"FF06B008";
    when 16#001B5# => romdata <= X"79708405";
    when 16#001B6# => romdata <= X"5B0C5652";
    when 16#001B7# => romdata <= X"555272E1";
    when 16#001B8# => romdata <= X"3872B00C";
    when 16#001B9# => romdata <= X"863D0D04";
    when 16#001BA# => romdata <= X"803D0D8C";
    when 16#001BB# => romdata <= X"5180D6F4";
    when 16#001BC# => romdata <= X"3F800BB0";
    when 16#001BD# => romdata <= X"0C823D0D";
    when 16#001BE# => romdata <= X"04FB3D0D";
    when 16#001BF# => romdata <= X"800B8199";
    when 16#001C0# => romdata <= X"FC525680";
    when 16#001C1# => romdata <= X"D6F83F75";
    when 16#001C2# => romdata <= X"55741081";
    when 16#001C3# => romdata <= X"FE065381";
    when 16#001C4# => romdata <= X"D05281B2";
    when 16#001C5# => romdata <= X"900851BD";
    when 16#001C6# => romdata <= X"983FB008";
    when 16#001C7# => romdata <= X"982B5480";
    when 16#001C8# => romdata <= X"7424A238";
    when 16#001C9# => romdata <= X"819A8851";
    when 16#001CA# => romdata <= X"80D6D33F";
    when 16#001CB# => romdata <= X"74528851";
    when 16#001CC# => romdata <= X"80D6EE3F";
    when 16#001CD# => romdata <= X"819A9451";
    when 16#001CE# => romdata <= X"80D6C33F";
    when 16#001CF# => romdata <= X"81167083";
    when 16#001D0# => romdata <= X"FFFF0657";
    when 16#001D1# => romdata <= X"54811570";
    when 16#001D2# => romdata <= X"81FF0670";
    when 16#001D3# => romdata <= X"982B5256";
    when 16#001D4# => romdata <= X"54738025";
    when 16#001D5# => romdata <= X"FFB33875";
    when 16#001D6# => romdata <= X"B00C873D";
    when 16#001D7# => romdata <= X"0D04F33D";
    when 16#001D8# => romdata <= X"0D7F0284";
    when 16#001D9# => romdata <= X"0580C305";
    when 16#001DA# => romdata <= X"33028805";
    when 16#001DB# => romdata <= X"80C60522";
    when 16#001DC# => romdata <= X"819AA454";
    when 16#001DD# => romdata <= X"5B555880";
    when 16#001DE# => romdata <= X"D6843F78";
    when 16#001DF# => romdata <= X"5180D7C8";
    when 16#001E0# => romdata <= X"3F819AB0";
    when 16#001E1# => romdata <= X"5180D5F6";
    when 16#001E2# => romdata <= X"3F735288";
    when 16#001E3# => romdata <= X"5180D691";
    when 16#001E4# => romdata <= X"3F819ACC";
    when 16#001E5# => romdata <= X"5180D5E6";
    when 16#001E6# => romdata <= X"3F805776";
    when 16#001E7# => romdata <= X"7927819C";
    when 16#001E8# => romdata <= X"3873108E";
    when 16#001E9# => romdata <= X"3D5D5A79";
    when 16#001EA# => romdata <= X"81FF0653";
    when 16#001EB# => romdata <= X"81905277";
    when 16#001EC# => romdata <= X"51BBFE3F";
    when 16#001ED# => romdata <= X"76882A53";
    when 16#001EE# => romdata <= X"90527751";
    when 16#001EF# => romdata <= X"BBF33F76";
    when 16#001F0# => romdata <= X"81FF0653";
    when 16#001F1# => romdata <= X"90527751";
    when 16#001F2# => romdata <= X"BBE73F81";
    when 16#001F3# => romdata <= X"1A7081FF";
    when 16#001F4# => romdata <= X"06545581";
    when 16#001F5# => romdata <= X"90527751";
    when 16#001F6# => romdata <= X"BBD73F80";
    when 16#001F7# => romdata <= X"5380E052";
    when 16#001F8# => romdata <= X"7751BBCD";
    when 16#001F9# => romdata <= X"3FB00898";
    when 16#001FA# => romdata <= X"2B548074";
    when 16#001FB# => romdata <= X"248A3888";
    when 16#001FC# => romdata <= X"18087081";
    when 16#001FD# => romdata <= X"FF065C56";
    when 16#001FE# => romdata <= X"7A81FF06";
    when 16#001FF# => romdata <= X"81A5F052";
    when 16#00200# => romdata <= X"5680D4FA";
    when 16#00201# => romdata <= X"3F755288";
    when 16#00202# => romdata <= X"5180D595";
    when 16#00203# => romdata <= X"3F819DEC";
    when 16#00204# => romdata <= X"5180D4EA";
    when 16#00205# => romdata <= X"3FE01654";
    when 16#00206# => romdata <= X"80DF7427";
    when 16#00207# => romdata <= X"B6387687";
    when 16#00208# => romdata <= X"06701D57";
    when 16#00209# => romdata <= X"55A07634";
    when 16#0020A# => romdata <= X"74872EB9";
    when 16#0020B# => romdata <= X"38811770";
    when 16#0020C# => romdata <= X"83FFFF06";
    when 16#0020D# => romdata <= X"58557877";
    when 16#0020E# => romdata <= X"26FEEC38";
    when 16#0020F# => romdata <= X"80E00B8C";
    when 16#00210# => romdata <= X"190C8C18";
    when 16#00211# => romdata <= X"0870812A";
    when 16#00212# => romdata <= X"8106585A";
    when 16#00213# => romdata <= X"76F4388F";
    when 16#00214# => romdata <= X"3D0D0476";
    when 16#00215# => romdata <= X"8706701D";
    when 16#00216# => romdata <= X"55557574";
    when 16#00217# => romdata <= X"3474872E";
    when 16#00218# => romdata <= X"098106C9";
    when 16#00219# => romdata <= X"387B5180";
    when 16#0021A# => romdata <= X"D4943F8A";
    when 16#0021B# => romdata <= X"5180D3F4";
    when 16#0021C# => romdata <= X"3F811770";
    when 16#0021D# => romdata <= X"83FFFF06";
    when 16#0021E# => romdata <= X"58557877";
    when 16#0021F# => romdata <= X"26FEA838";
    when 16#00220# => romdata <= X"FFBA39FB";
    when 16#00221# => romdata <= X"3D0D8151";
    when 16#00222# => romdata <= X"A5CE3FB0";
    when 16#00223# => romdata <= X"0881FF06";
    when 16#00224# => romdata <= X"548251A6";
    when 16#00225# => romdata <= X"F53FB008";
    when 16#00226# => romdata <= X"81FF0656";
    when 16#00227# => romdata <= X"8351A5B8";
    when 16#00228# => romdata <= X"3FB00883";
    when 16#00229# => romdata <= X"FFFF0655";
    when 16#0022A# => romdata <= X"739C3881";
    when 16#0022B# => romdata <= X"B2900854";
    when 16#0022C# => romdata <= X"74843881";
    when 16#0022D# => romdata <= X"80557453";
    when 16#0022E# => romdata <= X"75527351";
    when 16#0022F# => romdata <= X"FDA03F74";
    when 16#00230# => romdata <= X"B00C873D";
    when 16#00231# => romdata <= X"0D0481B2";
    when 16#00232# => romdata <= X"940854E4";
    when 16#00233# => romdata <= X"39F83D0D";
    when 16#00234# => romdata <= X"02AA0522";
    when 16#00235# => romdata <= X"81B1EC33";
    when 16#00236# => romdata <= X"81F70658";
    when 16#00237# => romdata <= X"587681B1";
    when 16#00238# => romdata <= X"EC3481B2";
    when 16#00239# => romdata <= X"90085580";
    when 16#0023A# => romdata <= X"C0538190";
    when 16#0023B# => romdata <= X"527451B9";
    when 16#0023C# => romdata <= X"C03F7451";
    when 16#0023D# => romdata <= X"B9ED3FB0";
    when 16#0023E# => romdata <= X"0881FF06";
    when 16#0023F# => romdata <= X"5473802E";
    when 16#00240# => romdata <= X"83FC3876";
    when 16#00241# => romdata <= X"5380D052";
    when 16#00242# => romdata <= X"7451B9A5";
    when 16#00243# => romdata <= X"3F80598F";
    when 16#00244# => romdata <= X"5781B1EC";
    when 16#00245# => romdata <= X"3381FE06";
    when 16#00246# => romdata <= X"547381B1";
    when 16#00247# => romdata <= X"EC3481B2";
    when 16#00248# => romdata <= X"90087457";
    when 16#00249# => romdata <= X"5580C053";
    when 16#0024A# => romdata <= X"81905274";
    when 16#0024B# => romdata <= X"51B9823F";
    when 16#0024C# => romdata <= X"7451B9AF";
    when 16#0024D# => romdata <= X"3FB00881";
    when 16#0024E# => romdata <= X"FF065473";
    when 16#0024F# => romdata <= X"802E83B3";
    when 16#00250# => romdata <= X"38755380";
    when 16#00251# => romdata <= X"D0527451";
    when 16#00252# => romdata <= X"B8E73F77";
    when 16#00253# => romdata <= X"772C8106";
    when 16#00254# => romdata <= X"5574802E";
    when 16#00255# => romdata <= X"83923881";
    when 16#00256# => romdata <= X"B1EC3382";
    when 16#00257# => romdata <= X"07547381";
    when 16#00258# => romdata <= X"B1EC3481";
    when 16#00259# => romdata <= X"B2900874";
    when 16#0025A# => romdata <= X"575580C0";
    when 16#0025B# => romdata <= X"53819052";
    when 16#0025C# => romdata <= X"7451B8BD";
    when 16#0025D# => romdata <= X"3F7451B8";
    when 16#0025E# => romdata <= X"EA3FB008";
    when 16#0025F# => romdata <= X"81FF0654";
    when 16#00260# => romdata <= X"73802E82";
    when 16#00261# => romdata <= X"D8387553";
    when 16#00262# => romdata <= X"80D05274";
    when 16#00263# => romdata <= X"51B8A23F";
    when 16#00264# => romdata <= X"81B29008";
    when 16#00265# => romdata <= X"5580C153";
    when 16#00266# => romdata <= X"81905274";
    when 16#00267# => romdata <= X"51B8923F";
    when 16#00268# => romdata <= X"7451B8BF";
    when 16#00269# => romdata <= X"3FB00881";
    when 16#0026A# => romdata <= X"FF065675";
    when 16#0026B# => romdata <= X"802E8281";
    when 16#0026C# => romdata <= X"38805380";
    when 16#0026D# => romdata <= X"E0527451";
    when 16#0026E# => romdata <= X"B7F73F74";
    when 16#0026F# => romdata <= X"51B8A43F";
    when 16#00270# => romdata <= X"B00881FF";
    when 16#00271# => romdata <= X"06547380";
    when 16#00272# => romdata <= X"2E81E638";
    when 16#00273# => romdata <= X"88150870";
    when 16#00274# => romdata <= X"902B7090";
    when 16#00275# => romdata <= X"2C565656";
    when 16#00276# => romdata <= X"73822A81";
    when 16#00277# => romdata <= X"06547380";
    when 16#00278# => romdata <= X"2E8D3881";
    when 16#00279# => romdata <= X"772B7907";
    when 16#0027A# => romdata <= X"7083FFFF";
    when 16#0027B# => romdata <= X"065A5681";
    when 16#0027C# => romdata <= X"B1EC3381";
    when 16#0027D# => romdata <= X"07547381";
    when 16#0027E# => romdata <= X"B1EC3481";
    when 16#0027F# => romdata <= X"B2900874";
    when 16#00280# => romdata <= X"575580C0";
    when 16#00281# => romdata <= X"53819052";
    when 16#00282# => romdata <= X"7451B7A5";
    when 16#00283# => romdata <= X"3F7451B7";
    when 16#00284# => romdata <= X"D23FB008";
    when 16#00285# => romdata <= X"81FF0654";
    when 16#00286# => romdata <= X"73802E81";
    when 16#00287# => romdata <= X"A1387553";
    when 16#00288# => romdata <= X"80D05274";
    when 16#00289# => romdata <= X"51B78A3F";
    when 16#0028A# => romdata <= X"7681800A";
    when 16#0028B# => romdata <= X"2981FF0A";
    when 16#0028C# => romdata <= X"0570982C";
    when 16#0028D# => romdata <= X"58567680";
    when 16#0028E# => romdata <= X"25FDD638";
    when 16#0028F# => romdata <= X"81B1EC33";
    when 16#00290# => romdata <= X"82075776";
    when 16#00291# => romdata <= X"81B1EC34";
    when 16#00292# => romdata <= X"81B29008";
    when 16#00293# => romdata <= X"5580C053";
    when 16#00294# => romdata <= X"81905274";
    when 16#00295# => romdata <= X"51B6DA3F";
    when 16#00296# => romdata <= X"7451B787";
    when 16#00297# => romdata <= X"3FB00881";
    when 16#00298# => romdata <= X"FF065877";
    when 16#00299# => romdata <= X"802E81B4";
    when 16#0029A# => romdata <= X"38765380";
    when 16#0029B# => romdata <= X"D0527451";
    when 16#0029C# => romdata <= X"B6BF3F81";
    when 16#0029D# => romdata <= X"B1EC3388";
    when 16#0029E# => romdata <= X"07577681";
    when 16#0029F# => romdata <= X"B1EC3481";
    when 16#002A0# => romdata <= X"B2900855";
    when 16#002A1# => romdata <= X"80C05381";
    when 16#002A2# => romdata <= X"90527451";
    when 16#002A3# => romdata <= X"B6A33F74";
    when 16#002A4# => romdata <= X"51B6D03F";
    when 16#002A5# => romdata <= X"B00881FF";
    when 16#002A6# => romdata <= X"06587780";
    when 16#002A7# => romdata <= X"2E80EE38";
    when 16#002A8# => romdata <= X"765380D0";
    when 16#002A9# => romdata <= X"527451B6";
    when 16#002AA# => romdata <= X"883F78B0";
    when 16#002AB# => romdata <= X"0C8A3D0D";
    when 16#002AC# => romdata <= X"04819AD0";
    when 16#002AD# => romdata <= X"5180CFC6";
    when 16#002AE# => romdata <= X"3FFF54FE";
    when 16#002AF# => romdata <= X"9B39819A";
    when 16#002B0# => romdata <= X"D05180CF";
    when 16#002B1# => romdata <= X"B93F7681";
    when 16#002B2# => romdata <= X"800A2981";
    when 16#002B3# => romdata <= X"FF0A0570";
    when 16#002B4# => romdata <= X"982C5856";
    when 16#002B5# => romdata <= X"768025FC";
    when 16#002B6# => romdata <= X"B838FEE0";
    when 16#002B7# => romdata <= X"39819AD0";
    when 16#002B8# => romdata <= X"5180CF9A";
    when 16#002B9# => romdata <= X"3FFDA939";
    when 16#002BA# => romdata <= X"81B1EC33";
    when 16#002BB# => romdata <= X"81FD0654";
    when 16#002BC# => romdata <= X"FCEC3981";
    when 16#002BD# => romdata <= X"9AD05180";
    when 16#002BE# => romdata <= X"CF843FFC";
    when 16#002BF# => romdata <= X"CE39819A";
    when 16#002C0# => romdata <= X"D05180CE";
    when 16#002C1# => romdata <= X"F93F8059";
    when 16#002C2# => romdata <= X"8F57FC85";
    when 16#002C3# => romdata <= X"39819AD0";
    when 16#002C4# => romdata <= X"5180CEEA";
    when 16#002C5# => romdata <= X"3F78B00C";
    when 16#002C6# => romdata <= X"8A3D0D04";
    when 16#002C7# => romdata <= X"819AD051";
    when 16#002C8# => romdata <= X"80CEDB3F";
    when 16#002C9# => romdata <= X"FECD39FF";
    when 16#002CA# => romdata <= X"3D0D8151";
    when 16#002CB# => romdata <= X"A0AA3FB0";
    when 16#002CC# => romdata <= X"0881FF06";
    when 16#002CD# => romdata <= X"52818051";
    when 16#002CE# => romdata <= X"FB933F82";
    when 16#002CF# => romdata <= X"8051FB8D";
    when 16#002D0# => romdata <= X"3F848351";
    when 16#002D1# => romdata <= X"FB873F86";
    when 16#002D2# => romdata <= X"F151FB81";
    when 16#002D3# => romdata <= X"3F71832B";
    when 16#002D4# => romdata <= X"88830751";
    when 16#002D5# => romdata <= X"FAF73F80";
    when 16#002D6# => romdata <= X"0BB00C83";
    when 16#002D7# => romdata <= X"3D0D04FE";
    when 16#002D8# => romdata <= X"3D0D0293";
    when 16#002D9# => romdata <= X"05330284";
    when 16#002DA# => romdata <= X"05970533";
    when 16#002DB# => romdata <= X"54527173";
    when 16#002DC# => romdata <= X"279438A0";
    when 16#002DD# => romdata <= X"5180CDEC";
    when 16#002DE# => romdata <= X"3F811270";
    when 16#002DF# => romdata <= X"81FF0651";
    when 16#002E0# => romdata <= X"52727226";
    when 16#002E1# => romdata <= X"EE38843D";
    when 16#002E2# => romdata <= X"0D04FD3D";
    when 16#002E3# => romdata <= X"0D819B88";
    when 16#002E4# => romdata <= X"5180CDEA";
    when 16#002E5# => romdata <= X"3F819BA8";
    when 16#002E6# => romdata <= X"5180CDE2";
    when 16#002E7# => romdata <= X"3F819BF0";
    when 16#002E8# => romdata <= X"5180CDDA";
    when 16#002E9# => romdata <= X"3F819CB8";
    when 16#002EA# => romdata <= X"5180CDD2";
    when 16#002EB# => romdata <= X"3F81B1E4";
    when 16#002EC# => romdata <= X"08700852";
    when 16#002ED# => romdata <= X"5380CF90";
    when 16#002EE# => romdata <= X"3FB00881";
    when 16#002EF# => romdata <= X"FF065372";
    when 16#002F0# => romdata <= X"8C279438";
    when 16#002F1# => romdata <= X"A05180CD";
    when 16#002F2# => romdata <= X"9B3F8113";
    when 16#002F3# => romdata <= X"7081FF06";
    when 16#002F4# => romdata <= X"54548C73";
    when 16#002F5# => romdata <= X"26EE3881";
    when 16#002F6# => romdata <= X"B1E40884";
    when 16#002F7# => romdata <= X"11085253";
    when 16#002F8# => romdata <= X"80CEE53F";
    when 16#002F9# => romdata <= X"B00881FF";
    when 16#002FA# => romdata <= X"0653728C";
    when 16#002FB# => romdata <= X"279438A0";
    when 16#002FC# => romdata <= X"5180CCF0";
    when 16#002FD# => romdata <= X"3F811370";
    when 16#002FE# => romdata <= X"81FF0654";
    when 16#002FF# => romdata <= X"548C7326";
    when 16#00300# => romdata <= X"EE3881B1";
    when 16#00301# => romdata <= X"E4088811";
    when 16#00302# => romdata <= X"08525380";
    when 16#00303# => romdata <= X"CEBA3FB0";
    when 16#00304# => romdata <= X"0881FF06";
    when 16#00305# => romdata <= X"53728C27";
    when 16#00306# => romdata <= X"9438A051";
    when 16#00307# => romdata <= X"80CCC53F";
    when 16#00308# => romdata <= X"81137081";
    when 16#00309# => romdata <= X"FF065454";
    when 16#0030A# => romdata <= X"8C7326EE";
    when 16#0030B# => romdata <= X"3881B1E4";
    when 16#0030C# => romdata <= X"088C1108";
    when 16#0030D# => romdata <= X"525380CE";
    when 16#0030E# => romdata <= X"8F3FB008";
    when 16#0030F# => romdata <= X"81FF0653";
    when 16#00310# => romdata <= X"728C2794";
    when 16#00311# => romdata <= X"38A05180";
    when 16#00312# => romdata <= X"CC9A3F81";
    when 16#00313# => romdata <= X"137081FF";
    when 16#00314# => romdata <= X"0654548C";
    when 16#00315# => romdata <= X"7326EE38";
    when 16#00316# => romdata <= X"819CD451";
    when 16#00317# => romdata <= X"80CC9F3F";
    when 16#00318# => romdata <= X"81B1E408";
    when 16#00319# => romdata <= X"90110852";
    when 16#0031A# => romdata <= X"5380CDDC";
    when 16#0031B# => romdata <= X"3FB00881";
    when 16#0031C# => romdata <= X"FF065372";
    when 16#0031D# => romdata <= X"8C279438";
    when 16#0031E# => romdata <= X"A05180CB";
    when 16#0031F# => romdata <= X"E73F8113";
    when 16#00320# => romdata <= X"7081FF06";
    when 16#00321# => romdata <= X"54548C73";
    when 16#00322# => romdata <= X"26EE3881";
    when 16#00323# => romdata <= X"B1E40894";
    when 16#00324# => romdata <= X"11085253";
    when 16#00325# => romdata <= X"80CDB13F";
    when 16#00326# => romdata <= X"B00881FF";
    when 16#00327# => romdata <= X"0653728C";
    when 16#00328# => romdata <= X"279438A0";
    when 16#00329# => romdata <= X"5180CBBC";
    when 16#0032A# => romdata <= X"3F811370";
    when 16#0032B# => romdata <= X"81FF0654";
    when 16#0032C# => romdata <= X"548C7326";
    when 16#0032D# => romdata <= X"EE3881B1";
    when 16#0032E# => romdata <= X"E4089811";
    when 16#0032F# => romdata <= X"08525380";
    when 16#00330# => romdata <= X"CD863FB0";
    when 16#00331# => romdata <= X"0881FF06";
    when 16#00332# => romdata <= X"53728C27";
    when 16#00333# => romdata <= X"9438A051";
    when 16#00334# => romdata <= X"80CB913F";
    when 16#00335# => romdata <= X"81137081";
    when 16#00336# => romdata <= X"FF065454";
    when 16#00337# => romdata <= X"8C7326EE";
    when 16#00338# => romdata <= X"3881B1E4";
    when 16#00339# => romdata <= X"089C1108";
    when 16#0033A# => romdata <= X"525380CC";
    when 16#0033B# => romdata <= X"DB3FB008";
    when 16#0033C# => romdata <= X"81FF0653";
    when 16#0033D# => romdata <= X"728C2794";
    when 16#0033E# => romdata <= X"38A05180";
    when 16#0033F# => romdata <= X"CAE63F81";
    when 16#00340# => romdata <= X"137081FF";
    when 16#00341# => romdata <= X"0654548C";
    when 16#00342# => romdata <= X"7326EE38";
    when 16#00343# => romdata <= X"819CF051";
    when 16#00344# => romdata <= X"80CAEB3F";
    when 16#00345# => romdata <= X"81B1E408";
    when 16#00346# => romdata <= X"54810BB0";
    when 16#00347# => romdata <= X"150CB014";
    when 16#00348# => romdata <= X"08537280";
    when 16#00349# => romdata <= X"25F838A0";
    when 16#0034A# => romdata <= X"14085180";
    when 16#0034B# => romdata <= X"CC9A3FB0";
    when 16#0034C# => romdata <= X"0881FF06";
    when 16#0034D# => romdata <= X"53728C27";
    when 16#0034E# => romdata <= X"9438A051";
    when 16#0034F# => romdata <= X"80CAA53F";
    when 16#00350# => romdata <= X"81137081";
    when 16#00351# => romdata <= X"FF065454";
    when 16#00352# => romdata <= X"8C7326EE";
    when 16#00353# => romdata <= X"3881B1E4";
    when 16#00354# => romdata <= X"08A41108";
    when 16#00355# => romdata <= X"525380CB";
    when 16#00356# => romdata <= X"EF3FB008";
    when 16#00357# => romdata <= X"81FF0653";
    when 16#00358# => romdata <= X"728C2794";
    when 16#00359# => romdata <= X"38A05180";
    when 16#0035A# => romdata <= X"C9FA3F81";
    when 16#0035B# => romdata <= X"137081FF";
    when 16#0035C# => romdata <= X"0654548C";
    when 16#0035D# => romdata <= X"7326EE38";
    when 16#0035E# => romdata <= X"81B1E408";
    when 16#0035F# => romdata <= X"A8110852";
    when 16#00360# => romdata <= X"5380CBC4";
    when 16#00361# => romdata <= X"3FB00881";
    when 16#00362# => romdata <= X"FF065372";
    when 16#00363# => romdata <= X"8C279438";
    when 16#00364# => romdata <= X"A05180C9";
    when 16#00365# => romdata <= X"CF3F8113";
    when 16#00366# => romdata <= X"7081FF06";
    when 16#00367# => romdata <= X"54548C73";
    when 16#00368# => romdata <= X"26EE3881";
    when 16#00369# => romdata <= X"B1E408AC";
    when 16#0036A# => romdata <= X"11085253";
    when 16#0036B# => romdata <= X"80CB993F";
    when 16#0036C# => romdata <= X"B00881FF";
    when 16#0036D# => romdata <= X"0653728C";
    when 16#0036E# => romdata <= X"279438A0";
    when 16#0036F# => romdata <= X"5180C9A4";
    when 16#00370# => romdata <= X"3F811370";
    when 16#00371# => romdata <= X"81FF0654";
    when 16#00372# => romdata <= X"548C7326";
    when 16#00373# => romdata <= X"EE38819D";
    when 16#00374# => romdata <= X"8C5180C9";
    when 16#00375# => romdata <= X"A93F81B1";
    when 16#00376# => romdata <= X"E408B011";
    when 16#00377# => romdata <= X"08FE0A06";
    when 16#00378# => romdata <= X"525480CA";
    when 16#00379# => romdata <= X"E33F81B1";
    when 16#0037A# => romdata <= X"E4085480";
    when 16#0037B# => romdata <= X"0BB0150C";
    when 16#0037C# => romdata <= X"819DA051";
    when 16#0037D# => romdata <= X"80C9873F";
    when 16#0037E# => romdata <= X"819DB851";
    when 16#0037F# => romdata <= X"80C8FF3F";
    when 16#00380# => romdata <= X"81B1E408";
    when 16#00381# => romdata <= X"80C01108";
    when 16#00382# => romdata <= X"525380CA";
    when 16#00383# => romdata <= X"BB3FB008";
    when 16#00384# => romdata <= X"81FF0653";
    when 16#00385# => romdata <= X"72982794";
    when 16#00386# => romdata <= X"38A05180";
    when 16#00387# => romdata <= X"C8C63F81";
    when 16#00388# => romdata <= X"137081FF";
    when 16#00389# => romdata <= X"06515398";
    when 16#0038A# => romdata <= X"7326EE38";
    when 16#0038B# => romdata <= X"81B1E408";
    when 16#0038C# => romdata <= X"80C81108";
    when 16#0038D# => romdata <= X"525480CA";
    when 16#0038E# => romdata <= X"8F3FB008";
    when 16#0038F# => romdata <= X"81FF0653";
    when 16#00390# => romdata <= X"72982794";
    when 16#00391# => romdata <= X"38A05180";
    when 16#00392# => romdata <= X"C89A3F81";
    when 16#00393# => romdata <= X"137081FF";
    when 16#00394# => romdata <= X"06515398";
    when 16#00395# => romdata <= X"7326EE38";
    when 16#00396# => romdata <= X"819DD451";
    when 16#00397# => romdata <= X"80C89F3F";
    when 16#00398# => romdata <= X"81B1E408";
    when 16#00399# => romdata <= X"80C41108";
    when 16#0039A# => romdata <= X"525480C9";
    when 16#0039B# => romdata <= X"DB3FB008";
    when 16#0039C# => romdata <= X"81FF0653";
    when 16#0039D# => romdata <= X"72982794";
    when 16#0039E# => romdata <= X"38A05180";
    when 16#0039F# => romdata <= X"C7E63F81";
    when 16#003A0# => romdata <= X"137081FF";
    when 16#003A1# => romdata <= X"06515398";
    when 16#003A2# => romdata <= X"7326EE38";
    when 16#003A3# => romdata <= X"81B1E408";
    when 16#003A4# => romdata <= X"80CC1108";
    when 16#003A5# => romdata <= X"525480C9";
    when 16#003A6# => romdata <= X"AF3FB008";
    when 16#003A7# => romdata <= X"81FF0653";
    when 16#003A8# => romdata <= X"72982794";
    when 16#003A9# => romdata <= X"38A05180";
    when 16#003AA# => romdata <= X"C7BA3F81";
    when 16#003AB# => romdata <= X"137081FF";
    when 16#003AC# => romdata <= X"06515398";
    when 16#003AD# => romdata <= X"7326EE38";
    when 16#003AE# => romdata <= X"8A5180C7";
    when 16#003AF# => romdata <= X"A73F81B1";
    when 16#003B0# => romdata <= X"E408B411";
    when 16#003B1# => romdata <= X"087081FF";
    when 16#003B2# => romdata <= X"06819DF0";
    when 16#003B3# => romdata <= X"54525553";
    when 16#003B4# => romdata <= X"80C7AB3F";
    when 16#003B5# => romdata <= X"725180C8";
    when 16#003B6# => romdata <= X"EF3FA051";
    when 16#003B7# => romdata <= X"80C7853F";
    when 16#003B8# => romdata <= X"72862694";
    when 16#003B9# => romdata <= X"38721010";
    when 16#003BA# => romdata <= X"81A2B005";
    when 16#003BB# => romdata <= X"54730804";
    when 16#003BC# => romdata <= X"819E8451";
    when 16#003BD# => romdata <= X"80C7873F";
    when 16#003BE# => romdata <= X"81B1E408";
    when 16#003BF# => romdata <= X"B8110870";
    when 16#003C0# => romdata <= X"81FF0681";
    when 16#003C1# => romdata <= X"9E905452";
    when 16#003C2# => romdata <= X"545480C6";
    when 16#003C3# => romdata <= X"F13F7352";
    when 16#003C4# => romdata <= X"885180C7";
    when 16#003C5# => romdata <= X"8C3F7381";
    when 16#003C6# => romdata <= X"06537280";
    when 16#003C7# => romdata <= X"F2387381";
    when 16#003C8# => romdata <= X"2A708106";
    when 16#003C9# => romdata <= X"51537280";
    when 16#003CA# => romdata <= X"CE387382";
    when 16#003CB# => romdata <= X"2A708106";
    when 16#003CC# => romdata <= X"515372AE";
    when 16#003CD# => romdata <= X"3873832A";
    when 16#003CE# => romdata <= X"81065473";
    when 16#003CF# => romdata <= X"8F388A51";
    when 16#003D0# => romdata <= X"80C6A13F";
    when 16#003D1# => romdata <= X"800BB00C";
    when 16#003D2# => romdata <= X"853D0D04";
    when 16#003D3# => romdata <= X"819EA451";
    when 16#003D4# => romdata <= X"80C6AB3F";
    when 16#003D5# => romdata <= X"8A5180C6";
    when 16#003D6# => romdata <= X"8B3F800B";
    when 16#003D7# => romdata <= X"B00C853D";
    when 16#003D8# => romdata <= X"0D04819E";
    when 16#003D9# => romdata <= X"B85180C6";
    when 16#003DA# => romdata <= X"953F7383";
    when 16#003DB# => romdata <= X"2A810654";
    when 16#003DC# => romdata <= X"73802ECA";
    when 16#003DD# => romdata <= X"38D63981";
    when 16#003DE# => romdata <= X"9ED85180";
    when 16#003DF# => romdata <= X"C6803F73";
    when 16#003E0# => romdata <= X"822A7081";
    when 16#003E1# => romdata <= X"06515372";
    when 16#003E2# => romdata <= X"802EFFA9";
    when 16#003E3# => romdata <= X"38D43981";
    when 16#003E4# => romdata <= X"9EF05180";
    when 16#003E5# => romdata <= X"C5E83F73";
    when 16#003E6# => romdata <= X"812A7081";
    when 16#003E7# => romdata <= X"06515372";
    when 16#003E8# => romdata <= X"802EFF86";
    when 16#003E9# => romdata <= X"38D13981";
    when 16#003EA# => romdata <= X"9F845180";
    when 16#003EB# => romdata <= X"C5D03FFE";
    when 16#003EC# => romdata <= X"C739819F";
    when 16#003ED# => romdata <= X"905180C5";
    when 16#003EE# => romdata <= X"C53FFEBC";
    when 16#003EF# => romdata <= X"39819F9C";
    when 16#003F0# => romdata <= X"5180C5BA";
    when 16#003F1# => romdata <= X"3FFEB139";
    when 16#003F2# => romdata <= X"819FA051";
    when 16#003F3# => romdata <= X"80C5AF3F";
    when 16#003F4# => romdata <= X"FEA63981";
    when 16#003F5# => romdata <= X"9FAC5180";
    when 16#003F6# => romdata <= X"C5A43FFE";
    when 16#003F7# => romdata <= X"9B39819F";
    when 16#003F8# => romdata <= X"B85180C5";
    when 16#003F9# => romdata <= X"993FFE90";
    when 16#003FA# => romdata <= X"39FE3D0D";
    when 16#003FB# => romdata <= X"880A5384";
    when 16#003FC# => romdata <= X"0A0B81B1";
    when 16#003FD# => romdata <= X"E0088C11";
    when 16#003FE# => romdata <= X"08515252";
    when 16#003FF# => romdata <= X"80712795";
    when 16#00400# => romdata <= X"38807370";
    when 16#00401# => romdata <= X"8405550C";
    when 16#00402# => romdata <= X"80727084";
    when 16#00403# => romdata <= X"05540CFF";
    when 16#00404# => romdata <= X"115170ED";
    when 16#00405# => romdata <= X"38800BB0";
    when 16#00406# => romdata <= X"0C843D0D";
    when 16#00407# => romdata <= X"04FA3D0D";
    when 16#00408# => romdata <= X"880A5784";
    when 16#00409# => romdata <= X"0A568151";
    when 16#0040A# => romdata <= X"96AE3FB0";
    when 16#0040B# => romdata <= X"0883FFFF";
    when 16#0040C# => romdata <= X"06547383";
    when 16#0040D# => romdata <= X"38905480";
    when 16#0040E# => romdata <= X"55747427";
    when 16#0040F# => romdata <= X"81C23875";
    when 16#00410# => romdata <= X"0870902C";
    when 16#00411# => romdata <= X"525380C5";
    when 16#00412# => romdata <= X"FF3FB008";
    when 16#00413# => romdata <= X"81FF0652";
    when 16#00414# => romdata <= X"718A2794";
    when 16#00415# => romdata <= X"38A05180";
    when 16#00416# => romdata <= X"C48A3F81";
    when 16#00417# => romdata <= X"127081FF";
    when 16#00418# => romdata <= X"0651528A";
    when 16#00419# => romdata <= X"7226EE38";
    when 16#0041A# => romdata <= X"72902B70";
    when 16#0041B# => romdata <= X"902C5252";
    when 16#0041C# => romdata <= X"80C5D53F";
    when 16#0041D# => romdata <= X"B00881FF";
    when 16#0041E# => romdata <= X"0652718A";
    when 16#0041F# => romdata <= X"279438A0";
    when 16#00420# => romdata <= X"5180C3E0";
    when 16#00421# => romdata <= X"3F811270";
    when 16#00422# => romdata <= X"81FF0653";
    when 16#00423# => romdata <= X"538A7226";
    when 16#00424# => romdata <= X"EE387608";
    when 16#00425# => romdata <= X"70902C52";
    when 16#00426# => romdata <= X"5380C5AC";
    when 16#00427# => romdata <= X"3FB00881";
    when 16#00428# => romdata <= X"FF065271";
    when 16#00429# => romdata <= X"8A279438";
    when 16#0042A# => romdata <= X"A05180C3";
    when 16#0042B# => romdata <= X"B73F8112";
    when 16#0042C# => romdata <= X"7081FF06";
    when 16#0042D# => romdata <= X"51528A72";
    when 16#0042E# => romdata <= X"26EE3872";
    when 16#0042F# => romdata <= X"902B7090";
    when 16#00430# => romdata <= X"2C525280";
    when 16#00431# => romdata <= X"C5823FB0";
    when 16#00432# => romdata <= X"0881FF06";
    when 16#00433# => romdata <= X"52718A27";
    when 16#00434# => romdata <= X"9438A051";
    when 16#00435# => romdata <= X"80C38D3F";
    when 16#00436# => romdata <= X"81127081";
    when 16#00437# => romdata <= X"FF065353";
    when 16#00438# => romdata <= X"8A7226EE";
    when 16#00439# => romdata <= X"388A5180";
    when 16#0043A# => romdata <= X"C2FA3F84";
    when 16#0043B# => romdata <= X"17841781";
    when 16#0043C# => romdata <= X"177083FF";
    when 16#0043D# => romdata <= X"FF065854";
    when 16#0043E# => romdata <= X"57577375";
    when 16#0043F# => romdata <= X"26FEC038";
    when 16#00440# => romdata <= X"73B00C88";
    when 16#00441# => romdata <= X"3D0D04FD";
    when 16#00442# => romdata <= X"3D0D81B1";
    when 16#00443# => romdata <= X"E0088C11";
    when 16#00444# => romdata <= X"0870822B";
    when 16#00445# => romdata <= X"83FFFC06";
    when 16#00446# => romdata <= X"819FC454";
    when 16#00447# => romdata <= X"51545480";
    when 16#00448# => romdata <= X"C2DC3F72";
    when 16#00449# => romdata <= X"52880A51";
    when 16#0044A# => romdata <= X"9AF63FB0";
    when 16#0044B# => romdata <= X"0854B008";
    when 16#0044C# => romdata <= X"FE2EAB38";
    when 16#0044D# => romdata <= X"B008FF2E";
    when 16#0044E# => romdata <= X"96387251";
    when 16#0044F# => romdata <= X"80C4893F";
    when 16#00450# => romdata <= X"819FD851";
    when 16#00451# => romdata <= X"80C2B73F";
    when 16#00452# => romdata <= X"73B00C85";
    when 16#00453# => romdata <= X"3D0D0481";
    when 16#00454# => romdata <= X"9FEC5180";
    when 16#00455# => romdata <= X"C2A83F73";
    when 16#00456# => romdata <= X"B00C853D";
    when 16#00457# => romdata <= X"0D04819F";
    when 16#00458# => romdata <= X"F45180C2";
    when 16#00459# => romdata <= X"993F73B0";
    when 16#0045A# => romdata <= X"0C853D0D";
    when 16#0045B# => romdata <= X"04FC3D0D";
    when 16#0045C# => romdata <= X"81B1E008";
    when 16#0045D# => romdata <= X"8C110870";
    when 16#0045E# => romdata <= X"822B83FF";
    when 16#0045F# => romdata <= X"FC0681A0";
    when 16#00460# => romdata <= X"80545155";
    when 16#00461# => romdata <= X"5580C1F6";
    when 16#00462# => romdata <= X"3F81B2A4";
    when 16#00463# => romdata <= X"08881108";
    when 16#00464# => romdata <= X"7080C007";
    when 16#00465# => romdata <= X"88130C54";
    when 16#00466# => romdata <= X"55735288";
    when 16#00467# => romdata <= X"0A519D82";
    when 16#00468# => romdata <= X"3FB00881";
    when 16#00469# => romdata <= X"B2A40888";
    when 16#0046A# => romdata <= X"110870FF";
    when 16#0046B# => romdata <= X"BF068813";
    when 16#0046C# => romdata <= X"0C555555";
    when 16#0046D# => romdata <= X"B008FE2E";
    when 16#0046E# => romdata <= X"80C938B0";
    when 16#0046F# => romdata <= X"08FE249C";
    when 16#00470# => romdata <= X"38B008FD";
    when 16#00471# => romdata <= X"2EAE3874";
    when 16#00472# => romdata <= X"5180C2FC";
    when 16#00473# => romdata <= X"3F81A094";
    when 16#00474# => romdata <= X"5180C1AA";
    when 16#00475# => romdata <= X"3F74B00C";
    when 16#00476# => romdata <= X"863D0D04";
    when 16#00477# => romdata <= X"B008FF2E";
    when 16#00478# => romdata <= X"098106E3";
    when 16#00479# => romdata <= X"38819FEC";
    when 16#0047A# => romdata <= X"5180C192";
    when 16#0047B# => romdata <= X"3F74B00C";
    when 16#0047C# => romdata <= X"863D0D04";
    when 16#0047D# => romdata <= X"81A0A851";
    when 16#0047E# => romdata <= X"80C1833F";
    when 16#0047F# => romdata <= X"74B00C86";
    when 16#00480# => romdata <= X"3D0D0481";
    when 16#00481# => romdata <= X"A0B85180";
    when 16#00482# => romdata <= X"C0F43F74";
    when 16#00483# => romdata <= X"B00C863D";
    when 16#00484# => romdata <= X"0D04FD3D";
    when 16#00485# => romdata <= X"0D815192";
    when 16#00486# => romdata <= X"BF3FB008";
    when 16#00487# => romdata <= X"81FF0654";
    when 16#00488# => romdata <= X"73802EA4";
    when 16#00489# => romdata <= X"38738426";
    when 16#0048A# => romdata <= X"903881B1";
    when 16#0048B# => romdata <= X"E0087471";
    when 16#0048C# => romdata <= X"0C5373B0";
    when 16#0048D# => romdata <= X"0C853D0D";
    when 16#0048E# => romdata <= X"0481B1E0";
    when 16#0048F# => romdata <= X"08538073";
    when 16#00490# => romdata <= X"0C73B00C";
    when 16#00491# => romdata <= X"853D0D04";
    when 16#00492# => romdata <= X"81A0C451";
    when 16#00493# => romdata <= X"80C0AF3F";
    when 16#00494# => romdata <= X"81A0D451";
    when 16#00495# => romdata <= X"80C0A73F";
    when 16#00496# => romdata <= X"81B1E008";
    when 16#00497# => romdata <= X"70085253";
    when 16#00498# => romdata <= X"80C1E53F";
    when 16#00499# => romdata <= X"81A0E451";
    when 16#0049A# => romdata <= X"80C0933F";
    when 16#0049B# => romdata <= X"81B1E008";
    when 16#0049C# => romdata <= X"84110853";
    when 16#0049D# => romdata <= X"53A05180";
    when 16#0049E# => romdata <= X"C0A73F81";
    when 16#0049F# => romdata <= X"A0F851BF";
    when 16#004A0# => romdata <= X"FD3F81B1";
    when 16#004A1# => romdata <= X"E0088811";
    when 16#004A2# => romdata <= X"085353A0";
    when 16#004A3# => romdata <= X"5180C091";
    when 16#004A4# => romdata <= X"3F81A18C";
    when 16#004A5# => romdata <= X"51BFE73F";
    when 16#004A6# => romdata <= X"81B1E008";
    when 16#004A7# => romdata <= X"8C110852";
    when 16#004A8# => romdata <= X"5380C1A4";
    when 16#004A9# => romdata <= X"3F8A51BF";
    when 16#004AA# => romdata <= X"BB3F73B0";
    when 16#004AB# => romdata <= X"0C853D0D";
    when 16#004AC# => romdata <= X"04F63D0D";
    when 16#004AD# => romdata <= X"880A5681";
    when 16#004AE# => romdata <= X"51919D3F";
    when 16#004AF# => romdata <= X"B0088B3D";
    when 16#004B0# => romdata <= X"23825191";
    when 16#004B1# => romdata <= X"933FB008";
    when 16#004B2# => romdata <= X"028405A6";
    when 16#004B3# => romdata <= X"05238351";
    when 16#004B4# => romdata <= X"91863FB0";
    when 16#004B5# => romdata <= X"088C3D23";
    when 16#004B6# => romdata <= X"845190FC";
    when 16#004B7# => romdata <= X"3FB00889";
    when 16#004B8# => romdata <= X"3D238551";
    when 16#004B9# => romdata <= X"90F23FB0";
    when 16#004BA# => romdata <= X"08028405";
    when 16#004BB# => romdata <= X"9E052386";
    when 16#004BC# => romdata <= X"5190E53F";
    when 16#004BD# => romdata <= X"B0088A3D";
    when 16#004BE# => romdata <= X"23800B81";
    when 16#004BF# => romdata <= X"B1E0088C";
    when 16#004C0# => romdata <= X"11085153";
    when 16#004C1# => romdata <= X"55747227";
    when 16#004C2# => romdata <= X"B8387154";
    when 16#004C3# => romdata <= X"8C3D7510";
    when 16#004C4# => romdata <= X"05F81122";
    when 16#004C5# => romdata <= X"70902BF0";
    when 16#004C6# => romdata <= X"13227084";
    when 16#004C7# => romdata <= X"80802972";
    when 16#004C8# => romdata <= X"902C057A";
    when 16#004C9# => romdata <= X"0C525558";
    when 16#004CA# => romdata <= X"81167081";
    when 16#004CB# => romdata <= X"FF065254";
    when 16#004CC# => romdata <= X"5274822E";
    when 16#004CD# => romdata <= X"94387184";
    when 16#004CE# => romdata <= X"17FF1656";
    when 16#004CF# => romdata <= X"575573CC";
    when 16#004D0# => romdata <= X"38800BB0";
    when 16#004D1# => romdata <= X"0C8C3D0D";
    when 16#004D2# => romdata <= X"04800B84";
    when 16#004D3# => romdata <= X"17FF1656";
    when 16#004D4# => romdata <= X"575573FF";
    when 16#004D5# => romdata <= X"B738EA39";
    when 16#004D6# => romdata <= X"FE3D0D81";
    when 16#004D7# => romdata <= X"518FF93F";
    when 16#004D8# => romdata <= X"B00881FF";
    when 16#004D9# => romdata <= X"0681B1DC";
    when 16#004DA# => romdata <= X"08718812";
    when 16#004DB# => romdata <= X"0C53B00C";
    when 16#004DC# => romdata <= X"843D0D04";
    when 16#004DD# => romdata <= X"803D0D81";
    when 16#004DE# => romdata <= X"51918F3F";
    when 16#004DF# => romdata <= X"B00883FF";
    when 16#004E0# => romdata <= X"FF0651EA";
    when 16#004E1# => romdata <= X"C83FB008";
    when 16#004E2# => romdata <= X"83FFFF06";
    when 16#004E3# => romdata <= X"B00C823D";
    when 16#004E4# => romdata <= X"0D04803D";
    when 16#004E5# => romdata <= X"0D81518F";
    when 16#004E6# => romdata <= X"BF3FB008";
    when 16#004E7# => romdata <= X"81FF0651";
    when 16#004E8# => romdata <= X"A0B93F80";
    when 16#004E9# => romdata <= X"0BB00C82";
    when 16#004EA# => romdata <= X"3D0D0480";
    when 16#004EB# => romdata <= X"3D0D81B2";
    when 16#004EC# => romdata <= X"A80851F8";
    when 16#004ED# => romdata <= X"BB9586A1";
    when 16#004EE# => romdata <= X"710C810B";
    when 16#004EF# => romdata <= X"B00C823D";
    when 16#004F0# => romdata <= X"0D04FC3D";
    when 16#004F1# => romdata <= X"0D81518F";
    when 16#004F2# => romdata <= X"8F3FB008";
    when 16#004F3# => romdata <= X"81FF0654";
    when 16#004F4# => romdata <= X"82518F84";
    when 16#004F5# => romdata <= X"3FB00881";
    when 16#004F6# => romdata <= X"FF0681B2";
    when 16#004F7# => romdata <= X"9C088411";
    when 16#004F8# => romdata <= X"0870FE8F";
    when 16#004F9# => romdata <= X"0A067798";
    when 16#004FA# => romdata <= X"2B075154";
    when 16#004FB# => romdata <= X"56537280";
    when 16#004FC# => romdata <= X"2E863871";
    when 16#004FD# => romdata <= X"810A0752";
    when 16#004FE# => romdata <= X"7184160C";
    when 16#004FF# => romdata <= X"71B00C86";
    when 16#00500# => romdata <= X"3D0D04FD";
    when 16#00501# => romdata <= X"3D0D81B2";
    when 16#00502# => romdata <= X"9C088411";
    when 16#00503# => romdata <= X"08555381";
    when 16#00504# => romdata <= X"518EC53F";
    when 16#00505# => romdata <= X"B00881FF";
    when 16#00506# => romdata <= X"0674DFFF";
    when 16#00507# => romdata <= X"FF065452";
    when 16#00508# => romdata <= X"71802E87";
    when 16#00509# => romdata <= X"3873A080";
    when 16#0050A# => romdata <= X"80075382";
    when 16#0050B# => romdata <= X"518EA93F";
    when 16#0050C# => romdata <= X"B00881FF";
    when 16#0050D# => romdata <= X"0673EFFF";
    when 16#0050E# => romdata <= X"0A065552";
    when 16#0050F# => romdata <= X"71802E87";
    when 16#00510# => romdata <= X"38729080";
    when 16#00511# => romdata <= X"0A075483";
    when 16#00512# => romdata <= X"518E8D3F";
    when 16#00513# => romdata <= X"B00881FF";
    when 16#00514# => romdata <= X"0674F7FF";
    when 16#00515# => romdata <= X"0A065452";
    when 16#00516# => romdata <= X"71802E87";
    when 16#00517# => romdata <= X"38738880";
    when 16#00518# => romdata <= X"0A075384";
    when 16#00519# => romdata <= X"518DF13F";
    when 16#0051A# => romdata <= X"B00881FF";
    when 16#0051B# => romdata <= X"0673FBFF";
    when 16#0051C# => romdata <= X"0A065552";
    when 16#0051D# => romdata <= X"71802E87";
    when 16#0051E# => romdata <= X"38728480";
    when 16#0051F# => romdata <= X"0A075485";
    when 16#00520# => romdata <= X"518DD53F";
    when 16#00521# => romdata <= X"B00881FF";
    when 16#00522# => romdata <= X"0674FDFF";
    when 16#00523# => romdata <= X"0A065452";
    when 16#00524# => romdata <= X"71802E87";
    when 16#00525# => romdata <= X"38738280";
    when 16#00526# => romdata <= X"0A075381";
    when 16#00527# => romdata <= X"B29C0873";
    when 16#00528# => romdata <= X"84120C54";
    when 16#00529# => romdata <= X"72B00C85";
    when 16#0052A# => romdata <= X"3D0D04FC";
    when 16#0052B# => romdata <= X"3D0D81B2";
    when 16#0052C# => romdata <= X"9C087008";
    when 16#0052D# => romdata <= X"81A19C53";
    when 16#0052E# => romdata <= X"5555BBC2";
    when 16#0052F# => romdata <= X"3F739E2A";
    when 16#00530# => romdata <= X"81065271";
    when 16#00531# => romdata <= X"802EB638";
    when 16#00532# => romdata <= X"81A1AC51";
    when 16#00533# => romdata <= X"BBB03F81";
    when 16#00534# => romdata <= X"518D853F";
    when 16#00535# => romdata <= X"B00881FF";
    when 16#00536# => romdata <= X"0681B29C";
    when 16#00537# => romdata <= X"08841108";
    when 16#00538# => romdata <= X"70FD0A06";
    when 16#00539# => romdata <= X"56565652";
    when 16#0053A# => romdata <= X"71802E86";
    when 16#0053B# => romdata <= X"3873820A";
    when 16#0053C# => romdata <= X"07537284";
    when 16#0053D# => romdata <= X"160C72B0";
    when 16#0053E# => romdata <= X"0C863D0D";
    when 16#0053F# => romdata <= X"0481A1B4";
    when 16#00540# => romdata <= X"51BAFB3F";
    when 16#00541# => romdata <= X"C339FD3D";
    when 16#00542# => romdata <= X"0D81C1F4";
    when 16#00543# => romdata <= X"0852F881";
    when 16#00544# => romdata <= X"C08E800B";
    when 16#00545# => romdata <= X"81B29C08";
    when 16#00546# => romdata <= X"55537180";
    when 16#00547# => romdata <= X"2E80F738";
    when 16#00548# => romdata <= X"7281FF06";
    when 16#00549# => romdata <= X"84150C81";
    when 16#0054A# => romdata <= X"B1D83370";
    when 16#0054B# => romdata <= X"81FF0651";
    when 16#0054C# => romdata <= X"5271802E";
    when 16#0054D# => romdata <= X"80C23872";
    when 16#0054E# => romdata <= X"9F2A7310";
    when 16#0054F# => romdata <= X"075381C1";
    when 16#00550# => romdata <= X"F8337081";
    when 16#00551# => romdata <= X"FF065152";
    when 16#00552# => romdata <= X"71802ED4";
    when 16#00553# => romdata <= X"38800B81";
    when 16#00554# => romdata <= X"C1F83490";
    when 16#00555# => romdata <= X"883F81B1";
    when 16#00556# => romdata <= X"E8335473";
    when 16#00557# => romdata <= X"80E23881";
    when 16#00558# => romdata <= X"B29C0873";
    when 16#00559# => romdata <= X"81FF0684";
    when 16#0055A# => romdata <= X"120C81B1";
    when 16#0055B# => romdata <= X"D8337081";
    when 16#0055C# => romdata <= X"FF065153";
    when 16#0055D# => romdata <= X"5471C038";
    when 16#0055E# => romdata <= X"72812A73";
    when 16#0055F# => romdata <= X"9F2B0753";
    when 16#00560# => romdata <= X"FFBC3972";
    when 16#00561# => romdata <= X"812A739F";
    when 16#00562# => romdata <= X"2B075380";
    when 16#00563# => romdata <= X"FD51BD81";
    when 16#00564# => romdata <= X"3F81B29C";
    when 16#00565# => romdata <= X"08547281";
    when 16#00566# => romdata <= X"FF068415";
    when 16#00567# => romdata <= X"0C81B1D8";
    when 16#00568# => romdata <= X"337081FF";
    when 16#00569# => romdata <= X"06535471";
    when 16#0056A# => romdata <= X"802ED838";
    when 16#0056B# => romdata <= X"729F2A73";
    when 16#0056C# => romdata <= X"10075380";
    when 16#0056D# => romdata <= X"FD51BCD9";
    when 16#0056E# => romdata <= X"3F81B29C";
    when 16#0056F# => romdata <= X"0854D739";
    when 16#00570# => romdata <= X"800BB00C";
    when 16#00571# => romdata <= X"853D0D04";
    when 16#00572# => romdata <= X"F73D0D85";
    when 16#00573# => romdata <= X"3D549653";
    when 16#00574# => romdata <= X"81A1BC52";
    when 16#00575# => romdata <= X"735180C0";
    when 16#00576# => romdata <= X"BD3FA3B8";
    when 16#00577# => romdata <= X"3F81518A";
    when 16#00578# => romdata <= X"F73F8052";
    when 16#00579# => romdata <= X"8051A289";
    when 16#0057A# => romdata <= X"3F735380";
    when 16#0057B# => romdata <= X"5281A6BC";
    when 16#0057C# => romdata <= X"51B4F43F";
    when 16#0057D# => romdata <= X"80528151";
    when 16#0057E# => romdata <= X"A1F73F73";
    when 16#0057F# => romdata <= X"53825281";
    when 16#00580# => romdata <= X"A6BC51B4";
    when 16#00581# => romdata <= X"E23F8052";
    when 16#00582# => romdata <= X"8251A1E5";
    when 16#00583# => romdata <= X"3F735381";
    when 16#00584# => romdata <= X"5281A6BC";
    when 16#00585# => romdata <= X"51B4D03F";
    when 16#00586# => romdata <= X"80528451";
    when 16#00587# => romdata <= X"A1D33F73";
    when 16#00588# => romdata <= X"53845281";
    when 16#00589# => romdata <= X"A6BC51B4";
    when 16#0058A# => romdata <= X"BE3F8052";
    when 16#0058B# => romdata <= X"8551A1C1";
    when 16#0058C# => romdata <= X"3F735390";
    when 16#0058D# => romdata <= X"5281A6BC";
    when 16#0058E# => romdata <= X"51B4AC3F";
    when 16#0058F# => romdata <= X"80528651";
    when 16#00590# => romdata <= X"A1AF3F73";
    when 16#00591# => romdata <= X"53835281";
    when 16#00592# => romdata <= X"A6BC51B4";
    when 16#00593# => romdata <= X"9A3F8B3D";
    when 16#00594# => romdata <= X"0D04FEF4";
    when 16#00595# => romdata <= X"3F800BB0";
    when 16#00596# => romdata <= X"0C04FC3D";
    when 16#00597# => romdata <= X"0D818DEC";
    when 16#00598# => romdata <= X"54805584";
    when 16#00599# => romdata <= X"527451A1";
    when 16#0059A# => romdata <= X"883F8053";
    when 16#0059B# => romdata <= X"73708105";
    when 16#0059C# => romdata <= X"553351A2";
    when 16#0059D# => romdata <= X"823F8113";
    when 16#0059E# => romdata <= X"7081FF06";
    when 16#0059F# => romdata <= X"515380DC";
    when 16#005A0# => romdata <= X"7327E938";
    when 16#005A1# => romdata <= X"81157081";
    when 16#005A2# => romdata <= X"FF065653";
    when 16#005A3# => romdata <= X"877527D3";
    when 16#005A4# => romdata <= X"38800BB0";
    when 16#005A5# => romdata <= X"0C863D0D";
    when 16#005A6# => romdata <= X"04FD3D0D";
    when 16#005A7# => romdata <= X"81B1D833";
    when 16#005A8# => romdata <= X"7081FF06";
    when 16#005A9# => romdata <= X"5454729F";
    when 16#005AA# => romdata <= X"26AB3881";
    when 16#005AB# => romdata <= X"B1D83370";
    when 16#005AC# => romdata <= X"81FF0681";
    when 16#005AD# => romdata <= X"B1DC0852";
    when 16#005AE# => romdata <= X"88120C54";
    when 16#005AF# => romdata <= X"80E452AD";
    when 16#005B0# => romdata <= X"99518DF9";
    when 16#005B1# => romdata <= X"3F81B1D8";
    when 16#005B2# => romdata <= X"33810553";
    when 16#005B3# => romdata <= X"7281B1D8";
    when 16#005B4# => romdata <= X"34853D0D";
    when 16#005B5# => romdata <= X"0480E452";
    when 16#005B6# => romdata <= X"ADEE518D";
    when 16#005B7# => romdata <= X"E03F81B1";
    when 16#005B8# => romdata <= X"D8338105";
    when 16#005B9# => romdata <= X"537281B1";
    when 16#005BA# => romdata <= X"D834853D";
    when 16#005BB# => romdata <= X"0D04FD3D";
    when 16#005BC# => romdata <= X"0D81B1D8";
    when 16#005BD# => romdata <= X"337081FF";
    when 16#005BE# => romdata <= X"06545472";
    when 16#005BF# => romdata <= X"9F26B738";
    when 16#005C0# => romdata <= X"81B1D833";
    when 16#005C1# => romdata <= X"7081FF06";
    when 16#005C2# => romdata <= X"81B1DC08";
    when 16#005C3# => romdata <= X"5688160C";
    when 16#005C4# => romdata <= X"5381B1D8";
    when 16#005C5# => romdata <= X"33810554";
    when 16#005C6# => romdata <= X"7381B1D8";
    when 16#005C7# => romdata <= X"3481B1D8";
    when 16#005C8# => romdata <= X"33BF0654";
    when 16#005C9# => romdata <= X"7381B1D8";
    when 16#005CA# => romdata <= X"3480E452";
    when 16#005CB# => romdata <= X"ADEE518D";
    when 16#005CC# => romdata <= X"8C3F853D";
    when 16#005CD# => romdata <= X"0D0481B1";
    when 16#005CE# => romdata <= X"D8337081";
    when 16#005CF# => romdata <= X"FF06BF71";
    when 16#005D0# => romdata <= X"3181B1DC";
    when 16#005D1# => romdata <= X"08528812";
    when 16#005D2# => romdata <= X"0C555381";
    when 16#005D3# => romdata <= X"B1D83381";
    when 16#005D4# => romdata <= X"05547381";
    when 16#005D5# => romdata <= X"B1D83481";
    when 16#005D6# => romdata <= X"B1D833BF";
    when 16#005D7# => romdata <= X"06547381";
    when 16#005D8# => romdata <= X"B1D83480";
    when 16#005D9# => romdata <= X"E452ADEE";
    when 16#005DA# => romdata <= X"518CD23F";
    when 16#005DB# => romdata <= X"853D0D04";
    when 16#005DC# => romdata <= X"810B81B1";
    when 16#005DD# => romdata <= X"E83404FE";
    when 16#005DE# => romdata <= X"3D0D81B2";
    when 16#005DF# => romdata <= X"A0089811";
    when 16#005E0# => romdata <= X"0870842A";
    when 16#005E1# => romdata <= X"70810651";
    when 16#005E2# => romdata <= X"53535370";
    when 16#005E3# => romdata <= X"802E8D38";
    when 16#005E4# => romdata <= X"71EF0698";
    when 16#005E5# => romdata <= X"140C810B";
    when 16#005E6# => romdata <= X"81C1F834";
    when 16#005E7# => romdata <= X"843D0D04";
    when 16#005E8# => romdata <= X"FC3D0D81";
    when 16#005E9# => romdata <= X"B29C0870";
    when 16#005EA# => romdata <= X"08810A06";
    when 16#005EB# => romdata <= X"81C1F40C";
    when 16#005EC# => romdata <= X"53B9813F";
    when 16#005ED# => romdata <= X"B9A43F8D";
    when 16#005EE# => romdata <= X"C13F81B2";
    when 16#005EF# => romdata <= X"A0089811";
    when 16#005F0# => romdata <= X"08880798";
    when 16#005F1# => romdata <= X"120C5481";
    when 16#005F2# => romdata <= X"C1F40880";
    when 16#005F3# => romdata <= X"E4CE5553";
    when 16#005F4# => romdata <= X"72843888";
    when 16#005F5# => romdata <= X"80547381";
    when 16#005F6# => romdata <= X"D5F40C72";
    when 16#005F7# => romdata <= X"802E82E4";
    when 16#005F8# => romdata <= X"38819ACC";
    when 16#005F9# => romdata <= X"51B5973F";
    when 16#005FA# => romdata <= X"8C51B4F8";
    when 16#005FB# => romdata <= X"3F81A1BC";
    when 16#005FC# => romdata <= X"51B58B3F";
    when 16#005FD# => romdata <= X"81C1F408";
    when 16#005FE# => romdata <= X"802E81B7";
    when 16#005FF# => romdata <= X"3881A1D4";
    when 16#00600# => romdata <= X"51B4FB3F";
    when 16#00601# => romdata <= X"81C1F408";
    when 16#00602# => romdata <= X"802E8295";
    when 16#00603# => romdata <= X"3881B29C";
    when 16#00604# => romdata <= X"08841108";
    when 16#00605# => romdata <= X"55558053";
    when 16#00606# => romdata <= X"73FE8F0A";
    when 16#00607# => romdata <= X"0673982B";
    when 16#00608# => romdata <= X"07708417";
    when 16#00609# => romdata <= X"0C811470";
    when 16#0060A# => romdata <= X"81FF0651";
    when 16#0060B# => romdata <= X"54548F73";
    when 16#0060C# => romdata <= X"27E63883";
    when 16#0060D# => romdata <= X"52AEF051";
    when 16#0060E# => romdata <= X"8B833FF8";
    when 16#0060F# => romdata <= X"81C08E80";
    when 16#00610# => romdata <= X"0B81B29C";
    when 16#00611# => romdata <= X"08565481";
    when 16#00612# => romdata <= X"C1F40880";
    when 16#00613# => romdata <= X"2E81A838";
    when 16#00614# => romdata <= X"7381FF06";
    when 16#00615# => romdata <= X"84160C81";
    when 16#00616# => romdata <= X"B1D83370";
    when 16#00617# => romdata <= X"81FF0651";
    when 16#00618# => romdata <= X"5372802E";
    when 16#00619# => romdata <= X"80C23873";
    when 16#0061A# => romdata <= X"9F2A7410";
    when 16#0061B# => romdata <= X"075481C1";
    when 16#0061C# => romdata <= X"F8337081";
    when 16#0061D# => romdata <= X"FF065153";
    when 16#0061E# => romdata <= X"72802ED4";
    when 16#0061F# => romdata <= X"38800B81";
    when 16#00620# => romdata <= X"C1F83489";
    when 16#00621# => romdata <= X"D83F81B1";
    when 16#00622# => romdata <= X"E8335574";
    when 16#00623# => romdata <= X"81C23881";
    when 16#00624# => romdata <= X"B29C0874";
    when 16#00625# => romdata <= X"81FF0684";
    when 16#00626# => romdata <= X"120C81B1";
    when 16#00627# => romdata <= X"D8337081";
    when 16#00628# => romdata <= X"FF065154";
    when 16#00629# => romdata <= X"5572C038";
    when 16#0062A# => romdata <= X"73812A74";
    when 16#0062B# => romdata <= X"9F2B0754";
    when 16#0062C# => romdata <= X"FFBC3981";
    when 16#0062D# => romdata <= X"A1E051B3";
    when 16#0062E# => romdata <= X"C53F81A2";
    when 16#0062F# => romdata <= X"8451B3BE";
    when 16#00630# => romdata <= X"3FB451B5";
    when 16#00631# => romdata <= X"833F81A2";
    when 16#00632# => romdata <= X"9451B3B2";
    when 16#00633# => romdata <= X"3F81A29C";
    when 16#00634# => romdata <= X"51B3AB3F";
    when 16#00635# => romdata <= X"81A2A851";
    when 16#00636# => romdata <= X"B3A43F81";
    when 16#00637# => romdata <= X"C1F408FE";
    when 16#00638# => romdata <= X"AC38BE39";
    when 16#00639# => romdata <= X"73812A74";
    when 16#0063A# => romdata <= X"9F2B0754";
    when 16#0063B# => romdata <= X"80FD51B6";
    when 16#0063C# => romdata <= X"A03F81B2";
    when 16#0063D# => romdata <= X"9C085573";
    when 16#0063E# => romdata <= X"81FF0684";
    when 16#0063F# => romdata <= X"160C81B1";
    when 16#00640# => romdata <= X"D8337081";
    when 16#00641# => romdata <= X"FF065653";
    when 16#00642# => romdata <= X"74802ED8";
    when 16#00643# => romdata <= X"38739F2A";
    when 16#00644# => romdata <= X"74100754";
    when 16#00645# => romdata <= X"80FD51B5";
    when 16#00646# => romdata <= X"F83F81B2";
    when 16#00647# => romdata <= X"9C0855D7";
    when 16#00648# => romdata <= X"39B6D852";
    when 16#00649# => romdata <= X"ACDA5189";
    when 16#0064A# => romdata <= X"943F87E8";
    when 16#0064B# => romdata <= X"52AD9951";
    when 16#0064C# => romdata <= X"898B3FD5";
    when 16#0064D# => romdata <= X"E63F81B2";
    when 16#0064E# => romdata <= X"9C088411";
    when 16#0064F# => romdata <= X"08555580";
    when 16#00650# => romdata <= X"53FDD539";
    when 16#00651# => romdata <= X"B7D23F99";
    when 16#00652# => romdata <= X"B03F9CC8";
    when 16#00653# => romdata <= X"3FFD9239";
    when 16#00654# => romdata <= X"B9B73F80";
    when 16#00655# => romdata <= X"0B81D590";
    when 16#00656# => romdata <= X"34800B81";
    when 16#00657# => romdata <= X"D58C3480";
    when 16#00658# => romdata <= X"0B81D594";
    when 16#00659# => romdata <= X"0C04FC3D";
    when 16#0065A# => romdata <= X"0D765281";
    when 16#0065B# => romdata <= X"D58C3370";
    when 16#0065C# => romdata <= X"10101071";
    when 16#0065D# => romdata <= X"100581C1";
    when 16#0065E# => romdata <= X"FC055254";
    when 16#0065F# => romdata <= X"BEA63F77";
    when 16#00660# => romdata <= X"5281D58C";
    when 16#00661# => romdata <= X"33709029";
    when 16#00662# => romdata <= X"71317010";
    when 16#00663# => romdata <= X"1081C4BC";
    when 16#00664# => romdata <= X"05535555";
    when 16#00665# => romdata <= X"BE8E3F81";
    when 16#00666# => romdata <= X"D58C3370";
    when 16#00667# => romdata <= X"101081D3";
    when 16#00668# => romdata <= X"BC057A71";
    when 16#00669# => romdata <= X"0C548105";
    when 16#0066A# => romdata <= X"537281D5";
    when 16#0066B# => romdata <= X"8C34863D";
    when 16#0066C# => romdata <= X"0D04803D";
    when 16#0066D# => romdata <= X"0D81A2DC";
    when 16#0066E# => romdata <= X"51B1C33F";
    when 16#0066F# => romdata <= X"823D0D04";
    when 16#00670# => romdata <= X"FE3D0D81";
    when 16#00671# => romdata <= X"D5940853";
    when 16#00672# => romdata <= X"72853884";
    when 16#00673# => romdata <= X"3D0D0472";
    when 16#00674# => romdata <= X"2DB00853";
    when 16#00675# => romdata <= X"800B81D5";
    when 16#00676# => romdata <= X"940CB008";
    when 16#00677# => romdata <= X"8C3881A2";
    when 16#00678# => romdata <= X"DC51B19A";
    when 16#00679# => romdata <= X"3F843D0D";
    when 16#0067A# => romdata <= X"0481A5F0";
    when 16#0067B# => romdata <= X"51B18F3F";
    when 16#0067C# => romdata <= X"7283FFFF";
    when 16#0067D# => romdata <= X"26AA3881";
    when 16#0067E# => romdata <= X"FF732796";
    when 16#0067F# => romdata <= X"38725290";
    when 16#00680# => romdata <= X"51B19E3F";
    when 16#00681# => romdata <= X"8A51B0DC";
    when 16#00682# => romdata <= X"3F81A2DC";
    when 16#00683# => romdata <= X"51B0EF3F";
    when 16#00684# => romdata <= X"D4397252";
    when 16#00685# => romdata <= X"8851B189";
    when 16#00686# => romdata <= X"3F8A51B0";
    when 16#00687# => romdata <= X"C73FEA39";
    when 16#00688# => romdata <= X"7252A051";
    when 16#00689# => romdata <= X"B0FB3F8A";
    when 16#0068A# => romdata <= X"51B0B93F";
    when 16#0068B# => romdata <= X"DC39FA3D";
    when 16#0068C# => romdata <= X"0D02A305";
    when 16#0068D# => romdata <= X"3356758D";
    when 16#0068E# => romdata <= X"2E80F438";
    when 16#0068F# => romdata <= X"75883270";
    when 16#00690# => romdata <= X"307780FF";
    when 16#00691# => romdata <= X"32703072";
    when 16#00692# => romdata <= X"80257180";
    when 16#00693# => romdata <= X"25075451";
    when 16#00694# => romdata <= X"56585574";
    when 16#00695# => romdata <= X"95389F76";
    when 16#00696# => romdata <= X"278C3881";
    when 16#00697# => romdata <= X"D5903355";
    when 16#00698# => romdata <= X"80CE7527";
    when 16#00699# => romdata <= X"AE38883D";
    when 16#0069A# => romdata <= X"0D0481D5";
    when 16#0069B# => romdata <= X"90335675";
    when 16#0069C# => romdata <= X"802EF338";
    when 16#0069D# => romdata <= X"8851AFEC";
    when 16#0069E# => romdata <= X"3FA051AF";
    when 16#0069F# => romdata <= X"E73F8851";
    when 16#006A0# => romdata <= X"AFE23F81";
    when 16#006A1# => romdata <= X"D59033FF";
    when 16#006A2# => romdata <= X"05577681";
    when 16#006A3# => romdata <= X"D5903488";
    when 16#006A4# => romdata <= X"3D0D0475";
    when 16#006A5# => romdata <= X"51AFCD3F";
    when 16#006A6# => romdata <= X"81D59033";
    when 16#006A7# => romdata <= X"81115557";
    when 16#006A8# => romdata <= X"7381D590";
    when 16#006A9# => romdata <= X"347581D4";
    when 16#006AA# => romdata <= X"BC183488";
    when 16#006AB# => romdata <= X"3D0D048A";
    when 16#006AC# => romdata <= X"51AFB13F";
    when 16#006AD# => romdata <= X"81D59033";
    when 16#006AE# => romdata <= X"81115654";
    when 16#006AF# => romdata <= X"7481D590";
    when 16#006B0# => romdata <= X"34800B81";
    when 16#006B1# => romdata <= X"D4BC1534";
    when 16#006B2# => romdata <= X"8056800B";
    when 16#006B3# => romdata <= X"81D4BC17";
    when 16#006B4# => romdata <= X"33565474";
    when 16#006B5# => romdata <= X"A02E8338";
    when 16#006B6# => romdata <= X"81547480";
    when 16#006B7# => romdata <= X"2E903873";
    when 16#006B8# => romdata <= X"802E8B38";
    when 16#006B9# => romdata <= X"81167081";
    when 16#006BA# => romdata <= X"FF065757";
    when 16#006BB# => romdata <= X"DD397580";
    when 16#006BC# => romdata <= X"2EBF3880";
    when 16#006BD# => romdata <= X"0B81D58C";
    when 16#006BE# => romdata <= X"33555574";
    when 16#006BF# => romdata <= X"7427AB38";
    when 16#006C0# => romdata <= X"73577410";
    when 16#006C1# => romdata <= X"10107510";
    when 16#006C2# => romdata <= X"05765481";
    when 16#006C3# => romdata <= X"D4BC5381";
    when 16#006C4# => romdata <= X"C1FC0551";
    when 16#006C5# => romdata <= X"BCDA3FB0";
    when 16#006C6# => romdata <= X"08802EA6";
    when 16#006C7# => romdata <= X"38811570";
    when 16#006C8# => romdata <= X"81FF0656";
    when 16#006C9# => romdata <= X"54767526";
    when 16#006CA# => romdata <= X"D93881A2";
    when 16#006CB# => romdata <= X"E051AECE";
    when 16#006CC# => romdata <= X"3F81A2DC";
    when 16#006CD# => romdata <= X"51AEC73F";
    when 16#006CE# => romdata <= X"800B81D5";
    when 16#006CF# => romdata <= X"9034883D";
    when 16#006D0# => romdata <= X"0D047410";
    when 16#006D1# => romdata <= X"1081D3BC";
    when 16#006D2# => romdata <= X"05700881";
    when 16#006D3# => romdata <= X"D5940C56";
    when 16#006D4# => romdata <= X"800B81D5";
    when 16#006D5# => romdata <= X"9034E739";
    when 16#006D6# => romdata <= X"F73D0D02";
    when 16#006D7# => romdata <= X"AF053359";
    when 16#006D8# => romdata <= X"800B81D4";
    when 16#006D9# => romdata <= X"BC3381D4";
    when 16#006DA# => romdata <= X"BC595556";
    when 16#006DB# => romdata <= X"73A02E09";
    when 16#006DC# => romdata <= X"81069638";
    when 16#006DD# => romdata <= X"81167081";
    when 16#006DE# => romdata <= X"FF0681D4";
    when 16#006DF# => romdata <= X"BC117033";
    when 16#006E0# => romdata <= X"53595754";
    when 16#006E1# => romdata <= X"73A02EEC";
    when 16#006E2# => romdata <= X"38805877";
    when 16#006E3# => romdata <= X"792780EA";
    when 16#006E4# => romdata <= X"38807733";
    when 16#006E5# => romdata <= X"56547474";
    when 16#006E6# => romdata <= X"2E833881";
    when 16#006E7# => romdata <= X"5474A02E";
    when 16#006E8# => romdata <= X"9A387380";
    when 16#006E9# => romdata <= X"C53874A0";
    when 16#006EA# => romdata <= X"2E913881";
    when 16#006EB# => romdata <= X"187081FF";
    when 16#006EC# => romdata <= X"06595578";
    when 16#006ED# => romdata <= X"7826DA38";
    when 16#006EE# => romdata <= X"80C03981";
    when 16#006EF# => romdata <= X"167081FF";
    when 16#006F0# => romdata <= X"0681D4BC";
    when 16#006F1# => romdata <= X"11703357";
    when 16#006F2# => romdata <= X"52575773";
    when 16#006F3# => romdata <= X"A02E0981";
    when 16#006F4# => romdata <= X"06D93881";
    when 16#006F5# => romdata <= X"167081FF";
    when 16#006F6# => romdata <= X"0681D4BC";
    when 16#006F7# => romdata <= X"11703357";
    when 16#006F8# => romdata <= X"52575773";
    when 16#006F9# => romdata <= X"A02ED438";
    when 16#006FA# => romdata <= X"C2398116";
    when 16#006FB# => romdata <= X"7081FF06";
    when 16#006FC# => romdata <= X"81D4BC11";
    when 16#006FD# => romdata <= X"595755FF";
    when 16#006FE# => romdata <= X"98398A53";
    when 16#006FF# => romdata <= X"8B3DFC05";
    when 16#00700# => romdata <= X"527651BF";
    when 16#00701# => romdata <= X"B03F8B3D";
    when 16#00702# => romdata <= X"0D04F73D";
    when 16#00703# => romdata <= X"0D02AF05";
    when 16#00704# => romdata <= X"3359800B";
    when 16#00705# => romdata <= X"81D4BC33";
    when 16#00706# => romdata <= X"81D4BC59";
    when 16#00707# => romdata <= X"555673A0";
    when 16#00708# => romdata <= X"2E098106";
    when 16#00709# => romdata <= X"96388116";
    when 16#0070A# => romdata <= X"7081FF06";
    when 16#0070B# => romdata <= X"81D4BC11";
    when 16#0070C# => romdata <= X"70335359";
    when 16#0070D# => romdata <= X"575473A0";
    when 16#0070E# => romdata <= X"2EEC3880";
    when 16#0070F# => romdata <= X"58777927";
    when 16#00710# => romdata <= X"80EA3880";
    when 16#00711# => romdata <= X"77335654";
    when 16#00712# => romdata <= X"74742E83";
    when 16#00713# => romdata <= X"38815474";
    when 16#00714# => romdata <= X"A02E9A38";
    when 16#00715# => romdata <= X"7380C538";
    when 16#00716# => romdata <= X"74A02E91";
    when 16#00717# => romdata <= X"38811870";
    when 16#00718# => romdata <= X"81FF0659";
    when 16#00719# => romdata <= X"55787826";
    when 16#0071A# => romdata <= X"DA3880C0";
    when 16#0071B# => romdata <= X"39811670";
    when 16#0071C# => romdata <= X"81FF0681";
    when 16#0071D# => romdata <= X"D4BC1170";
    when 16#0071E# => romdata <= X"33575257";
    when 16#0071F# => romdata <= X"5773A02E";
    when 16#00720# => romdata <= X"098106D9";
    when 16#00721# => romdata <= X"38811670";
    when 16#00722# => romdata <= X"81FF0681";
    when 16#00723# => romdata <= X"D4BC1170";
    when 16#00724# => romdata <= X"33575257";
    when 16#00725# => romdata <= X"5773A02E";
    when 16#00726# => romdata <= X"D438C239";
    when 16#00727# => romdata <= X"81167081";
    when 16#00728# => romdata <= X"FF0681D4";
    when 16#00729# => romdata <= X"BC115957";
    when 16#0072A# => romdata <= X"55FF9839";
    when 16#0072B# => romdata <= X"90538B3D";
    when 16#0072C# => romdata <= X"FC055276";
    when 16#0072D# => romdata <= X"5180C19A";
    when 16#0072E# => romdata <= X"3F8B3D0D";
    when 16#0072F# => romdata <= X"04FC3D0D";
    when 16#00730# => romdata <= X"8A51ABA0";
    when 16#00731# => romdata <= X"3F81A2F4";
    when 16#00732# => romdata <= X"51ABB33F";
    when 16#00733# => romdata <= X"800B81D5";
    when 16#00734# => romdata <= X"8C335353";
    when 16#00735# => romdata <= X"72722780";
    when 16#00736# => romdata <= X"F5387210";
    when 16#00737# => romdata <= X"10107310";
    when 16#00738# => romdata <= X"0581C1FC";
    when 16#00739# => romdata <= X"05705254";
    when 16#0073A# => romdata <= X"AB943F72";
    when 16#0073B# => romdata <= X"842B7074";
    when 16#0073C# => romdata <= X"31822B81";
    when 16#0073D# => romdata <= X"C4BC1133";
    when 16#0073E# => romdata <= X"51535571";
    when 16#0073F# => romdata <= X"802EB738";
    when 16#00740# => romdata <= X"7351B88D";
    when 16#00741# => romdata <= X"3FB00881";
    when 16#00742# => romdata <= X"FF065271";
    when 16#00743# => romdata <= X"89269338";
    when 16#00744# => romdata <= X"A051AAD0";
    when 16#00745# => romdata <= X"3F811270";
    when 16#00746# => romdata <= X"81FF0653";
    when 16#00747# => romdata <= X"54897227";
    when 16#00748# => romdata <= X"EF3881A3";
    when 16#00749# => romdata <= X"8C51AAD6";
    when 16#0074A# => romdata <= X"3F747331";
    when 16#0074B# => romdata <= X"822B81C4";
    when 16#0074C# => romdata <= X"BC0551AA";
    when 16#0074D# => romdata <= X"C93F8A51";
    when 16#0074E# => romdata <= X"AAAA3F81";
    when 16#0074F# => romdata <= X"137081FF";
    when 16#00750# => romdata <= X"0681D58C";
    when 16#00751# => romdata <= X"33545455";
    when 16#00752# => romdata <= X"717326FF";
    when 16#00753# => romdata <= X"8D388A51";
    when 16#00754# => romdata <= X"AA923F81";
    when 16#00755# => romdata <= X"D58C33B0";
    when 16#00756# => romdata <= X"0C863D0D";
    when 16#00757# => romdata <= X"04FE3D0D";
    when 16#00758# => romdata <= X"81D5EC22";
    when 16#00759# => romdata <= X"FF055170";
    when 16#0075A# => romdata <= X"81D5EC23";
    when 16#0075B# => romdata <= X"7083FFFF";
    when 16#0075C# => romdata <= X"06517080";
    when 16#0075D# => romdata <= X"C43881D5";
    when 16#0075E# => romdata <= X"F0335170";
    when 16#0075F# => romdata <= X"81FF2EB9";
    when 16#00760# => romdata <= X"38701010";
    when 16#00761# => romdata <= X"1081D59C";
    when 16#00762# => romdata <= X"05527133";
    when 16#00763# => romdata <= X"81D5F034";
    when 16#00764# => romdata <= X"FE723481";
    when 16#00765# => romdata <= X"D5F03370";
    when 16#00766# => romdata <= X"10101081";
    when 16#00767# => romdata <= X"D59C0552";
    when 16#00768# => romdata <= X"53821122";
    when 16#00769# => romdata <= X"81D5EC23";
    when 16#0076A# => romdata <= X"84120853";
    when 16#0076B# => romdata <= X"722D81D5";
    when 16#0076C# => romdata <= X"EC225170";
    when 16#0076D# => romdata <= X"802EFFBE";
    when 16#0076E# => romdata <= X"38843D0D";
    when 16#0076F# => romdata <= X"04F93D0D";
    when 16#00770# => romdata <= X"02AA0522";
    when 16#00771# => romdata <= X"56805574";
    when 16#00772# => romdata <= X"10101081";
    when 16#00773# => romdata <= X"D59C0570";
    when 16#00774# => romdata <= X"33525270";
    when 16#00775# => romdata <= X"81FE2E99";
    when 16#00776# => romdata <= X"38811570";
    when 16#00777# => romdata <= X"81FF0656";
    when 16#00778# => romdata <= X"52748A2E";
    when 16#00779# => romdata <= X"098106DF";
    when 16#0077A# => romdata <= X"38810BB0";
    when 16#0077B# => romdata <= X"0C893D0D";
    when 16#0077C# => romdata <= X"0481D5F0";
    when 16#0077D# => romdata <= X"337081FF";
    when 16#0077E# => romdata <= X"0681D5EC";
    when 16#0077F# => romdata <= X"22535458";
    when 16#00780# => romdata <= X"7281FF2E";
    when 16#00781# => romdata <= X"B0387283";
    when 16#00782# => romdata <= X"2B547076";
    when 16#00783# => romdata <= X"2780DE38";
    when 16#00784# => romdata <= X"75713170";
    when 16#00785# => romdata <= X"83FFFF06";
    when 16#00786# => romdata <= X"7481D59C";
    when 16#00787# => romdata <= X"17337083";
    when 16#00788# => romdata <= X"2B81D59E";
    when 16#00789# => romdata <= X"11225658";
    when 16#0078A# => romdata <= X"56525757";
    when 16#0078B# => romdata <= X"7281FF2E";
    when 16#0078C# => romdata <= X"098106D6";
    when 16#0078D# => romdata <= X"38727234";
    when 16#0078E# => romdata <= X"75821323";
    when 16#0078F# => romdata <= X"7984130C";
    when 16#00790# => romdata <= X"7781FF06";
    when 16#00791# => romdata <= X"5473732E";
    when 16#00792# => romdata <= X"96387610";
    when 16#00793# => romdata <= X"101081D5";
    when 16#00794# => romdata <= X"9C055374";
    when 16#00795# => romdata <= X"73348051";
    when 16#00796# => romdata <= X"70B00C89";
    when 16#00797# => romdata <= X"3D0D0474";
    when 16#00798# => romdata <= X"81D5F034";
    when 16#00799# => romdata <= X"7581D5EC";
    when 16#0079A# => romdata <= X"238051EC";
    when 16#0079B# => romdata <= X"39707631";
    when 16#0079C# => romdata <= X"517081D5";
    when 16#0079D# => romdata <= X"9E1523FF";
    when 16#0079E# => romdata <= X"BC39FF3D";
    when 16#0079F# => romdata <= X"0D8A5271";
    when 16#007A0# => romdata <= X"10101081";
    when 16#007A1# => romdata <= X"D5940551";
    when 16#007A2# => romdata <= X"FE7134FF";
    when 16#007A3# => romdata <= X"127081FF";
    when 16#007A4# => romdata <= X"06535171";
    when 16#007A5# => romdata <= X"EA38FF0B";
    when 16#007A6# => romdata <= X"81D5F034";
    when 16#007A7# => romdata <= X"833D0D04";
    when 16#007A8# => romdata <= X"F53D0D7D";
    when 16#007A9# => romdata <= X"598A5481";
    when 16#007AA# => romdata <= X"028405BA";
    when 16#007AB# => romdata <= X"0522575C";
    when 16#007AC# => romdata <= X"80E45380";
    when 16#007AD# => romdata <= X"52ABB93F";
    when 16#007AE# => romdata <= X"B008722E";
    when 16#007AF# => romdata <= X"09810683";
    when 16#007B0# => romdata <= X"38815272";
    when 16#007B1# => romdata <= X"802EB138";
    when 16#007B2# => romdata <= X"71802E91";
    when 16#007B3# => romdata <= X"3880E451";
    when 16#007B4# => romdata <= X"AABF3FFF";
    when 16#007B5# => romdata <= X"137081FF";
    when 16#007B6# => romdata <= X"065452D7";
    when 16#007B7# => romdata <= X"3972802E";
    when 16#007B8# => romdata <= X"9738AB9F";
    when 16#007B9# => romdata <= X"3FB00881";
    when 16#007BA# => romdata <= X"FF065271";
    when 16#007BB# => romdata <= X"952E829A";
    when 16#007BC# => romdata <= X"387180C3";
    when 16#007BD# => romdata <= X"2E81EC38";
    when 16#007BE# => romdata <= X"FF147081";
    when 16#007BF# => romdata <= X"FF065553";
    when 16#007C0# => romdata <= X"73FFAD38";
    when 16#007C1# => romdata <= X"75802E81";
    when 16#007C2# => romdata <= X"CC388A7C";
    when 16#007C3# => romdata <= X"095C5A81";
    when 16#007C4# => romdata <= X"51AB923F";
    when 16#007C5# => romdata <= X"7B51AB8D";
    when 16#007C6# => romdata <= X"3F7A51AB";
    when 16#007C7# => romdata <= X"883F8070";
    when 16#007C8# => romdata <= X"55578180";
    when 16#007C9# => romdata <= X"55FF1570";
    when 16#007CA# => romdata <= X"81FF0656";
    when 16#007CB# => romdata <= X"529A5375";
    when 16#007CC# => romdata <= X"802E9138";
    when 16#007CD# => romdata <= X"78708105";
    when 16#007CE# => romdata <= X"5A33FF17";
    when 16#007CF# => romdata <= X"7083FFFF";
    when 16#007D0# => romdata <= X"06585353";
    when 16#007D1# => romdata <= X"7251AADD";
    when 16#007D2# => romdata <= X"3F77802E";
    when 16#007D3# => romdata <= X"81A93872";
    when 16#007D4# => romdata <= X"882B7432";
    when 16#007D5# => romdata <= X"53875472";
    when 16#007D6# => romdata <= X"902B5280";
    when 16#007D7# => romdata <= X"72248188";
    when 16#007D8# => romdata <= X"38721083";
    when 16#007D9# => romdata <= X"FFFE0653";
    when 16#007DA# => romdata <= X"FF145473";
    when 16#007DB# => romdata <= X"8025E838";
    when 16#007DC# => romdata <= X"7283FFFF";
    when 16#007DD# => romdata <= X"065474FF";
    when 16#007DE# => romdata <= X"AC387780";
    when 16#007DF# => romdata <= X"2E818338";
    when 16#007E0# => romdata <= X"73882A51";
    when 16#007E1# => romdata <= X"AA9F3F73";
    when 16#007E2# => romdata <= X"81FF0651";
    when 16#007E3# => romdata <= X"AA973FA9";
    when 16#007E4# => romdata <= X"DF3FB008";
    when 16#007E5# => romdata <= X"FA38A9EB";
    when 16#007E6# => romdata <= X"3FB00881";
    when 16#007E7# => romdata <= X"FF065271";
    when 16#007E8# => romdata <= X"862E80EB";
    when 16#007E9# => romdata <= X"3871982E";
    when 16#007EA# => romdata <= X"80F038FF";
    when 16#007EB# => romdata <= X"1A7081FF";
    when 16#007EC# => romdata <= X"065B5479";
    when 16#007ED# => romdata <= X"FED938FE";
    when 16#007EE# => romdata <= X"5271B00C";
    when 16#007EF# => romdata <= X"8D3D0D04";
    when 16#007F0# => romdata <= X"A9AE3FB0";
    when 16#007F1# => romdata <= X"08FA38A9";
    when 16#007F2# => romdata <= X"BA3FB008";
    when 16#007F3# => romdata <= X"81FF0652";
    when 16#007F4# => romdata <= X"71862EE5";
    when 16#007F5# => romdata <= X"388451A9";
    when 16#007F6# => romdata <= X"CC3FA994";
    when 16#007F7# => romdata <= X"3FB008E0";
    when 16#007F8# => romdata <= X"38E53981";
    when 16#007F9# => romdata <= X"58FE9D39";
    when 16#007FA# => romdata <= X"7210A0A1";
    when 16#007FB# => romdata <= X"327083FF";
    when 16#007FC# => romdata <= X"FF065452";
    when 16#007FD# => romdata <= X"FEF23972";
    when 16#007FE# => romdata <= X"177081FF";
    when 16#007FF# => romdata <= X"065852FE";
    when 16#00800# => romdata <= X"F5397651";
    when 16#00801# => romdata <= X"A99F3FFF";
    when 16#00802# => romdata <= X"86398058";
    when 16#00803# => romdata <= X"FDF63981";
    when 16#00804# => romdata <= X"1C7081FF";
    when 16#00805# => romdata <= X"065D55FD";
    when 16#00806# => romdata <= X"EB39FF0B";
    when 16#00807# => romdata <= X"B00C8D3D";
    when 16#00808# => romdata <= X"0D04F63D";
    when 16#00809# => romdata <= X"0D7C7E5B";
    when 16#0080A# => romdata <= X"5980C357";
    when 16#0080B# => romdata <= X"8A55815B";
    when 16#0080C# => romdata <= X"805880E4";
    when 16#0080D# => romdata <= X"53805477";
    when 16#0080E# => romdata <= X"7A2482AA";
    when 16#0080F# => romdata <= X"387651A8";
    when 16#00810# => romdata <= X"E43F8052";
    when 16#00811# => romdata <= X"A8AA3FB0";
    when 16#00812# => romdata <= X"08722E09";
    when 16#00813# => romdata <= X"81068338";
    when 16#00814# => romdata <= X"81527280";
    when 16#00815# => romdata <= X"2E81E638";
    when 16#00816# => romdata <= X"71802E91";
    when 16#00817# => romdata <= X"3880E451";
    when 16#00818# => romdata <= X"A7AF3FFF";
    when 16#00819# => romdata <= X"137081FF";
    when 16#0081A# => romdata <= X"065452D6";
    when 16#0081B# => romdata <= X"3972802E";
    when 16#0081C# => romdata <= X"81CB38A8";
    when 16#0081D# => romdata <= X"8E3FB008";
    when 16#0081E# => romdata <= X"81FF0652";
    when 16#0081F# => romdata <= X"71842E82";
    when 16#00820# => romdata <= X"81387184";
    when 16#00821# => romdata <= X"2481CA38";
    when 16#00822# => romdata <= X"71812E09";
    when 16#00823# => romdata <= X"810681AD";
    when 16#00824# => romdata <= X"388657A7";
    when 16#00825# => romdata <= X"EE3FB008";
    when 16#00826# => romdata <= X"81FF0653";
    when 16#00827# => romdata <= X"7A732E83";
    when 16#00828# => romdata <= X"389557A7";
    when 16#00829# => romdata <= X"DE3FB008";
    when 16#0082A# => romdata <= X"097081FF";
    when 16#0082B# => romdata <= X"0657527A";
    when 16#0082C# => romdata <= X"762E8338";
    when 16#0082D# => romdata <= X"95578053";
    when 16#0082E# => romdata <= X"A7C93F78";
    when 16#0082F# => romdata <= X"1356B008";
    when 16#00830# => romdata <= X"76348113";
    when 16#00831# => romdata <= X"7081FF06";
    when 16#00832# => romdata <= X"70982B58";
    when 16#00833# => romdata <= X"54527580";
    when 16#00834# => romdata <= X"25E63880";
    when 16#00835# => romdata <= X"56781670";
    when 16#00836# => romdata <= X"3370882B";
    when 16#00837# => romdata <= X"76325253";
    when 16#00838# => romdata <= X"53875472";
    when 16#00839# => romdata <= X"902B5280";
    when 16#0083A# => romdata <= X"72248187";
    when 16#0083B# => romdata <= X"38721083";
    when 16#0083C# => romdata <= X"FFFE0653";
    when 16#0083D# => romdata <= X"FF145473";
    when 16#0083E# => romdata <= X"8025E838";
    when 16#0083F# => romdata <= X"7283FFFF";
    when 16#00840# => romdata <= X"06811770";
    when 16#00841# => romdata <= X"81FF0670";
    when 16#00842# => romdata <= X"982B5658";
    when 16#00843# => romdata <= X"53547280";
    when 16#00844# => romdata <= X"25C338A6";
    when 16#00845# => romdata <= X"EE3FB008";
    when 16#00846# => romdata <= X"81FF0674";
    when 16#00847# => romdata <= X"882A5753";
    when 16#00848# => romdata <= X"72762E83";
    when 16#00849# => romdata <= X"389557A6";
    when 16#0084A# => romdata <= X"DA3FB008";
    when 16#0084B# => romdata <= X"81FF0674";
    when 16#0084C# => romdata <= X"81FF0653";
    when 16#0084D# => romdata <= X"5675722E";
    when 16#0084E# => romdata <= X"80D43895";
    when 16#0084F# => romdata <= X"57FF1570";
    when 16#00850# => romdata <= X"81FF0656";
    when 16#00851# => romdata <= X"5274FDEA";
    when 16#00852# => romdata <= X"38FE0BB0";
    when 16#00853# => romdata <= X"0C8C3D0D";
    when 16#00854# => romdata <= X"0471982E";
    when 16#00855# => romdata <= X"098106E5";
    when 16#00856# => romdata <= X"388651A6";
    when 16#00857# => romdata <= X"C83FFF0B";
    when 16#00858# => romdata <= X"B00C8C3D";
    when 16#00859# => romdata <= X"0D049851";
    when 16#0085A# => romdata <= X"A6BB3FFD";
    when 16#0085B# => romdata <= X"0BB00C8C";
    when 16#0085C# => romdata <= X"3D0D0472";
    when 16#0085D# => romdata <= X"10A0A132";
    when 16#0085E# => romdata <= X"7083FFFF";
    when 16#0085F# => romdata <= X"065452FE";
    when 16#00860# => romdata <= X"F3398651";
    when 16#00861# => romdata <= X"A69F3F77";
    when 16#00862# => romdata <= X"B00C8C3D";
    when 16#00863# => romdata <= X"0D047686";
    when 16#00864# => romdata <= X"2E098106";
    when 16#00865# => romdata <= X"FFA73877";
    when 16#00866# => romdata <= X"84808029";
    when 16#00867# => romdata <= X"82800A05";
    when 16#00868# => romdata <= X"70902C81";
    when 16#00869# => romdata <= X"801B811E";
    when 16#0086A# => romdata <= X"7081FF06";
    when 16#0086B# => romdata <= X"5F575B59";
    when 16#0086C# => romdata <= X"5374FCFE";
    when 16#0086D# => romdata <= X"38FF9239";
    when 16#0086E# => romdata <= X"FE3D0D02";
    when 16#0086F# => romdata <= X"93053302";
    when 16#00870# => romdata <= X"84059705";
    when 16#00871# => romdata <= X"33545271";
    when 16#00872# => romdata <= X"812E9238";
    when 16#00873# => romdata <= X"7180D52E";
    when 16#00874# => romdata <= X"BB3881A3";
    when 16#00875# => romdata <= X"9051A1A6";
    when 16#00876# => romdata <= X"3F843D0D";
    when 16#00877# => romdata <= X"0481A39C";
    when 16#00878# => romdata <= X"51A19B3F";
    when 16#00879# => romdata <= X"72912E81";
    when 16#0087A# => romdata <= X"D9387291";
    when 16#0087B# => romdata <= X"24B53872";
    when 16#0087C# => romdata <= X"8C2E81E4";
    when 16#0087D# => romdata <= X"38728C24";
    when 16#0087E# => romdata <= X"80DC3872";
    when 16#0087F# => romdata <= X"862E81B7";
    when 16#00880# => romdata <= X"3881A3A8";
    when 16#00881# => romdata <= X"51A0F73F";
    when 16#00882# => romdata <= X"843D0D04";
    when 16#00883# => romdata <= X"81A3B851";
    when 16#00884# => romdata <= X"A0EC3F72";
    when 16#00885# => romdata <= X"8726EA38";
    when 16#00886# => romdata <= X"72101081";
    when 16#00887# => romdata <= X"A69C0552";
    when 16#00888# => romdata <= X"71080472";
    when 16#00889# => romdata <= X"A82E81A5";
    when 16#0088A# => romdata <= X"3872A824";
    when 16#0088B# => romdata <= X"9438729A";
    when 16#0088C# => romdata <= X"2E098106";
    when 16#0088D# => romdata <= X"CC3881A3";
    when 16#0088E# => romdata <= X"C451A0C2";
    when 16#0088F# => romdata <= X"3F843D0D";
    when 16#00890# => romdata <= X"047280E1";
    when 16#00891# => romdata <= X"2E098106";
    when 16#00892# => romdata <= X"FFB73881";
    when 16#00893# => romdata <= X"A3E051A0";
    when 16#00894# => romdata <= X"AD3F843D";
    when 16#00895# => romdata <= X"0D04728F";
    when 16#00896# => romdata <= X"2E098106";
    when 16#00897# => romdata <= X"FFA33881";
    when 16#00898# => romdata <= X"A3F051A0";
    when 16#00899# => romdata <= X"993F843D";
    when 16#0089A# => romdata <= X"0D0481A4";
    when 16#0089B# => romdata <= X"8C51A08E";
    when 16#0089C# => romdata <= X"3F843D0D";
    when 16#0089D# => romdata <= X"0481A1BC";
    when 16#0089E# => romdata <= X"51A0833F";
    when 16#0089F# => romdata <= X"843D0D04";
    when 16#008A0# => romdata <= X"81A4A451";
    when 16#008A1# => romdata <= X"9FF83F84";
    when 16#008A2# => romdata <= X"3D0D0481";
    when 16#008A3# => romdata <= X"A4B8519F";
    when 16#008A4# => romdata <= X"ED3F843D";
    when 16#008A5# => romdata <= X"0D0481A4";
    when 16#008A6# => romdata <= X"C8519FE2";
    when 16#008A7# => romdata <= X"3F843D0D";
    when 16#008A8# => romdata <= X"0481A4E0";
    when 16#008A9# => romdata <= X"519FD73F";
    when 16#008AA# => romdata <= X"843D0D04";
    when 16#008AB# => romdata <= X"81A4F451";
    when 16#008AC# => romdata <= X"9FCC3F84";
    when 16#008AD# => romdata <= X"3D0D0481";
    when 16#008AE# => romdata <= X"A584519F";
    when 16#008AF# => romdata <= X"C13F843D";
    when 16#008B0# => romdata <= X"0D0481A5";
    when 16#008B1# => romdata <= X"94519FB6";
    when 16#008B2# => romdata <= X"3F843D0D";
    when 16#008B3# => romdata <= X"0481A5A8";
    when 16#008B4# => romdata <= X"519FAB3F";
    when 16#008B5# => romdata <= X"843D0D04";
    when 16#008B6# => romdata <= X"81A5C851";
    when 16#008B7# => romdata <= X"9FA03F84";
    when 16#008B8# => romdata <= X"3D0D04F7";
    when 16#008B9# => romdata <= X"3D0D02B3";
    when 16#008BA# => romdata <= X"05337C70";
    when 16#008BB# => romdata <= X"08C08080";
    when 16#008BC# => romdata <= X"0659545A";
    when 16#008BD# => romdata <= X"80567583";
    when 16#008BE# => romdata <= X"2B7707BF";
    when 16#008BF# => romdata <= X"E0800770";
    when 16#008C0# => romdata <= X"70840552";
    when 16#008C1# => romdata <= X"0871088C";
    when 16#008C2# => romdata <= X"2ABFFE80";
    when 16#008C3# => romdata <= X"06790771";
    when 16#008C4# => romdata <= X"982A728C";
    when 16#008C5# => romdata <= X"2A9FFF06";
    when 16#008C6# => romdata <= X"73852A70";
    when 16#008C7# => romdata <= X"8F06759F";
    when 16#008C8# => romdata <= X"06565158";
    when 16#008C9# => romdata <= X"5D585255";
    when 16#008CA# => romdata <= X"58748D38";
    when 16#008CB# => romdata <= X"8116568F";
    when 16#008CC# => romdata <= X"7627C338";
    when 16#008CD# => romdata <= X"8B3D0D04";
    when 16#008CE# => romdata <= X"81A5D851";
    when 16#008CF# => romdata <= X"9EC03F75";
    when 16#008D0# => romdata <= X"51A0853F";
    when 16#008D1# => romdata <= X"8452B008";
    when 16#008D2# => romdata <= X"51D0943F";
    when 16#008D3# => romdata <= X"81A5E451";
    when 16#008D4# => romdata <= X"9EAC3F74";
    when 16#008D5# => romdata <= X"5288519E";
    when 16#008D6# => romdata <= X"C83F8452";
    when 16#008D7# => romdata <= X"B00851CF";
    when 16#008D8# => romdata <= X"FE3F81A5";
    when 16#008D9# => romdata <= X"EC519E96";
    when 16#008DA# => romdata <= X"3F785290";
    when 16#008DB# => romdata <= X"519EB23F";
    when 16#008DC# => romdata <= X"8652B008";
    when 16#008DD# => romdata <= X"51CFE83F";
    when 16#008DE# => romdata <= X"81A5F451";
    when 16#008DF# => romdata <= X"9E803F72";
    when 16#008E0# => romdata <= X"519FC53F";
    when 16#008E1# => romdata <= X"8452B008";
    when 16#008E2# => romdata <= X"51CFD43F";
    when 16#008E3# => romdata <= X"81A5FC51";
    when 16#008E4# => romdata <= X"9DEC3F73";
    when 16#008E5# => romdata <= X"519FB13F";
    when 16#008E6# => romdata <= X"8452B008";
    when 16#008E7# => romdata <= X"51CFC03F";
    when 16#008E8# => romdata <= X"81A68451";
    when 16#008E9# => romdata <= X"9DD83F77";
    when 16#008EA# => romdata <= X"52A0519D";
    when 16#008EB# => romdata <= X"F43F8A52";
    when 16#008EC# => romdata <= X"B00851CF";
    when 16#008ED# => romdata <= X"AA3F7992";
    when 16#008EE# => romdata <= X"388A519D";
    when 16#008EF# => romdata <= X"A73F8116";
    when 16#008F0# => romdata <= X"568F7627";
    when 16#008F1# => romdata <= X"FEB038FE";
    when 16#008F2# => romdata <= X"EB397881";
    when 16#008F3# => romdata <= X"FF065274";
    when 16#008F4# => romdata <= X"51FBE53F";
    when 16#008F5# => romdata <= X"8A519D8C";
    when 16#008F6# => romdata <= X"3FE439F8";
    when 16#008F7# => romdata <= X"3D0D02AB";
    when 16#008F8# => romdata <= X"05335980";
    when 16#008F9# => romdata <= X"5675852B";
    when 16#008FA# => romdata <= X"E09011E0";
    when 16#008FB# => romdata <= X"80120870";
    when 16#008FC# => romdata <= X"982A718C";
    when 16#008FD# => romdata <= X"2A9FFF06";
    when 16#008FE# => romdata <= X"72852A70";
    when 16#008FF# => romdata <= X"8F06749F";
    when 16#00900# => romdata <= X"06555158";
    when 16#00901# => romdata <= X"5B535659";
    when 16#00902# => romdata <= X"5574802E";
    when 16#00903# => romdata <= X"81A13875";
    when 16#00904# => romdata <= X"BF2681A9";
    when 16#00905# => romdata <= X"3881A68C";
    when 16#00906# => romdata <= X"519CE33F";
    when 16#00907# => romdata <= X"75519EA8";
    when 16#00908# => romdata <= X"3F8652B0";
    when 16#00909# => romdata <= X"0851CEB7";
    when 16#0090A# => romdata <= X"3F81A5E4";
    when 16#0090B# => romdata <= X"519CCF3F";
    when 16#0090C# => romdata <= X"74528851";
    when 16#0090D# => romdata <= X"9CEB3F84";
    when 16#0090E# => romdata <= X"52B00851";
    when 16#0090F# => romdata <= X"CEA13F81";
    when 16#00910# => romdata <= X"A5EC519C";
    when 16#00911# => romdata <= X"B93F7652";
    when 16#00912# => romdata <= X"90519CD5";
    when 16#00913# => romdata <= X"3F8652B0";
    when 16#00914# => romdata <= X"0851CE8B";
    when 16#00915# => romdata <= X"3F81A5F4";
    when 16#00916# => romdata <= X"519CA33F";
    when 16#00917# => romdata <= X"72519DE8";
    when 16#00918# => romdata <= X"3F8452B0";
    when 16#00919# => romdata <= X"0851CDF7";
    when 16#0091A# => romdata <= X"3F81A5FC";
    when 16#0091B# => romdata <= X"519C8F3F";
    when 16#0091C# => romdata <= X"73519DD4";
    when 16#0091D# => romdata <= X"3F8452B0";
    when 16#0091E# => romdata <= X"0851CDE3";
    when 16#0091F# => romdata <= X"3F81A684";
    when 16#00920# => romdata <= X"519BFB3F";
    when 16#00921# => romdata <= X"7708C080";
    when 16#00922# => romdata <= X"800652A0";
    when 16#00923# => romdata <= X"519C923F";
    when 16#00924# => romdata <= X"8A52B008";
    when 16#00925# => romdata <= X"51CDC83F";
    when 16#00926# => romdata <= X"7881AC38";
    when 16#00927# => romdata <= X"8A519BC4";
    when 16#00928# => romdata <= X"3F805374";
    when 16#00929# => romdata <= X"812E81D9";
    when 16#0092A# => romdata <= X"3876862E";
    when 16#0092B# => romdata <= X"81B53881";
    when 16#0092C# => romdata <= X"165680FF";
    when 16#0092D# => romdata <= X"7627FEAD";
    when 16#0092E# => romdata <= X"388A3D0D";
    when 16#0092F# => romdata <= X"0481A694";
    when 16#00930# => romdata <= X"519BBB3F";
    when 16#00931# => romdata <= X"C016519C";
    when 16#00932# => romdata <= X"FF3F8652";
    when 16#00933# => romdata <= X"B00851CD";
    when 16#00934# => romdata <= X"8E3F81A5";
    when 16#00935# => romdata <= X"E4519BA6";
    when 16#00936# => romdata <= X"3F745288";
    when 16#00937# => romdata <= X"519BC23F";
    when 16#00938# => romdata <= X"8452B008";
    when 16#00939# => romdata <= X"51CCF83F";
    when 16#0093A# => romdata <= X"81A5EC51";
    when 16#0093B# => romdata <= X"9B903F76";
    when 16#0093C# => romdata <= X"5290519B";
    when 16#0093D# => romdata <= X"AC3F8652";
    when 16#0093E# => romdata <= X"B00851CC";
    when 16#0093F# => romdata <= X"E23F81A5";
    when 16#00940# => romdata <= X"F4519AFA";
    when 16#00941# => romdata <= X"3F72519C";
    when 16#00942# => romdata <= X"BF3F8452";
    when 16#00943# => romdata <= X"B00851CC";
    when 16#00944# => romdata <= X"CE3F81A5";
    when 16#00945# => romdata <= X"FC519AE6";
    when 16#00946# => romdata <= X"3F73519C";
    when 16#00947# => romdata <= X"AB3F8452";
    when 16#00948# => romdata <= X"B00851CC";
    when 16#00949# => romdata <= X"BA3F81A6";
    when 16#0094A# => romdata <= X"84519AD2";
    when 16#0094B# => romdata <= X"3F7708C0";
    when 16#0094C# => romdata <= X"80800652";
    when 16#0094D# => romdata <= X"A0519AE9";
    when 16#0094E# => romdata <= X"3F8A52B0";
    when 16#0094F# => romdata <= X"0851CC9F";
    when 16#00950# => romdata <= X"3F78802E";
    when 16#00951# => romdata <= X"FED63876";
    when 16#00952# => romdata <= X"81FF0652";
    when 16#00953# => romdata <= X"7451F8E8";
    when 16#00954# => romdata <= X"3F8A519A";
    when 16#00955# => romdata <= X"8F3F8053";
    when 16#00956# => romdata <= X"74812E09";
    when 16#00957# => romdata <= X"8106FEC9";
    when 16#00958# => romdata <= X"389F3972";
    when 16#00959# => romdata <= X"81065776";
    when 16#0095A# => romdata <= X"802EFEC3";
    when 16#0095B# => romdata <= X"38785277";
    when 16#0095C# => romdata <= X"51FAF03F";
    when 16#0095D# => romdata <= X"81165680";
    when 16#0095E# => romdata <= X"FF7627FC";
    when 16#0095F# => romdata <= X"E838FEB9";
    when 16#00960# => romdata <= X"39745376";
    when 16#00961# => romdata <= X"862E0981";
    when 16#00962# => romdata <= X"06FEA438";
    when 16#00963# => romdata <= X"D639803D";
    when 16#00964# => romdata <= X"0D81B294";
    when 16#00965# => romdata <= X"08519971";
    when 16#00966# => romdata <= X"0C81800B";
    when 16#00967# => romdata <= X"84120C81";
    when 16#00968# => romdata <= X"B2900851";
    when 16#00969# => romdata <= X"99710C81";
    when 16#0096A# => romdata <= X"800B8412";
    when 16#0096B# => romdata <= X"0C823D0D";
    when 16#0096C# => romdata <= X"04FE3D0D";
    when 16#0096D# => romdata <= X"74028405";
    when 16#0096E# => romdata <= X"97053302";
    when 16#0096F# => romdata <= X"88059B05";
    when 16#00970# => romdata <= X"3388130C";
    when 16#00971# => romdata <= X"8C120C53";
    when 16#00972# => romdata <= X"8C130870";
    when 16#00973# => romdata <= X"812A8106";
    when 16#00974# => romdata <= X"515271F4";
    when 16#00975# => romdata <= X"388C1308";
    when 16#00976# => romdata <= X"7081FF06";
    when 16#00977# => romdata <= X"B00C5184";
    when 16#00978# => romdata <= X"3D0D0480";
    when 16#00979# => romdata <= X"3D0D728C";
    when 16#0097A# => romdata <= X"11087087";
    when 16#0097B# => romdata <= X"2A813281";
    when 16#0097C# => romdata <= X"06B00C51";
    when 16#0097D# => romdata <= X"51823D0D";
    when 16#0097E# => romdata <= X"04FE3D0D";
    when 16#0097F# => romdata <= X"FF903F81";
    when 16#00980# => romdata <= X"EC538190";
    when 16#00981# => romdata <= X"5281B294";
    when 16#00982# => romdata <= X"0851FFA5";
    when 16#00983# => romdata <= X"3F9D5390";
    when 16#00984# => romdata <= X"5281B294";
    when 16#00985# => romdata <= X"0851FF99";
    when 16#00986# => romdata <= X"3F80C553";
    when 16#00987# => romdata <= X"80D05281";
    when 16#00988# => romdata <= X"B2940851";
    when 16#00989# => romdata <= X"FF8B3F81";
    when 16#0098A# => romdata <= X"EC538190";
    when 16#0098B# => romdata <= X"5281B294";
    when 16#0098C# => romdata <= X"0851FEFD";
    when 16#0098D# => romdata <= X"3FA15390";
    when 16#0098E# => romdata <= X"5281B294";
    when 16#0098F# => romdata <= X"0851FEF1";
    when 16#00990# => romdata <= X"3F895380";
    when 16#00991# => romdata <= X"D05281B2";
    when 16#00992# => romdata <= X"940851FE";
    when 16#00993# => romdata <= X"E43F81EC";
    when 16#00994# => romdata <= X"53819052";
    when 16#00995# => romdata <= X"81B29408";
    when 16#00996# => romdata <= X"51FED63F";
    when 16#00997# => romdata <= X"B3539052";
    when 16#00998# => romdata <= X"81B29408";
    when 16#00999# => romdata <= X"51FECA3F";
    when 16#0099A# => romdata <= X"885380D0";
    when 16#0099B# => romdata <= X"5281B294";
    when 16#0099C# => romdata <= X"0851FEBD";
    when 16#0099D# => romdata <= X"3F81EC53";
    when 16#0099E# => romdata <= X"81905281";
    when 16#0099F# => romdata <= X"B2940851";
    when 16#009A0# => romdata <= X"FEAF3FB4";
    when 16#009A1# => romdata <= X"53905281";
    when 16#009A2# => romdata <= X"B2940851";
    when 16#009A3# => romdata <= X"FEA33F96";
    when 16#009A4# => romdata <= X"5380D052";
    when 16#009A5# => romdata <= X"81B29408";
    when 16#009A6# => romdata <= X"51FE963F";
    when 16#009A7# => romdata <= X"81EC5381";
    when 16#009A8# => romdata <= X"905281B2";
    when 16#009A9# => romdata <= X"940851FE";
    when 16#009AA# => romdata <= X"883FB653";
    when 16#009AB# => romdata <= X"905281B2";
    when 16#009AC# => romdata <= X"940851FD";
    when 16#009AD# => romdata <= X"FC3F80E0";
    when 16#009AE# => romdata <= X"5380D052";
    when 16#009AF# => romdata <= X"81B29408";
    when 16#009B0# => romdata <= X"51FDEE3F";
    when 16#009B1# => romdata <= X"81EC5381";
    when 16#009B2# => romdata <= X"905281B2";
    when 16#009B3# => romdata <= X"940851FD";
    when 16#009B4# => romdata <= X"E03F80C9";
    when 16#009B5# => romdata <= X"53905281";
    when 16#009B6# => romdata <= X"B2940851";
    when 16#009B7# => romdata <= X"FDD33F81";
    when 16#009B8# => romdata <= X"C05380D0";
    when 16#009B9# => romdata <= X"5281B294";
    when 16#009BA# => romdata <= X"0851FDC5";
    when 16#009BB# => romdata <= X"3F843D0D";
    when 16#009BC# => romdata <= X"04FD3D0D";
    when 16#009BD# => romdata <= X"02970533";
    when 16#009BE# => romdata <= X"0284059B";
    when 16#009BF# => romdata <= X"05337181";
    when 16#009C0# => romdata <= X"B00781BF";
    when 16#009C1# => romdata <= X"06535454";
    when 16#009C2# => romdata <= X"F8808098";
    when 16#009C3# => romdata <= X"8071710C";
    when 16#009C4# => romdata <= X"73842A90";
    when 16#009C5# => romdata <= X"07710C73";
    when 16#009C6# => romdata <= X"8F06710C";
    when 16#009C7# => romdata <= X"527281B1";
    when 16#009C8# => romdata <= X"F0347381";
    when 16#009C9# => romdata <= X"B1F43485";
    when 16#009CA# => romdata <= X"3D0D04FD";
    when 16#009CB# => romdata <= X"3D0D0297";
    when 16#009CC# => romdata <= X"053381B1";
    when 16#009CD# => romdata <= X"F4335473";
    when 16#009CE# => romdata <= X"05870602";
    when 16#009CF# => romdata <= X"84059A05";
    when 16#009D0# => romdata <= X"2281B1F0";
    when 16#009D1# => romdata <= X"33547305";
    when 16#009D2# => romdata <= X"7081FF06";
    when 16#009D3# => romdata <= X"7281B007";
    when 16#009D4# => romdata <= X"54515454";
    when 16#009D5# => romdata <= X"F8808098";
    when 16#009D6# => romdata <= X"8071710C";
    when 16#009D7# => romdata <= X"73842A90";
    when 16#009D8# => romdata <= X"07710C73";
    when 16#009D9# => romdata <= X"8F06710C";
    when 16#009DA# => romdata <= X"527281B1";
    when 16#009DB# => romdata <= X"F0347381";
    when 16#009DC# => romdata <= X"B1F43485";
    when 16#009DD# => romdata <= X"3D0D04FF";
    when 16#009DE# => romdata <= X"3D0D028F";
    when 16#009DF# => romdata <= X"0533F880";
    when 16#009E0# => romdata <= X"8098840C";
    when 16#009E1# => romdata <= X"81B1F033";
    when 16#009E2# => romdata <= X"81055170";
    when 16#009E3# => romdata <= X"81B1F034";
    when 16#009E4# => romdata <= X"833D0D04";
    when 16#009E5# => romdata <= X"FF3D0D80";
    when 16#009E6# => romdata <= X"C00BF880";
    when 16#009E7# => romdata <= X"8098800C";
    when 16#009E8# => romdata <= X"81A10BF8";
    when 16#009E9# => romdata <= X"80809880";
    when 16#009EA# => romdata <= X"0C81C00B";
    when 16#009EB# => romdata <= X"F8808098";
    when 16#009EC# => romdata <= X"800C81A4";
    when 16#009ED# => romdata <= X"0BF88080";
    when 16#009EE# => romdata <= X"98800C81";
    when 16#009EF# => romdata <= X"A60BF880";
    when 16#009F0# => romdata <= X"8098800C";
    when 16#009F1# => romdata <= X"81A20BF8";
    when 16#009F2# => romdata <= X"80809880";
    when 16#009F3# => romdata <= X"0CAF0BF8";
    when 16#009F4# => romdata <= X"80809880";
    when 16#009F5# => romdata <= X"0CA50BF8";
    when 16#009F6# => romdata <= X"80809880";
    when 16#009F7# => romdata <= X"0C81810B";
    when 16#009F8# => romdata <= X"F8808098";
    when 16#009F9# => romdata <= X"800C9D0B";
    when 16#009FA# => romdata <= X"F8808098";
    when 16#009FB# => romdata <= X"800C81FA";
    when 16#009FC# => romdata <= X"0BF88080";
    when 16#009FD# => romdata <= X"98800C80";
    when 16#009FE# => romdata <= X"0BF88080";
    when 16#009FF# => romdata <= X"98800C80";
    when 16#00A00# => romdata <= X"527181B0";
    when 16#00A01# => romdata <= X"0781BF06";
    when 16#00A02# => romdata <= X"F8808098";
    when 16#00A03# => romdata <= X"800C900B";
    when 16#00A04# => romdata <= X"F8808098";
    when 16#00A05# => romdata <= X"800C800B";
    when 16#00A06# => romdata <= X"F8808098";
    when 16#00A07# => romdata <= X"800C8051";
    when 16#00A08# => romdata <= X"800BF880";
    when 16#00A09# => romdata <= X"8098840C";
    when 16#00A0A# => romdata <= X"81117081";
    when 16#00A0B# => romdata <= X"FF065151";
    when 16#00A0C# => romdata <= X"80E57127";
    when 16#00A0D# => romdata <= X"EB388112";
    when 16#00A0E# => romdata <= X"7081FF06";
    when 16#00A0F# => romdata <= X"53518772";
    when 16#00A10# => romdata <= X"27FFBE38";
    when 16#00A11# => romdata <= X"81B00BF8";
    when 16#00A12# => romdata <= X"80809880";
    when 16#00A13# => romdata <= X"0C900BF8";
    when 16#00A14# => romdata <= X"80809880";
    when 16#00A15# => romdata <= X"0C800BF8";
    when 16#00A16# => romdata <= X"80809880";
    when 16#00A17# => romdata <= X"0C800B81";
    when 16#00A18# => romdata <= X"B1F03480";
    when 16#00A19# => romdata <= X"0B81B1F4";
    when 16#00A1A# => romdata <= X"3481AF0B";
    when 16#00A1B# => romdata <= X"F8808098";
    when 16#00A1C# => romdata <= X"800C833D";
    when 16#00A1D# => romdata <= X"0D04ED3D";
    when 16#00A1E# => romdata <= X"0D650284";
    when 16#00A1F# => romdata <= X"0580DB05";
    when 16#00A20# => romdata <= X"33028805";
    when 16#00A21# => romdata <= X"80DF0533";
    when 16#00A22# => romdata <= X"5F5A5680";
    when 16#00A23# => romdata <= X"7981067A";
    when 16#00A24# => romdata <= X"812A8106";
    when 16#00A25# => romdata <= X"7B832B81";
    when 16#00A26# => romdata <= X"80067C82";
    when 16#00A27# => romdata <= X"2A810657";
    when 16#00A28# => romdata <= X"5E435F5C";
    when 16#00A29# => romdata <= X"81FF4272";
    when 16#00A2A# => romdata <= X"7C2E0981";
    when 16#00A2B# => romdata <= X"0683387B";
    when 16#00A2C# => romdata <= X"42881608";
    when 16#00A2D# => romdata <= X"5574802E";
    when 16#00A2E# => romdata <= X"839F3885";
    when 16#00A2F# => romdata <= X"16335AFF";
    when 16#00A30# => romdata <= X"537C7A26";
    when 16#00A31# => romdata <= X"8E388416";
    when 16#00A32# => romdata <= X"3354737D";
    when 16#00A33# => romdata <= X"2685387C";
    when 16#00A34# => romdata <= X"74315374";
    when 16#00A35# => romdata <= X"13703354";
    when 16#00A36# => romdata <= X"577281FF";
    when 16#00A37# => romdata <= X"06831733";
    when 16#00A38# => romdata <= X"70982B81";
    when 16#00A39# => romdata <= X"FF0A119B";
    when 16#00A3A# => romdata <= X"2A810551";
    when 16#00A3B# => romdata <= X"5A404081";
    when 16#00A3C# => romdata <= X"53748338";
    when 16#00A3D# => romdata <= X"74537281";
    when 16#00A3E# => romdata <= X"FF064380";
    when 16#00A3F# => romdata <= X"7A81FF06";
    when 16#00A40# => romdata <= X"4557FF54";
    when 16#00A41# => romdata <= X"7C64268B";
    when 16#00A42# => romdata <= X"38841633";
    when 16#00A43# => romdata <= X"537C7327";
    when 16#00A44# => romdata <= X"83CE3873";
    when 16#00A45# => romdata <= X"7481FF06";
    when 16#00A46# => romdata <= X"5553805A";
    when 16#00A47# => romdata <= X"797324AB";
    when 16#00A48# => romdata <= X"38747A2E";
    when 16#00A49# => romdata <= X"09810682";
    when 16#00A4A# => romdata <= X"BB387E98";
    when 16#00A4B# => romdata <= X"2B81FF0A";
    when 16#00A4C# => romdata <= X"119B2A82";
    when 16#00A4D# => romdata <= X"18337171";
    when 16#00A4E# => romdata <= X"29117081";
    when 16#00A4F# => romdata <= X"FF067871";
    when 16#00A50# => romdata <= X"298C1C08";
    when 16#00A51# => romdata <= X"0552435D";
    when 16#00A52# => romdata <= X"5758447F";
    when 16#00A53# => romdata <= X"63057081";
    when 16#00A54# => romdata <= X"FF067063";
    when 16#00A55# => romdata <= X"2B7081FF";
    when 16#00A56# => romdata <= X"067B622B";
    when 16#00A57# => romdata <= X"7081FF06";
    when 16#00A58# => romdata <= X"7E832A81";
    when 16#00A59# => romdata <= X"065C5557";
    when 16#00A5A# => romdata <= X"5256455F";
    when 16#00A5B# => romdata <= X"75802E8F";
    when 16#00A5C# => romdata <= X"3881B1F0";
    when 16#00A5D# => romdata <= X"33640559";
    when 16#00A5E# => romdata <= X"7880E624";
    when 16#00A5F# => romdata <= X"8DC6387F";
    when 16#00A60# => romdata <= X"78296430";
    when 16#00A61# => romdata <= X"5E577B7E";
    when 16#00A62# => romdata <= X"2C982B70";
    when 16#00A63# => romdata <= X"982C5540";
    when 16#00A64# => romdata <= X"73772580";
    when 16#00A65# => romdata <= X"FC38FF1F";
    when 16#00A66# => romdata <= X"7C81065A";
    when 16#00A67# => romdata <= X"537B732E";
    when 16#00A68# => romdata <= X"83843860";
    when 16#00A69# => romdata <= X"85DA3861";
    when 16#00A6A# => romdata <= X"84A5387D";
    when 16#00A6B# => romdata <= X"802E81FE";
    when 16#00A6C# => romdata <= X"38791470";
    when 16#00A6D# => romdata <= X"33705254";
    when 16#00A6E# => romdata <= X"56805578";
    when 16#00A6F# => romdata <= X"752E8538";
    when 16#00A70# => romdata <= X"72842A56";
    when 16#00A71# => romdata <= X"75832A81";
    when 16#00A72# => romdata <= X"06407F80";
    when 16#00A73# => romdata <= X"2E843881";
    when 16#00A74# => romdata <= X"C0557582";
    when 16#00A75# => romdata <= X"2A810640";
    when 16#00A76# => romdata <= X"7F802E85";
    when 16#00A77# => romdata <= X"3874B007";
    when 16#00A78# => romdata <= X"5575812A";
    when 16#00A79# => romdata <= X"8106407F";
    when 16#00A7A# => romdata <= X"802E8538";
    when 16#00A7B# => romdata <= X"748C0755";
    when 16#00A7C# => romdata <= X"75810653";
    when 16#00A7D# => romdata <= X"72802E85";
    when 16#00A7E# => romdata <= X"38748307";
    when 16#00A7F# => romdata <= X"557451FA";
    when 16#00A80# => romdata <= X"F63F7714";
    when 16#00A81# => romdata <= X"982B7098";
    when 16#00A82# => romdata <= X"2C555576";
    when 16#00A83# => romdata <= X"7424FFA1";
    when 16#00A84# => romdata <= X"3862802E";
    when 16#00A85# => romdata <= X"9638617F";
    when 16#00A86# => romdata <= X"FF055654";
    when 16#00A87# => romdata <= X"7B752E81";
    when 16#00A88# => romdata <= X"E3387351";
    when 16#00A89# => romdata <= X"FAD13F60";
    when 16#00A8A# => romdata <= X"81BD387C";
    when 16#00A8B# => romdata <= X"528151F9";
    when 16#00A8C# => romdata <= X"FA3F811C";
    when 16#00A8D# => romdata <= X"7081FF06";
    when 16#00A8E# => romdata <= X"5D547E7C";
    when 16#00A8F# => romdata <= X"26FEC738";
    when 16#00A90# => romdata <= X"63527E30";
    when 16#00A91# => romdata <= X"70982B70";
    when 16#00A92# => romdata <= X"982C535C";
    when 16#00A93# => romdata <= X"5CF9DC3F";
    when 16#00A94# => romdata <= X"635372B0";
    when 16#00A95# => romdata <= X"0C953D0D";
    when 16#00A96# => romdata <= X"04821633";
    when 16#00A97# => romdata <= X"8517335B";
    when 16#00A98# => romdata <= X"53FCF639";
    when 16#00A99# => romdata <= X"73802EAF";
    when 16#00A9A# => romdata <= X"38FF1470";
    when 16#00A9B# => romdata <= X"81FF0655";
    when 16#00A9C# => romdata <= X"537381FF";
    when 16#00A9D# => romdata <= X"2EA13874";
    when 16#00A9E# => romdata <= X"70810556";
    when 16#00A9F# => romdata <= X"33770570";
    when 16#00AA0# => romdata <= X"83FFFF06";
    when 16#00AA1# => romdata <= X"FF167081";
    when 16#00AA2# => romdata <= X"FF065755";
    when 16#00AA3# => romdata <= X"585A7381";
    when 16#00AA4# => romdata <= X"FF2E0981";
    when 16#00AA5# => romdata <= X"06E1387E";
    when 16#00AA6# => romdata <= X"982B81FF";
    when 16#00AA7# => romdata <= X"0A119B2A";
    when 16#00AA8# => romdata <= X"70792919";
    when 16#00AA9# => romdata <= X"8C190805";
    when 16#00AAA# => romdata <= X"5C4055FD";
    when 16#00AAB# => romdata <= X"9E397914";
    when 16#00AAC# => romdata <= X"70335259";
    when 16#00AAD# => romdata <= X"F9C13F77";
    when 16#00AAE# => romdata <= X"14982B70";
    when 16#00AAF# => romdata <= X"982C5553";
    when 16#00AB0# => romdata <= X"737725FE";
    when 16#00AB1# => romdata <= X"CC387914";
    when 16#00AB2# => romdata <= X"70335259";
    when 16#00AB3# => romdata <= X"F9A93F77";
    when 16#00AB4# => romdata <= X"14982B70";
    when 16#00AB5# => romdata <= X"982C5553";
    when 16#00AB6# => romdata <= X"767424D2";
    when 16#00AB7# => romdata <= X"38FEB239";
    when 16#00AB8# => romdata <= X"7C733154";
    when 16#00AB9# => romdata <= X"FCAD3973";
    when 16#00ABA# => romdata <= X"51F98C3F";
    when 16#00ABB# => romdata <= X"7C528151";
    when 16#00ABC# => romdata <= X"F8B93F81";
    when 16#00ABD# => romdata <= X"1C7081FF";
    when 16#00ABE# => romdata <= X"065D547E";
    when 16#00ABF# => romdata <= X"7C26FD86";
    when 16#00AC0# => romdata <= X"38FEBD39";
    when 16#00AC1# => romdata <= X"617B3270";
    when 16#00AC2# => romdata <= X"81FF0655";
    when 16#00AC3# => romdata <= X"567D802E";
    when 16#00AC4# => romdata <= X"FE90387A";
    when 16#00AC5# => romdata <= X"812A7432";
    when 16#00AC6# => romdata <= X"705254F8";
    when 16#00AC7# => romdata <= X"DA3F6080";
    when 16#00AC8# => romdata <= X"2EFE8838";
    when 16#00AC9# => romdata <= X"C2396087";
    when 16#00ACA# => romdata <= X"8F386185";
    when 16#00ACB# => romdata <= X"D3387D80";
    when 16#00ACC# => romdata <= X"2E80E638";
    when 16#00ACD# => romdata <= X"79147033";
    when 16#00ACE# => romdata <= X"7C077052";
    when 16#00ACF# => romdata <= X"54568055";
    when 16#00AD0# => romdata <= X"78752E85";
    when 16#00AD1# => romdata <= X"3872842A";
    when 16#00AD2# => romdata <= X"5675832A";
    when 16#00AD3# => romdata <= X"81065372";
    when 16#00AD4# => romdata <= X"802E8438";
    when 16#00AD5# => romdata <= X"81C05575";
    when 16#00AD6# => romdata <= X"822A8106";
    when 16#00AD7# => romdata <= X"5372802E";
    when 16#00AD8# => romdata <= X"853874B0";
    when 16#00AD9# => romdata <= X"07557581";
    when 16#00ADA# => romdata <= X"2A810653";
    when 16#00ADB# => romdata <= X"72802E85";
    when 16#00ADC# => romdata <= X"38748C07";
    when 16#00ADD# => romdata <= X"55758106";
    when 16#00ADE# => romdata <= X"407F802E";
    when 16#00ADF# => romdata <= X"85387483";
    when 16#00AE0# => romdata <= X"07557451";
    when 16#00AE1# => romdata <= X"F7F13F77";
    when 16#00AE2# => romdata <= X"14982B70";
    when 16#00AE3# => romdata <= X"982C5553";
    when 16#00AE4# => romdata <= X"767424FF";
    when 16#00AE5# => romdata <= X"9F38FCF9";
    when 16#00AE6# => romdata <= X"39791470";
    when 16#00AE7# => romdata <= X"337C0752";
    when 16#00AE8# => romdata <= X"55F7D43F";
    when 16#00AE9# => romdata <= X"7714982B";
    when 16#00AEA# => romdata <= X"70982C55";
    when 16#00AEB# => romdata <= X"59737725";
    when 16#00AEC# => romdata <= X"FCDF3879";
    when 16#00AED# => romdata <= X"1470337C";
    when 16#00AEE# => romdata <= X"075255F7";
    when 16#00AEF# => romdata <= X"BA3F7714";
    when 16#00AF0# => romdata <= X"982B7098";
    when 16#00AF1# => romdata <= X"2C555976";
    when 16#00AF2# => romdata <= X"7424CE38";
    when 16#00AF3# => romdata <= X"FCC3397D";
    when 16#00AF4# => romdata <= X"802E80EA";
    when 16#00AF5# => romdata <= X"38791470";
    when 16#00AF6# => romdata <= X"33705854";
    when 16#00AF7# => romdata <= X"55805578";
    when 16#00AF8# => romdata <= X"752E8538";
    when 16#00AF9# => romdata <= X"72842A56";
    when 16#00AFA# => romdata <= X"75832A81";
    when 16#00AFB# => romdata <= X"06537280";
    when 16#00AFC# => romdata <= X"2E843881";
    when 16#00AFD# => romdata <= X"C0557582";
    when 16#00AFE# => romdata <= X"2A810653";
    when 16#00AFF# => romdata <= X"72802E85";
    when 16#00B00# => romdata <= X"3874B007";
    when 16#00B01# => romdata <= X"5575812A";
    when 16#00B02# => romdata <= X"81065372";
    when 16#00B03# => romdata <= X"802E8538";
    when 16#00B04# => romdata <= X"748C0755";
    when 16#00B05# => romdata <= X"75810640";
    when 16#00B06# => romdata <= X"7F802E85";
    when 16#00B07# => romdata <= X"38748307";
    when 16#00B08# => romdata <= X"55740970";
    when 16#00B09# => romdata <= X"81FF0652";
    when 16#00B0A# => romdata <= X"53F6CC3F";
    when 16#00B0B# => romdata <= X"7714982B";
    when 16#00B0C# => romdata <= X"70982C55";
    when 16#00B0D# => romdata <= X"56767424";
    when 16#00B0E# => romdata <= X"FF9B38FB";
    when 16#00B0F# => romdata <= X"D4397914";
    when 16#00B10# => romdata <= X"70337009";
    when 16#00B11# => romdata <= X"7081FF06";
    when 16#00B12# => romdata <= X"54585440";
    when 16#00B13# => romdata <= X"F6A93F77";
    when 16#00B14# => romdata <= X"14982B70";
    when 16#00B15# => romdata <= X"982C5559";
    when 16#00B16# => romdata <= X"737725FB";
    when 16#00B17# => romdata <= X"B4387914";
    when 16#00B18# => romdata <= X"70337009";
    when 16#00B19# => romdata <= X"7081FF06";
    when 16#00B1A# => romdata <= X"54585440";
    when 16#00B1B# => romdata <= X"F6893F77";
    when 16#00B1C# => romdata <= X"14982B70";
    when 16#00B1D# => romdata <= X"982C5559";
    when 16#00B1E# => romdata <= X"767424C2";
    when 16#00B1F# => romdata <= X"38FB9239";
    when 16#00B20# => romdata <= X"61802E81";
    when 16#00B21# => romdata <= X"C8387D80";
    when 16#00B22# => romdata <= X"2E80F138";
    when 16#00B23# => romdata <= X"79147033";
    when 16#00B24# => romdata <= X"70585455";
    when 16#00B25# => romdata <= X"80557875";
    when 16#00B26# => romdata <= X"2E853872";
    when 16#00B27# => romdata <= X"842A5675";
    when 16#00B28# => romdata <= X"832A8106";
    when 16#00B29# => romdata <= X"407F802E";
    when 16#00B2A# => romdata <= X"843881C0";
    when 16#00B2B# => romdata <= X"5575822A";
    when 16#00B2C# => romdata <= X"8106407F";
    when 16#00B2D# => romdata <= X"802E8538";
    when 16#00B2E# => romdata <= X"74B00755";
    when 16#00B2F# => romdata <= X"75812A81";
    when 16#00B30# => romdata <= X"06407F80";
    when 16#00B31# => romdata <= X"2E853874";
    when 16#00B32# => romdata <= X"8C075575";
    when 16#00B33# => romdata <= X"81065372";
    when 16#00B34# => romdata <= X"802E8538";
    when 16#00B35# => romdata <= X"74830755";
    when 16#00B36# => romdata <= X"74097081";
    when 16#00B37# => romdata <= X"FF067053";
    when 16#00B38# => romdata <= X"4156F593";
    when 16#00B39# => romdata <= X"3F7F51F5";
    when 16#00B3A# => romdata <= X"8E3F7714";
    when 16#00B3B# => romdata <= X"982B7098";
    when 16#00B3C# => romdata <= X"2C555376";
    when 16#00B3D# => romdata <= X"7424FF94";
    when 16#00B3E# => romdata <= X"38FA9639";
    when 16#00B3F# => romdata <= X"79147033";
    when 16#00B40# => romdata <= X"70097081";
    when 16#00B41# => romdata <= X"FF067055";
    when 16#00B42# => romdata <= X"59554155";
    when 16#00B43# => romdata <= X"F4E93F75";
    when 16#00B44# => romdata <= X"51F4E43F";
    when 16#00B45# => romdata <= X"7714982B";
    when 16#00B46# => romdata <= X"70982C55";
    when 16#00B47# => romdata <= X"59737725";
    when 16#00B48# => romdata <= X"F9EF3879";
    when 16#00B49# => romdata <= X"14703370";
    when 16#00B4A# => romdata <= X"097081FF";
    when 16#00B4B# => romdata <= X"06705559";
    when 16#00B4C# => romdata <= X"554155F4";
    when 16#00B4D# => romdata <= X"C23F7551";
    when 16#00B4E# => romdata <= X"F4BD3F77";
    when 16#00B4F# => romdata <= X"14982B70";
    when 16#00B50# => romdata <= X"982C5559";
    when 16#00B51# => romdata <= X"767424FF";
    when 16#00B52# => romdata <= X"B338F9C5";
    when 16#00B53# => romdata <= X"397D802E";
    when 16#00B54# => romdata <= X"80EE3879";
    when 16#00B55# => romdata <= X"14703370";
    when 16#00B56# => romdata <= X"58545580";
    when 16#00B57# => romdata <= X"5578752E";
    when 16#00B58# => romdata <= X"85387284";
    when 16#00B59# => romdata <= X"2A567583";
    when 16#00B5A# => romdata <= X"2A810653";
    when 16#00B5B# => romdata <= X"72802E84";
    when 16#00B5C# => romdata <= X"3881C055";
    when 16#00B5D# => romdata <= X"75822A81";
    when 16#00B5E# => romdata <= X"06537280";
    when 16#00B5F# => romdata <= X"2E853874";
    when 16#00B60# => romdata <= X"B0075575";
    when 16#00B61# => romdata <= X"812A8106";
    when 16#00B62# => romdata <= X"5372802E";
    when 16#00B63# => romdata <= X"8538748C";
    when 16#00B64# => romdata <= X"07557581";
    when 16#00B65# => romdata <= X"06407F80";
    when 16#00B66# => romdata <= X"2E853874";
    when 16#00B67# => romdata <= X"83075574";
    when 16#00B68# => romdata <= X"81FF0670";
    when 16#00B69# => romdata <= X"5256F3CF";
    when 16#00B6A# => romdata <= X"3F7551F3";
    when 16#00B6B# => romdata <= X"CA3F7714";
    when 16#00B6C# => romdata <= X"982B7098";
    when 16#00B6D# => romdata <= X"2C555376";
    when 16#00B6E# => romdata <= X"7424FF97";
    when 16#00B6F# => romdata <= X"38F8D239";
    when 16#00B70# => romdata <= X"79147033";
    when 16#00B71# => romdata <= X"70535740";
    when 16#00B72# => romdata <= X"F3AD3F75";
    when 16#00B73# => romdata <= X"51F3A83F";
    when 16#00B74# => romdata <= X"7714982B";
    when 16#00B75# => romdata <= X"70982C55";
    when 16#00B76# => romdata <= X"59737725";
    when 16#00B77# => romdata <= X"F8B33879";
    when 16#00B78# => romdata <= X"14703370";
    when 16#00B79# => romdata <= X"535740F3";
    when 16#00B7A# => romdata <= X"8E3F7551";
    when 16#00B7B# => romdata <= X"F3893F77";
    when 16#00B7C# => romdata <= X"14982B70";
    when 16#00B7D# => romdata <= X"982C5559";
    when 16#00B7E# => romdata <= X"767424C4";
    when 16#00B7F# => romdata <= X"38F89239";
    when 16#00B80# => romdata <= X"7D802E80";
    when 16#00B81# => romdata <= X"EC387914";
    when 16#00B82# => romdata <= X"70337C07";
    when 16#00B83# => romdata <= X"70525456";
    when 16#00B84# => romdata <= X"80557875";
    when 16#00B85# => romdata <= X"2E853872";
    when 16#00B86# => romdata <= X"842A5675";
    when 16#00B87# => romdata <= X"832A8106";
    when 16#00B88# => romdata <= X"5372802E";
    when 16#00B89# => romdata <= X"843881C0";
    when 16#00B8A# => romdata <= X"5575822A";
    when 16#00B8B# => romdata <= X"81065372";
    when 16#00B8C# => romdata <= X"802E8538";
    when 16#00B8D# => romdata <= X"74B00755";
    when 16#00B8E# => romdata <= X"75812A81";
    when 16#00B8F# => romdata <= X"06537280";
    when 16#00B90# => romdata <= X"2E853874";
    when 16#00B91# => romdata <= X"8C075575";
    when 16#00B92# => romdata <= X"8106407F";
    when 16#00B93# => romdata <= X"802E8538";
    when 16#00B94# => romdata <= X"74830755";
    when 16#00B95# => romdata <= X"74097081";
    when 16#00B96# => romdata <= X"FF065253";
    when 16#00B97# => romdata <= X"F2993F77";
    when 16#00B98# => romdata <= X"14982B70";
    when 16#00B99# => romdata <= X"982C5556";
    when 16#00B9A# => romdata <= X"767424FF";
    when 16#00B9B# => romdata <= X"9938F7A1";
    when 16#00B9C# => romdata <= X"39791470";
    when 16#00B9D# => romdata <= X"337C0770";
    when 16#00B9E# => romdata <= X"097081FF";
    when 16#00B9F# => romdata <= X"06545541";
    when 16#00BA0# => romdata <= X"56F1F43F";
    when 16#00BA1# => romdata <= X"7714982B";
    when 16#00BA2# => romdata <= X"70982C55";
    when 16#00BA3# => romdata <= X"59737725";
    when 16#00BA4# => romdata <= X"F6FF3879";
    when 16#00BA5# => romdata <= X"1470337C";
    when 16#00BA6# => romdata <= X"07700970";
    when 16#00BA7# => romdata <= X"81FF0654";
    when 16#00BA8# => romdata <= X"554156F1";
    when 16#00BA9# => romdata <= X"D23F7714";
    when 16#00BAA# => romdata <= X"982B7098";
    when 16#00BAB# => romdata <= X"2C555976";
    when 16#00BAC# => romdata <= X"7424FFBD";
    when 16#00BAD# => romdata <= X"38F6DA39";
    when 16#00BAE# => romdata <= X"61802E80";
    when 16#00BAF# => romdata <= X"F9387D80";
    when 16#00BB0# => romdata <= X"2E81E838";
    when 16#00BB1# => romdata <= X"79147033";
    when 16#00BB2# => romdata <= X"7C077052";
    when 16#00BB3# => romdata <= X"54568055";
    when 16#00BB4# => romdata <= X"78752E85";
    when 16#00BB5# => romdata <= X"3872842A";
    when 16#00BB6# => romdata <= X"5675832A";
    when 16#00BB7# => romdata <= X"81065372";
    when 16#00BB8# => romdata <= X"802E8438";
    when 16#00BB9# => romdata <= X"81C05575";
    when 16#00BBA# => romdata <= X"822A8106";
    when 16#00BBB# => romdata <= X"5372802E";
    when 16#00BBC# => romdata <= X"853874B0";
    when 16#00BBD# => romdata <= X"07557581";
    when 16#00BBE# => romdata <= X"2A810653";
    when 16#00BBF# => romdata <= X"72802E85";
    when 16#00BC0# => romdata <= X"38748C07";
    when 16#00BC1# => romdata <= X"55758106";
    when 16#00BC2# => romdata <= X"407F802E";
    when 16#00BC3# => romdata <= X"85387483";
    when 16#00BC4# => romdata <= X"07557409";
    when 16#00BC5# => romdata <= X"7081FF06";
    when 16#00BC6# => romdata <= X"70535456";
    when 16#00BC7# => romdata <= X"F0D93F72";
    when 16#00BC8# => romdata <= X"51F0D43F";
    when 16#00BC9# => romdata <= X"7714982B";
    when 16#00BCA# => romdata <= X"70982C55";
    when 16#00BCB# => romdata <= X"40767424";
    when 16#00BCC# => romdata <= X"FF9238F5";
    when 16#00BCD# => romdata <= X"DC397D80";
    when 16#00BCE# => romdata <= X"2E81C538";
    when 16#00BCF# => romdata <= X"79147033";
    when 16#00BD0# => romdata <= X"7C077052";
    when 16#00BD1# => romdata <= X"54568055";
    when 16#00BD2# => romdata <= X"78752E85";
    when 16#00BD3# => romdata <= X"3872842A";
    when 16#00BD4# => romdata <= X"5675832A";
    when 16#00BD5# => romdata <= X"81065372";
    when 16#00BD6# => romdata <= X"802E8438";
    when 16#00BD7# => romdata <= X"81C05575";
    when 16#00BD8# => romdata <= X"822A8106";
    when 16#00BD9# => romdata <= X"5372802E";
    when 16#00BDA# => romdata <= X"853874B0";
    when 16#00BDB# => romdata <= X"07557581";
    when 16#00BDC# => romdata <= X"2A810653";
    when 16#00BDD# => romdata <= X"72802E85";
    when 16#00BDE# => romdata <= X"38748C07";
    when 16#00BDF# => romdata <= X"55758106";
    when 16#00BE0# => romdata <= X"407F802E";
    when 16#00BE1# => romdata <= X"85387483";
    when 16#00BE2# => romdata <= X"07557481";
    when 16#00BE3# => romdata <= X"FF067052";
    when 16#00BE4# => romdata <= X"53EFE43F";
    when 16#00BE5# => romdata <= X"7251EFDF";
    when 16#00BE6# => romdata <= X"3F771498";
    when 16#00BE7# => romdata <= X"2B70982C";
    when 16#00BE8# => romdata <= X"55567674";
    when 16#00BE9# => romdata <= X"24FF9538";
    when 16#00BEA# => romdata <= X"F4E73979";
    when 16#00BEB# => romdata <= X"1470337C";
    when 16#00BEC# => romdata <= X"07700970";
    when 16#00BED# => romdata <= X"81FF0670";
    when 16#00BEE# => romdata <= X"55564256";
    when 16#00BEF# => romdata <= X"59EFB83F";
    when 16#00BF0# => romdata <= X"7251EFB3";
    when 16#00BF1# => romdata <= X"3F771498";
    when 16#00BF2# => romdata <= X"2B70982C";
    when 16#00BF3# => romdata <= X"55597377";
    when 16#00BF4# => romdata <= X"25F4BE38";
    when 16#00BF5# => romdata <= X"79147033";
    when 16#00BF6# => romdata <= X"7C077009";
    when 16#00BF7# => romdata <= X"7081FF06";
    when 16#00BF8# => romdata <= X"70555642";
    when 16#00BF9# => romdata <= X"5659EF8F";
    when 16#00BFA# => romdata <= X"3F7251EF";
    when 16#00BFB# => romdata <= X"8A3F7714";
    when 16#00BFC# => romdata <= X"982B7098";
    when 16#00BFD# => romdata <= X"2C555976";
    when 16#00BFE# => romdata <= X"7424FFAF";
    when 16#00BFF# => romdata <= X"38F49239";
    when 16#00C00# => romdata <= X"79147033";
    when 16#00C01# => romdata <= X"7C077053";
    when 16#00C02# => romdata <= X"5455EEEB";
    when 16#00C03# => romdata <= X"3F7251EE";
    when 16#00C04# => romdata <= X"E63F7714";
    when 16#00C05# => romdata <= X"982B7098";
    when 16#00C06# => romdata <= X"2C555973";
    when 16#00C07# => romdata <= X"7725F3F1";
    when 16#00C08# => romdata <= X"38791470";
    when 16#00C09# => romdata <= X"337C0770";
    when 16#00C0A# => romdata <= X"535455EE";
    when 16#00C0B# => romdata <= X"CA3F7251";
    when 16#00C0C# => romdata <= X"EEC53F77";
    when 16#00C0D# => romdata <= X"14982B70";
    when 16#00C0E# => romdata <= X"982C5559";
    when 16#00C0F# => romdata <= X"767424C0";
    when 16#00C10# => romdata <= X"38F3CE39";
    when 16#00C11# => romdata <= X"81B1F433";
    when 16#00C12# => romdata <= X"7F055680";
    when 16#00C13# => romdata <= X"527581FF";
    when 16#00C14# => romdata <= X"0651ED9D";
    when 16#00C15# => romdata <= X"3F80537C";
    when 16#00C16# => romdata <= X"A02EF3F6";
    when 16#00C17# => romdata <= X"387F7829";
    when 16#00C18# => romdata <= X"64305E57";
    when 16#00C19# => romdata <= X"F2A039F8";
    when 16#00C1A# => romdata <= X"3D0D7A7D";
    when 16#00C1B# => romdata <= X"028805AF";
    when 16#00C1C# => romdata <= X"05335A55";
    when 16#00C1D# => romdata <= X"59807470";
    when 16#00C1E# => romdata <= X"81055633";
    when 16#00C1F# => romdata <= X"75585657";
    when 16#00C20# => romdata <= X"74772E09";
    when 16#00C21# => romdata <= X"81068838";
    when 16#00C22# => romdata <= X"76B00C8A";
    when 16#00C23# => romdata <= X"3D0D0474";
    when 16#00C24# => romdata <= X"53775278";
    when 16#00C25# => romdata <= X"51EFDF3F";
    when 16#00C26# => romdata <= X"B00881FF";
    when 16#00C27# => romdata <= X"06770570";
    when 16#00C28# => romdata <= X"83FFFF06";
    when 16#00C29# => romdata <= X"77708105";
    when 16#00C2A# => romdata <= X"59335258";
    when 16#00C2B# => romdata <= X"5574802E";
    when 16#00C2C# => romdata <= X"D7387453";
    when 16#00C2D# => romdata <= X"77527851";
    when 16#00C2E# => romdata <= X"EFBC3FB0";
    when 16#00C2F# => romdata <= X"0881FF06";
    when 16#00C30# => romdata <= X"77057083";
    when 16#00C31# => romdata <= X"FFFF0677";
    when 16#00C32# => romdata <= X"70810559";
    when 16#00C33# => romdata <= X"33525855";
    when 16#00C34# => romdata <= X"74FFBC38";
    when 16#00C35# => romdata <= X"FFB239CD";
    when 16#00C36# => romdata <= X"C73F04FB";
    when 16#00C37# => romdata <= X"3D0D7779";
    when 16#00C38# => romdata <= X"55558056";
    when 16#00C39# => romdata <= X"757524AB";
    when 16#00C3A# => romdata <= X"38807424";
    when 16#00C3B# => romdata <= X"9D388053";
    when 16#00C3C# => romdata <= X"73527451";
    when 16#00C3D# => romdata <= X"80E13FB0";
    when 16#00C3E# => romdata <= X"08547580";
    when 16#00C3F# => romdata <= X"2E8538B0";
    when 16#00C40# => romdata <= X"08305473";
    when 16#00C41# => romdata <= X"B00C873D";
    when 16#00C42# => romdata <= X"0D047330";
    when 16#00C43# => romdata <= X"76813257";
    when 16#00C44# => romdata <= X"54DC3974";
    when 16#00C45# => romdata <= X"30558156";
    when 16#00C46# => romdata <= X"738025D2";
    when 16#00C47# => romdata <= X"38EC39FA";
    when 16#00C48# => romdata <= X"3D0D787A";
    when 16#00C49# => romdata <= X"57558057";
    when 16#00C4A# => romdata <= X"767524A4";
    when 16#00C4B# => romdata <= X"38759F2C";
    when 16#00C4C# => romdata <= X"54815375";
    when 16#00C4D# => romdata <= X"74327431";
    when 16#00C4E# => romdata <= X"5274519B";
    when 16#00C4F# => romdata <= X"3FB00854";
    when 16#00C50# => romdata <= X"76802E85";
    when 16#00C51# => romdata <= X"38B00830";
    when 16#00C52# => romdata <= X"5473B00C";
    when 16#00C53# => romdata <= X"883D0D04";
    when 16#00C54# => romdata <= X"74305581";
    when 16#00C55# => romdata <= X"57D739FC";
    when 16#00C56# => romdata <= X"3D0D7678";
    when 16#00C57# => romdata <= X"53548153";
    when 16#00C58# => romdata <= X"80747326";
    when 16#00C59# => romdata <= X"52557280";
    when 16#00C5A# => romdata <= X"2E983870";
    when 16#00C5B# => romdata <= X"802EA938";
    when 16#00C5C# => romdata <= X"807224A4";
    when 16#00C5D# => romdata <= X"38711073";
    when 16#00C5E# => romdata <= X"10757226";
    when 16#00C5F# => romdata <= X"53545272";
    when 16#00C60# => romdata <= X"EA387351";
    when 16#00C61# => romdata <= X"78833874";
    when 16#00C62# => romdata <= X"5170B00C";
    when 16#00C63# => romdata <= X"863D0D04";
    when 16#00C64# => romdata <= X"72812A72";
    when 16#00C65# => romdata <= X"812A5353";
    when 16#00C66# => romdata <= X"72802EE6";
    when 16#00C67# => romdata <= X"38717426";
    when 16#00C68# => romdata <= X"EF387372";
    when 16#00C69# => romdata <= X"31757407";
    when 16#00C6A# => romdata <= X"74812A74";
    when 16#00C6B# => romdata <= X"812A5555";
    when 16#00C6C# => romdata <= X"5654E539";
    when 16#00C6D# => romdata <= X"10101010";
    when 16#00C6E# => romdata <= X"10101010";
    when 16#00C6F# => romdata <= X"10101010";
    when 16#00C70# => romdata <= X"10101010";
    when 16#00C71# => romdata <= X"10101010";
    when 16#00C72# => romdata <= X"10101010";
    when 16#00C73# => romdata <= X"10101010";
    when 16#00C74# => romdata <= X"10101053";
    when 16#00C75# => romdata <= X"51047381";
    when 16#00C76# => romdata <= X"FF067383";
    when 16#00C77# => romdata <= X"06098105";
    when 16#00C78# => romdata <= X"83051010";
    when 16#00C79# => romdata <= X"102B0772";
    when 16#00C7A# => romdata <= X"FC060C51";
    when 16#00C7B# => romdata <= X"51043C04";
    when 16#00C7C# => romdata <= X"72728072";
    when 16#00C7D# => romdata <= X"8106FF05";
    when 16#00C7E# => romdata <= X"09720605";
    when 16#00C7F# => romdata <= X"71105272";
    when 16#00C80# => romdata <= X"0A100A53";
    when 16#00C81# => romdata <= X"72ED3851";
    when 16#00C82# => romdata <= X"51535104";
    when 16#00C83# => romdata <= X"B008B408";
    when 16#00C84# => romdata <= X"B8087575";
    when 16#00C85# => romdata <= X"80E29F2D";
    when 16#00C86# => romdata <= X"5050B008";
    when 16#00C87# => romdata <= X"56B80CB4";
    when 16#00C88# => romdata <= X"0CB00C51";
    when 16#00C89# => romdata <= X"04B008B4";
    when 16#00C8A# => romdata <= X"08B80875";
    when 16#00C8B# => romdata <= X"7580E1DB";
    when 16#00C8C# => romdata <= X"2D5050B0";
    when 16#00C8D# => romdata <= X"0856B80C";
    when 16#00C8E# => romdata <= X"B40CB00C";
    when 16#00C8F# => romdata <= X"5104B008";
    when 16#00C90# => romdata <= X"B408B808";
    when 16#00C91# => romdata <= X"AEF72DB8";
    when 16#00C92# => romdata <= X"0CB40CB0";
    when 16#00C93# => romdata <= X"0C04FF3D";
    when 16#00C94# => romdata <= X"0D028F05";
    when 16#00C95# => romdata <= X"3381B2AC";
    when 16#00C96# => romdata <= X"0852710C";
    when 16#00C97# => romdata <= X"800BB00C";
    when 16#00C98# => romdata <= X"833D0D04";
    when 16#00C99# => romdata <= X"FF3D0D02";
    when 16#00C9A# => romdata <= X"8F053351";
    when 16#00C9B# => romdata <= X"81D5F408";
    when 16#00C9C# => romdata <= X"52712DB0";
    when 16#00C9D# => romdata <= X"0881FF06";
    when 16#00C9E# => romdata <= X"B00C833D";
    when 16#00C9F# => romdata <= X"0D04FE3D";
    when 16#00CA0# => romdata <= X"0D747033";
    when 16#00CA1# => romdata <= X"53537180";
    when 16#00CA2# => romdata <= X"2E933881";
    when 16#00CA3# => romdata <= X"13725281";
    when 16#00CA4# => romdata <= X"D5F40853";
    when 16#00CA5# => romdata <= X"53712D72";
    when 16#00CA6# => romdata <= X"335271EF";
    when 16#00CA7# => romdata <= X"38843D0D";
    when 16#00CA8# => romdata <= X"04F43D0D";
    when 16#00CA9# => romdata <= X"7F028405";
    when 16#00CAA# => romdata <= X"BB053355";
    when 16#00CAB# => romdata <= X"57880B8C";
    when 16#00CAC# => romdata <= X"3D5B5989";
    when 16#00CAD# => romdata <= X"5381AFC4";
    when 16#00CAE# => romdata <= X"52795186";
    when 16#00CAF# => romdata <= X"D93F7379";
    when 16#00CB0# => romdata <= X"2E80FF38";
    when 16#00CB1# => romdata <= X"78567390";
    when 16#00CB2# => romdata <= X"2E80EC38";
    when 16#00CB3# => romdata <= X"02A70558";
    when 16#00CB4# => romdata <= X"768F0654";
    when 16#00CB5# => romdata <= X"73892680";
    when 16#00CB6# => romdata <= X"C2387518";
    when 16#00CB7# => romdata <= X"B0155555";
    when 16#00CB8# => romdata <= X"73753476";
    when 16#00CB9# => romdata <= X"842AFF17";
    when 16#00CBA# => romdata <= X"7081FF06";
    when 16#00CBB# => romdata <= X"58555775";
    when 16#00CBC# => romdata <= X"DF38781A";
    when 16#00CBD# => romdata <= X"55757534";
    when 16#00CBE# => romdata <= X"79703355";
    when 16#00CBF# => romdata <= X"5573802E";
    when 16#00CC0# => romdata <= X"93388115";
    when 16#00CC1# => romdata <= X"745281D5";
    when 16#00CC2# => romdata <= X"F4085755";
    when 16#00CC3# => romdata <= X"752D7433";
    when 16#00CC4# => romdata <= X"5473EF38";
    when 16#00CC5# => romdata <= X"78B00C8E";
    when 16#00CC6# => romdata <= X"3D0D0475";
    when 16#00CC7# => romdata <= X"18B71555";
    when 16#00CC8# => romdata <= X"55737534";
    when 16#00CC9# => romdata <= X"76842AFF";
    when 16#00CCA# => romdata <= X"177081FF";
    when 16#00CCB# => romdata <= X"06585557";
    when 16#00CCC# => romdata <= X"75FF9D38";
    when 16#00CCD# => romdata <= X"FFBC3984";
    when 16#00CCE# => romdata <= X"70575902";
    when 16#00CCF# => romdata <= X"A70558FF";
    when 16#00CD0# => romdata <= X"8F398270";
    when 16#00CD1# => romdata <= X"5759F439";
    when 16#00CD2# => romdata <= X"F13D0D61";
    when 16#00CD3# => romdata <= X"8D3D705B";
    when 16#00CD4# => romdata <= X"5C5A807A";
    when 16#00CD5# => romdata <= X"5657767A";
    when 16#00CD6# => romdata <= X"24818538";
    when 16#00CD7# => romdata <= X"7817548A";
    when 16#00CD8# => romdata <= X"52745184";
    when 16#00CD9# => romdata <= X"FF3FB008";
    when 16#00CDA# => romdata <= X"B0055372";
    when 16#00CDB# => romdata <= X"74348117";
    when 16#00CDC# => romdata <= X"578A5274";
    when 16#00CDD# => romdata <= X"5184C83F";
    when 16#00CDE# => romdata <= X"B00855B0";
    when 16#00CDF# => romdata <= X"08DE38B0";
    when 16#00CE0# => romdata <= X"08779F2A";
    when 16#00CE1# => romdata <= X"1870812C";
    when 16#00CE2# => romdata <= X"5A565680";
    when 16#00CE3# => romdata <= X"78259E38";
    when 16#00CE4# => romdata <= X"7817FF05";
    when 16#00CE5# => romdata <= X"55751970";
    when 16#00CE6# => romdata <= X"33555374";
    when 16#00CE7# => romdata <= X"33733473";
    when 16#00CE8# => romdata <= X"75348116";
    when 16#00CE9# => romdata <= X"FF165656";
    when 16#00CEA# => romdata <= X"777624E9";
    when 16#00CEB# => romdata <= X"38761958";
    when 16#00CEC# => romdata <= X"80783480";
    when 16#00CED# => romdata <= X"7A241770";
    when 16#00CEE# => romdata <= X"81FF067C";
    when 16#00CEF# => romdata <= X"70335657";
    when 16#00CF0# => romdata <= X"55567280";
    when 16#00CF1# => romdata <= X"2E933881";
    when 16#00CF2# => romdata <= X"15735281";
    when 16#00CF3# => romdata <= X"D5F40858";
    when 16#00CF4# => romdata <= X"55762D74";
    when 16#00CF5# => romdata <= X"335372EF";
    when 16#00CF6# => romdata <= X"3873B00C";
    when 16#00CF7# => romdata <= X"913D0D04";
    when 16#00CF8# => romdata <= X"AD7B3402";
    when 16#00CF9# => romdata <= X"AD057A30";
    when 16#00CFA# => romdata <= X"71195656";
    when 16#00CFB# => romdata <= X"598A5274";
    when 16#00CFC# => romdata <= X"5183F13F";
    when 16#00CFD# => romdata <= X"B008B005";
    when 16#00CFE# => romdata <= X"53727434";
    when 16#00CFF# => romdata <= X"8117578A";
    when 16#00D00# => romdata <= X"52745183";
    when 16#00D01# => romdata <= X"BA3FB008";
    when 16#00D02# => romdata <= X"55B008FE";
    when 16#00D03# => romdata <= X"CF38FEEF";
    when 16#00D04# => romdata <= X"39FD3D0D";
    when 16#00D05# => romdata <= X"81B2A008";
    when 16#00D06# => romdata <= X"76B2E429";
    when 16#00D07# => romdata <= X"94120C54";
    when 16#00D08# => romdata <= X"850B9815";
    when 16#00D09# => romdata <= X"0C981408";
    when 16#00D0A# => romdata <= X"70810651";
    when 16#00D0B# => romdata <= X"5372F638";
    when 16#00D0C# => romdata <= X"853D0D04";
    when 16#00D0D# => romdata <= X"803D0D81";
    when 16#00D0E# => romdata <= X"B2A00851";
    when 16#00D0F# => romdata <= X"870B8412";
    when 16#00D10# => romdata <= X"0CFF0BA4";
    when 16#00D11# => romdata <= X"120CA70B";
    when 16#00D12# => romdata <= X"A8120CB2";
    when 16#00D13# => romdata <= X"E40B9412";
    when 16#00D14# => romdata <= X"0C870B98";
    when 16#00D15# => romdata <= X"120C823D";
    when 16#00D16# => romdata <= X"0D04803D";
    when 16#00D17# => romdata <= X"0D81B2A4";
    when 16#00D18# => romdata <= X"0851B80B";
    when 16#00D19# => romdata <= X"8C120C83";
    when 16#00D1A# => romdata <= X"0B88120C";
    when 16#00D1B# => romdata <= X"823D0D04";
    when 16#00D1C# => romdata <= X"803D0D81";
    when 16#00D1D# => romdata <= X"B2A40884";
    when 16#00D1E# => romdata <= X"11088106";
    when 16#00D1F# => romdata <= X"B00C5182";
    when 16#00D20# => romdata <= X"3D0D04FF";
    when 16#00D21# => romdata <= X"3D0D81B2";
    when 16#00D22# => romdata <= X"A4085284";
    when 16#00D23# => romdata <= X"12087081";
    when 16#00D24# => romdata <= X"06515170";
    when 16#00D25# => romdata <= X"802EF438";
    when 16#00D26# => romdata <= X"71087081";
    when 16#00D27# => romdata <= X"FF06B00C";
    when 16#00D28# => romdata <= X"51833D0D";
    when 16#00D29# => romdata <= X"04FE3D0D";
    when 16#00D2A# => romdata <= X"02930533";
    when 16#00D2B# => romdata <= X"81B2A408";
    when 16#00D2C# => romdata <= X"53538412";
    when 16#00D2D# => romdata <= X"0870892A";
    when 16#00D2E# => romdata <= X"70810651";
    when 16#00D2F# => romdata <= X"515170F2";
    when 16#00D30# => romdata <= X"3872720C";
    when 16#00D31# => romdata <= X"843D0D04";
    when 16#00D32# => romdata <= X"FE3D0D02";
    when 16#00D33# => romdata <= X"93053353";
    when 16#00D34# => romdata <= X"728A2E9C";
    when 16#00D35# => romdata <= X"3881B2A4";
    when 16#00D36# => romdata <= X"08528412";
    when 16#00D37# => romdata <= X"0870892A";
    when 16#00D38# => romdata <= X"70810651";
    when 16#00D39# => romdata <= X"515170F2";
    when 16#00D3A# => romdata <= X"3872720C";
    when 16#00D3B# => romdata <= X"843D0D04";
    when 16#00D3C# => romdata <= X"81B2A408";
    when 16#00D3D# => romdata <= X"52841208";
    when 16#00D3E# => romdata <= X"70892A70";
    when 16#00D3F# => romdata <= X"81065151";
    when 16#00D40# => romdata <= X"5170F238";
    when 16#00D41# => romdata <= X"8D720C84";
    when 16#00D42# => romdata <= X"12087089";
    when 16#00D43# => romdata <= X"2A708106";
    when 16#00D44# => romdata <= X"51515170";
    when 16#00D45# => romdata <= X"C538D239";
    when 16#00D46# => romdata <= X"803D0D81";
    when 16#00D47# => romdata <= X"B2980851";
    when 16#00D48# => romdata <= X"800B8412";
    when 16#00D49# => romdata <= X"0C83FE80";
    when 16#00D4A# => romdata <= X"0B88120C";
    when 16#00D4B# => romdata <= X"800B81D5";
    when 16#00D4C# => romdata <= X"F834800B";
    when 16#00D4D# => romdata <= X"81D5FC34";
    when 16#00D4E# => romdata <= X"823D0D04";
    when 16#00D4F# => romdata <= X"FA3D0D02";
    when 16#00D50# => romdata <= X"A3053381";
    when 16#00D51# => romdata <= X"B2980881";
    when 16#00D52# => romdata <= X"D5F83370";
    when 16#00D53# => romdata <= X"81FF0670";
    when 16#00D54# => romdata <= X"10101181";
    when 16#00D55# => romdata <= X"D5FC3370";
    when 16#00D56# => romdata <= X"81FF0672";
    when 16#00D57# => romdata <= X"90291170";
    when 16#00D58# => romdata <= X"882B7807";
    when 16#00D59# => romdata <= X"770C535B";
    when 16#00D5A# => romdata <= X"5B555559";
    when 16#00D5B# => romdata <= X"5454738A";
    when 16#00D5C# => romdata <= X"2E983874";
    when 16#00D5D# => romdata <= X"80CF2E92";
    when 16#00D5E# => romdata <= X"38738C2E";
    when 16#00D5F# => romdata <= X"A4388116";
    when 16#00D60# => romdata <= X"537281D5";
    when 16#00D61# => romdata <= X"FC34883D";
    when 16#00D62# => romdata <= X"0D0471A3";
    when 16#00D63# => romdata <= X"26A33881";
    when 16#00D64# => romdata <= X"17527181";
    when 16#00D65# => romdata <= X"D5F83480";
    when 16#00D66# => romdata <= X"0B81D5FC";
    when 16#00D67# => romdata <= X"34883D0D";
    when 16#00D68# => romdata <= X"04805271";
    when 16#00D69# => romdata <= X"882B730C";
    when 16#00D6A# => romdata <= X"81125297";
    when 16#00D6B# => romdata <= X"907226F3";
    when 16#00D6C# => romdata <= X"38800B81";
    when 16#00D6D# => romdata <= X"D5F83480";
    when 16#00D6E# => romdata <= X"0B81D5FC";
    when 16#00D6F# => romdata <= X"34DF39BC";
    when 16#00D70# => romdata <= X"0802BC0C";
    when 16#00D71# => romdata <= X"FD3D0D80";
    when 16#00D72# => romdata <= X"53BC088C";
    when 16#00D73# => romdata <= X"050852BC";
    when 16#00D74# => romdata <= X"08880508";
    when 16#00D75# => romdata <= X"51F7803F";
    when 16#00D76# => romdata <= X"B00870B0";
    when 16#00D77# => romdata <= X"0C54853D";
    when 16#00D78# => romdata <= X"0DBC0C04";
    when 16#00D79# => romdata <= X"BC0802BC";
    when 16#00D7A# => romdata <= X"0CFD3D0D";
    when 16#00D7B# => romdata <= X"8153BC08";
    when 16#00D7C# => romdata <= X"8C050852";
    when 16#00D7D# => romdata <= X"BC088805";
    when 16#00D7E# => romdata <= X"0851F6DB";
    when 16#00D7F# => romdata <= X"3FB00870";
    when 16#00D80# => romdata <= X"B00C5485";
    when 16#00D81# => romdata <= X"3D0DBC0C";
    when 16#00D82# => romdata <= X"04803D0D";
    when 16#00D83# => romdata <= X"86518496";
    when 16#00D84# => romdata <= X"3F8151A1";
    when 16#00D85# => romdata <= X"D33FFC3D";
    when 16#00D86# => romdata <= X"0D767079";
    when 16#00D87# => romdata <= X"7B555555";
    when 16#00D88# => romdata <= X"558F7227";
    when 16#00D89# => romdata <= X"8C387275";
    when 16#00D8A# => romdata <= X"07830651";
    when 16#00D8B# => romdata <= X"70802EA7";
    when 16#00D8C# => romdata <= X"38FF1252";
    when 16#00D8D# => romdata <= X"71FF2E98";
    when 16#00D8E# => romdata <= X"38727081";
    when 16#00D8F# => romdata <= X"05543374";
    when 16#00D90# => romdata <= X"70810556";
    when 16#00D91# => romdata <= X"34FF1252";
    when 16#00D92# => romdata <= X"71FF2E09";
    when 16#00D93# => romdata <= X"8106EA38";
    when 16#00D94# => romdata <= X"74B00C86";
    when 16#00D95# => romdata <= X"3D0D0474";
    when 16#00D96# => romdata <= X"51727084";
    when 16#00D97# => romdata <= X"05540871";
    when 16#00D98# => romdata <= X"70840553";
    when 16#00D99# => romdata <= X"0C727084";
    when 16#00D9A# => romdata <= X"05540871";
    when 16#00D9B# => romdata <= X"70840553";
    when 16#00D9C# => romdata <= X"0C727084";
    when 16#00D9D# => romdata <= X"05540871";
    when 16#00D9E# => romdata <= X"70840553";
    when 16#00D9F# => romdata <= X"0C727084";
    when 16#00DA0# => romdata <= X"05540871";
    when 16#00DA1# => romdata <= X"70840553";
    when 16#00DA2# => romdata <= X"0CF01252";
    when 16#00DA3# => romdata <= X"718F26C9";
    when 16#00DA4# => romdata <= X"38837227";
    when 16#00DA5# => romdata <= X"95387270";
    when 16#00DA6# => romdata <= X"84055408";
    when 16#00DA7# => romdata <= X"71708405";
    when 16#00DA8# => romdata <= X"530CFC12";
    when 16#00DA9# => romdata <= X"52718326";
    when 16#00DAA# => romdata <= X"ED387054";
    when 16#00DAB# => romdata <= X"FF8339FD";
    when 16#00DAC# => romdata <= X"3D0D7553";
    when 16#00DAD# => romdata <= X"84D81308";
    when 16#00DAE# => romdata <= X"802E8A38";
    when 16#00DAF# => romdata <= X"805372B0";
    when 16#00DB0# => romdata <= X"0C853D0D";
    when 16#00DB1# => romdata <= X"04818052";
    when 16#00DB2# => romdata <= X"72518D9B";
    when 16#00DB3# => romdata <= X"3FB00884";
    when 16#00DB4# => romdata <= X"D8140CFF";
    when 16#00DB5# => romdata <= X"53B00880";
    when 16#00DB6# => romdata <= X"2EE438B0";
    when 16#00DB7# => romdata <= X"08549F53";
    when 16#00DB8# => romdata <= X"80747084";
    when 16#00DB9# => romdata <= X"05560CFF";
    when 16#00DBA# => romdata <= X"13538073";
    when 16#00DBB# => romdata <= X"24CE3880";
    when 16#00DBC# => romdata <= X"74708405";
    when 16#00DBD# => romdata <= X"560CFF13";
    when 16#00DBE# => romdata <= X"53728025";
    when 16#00DBF# => romdata <= X"E338FFBC";
    when 16#00DC0# => romdata <= X"39FD3D0D";
    when 16#00DC1# => romdata <= X"75775553";
    when 16#00DC2# => romdata <= X"9F74278D";
    when 16#00DC3# => romdata <= X"3896730C";
    when 16#00DC4# => romdata <= X"FF5271B0";
    when 16#00DC5# => romdata <= X"0C853D0D";
    when 16#00DC6# => romdata <= X"0484D813";
    when 16#00DC7# => romdata <= X"08527180";
    when 16#00DC8# => romdata <= X"2E933873";
    when 16#00DC9# => romdata <= X"10101270";
    when 16#00DCA# => romdata <= X"0879720C";
    when 16#00DCB# => romdata <= X"515271B0";
    when 16#00DCC# => romdata <= X"0C853D0D";
    when 16#00DCD# => romdata <= X"047251FE";
    when 16#00DCE# => romdata <= X"F63FFF52";
    when 16#00DCF# => romdata <= X"B008D338";
    when 16#00DD0# => romdata <= X"84D81308";
    when 16#00DD1# => romdata <= X"74101011";
    when 16#00DD2# => romdata <= X"70087A72";
    when 16#00DD3# => romdata <= X"0C515152";
    when 16#00DD4# => romdata <= X"DD39F93D";
    when 16#00DD5# => romdata <= X"0D797B58";
    when 16#00DD6# => romdata <= X"56769F26";
    when 16#00DD7# => romdata <= X"80E83884";
    when 16#00DD8# => romdata <= X"D8160854";
    when 16#00DD9# => romdata <= X"73802EAA";
    when 16#00DDA# => romdata <= X"38761010";
    when 16#00DDB# => romdata <= X"14700855";
    when 16#00DDC# => romdata <= X"5573802E";
    when 16#00DDD# => romdata <= X"BA388058";
    when 16#00DDE# => romdata <= X"73812E8F";
    when 16#00DDF# => romdata <= X"3873FF2E";
    when 16#00DE0# => romdata <= X"A3388075";
    when 16#00DE1# => romdata <= X"0C765173";
    when 16#00DE2# => romdata <= X"2D805877";
    when 16#00DE3# => romdata <= X"B00C893D";
    when 16#00DE4# => romdata <= X"0D047551";
    when 16#00DE5# => romdata <= X"FE993FFF";
    when 16#00DE6# => romdata <= X"58B008EF";
    when 16#00DE7# => romdata <= X"3884D816";
    when 16#00DE8# => romdata <= X"0854C639";
    when 16#00DE9# => romdata <= X"96760C81";
    when 16#00DEA# => romdata <= X"0BB00C89";
    when 16#00DEB# => romdata <= X"3D0D0475";
    when 16#00DEC# => romdata <= X"5181ED3F";
    when 16#00DED# => romdata <= X"7653B008";
    when 16#00DEE# => romdata <= X"52755181";
    when 16#00DEF# => romdata <= X"AD3FB008";
    when 16#00DF0# => romdata <= X"B00C893D";
    when 16#00DF1# => romdata <= X"0D049676";
    when 16#00DF2# => romdata <= X"0CFF0BB0";
    when 16#00DF3# => romdata <= X"0C893D0D";
    when 16#00DF4# => romdata <= X"04FC3D0D";
    when 16#00DF5# => romdata <= X"76785653";
    when 16#00DF6# => romdata <= X"FF54749F";
    when 16#00DF7# => romdata <= X"26B13884";
    when 16#00DF8# => romdata <= X"D8130852";
    when 16#00DF9# => romdata <= X"71802EAE";
    when 16#00DFA# => romdata <= X"38741010";
    when 16#00DFB# => romdata <= X"12700853";
    when 16#00DFC# => romdata <= X"53815471";
    when 16#00DFD# => romdata <= X"802E9838";
    when 16#00DFE# => romdata <= X"825471FF";
    when 16#00DFF# => romdata <= X"2E913883";
    when 16#00E00# => romdata <= X"5471812E";
    when 16#00E01# => romdata <= X"8A388073";
    when 16#00E02# => romdata <= X"0C745171";
    when 16#00E03# => romdata <= X"2D805473";
    when 16#00E04# => romdata <= X"B00C863D";
    when 16#00E05# => romdata <= X"0D047251";
    when 16#00E06# => romdata <= X"FD953FB0";
    when 16#00E07# => romdata <= X"08F13884";
    when 16#00E08# => romdata <= X"D8130852";
    when 16#00E09# => romdata <= X"C439FF3D";
    when 16#00E0A# => romdata <= X"0D735281";
    when 16#00E0B# => romdata <= X"B2B00851";
    when 16#00E0C# => romdata <= X"FEA03F83";
    when 16#00E0D# => romdata <= X"3D0D04FE";
    when 16#00E0E# => romdata <= X"3D0D7553";
    when 16#00E0F# => romdata <= X"745281B2";
    when 16#00E10# => romdata <= X"B00851FD";
    when 16#00E11# => romdata <= X"BC3F843D";
    when 16#00E12# => romdata <= X"0D04803D";
    when 16#00E13# => romdata <= X"0D81B2B0";
    when 16#00E14# => romdata <= X"0851FCDB";
    when 16#00E15# => romdata <= X"3F823D0D";
    when 16#00E16# => romdata <= X"04FF3D0D";
    when 16#00E17# => romdata <= X"735281B2";
    when 16#00E18# => romdata <= X"B00851FE";
    when 16#00E19# => romdata <= X"EC3F833D";
    when 16#00E1A# => romdata <= X"0D04FC3D";
    when 16#00E1B# => romdata <= X"0D800B81";
    when 16#00E1C# => romdata <= X"D6840C78";
    when 16#00E1D# => romdata <= X"5277519C";
    when 16#00E1E# => romdata <= X"AA3FB008";
    when 16#00E1F# => romdata <= X"54B008FF";
    when 16#00E20# => romdata <= X"2E883873";
    when 16#00E21# => romdata <= X"B00C863D";
    when 16#00E22# => romdata <= X"0D0481D6";
    when 16#00E23# => romdata <= X"84085574";
    when 16#00E24# => romdata <= X"802EF038";
    when 16#00E25# => romdata <= X"7675710C";
    when 16#00E26# => romdata <= X"5373B00C";
    when 16#00E27# => romdata <= X"863D0D04";
    when 16#00E28# => romdata <= X"9BFC3F04";
    when 16#00E29# => romdata <= X"FC3D0D76";
    when 16#00E2A# => romdata <= X"70797073";
    when 16#00E2B# => romdata <= X"07830654";
    when 16#00E2C# => romdata <= X"54545570";
    when 16#00E2D# => romdata <= X"80C33871";
    when 16#00E2E# => romdata <= X"70087009";
    when 16#00E2F# => romdata <= X"70F7FBFD";
    when 16#00E30# => romdata <= X"FF130670";
    when 16#00E31# => romdata <= X"F8848281";
    when 16#00E32# => romdata <= X"80065151";
    when 16#00E33# => romdata <= X"53535470";
    when 16#00E34# => romdata <= X"A6388414";
    when 16#00E35# => romdata <= X"72747084";
    when 16#00E36# => romdata <= X"05560C70";
    when 16#00E37# => romdata <= X"08700970";
    when 16#00E38# => romdata <= X"F7FBFDFF";
    when 16#00E39# => romdata <= X"130670F8";
    when 16#00E3A# => romdata <= X"84828180";
    when 16#00E3B# => romdata <= X"06515153";
    when 16#00E3C# => romdata <= X"53547080";
    when 16#00E3D# => romdata <= X"2EDC3873";
    when 16#00E3E# => romdata <= X"52717081";
    when 16#00E3F# => romdata <= X"05533351";
    when 16#00E40# => romdata <= X"70737081";
    when 16#00E41# => romdata <= X"05553470";
    when 16#00E42# => romdata <= X"F03874B0";
    when 16#00E43# => romdata <= X"0C863D0D";
    when 16#00E44# => romdata <= X"04FD3D0D";
    when 16#00E45# => romdata <= X"75707183";
    when 16#00E46# => romdata <= X"06535552";
    when 16#00E47# => romdata <= X"70B83871";
    when 16#00E48# => romdata <= X"70087009";
    when 16#00E49# => romdata <= X"F7FBFDFF";
    when 16#00E4A# => romdata <= X"120670F8";
    when 16#00E4B# => romdata <= X"84828180";
    when 16#00E4C# => romdata <= X"06515152";
    when 16#00E4D# => romdata <= X"53709D38";
    when 16#00E4E# => romdata <= X"84137008";
    when 16#00E4F# => romdata <= X"7009F7FB";
    when 16#00E50# => romdata <= X"FDFF1206";
    when 16#00E51# => romdata <= X"70F88482";
    when 16#00E52# => romdata <= X"81800651";
    when 16#00E53# => romdata <= X"51525370";
    when 16#00E54# => romdata <= X"802EE538";
    when 16#00E55# => romdata <= X"72527133";
    when 16#00E56# => romdata <= X"5170802E";
    when 16#00E57# => romdata <= X"8A388112";
    when 16#00E58# => romdata <= X"70335252";
    when 16#00E59# => romdata <= X"70F83871";
    when 16#00E5A# => romdata <= X"7431B00C";
    when 16#00E5B# => romdata <= X"853D0D04";
    when 16#00E5C# => romdata <= X"FA3D0D78";
    when 16#00E5D# => romdata <= X"7A7C7054";
    when 16#00E5E# => romdata <= X"55555272";
    when 16#00E5F# => romdata <= X"802E80D9";
    when 16#00E60# => romdata <= X"38717407";
    when 16#00E61# => romdata <= X"83065170";
    when 16#00E62# => romdata <= X"802E80D4";
    when 16#00E63# => romdata <= X"38FF1353";
    when 16#00E64# => romdata <= X"72FF2EB1";
    when 16#00E65# => romdata <= X"38713374";
    when 16#00E66# => romdata <= X"33565174";
    when 16#00E67# => romdata <= X"712E0981";
    when 16#00E68# => romdata <= X"06A93872";
    when 16#00E69# => romdata <= X"802E8187";
    when 16#00E6A# => romdata <= X"387081FF";
    when 16#00E6B# => romdata <= X"06517080";
    when 16#00E6C# => romdata <= X"2E80FC38";
    when 16#00E6D# => romdata <= X"81128115";
    when 16#00E6E# => romdata <= X"FF155555";
    when 16#00E6F# => romdata <= X"5272FF2E";
    when 16#00E70# => romdata <= X"098106D1";
    when 16#00E71# => romdata <= X"38713374";
    when 16#00E72# => romdata <= X"33565170";
    when 16#00E73# => romdata <= X"81FF0675";
    when 16#00E74# => romdata <= X"81FF0671";
    when 16#00E75# => romdata <= X"71315152";
    when 16#00E76# => romdata <= X"5270B00C";
    when 16#00E77# => romdata <= X"883D0D04";
    when 16#00E78# => romdata <= X"71745755";
    when 16#00E79# => romdata <= X"83732788";
    when 16#00E7A# => romdata <= X"38710874";
    when 16#00E7B# => romdata <= X"082E8838";
    when 16#00E7C# => romdata <= X"74765552";
    when 16#00E7D# => romdata <= X"FF9739FC";
    when 16#00E7E# => romdata <= X"13537280";
    when 16#00E7F# => romdata <= X"2EB13874";
    when 16#00E80# => romdata <= X"087009F7";
    when 16#00E81# => romdata <= X"FBFDFF12";
    when 16#00E82# => romdata <= X"0670F884";
    when 16#00E83# => romdata <= X"82818006";
    when 16#00E84# => romdata <= X"51515170";
    when 16#00E85# => romdata <= X"9A388415";
    when 16#00E86# => romdata <= X"84175755";
    when 16#00E87# => romdata <= X"837327D0";
    when 16#00E88# => romdata <= X"38740876";
    when 16#00E89# => romdata <= X"082ED038";
    when 16#00E8A# => romdata <= X"74765552";
    when 16#00E8B# => romdata <= X"FEDF3980";
    when 16#00E8C# => romdata <= X"0BB00C88";
    when 16#00E8D# => romdata <= X"3D0D04F3";
    when 16#00E8E# => romdata <= X"3D0D6062";
    when 16#00E8F# => romdata <= X"64725A5A";
    when 16#00E90# => romdata <= X"5E5E805C";
    when 16#00E91# => romdata <= X"76708105";
    when 16#00E92# => romdata <= X"583381AF";
    when 16#00E93# => romdata <= X"D1113370";
    when 16#00E94# => romdata <= X"832A7081";
    when 16#00E95# => romdata <= X"06515555";
    when 16#00E96# => romdata <= X"5672E938";
    when 16#00E97# => romdata <= X"75AD2E82";
    when 16#00E98# => romdata <= X"883875AB";
    when 16#00E99# => romdata <= X"2E828438";
    when 16#00E9A# => romdata <= X"77307079";
    when 16#00E9B# => romdata <= X"07802579";
    when 16#00E9C# => romdata <= X"90327030";
    when 16#00E9D# => romdata <= X"70720780";
    when 16#00E9E# => romdata <= X"25730753";
    when 16#00E9F# => romdata <= X"57575153";
    when 16#00EA0# => romdata <= X"72802E87";
    when 16#00EA1# => romdata <= X"3875B02E";
    when 16#00EA2# => romdata <= X"81EB3877";
    when 16#00EA3# => romdata <= X"8A388858";
    when 16#00EA4# => romdata <= X"75B02E83";
    when 16#00EA5# => romdata <= X"388A5881";
    when 16#00EA6# => romdata <= X"0A5A7B84";
    when 16#00EA7# => romdata <= X"38FE0A5A";
    when 16#00EA8# => romdata <= X"77527951";
    when 16#00EA9# => romdata <= X"F6BE3FB0";
    when 16#00EAA# => romdata <= X"0878537A";
    when 16#00EAB# => romdata <= X"525BF68F";
    when 16#00EAC# => romdata <= X"3FB0085A";
    when 16#00EAD# => romdata <= X"807081AF";
    when 16#00EAE# => romdata <= X"D1183370";
    when 16#00EAF# => romdata <= X"822A7081";
    when 16#00EB0# => romdata <= X"06515656";
    when 16#00EB1# => romdata <= X"5A557280";
    when 16#00EB2# => romdata <= X"2E80C138";
    when 16#00EB3# => romdata <= X"D0165675";
    when 16#00EB4# => romdata <= X"782580D7";
    when 16#00EB5# => romdata <= X"38807924";
    when 16#00EB6# => romdata <= X"757B2607";
    when 16#00EB7# => romdata <= X"53729338";
    when 16#00EB8# => romdata <= X"747A2E80";
    when 16#00EB9# => romdata <= X"EB387A76";
    when 16#00EBA# => romdata <= X"2580ED38";
    when 16#00EBB# => romdata <= X"72802E80";
    when 16#00EBC# => romdata <= X"E738FF77";
    when 16#00EBD# => romdata <= X"70810559";
    when 16#00EBE# => romdata <= X"33575981";
    when 16#00EBF# => romdata <= X"AFD11633";
    when 16#00EC0# => romdata <= X"70822A70";
    when 16#00EC1# => romdata <= X"81065154";
    when 16#00EC2# => romdata <= X"5472C138";
    when 16#00EC3# => romdata <= X"73830653";
    when 16#00EC4# => romdata <= X"72802E97";
    when 16#00EC5# => romdata <= X"38738106";
    when 16#00EC6# => romdata <= X"C9175553";
    when 16#00EC7# => romdata <= X"728538FF";
    when 16#00EC8# => romdata <= X"A9165473";
    when 16#00EC9# => romdata <= X"56777624";
    when 16#00ECA# => romdata <= X"FFAB3880";
    when 16#00ECB# => romdata <= X"792480F0";
    when 16#00ECC# => romdata <= X"387B802E";
    when 16#00ECD# => romdata <= X"84387430";
    when 16#00ECE# => romdata <= X"557C802E";
    when 16#00ECF# => romdata <= X"8C38FF17";
    when 16#00ED0# => romdata <= X"53788338";
    when 16#00ED1# => romdata <= X"7D53727D";
    when 16#00ED2# => romdata <= X"0C74B00C";
    when 16#00ED3# => romdata <= X"8F3D0D04";
    when 16#00ED4# => romdata <= X"8153757B";
    when 16#00ED5# => romdata <= X"24FF9538";
    when 16#00ED6# => romdata <= X"81757929";
    when 16#00ED7# => romdata <= X"17787081";
    when 16#00ED8# => romdata <= X"055A3358";
    when 16#00ED9# => romdata <= X"5659FF93";
    when 16#00EDA# => romdata <= X"39815C76";
    when 16#00EDB# => romdata <= X"70810558";
    when 16#00EDC# => romdata <= X"3356FDF4";
    when 16#00EDD# => romdata <= X"39807733";
    when 16#00EDE# => romdata <= X"54547280";
    when 16#00EDF# => romdata <= X"F82EB238";
    when 16#00EE0# => romdata <= X"7280D832";
    when 16#00EE1# => romdata <= X"70307080";
    when 16#00EE2# => romdata <= X"25760751";
    when 16#00EE3# => romdata <= X"51537280";
    when 16#00EE4# => romdata <= X"2EFDF838";
    when 16#00EE5# => romdata <= X"81173382";
    when 16#00EE6# => romdata <= X"18585690";
    when 16#00EE7# => romdata <= X"58FDF839";
    when 16#00EE8# => romdata <= X"810A557B";
    when 16#00EE9# => romdata <= X"8438FE0A";
    when 16#00EEA# => romdata <= X"557F53A2";
    when 16#00EEB# => romdata <= X"730CFF89";
    when 16#00EEC# => romdata <= X"398154CC";
    when 16#00EED# => romdata <= X"39FD3D0D";
    when 16#00EEE# => romdata <= X"77547653";
    when 16#00EEF# => romdata <= X"755281B2";
    when 16#00EF0# => romdata <= X"B00851FC";
    when 16#00EF1# => romdata <= X"F23F853D";
    when 16#00EF2# => romdata <= X"0D04F33D";
    when 16#00EF3# => romdata <= X"0D606264";
    when 16#00EF4# => romdata <= X"725A5A5D";
    when 16#00EF5# => romdata <= X"5D805E76";
    when 16#00EF6# => romdata <= X"70810558";
    when 16#00EF7# => romdata <= X"3381AFD1";
    when 16#00EF8# => romdata <= X"11337083";
    when 16#00EF9# => romdata <= X"2A708106";
    when 16#00EFA# => romdata <= X"51555556";
    when 16#00EFB# => romdata <= X"72E93875";
    when 16#00EFC# => romdata <= X"AD2E81FF";
    when 16#00EFD# => romdata <= X"3875AB2E";
    when 16#00EFE# => romdata <= X"81FB3877";
    when 16#00EFF# => romdata <= X"30707907";
    when 16#00F00# => romdata <= X"80257990";
    when 16#00F01# => romdata <= X"32703070";
    when 16#00F02# => romdata <= X"72078025";
    when 16#00F03# => romdata <= X"73075357";
    when 16#00F04# => romdata <= X"57515372";
    when 16#00F05# => romdata <= X"802E8738";
    when 16#00F06# => romdata <= X"75B02E81";
    when 16#00F07# => romdata <= X"E238778A";
    when 16#00F08# => romdata <= X"38885875";
    when 16#00F09# => romdata <= X"B02E8338";
    when 16#00F0A# => romdata <= X"8A587752";
    when 16#00F0B# => romdata <= X"FF51F38F";
    when 16#00F0C# => romdata <= X"3FB00878";
    when 16#00F0D# => romdata <= X"535AFF51";
    when 16#00F0E# => romdata <= X"F3AA3FB0";
    when 16#00F0F# => romdata <= X"085B8070";
    when 16#00F10# => romdata <= X"5A5581AF";
    when 16#00F11# => romdata <= X"D1163370";
    when 16#00F12# => romdata <= X"822A7081";
    when 16#00F13# => romdata <= X"06515454";
    when 16#00F14# => romdata <= X"72802E80";
    when 16#00F15# => romdata <= X"C138D016";
    when 16#00F16# => romdata <= X"56757825";
    when 16#00F17# => romdata <= X"80D73880";
    when 16#00F18# => romdata <= X"7924757B";
    when 16#00F19# => romdata <= X"26075372";
    when 16#00F1A# => romdata <= X"9338747A";
    when 16#00F1B# => romdata <= X"2E80EB38";
    when 16#00F1C# => romdata <= X"7A762580";
    when 16#00F1D# => romdata <= X"ED387280";
    when 16#00F1E# => romdata <= X"2E80E738";
    when 16#00F1F# => romdata <= X"FF777081";
    when 16#00F20# => romdata <= X"05593357";
    when 16#00F21# => romdata <= X"5981AFD1";
    when 16#00F22# => romdata <= X"16337082";
    when 16#00F23# => romdata <= X"2A708106";
    when 16#00F24# => romdata <= X"51545472";
    when 16#00F25# => romdata <= X"C1387383";
    when 16#00F26# => romdata <= X"06537280";
    when 16#00F27# => romdata <= X"2E973873";
    when 16#00F28# => romdata <= X"8106C917";
    when 16#00F29# => romdata <= X"55537285";
    when 16#00F2A# => romdata <= X"38FFA916";
    when 16#00F2B# => romdata <= X"54735677";
    when 16#00F2C# => romdata <= X"7624FFAB";
    when 16#00F2D# => romdata <= X"38807924";
    when 16#00F2E# => romdata <= X"8189387D";
    when 16#00F2F# => romdata <= X"802E8438";
    when 16#00F30# => romdata <= X"7430557B";
    when 16#00F31# => romdata <= X"802E8C38";
    when 16#00F32# => romdata <= X"FF175378";
    when 16#00F33# => romdata <= X"83387C53";
    when 16#00F34# => romdata <= X"727C0C74";
    when 16#00F35# => romdata <= X"B00C8F3D";
    when 16#00F36# => romdata <= X"0D048153";
    when 16#00F37# => romdata <= X"757B24FF";
    when 16#00F38# => romdata <= X"95388175";
    when 16#00F39# => romdata <= X"79291778";
    when 16#00F3A# => romdata <= X"7081055A";
    when 16#00F3B# => romdata <= X"33585659";
    when 16#00F3C# => romdata <= X"FF933981";
    when 16#00F3D# => romdata <= X"5E767081";
    when 16#00F3E# => romdata <= X"05583356";
    when 16#00F3F# => romdata <= X"FDFD3980";
    when 16#00F40# => romdata <= X"77335454";
    when 16#00F41# => romdata <= X"7280F82E";
    when 16#00F42# => romdata <= X"80C33872";
    when 16#00F43# => romdata <= X"80D83270";
    when 16#00F44# => romdata <= X"30708025";
    when 16#00F45# => romdata <= X"76075151";
    when 16#00F46# => romdata <= X"5372802E";
    when 16#00F47# => romdata <= X"FE803881";
    when 16#00F48# => romdata <= X"17338218";
    when 16#00F49# => romdata <= X"58569070";
    when 16#00F4A# => romdata <= X"5358FF51";
    when 16#00F4B# => romdata <= X"F1913FB0";
    when 16#00F4C# => romdata <= X"0878535A";
    when 16#00F4D# => romdata <= X"FF51F1AC";
    when 16#00F4E# => romdata <= X"3FB0085B";
    when 16#00F4F# => romdata <= X"80705A55";
    when 16#00F50# => romdata <= X"FE8039FF";
    when 16#00F51# => romdata <= X"605455A2";
    when 16#00F52# => romdata <= X"730CFEF7";
    when 16#00F53# => romdata <= X"398154FF";
    when 16#00F54# => romdata <= X"BA39FD3D";
    when 16#00F55# => romdata <= X"0D775476";
    when 16#00F56# => romdata <= X"53755281";
    when 16#00F57# => romdata <= X"B2B00851";
    when 16#00F58# => romdata <= X"FCE83F85";
    when 16#00F59# => romdata <= X"3D0D04F3";
    when 16#00F5A# => romdata <= X"3D0D7F61";
    when 16#00F5B# => romdata <= X"8B1170F8";
    when 16#00F5C# => romdata <= X"065C5555";
    when 16#00F5D# => romdata <= X"5E729626";
    when 16#00F5E# => romdata <= X"83389059";
    when 16#00F5F# => romdata <= X"80792474";
    when 16#00F60# => romdata <= X"7A260753";
    when 16#00F61# => romdata <= X"80547274";
    when 16#00F62# => romdata <= X"2E098106";
    when 16#00F63# => romdata <= X"80CB387D";
    when 16#00F64# => romdata <= X"518BCA3F";
    when 16#00F65# => romdata <= X"7883F726";
    when 16#00F66# => romdata <= X"80C63878";
    when 16#00F67# => romdata <= X"832A7010";
    when 16#00F68# => romdata <= X"101081B9";
    when 16#00F69# => romdata <= X"EC058C11";
    when 16#00F6A# => romdata <= X"0859595A";
    when 16#00F6B# => romdata <= X"76782E83";
    when 16#00F6C# => romdata <= X"B0388417";
    when 16#00F6D# => romdata <= X"08FC0656";
    when 16#00F6E# => romdata <= X"8C170888";
    when 16#00F6F# => romdata <= X"1808718C";
    when 16#00F70# => romdata <= X"120C8812";
    when 16#00F71# => romdata <= X"0C587517";
    when 16#00F72# => romdata <= X"84110881";
    when 16#00F73# => romdata <= X"0784120C";
    when 16#00F74# => romdata <= X"537D518B";
    when 16#00F75# => romdata <= X"893F8817";
    when 16#00F76# => romdata <= X"5473B00C";
    when 16#00F77# => romdata <= X"8F3D0D04";
    when 16#00F78# => romdata <= X"78892A79";
    when 16#00F79# => romdata <= X"832A5B53";
    when 16#00F7A# => romdata <= X"72802EBF";
    when 16#00F7B# => romdata <= X"3878862A";
    when 16#00F7C# => romdata <= X"B8055A84";
    when 16#00F7D# => romdata <= X"7327B438";
    when 16#00F7E# => romdata <= X"80DB135A";
    when 16#00F7F# => romdata <= X"947327AB";
    when 16#00F80# => romdata <= X"38788C2A";
    when 16#00F81# => romdata <= X"80EE055A";
    when 16#00F82# => romdata <= X"80D47327";
    when 16#00F83# => romdata <= X"9E38788F";
    when 16#00F84# => romdata <= X"2A80F705";
    when 16#00F85# => romdata <= X"5A82D473";
    when 16#00F86# => romdata <= X"27913878";
    when 16#00F87# => romdata <= X"922A80FC";
    when 16#00F88# => romdata <= X"055A8AD4";
    when 16#00F89# => romdata <= X"73278438";
    when 16#00F8A# => romdata <= X"80FE5A79";
    when 16#00F8B# => romdata <= X"10101081";
    when 16#00F8C# => romdata <= X"B9EC058C";
    when 16#00F8D# => romdata <= X"11085855";
    when 16#00F8E# => romdata <= X"76752EA3";
    when 16#00F8F# => romdata <= X"38841708";
    when 16#00F90# => romdata <= X"FC06707A";
    when 16#00F91# => romdata <= X"31555673";
    when 16#00F92# => romdata <= X"8F2488D5";
    when 16#00F93# => romdata <= X"38738025";
    when 16#00F94# => romdata <= X"FEE6388C";
    when 16#00F95# => romdata <= X"17085776";
    when 16#00F96# => romdata <= X"752E0981";
    when 16#00F97# => romdata <= X"06DF3881";
    when 16#00F98# => romdata <= X"1A5A81B9";
    when 16#00F99# => romdata <= X"FC085776";
    when 16#00F9A# => romdata <= X"81B9F42E";
    when 16#00F9B# => romdata <= X"82C03884";
    when 16#00F9C# => romdata <= X"1708FC06";
    when 16#00F9D# => romdata <= X"707A3155";
    when 16#00F9E# => romdata <= X"56738F24";
    when 16#00F9F# => romdata <= X"81F93881";
    when 16#00FA0# => romdata <= X"B9F40B81";
    when 16#00FA1# => romdata <= X"BA800C81";
    when 16#00FA2# => romdata <= X"B9F40B81";
    when 16#00FA3# => romdata <= X"B9FC0C73";
    when 16#00FA4# => romdata <= X"8025FEB2";
    when 16#00FA5# => romdata <= X"3883FF76";
    when 16#00FA6# => romdata <= X"2783DF38";
    when 16#00FA7# => romdata <= X"75892A76";
    when 16#00FA8# => romdata <= X"832A5553";
    when 16#00FA9# => romdata <= X"72802EBF";
    when 16#00FAA# => romdata <= X"3875862A";
    when 16#00FAB# => romdata <= X"B8055484";
    when 16#00FAC# => romdata <= X"7327B438";
    when 16#00FAD# => romdata <= X"80DB1354";
    when 16#00FAE# => romdata <= X"947327AB";
    when 16#00FAF# => romdata <= X"38758C2A";
    when 16#00FB0# => romdata <= X"80EE0554";
    when 16#00FB1# => romdata <= X"80D47327";
    when 16#00FB2# => romdata <= X"9E38758F";
    when 16#00FB3# => romdata <= X"2A80F705";
    when 16#00FB4# => romdata <= X"5482D473";
    when 16#00FB5# => romdata <= X"27913875";
    when 16#00FB6# => romdata <= X"922A80FC";
    when 16#00FB7# => romdata <= X"05548AD4";
    when 16#00FB8# => romdata <= X"73278438";
    when 16#00FB9# => romdata <= X"80FE5473";
    when 16#00FBA# => romdata <= X"10101081";
    when 16#00FBB# => romdata <= X"B9EC0588";
    when 16#00FBC# => romdata <= X"11085658";
    when 16#00FBD# => romdata <= X"74782E86";
    when 16#00FBE# => romdata <= X"CF388415";
    when 16#00FBF# => romdata <= X"08FC0653";
    when 16#00FC0# => romdata <= X"7573278D";
    when 16#00FC1# => romdata <= X"38881508";
    when 16#00FC2# => romdata <= X"5574782E";
    when 16#00FC3# => romdata <= X"098106EA";
    when 16#00FC4# => romdata <= X"388C1508";
    when 16#00FC5# => romdata <= X"81B9EC0B";
    when 16#00FC6# => romdata <= X"84050871";
    when 16#00FC7# => romdata <= X"8C1A0C76";
    when 16#00FC8# => romdata <= X"881A0C78";
    when 16#00FC9# => romdata <= X"88130C78";
    when 16#00FCA# => romdata <= X"8C180C5D";
    when 16#00FCB# => romdata <= X"58795380";
    when 16#00FCC# => romdata <= X"7A2483E6";
    when 16#00FCD# => romdata <= X"3872822C";
    when 16#00FCE# => romdata <= X"81712B5C";
    when 16#00FCF# => romdata <= X"537A7C26";
    when 16#00FD0# => romdata <= X"8198387B";
    when 16#00FD1# => romdata <= X"7B065372";
    when 16#00FD2# => romdata <= X"82F13879";
    when 16#00FD3# => romdata <= X"FC068405";
    when 16#00FD4# => romdata <= X"5A7A1070";
    when 16#00FD5# => romdata <= X"7D06545B";
    when 16#00FD6# => romdata <= X"7282E038";
    when 16#00FD7# => romdata <= X"841A5AF1";
    when 16#00FD8# => romdata <= X"3988178C";
    when 16#00FD9# => romdata <= X"11085858";
    when 16#00FDA# => romdata <= X"76782E09";
    when 16#00FDB# => romdata <= X"8106FCC2";
    when 16#00FDC# => romdata <= X"38821A5A";
    when 16#00FDD# => romdata <= X"FDEC3978";
    when 16#00FDE# => romdata <= X"17798107";
    when 16#00FDF# => romdata <= X"84190C70";
    when 16#00FE0# => romdata <= X"81BA800C";
    when 16#00FE1# => romdata <= X"7081B9FC";
    when 16#00FE2# => romdata <= X"0C81B9F4";
    when 16#00FE3# => romdata <= X"0B8C120C";
    when 16#00FE4# => romdata <= X"8C110888";
    when 16#00FE5# => romdata <= X"120C7481";
    when 16#00FE6# => romdata <= X"0784120C";
    when 16#00FE7# => romdata <= X"74117571";
    when 16#00FE8# => romdata <= X"0C51537D";
    when 16#00FE9# => romdata <= X"5187B73F";
    when 16#00FEA# => romdata <= X"881754FC";
    when 16#00FEB# => romdata <= X"AC3981B9";
    when 16#00FEC# => romdata <= X"EC0B8405";
    when 16#00FED# => romdata <= X"087A545C";
    when 16#00FEE# => romdata <= X"798025FE";
    when 16#00FEF# => romdata <= X"F83882DA";
    when 16#00FF0# => romdata <= X"397A097C";
    when 16#00FF1# => romdata <= X"067081B9";
    when 16#00FF2# => romdata <= X"EC0B8405";
    when 16#00FF3# => romdata <= X"0C5C7A10";
    when 16#00FF4# => romdata <= X"5B7A7C26";
    when 16#00FF5# => romdata <= X"85387A85";
    when 16#00FF6# => romdata <= X"B83881B9";
    when 16#00FF7# => romdata <= X"EC0B8805";
    when 16#00FF8# => romdata <= X"08708412";
    when 16#00FF9# => romdata <= X"08FC0670";
    when 16#00FFA# => romdata <= X"7C317C72";
    when 16#00FFB# => romdata <= X"268F7225";
    when 16#00FFC# => romdata <= X"0757575C";
    when 16#00FFD# => romdata <= X"5D557280";
    when 16#00FFE# => romdata <= X"2E80DB38";
    when 16#00FFF# => romdata <= X"797A1681";
    when 16#01000# => romdata <= X"B9E4081B";
    when 16#01001# => romdata <= X"90115A55";
    when 16#01002# => romdata <= X"575B81B9";
    when 16#01003# => romdata <= X"E008FF2E";
    when 16#01004# => romdata <= X"8838A08F";
    when 16#01005# => romdata <= X"13E08006";
    when 16#01006# => romdata <= X"5776527D";
    when 16#01007# => romdata <= X"5186C03F";
    when 16#01008# => romdata <= X"B00854B0";
    when 16#01009# => romdata <= X"08FF2E90";
    when 16#0100A# => romdata <= X"38B00876";
    when 16#0100B# => romdata <= X"27829938";
    when 16#0100C# => romdata <= X"7481B9EC";
    when 16#0100D# => romdata <= X"2E829138";
    when 16#0100E# => romdata <= X"81B9EC0B";
    when 16#0100F# => romdata <= X"88050855";
    when 16#01010# => romdata <= X"841508FC";
    when 16#01011# => romdata <= X"06707A31";
    when 16#01012# => romdata <= X"7A72268F";
    when 16#01013# => romdata <= X"72250752";
    when 16#01014# => romdata <= X"55537283";
    when 16#01015# => romdata <= X"E6387479";
    when 16#01016# => romdata <= X"81078417";
    when 16#01017# => romdata <= X"0C791670";
    when 16#01018# => romdata <= X"81B9EC0B";
    when 16#01019# => romdata <= X"88050C75";
    when 16#0101A# => romdata <= X"81078412";
    when 16#0101B# => romdata <= X"0C547E52";
    when 16#0101C# => romdata <= X"5785EB3F";
    when 16#0101D# => romdata <= X"881754FA";
    when 16#0101E# => romdata <= X"E0397583";
    when 16#0101F# => romdata <= X"2A705454";
    when 16#01020# => romdata <= X"80742481";
    when 16#01021# => romdata <= X"9B387282";
    when 16#01022# => romdata <= X"2C81712B";
    when 16#01023# => romdata <= X"81B9F008";
    when 16#01024# => romdata <= X"077081B9";
    when 16#01025# => romdata <= X"EC0B8405";
    when 16#01026# => romdata <= X"0C751010";
    when 16#01027# => romdata <= X"1081B9EC";
    when 16#01028# => romdata <= X"05881108";
    when 16#01029# => romdata <= X"585A5D53";
    when 16#0102A# => romdata <= X"778C180C";
    when 16#0102B# => romdata <= X"7488180C";
    when 16#0102C# => romdata <= X"7688190C";
    when 16#0102D# => romdata <= X"768C160C";
    when 16#0102E# => romdata <= X"FCF33979";
    when 16#0102F# => romdata <= X"7A101010";
    when 16#01030# => romdata <= X"81B9EC05";
    when 16#01031# => romdata <= X"7057595D";
    when 16#01032# => romdata <= X"8C150857";
    when 16#01033# => romdata <= X"76752EA3";
    when 16#01034# => romdata <= X"38841708";
    when 16#01035# => romdata <= X"FC06707A";
    when 16#01036# => romdata <= X"31555673";
    when 16#01037# => romdata <= X"8F2483CA";
    when 16#01038# => romdata <= X"38738025";
    when 16#01039# => romdata <= X"8481388C";
    when 16#0103A# => romdata <= X"17085776";
    when 16#0103B# => romdata <= X"752E0981";
    when 16#0103C# => romdata <= X"06DF3888";
    when 16#0103D# => romdata <= X"15811B70";
    when 16#0103E# => romdata <= X"8306555B";
    when 16#0103F# => romdata <= X"5572C938";
    when 16#01040# => romdata <= X"7C830653";
    when 16#01041# => romdata <= X"72802EFD";
    when 16#01042# => romdata <= X"B838FF1D";
    when 16#01043# => romdata <= X"F819595D";
    when 16#01044# => romdata <= X"88180878";
    when 16#01045# => romdata <= X"2EEA38FD";
    when 16#01046# => romdata <= X"B539831A";
    when 16#01047# => romdata <= X"53FC9639";
    when 16#01048# => romdata <= X"83147082";
    when 16#01049# => romdata <= X"2C81712B";
    when 16#0104A# => romdata <= X"81B9F008";
    when 16#0104B# => romdata <= X"077081B9";
    when 16#0104C# => romdata <= X"EC0B8405";
    when 16#0104D# => romdata <= X"0C761010";
    when 16#0104E# => romdata <= X"1081B9EC";
    when 16#0104F# => romdata <= X"05881108";
    when 16#01050# => romdata <= X"595B5E51";
    when 16#01051# => romdata <= X"53FEE139";
    when 16#01052# => romdata <= X"81B9B008";
    when 16#01053# => romdata <= X"1758B008";
    when 16#01054# => romdata <= X"762E818D";
    when 16#01055# => romdata <= X"3881B9E0";
    when 16#01056# => romdata <= X"08FF2E83";
    when 16#01057# => romdata <= X"EC387376";
    when 16#01058# => romdata <= X"311881B9";
    when 16#01059# => romdata <= X"B00C7387";
    when 16#0105A# => romdata <= X"06705753";
    when 16#0105B# => romdata <= X"72802E88";
    when 16#0105C# => romdata <= X"38887331";
    when 16#0105D# => romdata <= X"70155556";
    when 16#0105E# => romdata <= X"76149FFF";
    when 16#0105F# => romdata <= X"06A08071";
    when 16#01060# => romdata <= X"31177054";
    when 16#01061# => romdata <= X"7F535753";
    when 16#01062# => romdata <= X"83D53FB0";
    when 16#01063# => romdata <= X"0853B008";
    when 16#01064# => romdata <= X"FF2E81A0";
    when 16#01065# => romdata <= X"3881B9B0";
    when 16#01066# => romdata <= X"08167081";
    when 16#01067# => romdata <= X"B9B00C74";
    when 16#01068# => romdata <= X"7581B9EC";
    when 16#01069# => romdata <= X"0B88050C";
    when 16#0106A# => romdata <= X"74763118";
    when 16#0106B# => romdata <= X"70810751";
    when 16#0106C# => romdata <= X"5556587B";
    when 16#0106D# => romdata <= X"81B9EC2E";
    when 16#0106E# => romdata <= X"839C3879";
    when 16#0106F# => romdata <= X"8F2682CB";
    when 16#01070# => romdata <= X"38810B84";
    when 16#01071# => romdata <= X"150C8415";
    when 16#01072# => romdata <= X"08FC0670";
    when 16#01073# => romdata <= X"7A317A72";
    when 16#01074# => romdata <= X"268F7225";
    when 16#01075# => romdata <= X"07525553";
    when 16#01076# => romdata <= X"72802EFC";
    when 16#01077# => romdata <= X"F93880DB";
    when 16#01078# => romdata <= X"39B0089F";
    when 16#01079# => romdata <= X"FF065372";
    when 16#0107A# => romdata <= X"FEEB3877";
    when 16#0107B# => romdata <= X"81B9B00C";
    when 16#0107C# => romdata <= X"81B9EC0B";
    when 16#0107D# => romdata <= X"8805087B";
    when 16#0107E# => romdata <= X"18810784";
    when 16#0107F# => romdata <= X"120C5581";
    when 16#01080# => romdata <= X"B9DC0878";
    when 16#01081# => romdata <= X"27863877";
    when 16#01082# => romdata <= X"81B9DC0C";
    when 16#01083# => romdata <= X"81B9D808";
    when 16#01084# => romdata <= X"7827FCAC";
    when 16#01085# => romdata <= X"387781B9";
    when 16#01086# => romdata <= X"D80C8415";
    when 16#01087# => romdata <= X"08FC0670";
    when 16#01088# => romdata <= X"7A317A72";
    when 16#01089# => romdata <= X"268F7225";
    when 16#0108A# => romdata <= X"07525553";
    when 16#0108B# => romdata <= X"72802EFC";
    when 16#0108C# => romdata <= X"A5388839";
    when 16#0108D# => romdata <= X"80745456";
    when 16#0108E# => romdata <= X"FEDB397D";
    when 16#0108F# => romdata <= X"51829F3F";
    when 16#01090# => romdata <= X"800BB00C";
    when 16#01091# => romdata <= X"8F3D0D04";
    when 16#01092# => romdata <= X"73538074";
    when 16#01093# => romdata <= X"24A93872";
    when 16#01094# => romdata <= X"822C8171";
    when 16#01095# => romdata <= X"2B81B9F0";
    when 16#01096# => romdata <= X"08077081";
    when 16#01097# => romdata <= X"B9EC0B84";
    when 16#01098# => romdata <= X"050C5D53";
    when 16#01099# => romdata <= X"778C180C";
    when 16#0109A# => romdata <= X"7488180C";
    when 16#0109B# => romdata <= X"7688190C";
    when 16#0109C# => romdata <= X"768C160C";
    when 16#0109D# => romdata <= X"F9B73983";
    when 16#0109E# => romdata <= X"1470822C";
    when 16#0109F# => romdata <= X"81712B81";
    when 16#010A0# => romdata <= X"B9F00807";
    when 16#010A1# => romdata <= X"7081B9EC";
    when 16#010A2# => romdata <= X"0B84050C";
    when 16#010A3# => romdata <= X"5E5153D4";
    when 16#010A4# => romdata <= X"397B7B06";
    when 16#010A5# => romdata <= X"5372FCA3";
    when 16#010A6# => romdata <= X"38841A7B";
    when 16#010A7# => romdata <= X"105C5AF1";
    when 16#010A8# => romdata <= X"39FF1A81";
    when 16#010A9# => romdata <= X"11515AF7";
    when 16#010AA# => romdata <= X"B9397817";
    when 16#010AB# => romdata <= X"79810784";
    when 16#010AC# => romdata <= X"190C8C18";
    when 16#010AD# => romdata <= X"08881908";
    when 16#010AE# => romdata <= X"718C120C";
    when 16#010AF# => romdata <= X"88120C59";
    when 16#010B0# => romdata <= X"7081BA80";
    when 16#010B1# => romdata <= X"0C7081B9";
    when 16#010B2# => romdata <= X"FC0C81B9";
    when 16#010B3# => romdata <= X"F40B8C12";
    when 16#010B4# => romdata <= X"0C8C1108";
    when 16#010B5# => romdata <= X"88120C74";
    when 16#010B6# => romdata <= X"81078412";
    when 16#010B7# => romdata <= X"0C741175";
    when 16#010B8# => romdata <= X"710C5153";
    when 16#010B9# => romdata <= X"F9BD3975";
    when 16#010BA# => romdata <= X"17841108";
    when 16#010BB# => romdata <= X"81078412";
    when 16#010BC# => romdata <= X"0C538C17";
    when 16#010BD# => romdata <= X"08881808";
    when 16#010BE# => romdata <= X"718C120C";
    when 16#010BF# => romdata <= X"88120C58";
    when 16#010C0# => romdata <= X"7D5180DA";
    when 16#010C1# => romdata <= X"3F881754";
    when 16#010C2# => romdata <= X"F5CF3972";
    when 16#010C3# => romdata <= X"84150CF4";
    when 16#010C4# => romdata <= X"1AF80670";
    when 16#010C5# => romdata <= X"841E0881";
    when 16#010C6# => romdata <= X"0607841E";
    when 16#010C7# => romdata <= X"0C701D54";
    when 16#010C8# => romdata <= X"5B850B84";
    when 16#010C9# => romdata <= X"140C850B";
    when 16#010CA# => romdata <= X"88140C8F";
    when 16#010CB# => romdata <= X"7B27FDCF";
    when 16#010CC# => romdata <= X"38881C52";
    when 16#010CD# => romdata <= X"7D518290";
    when 16#010CE# => romdata <= X"3F81B9EC";
    when 16#010CF# => romdata <= X"0B880508";
    when 16#010D0# => romdata <= X"81B9B008";
    when 16#010D1# => romdata <= X"5955FDB7";
    when 16#010D2# => romdata <= X"397781B9";
    when 16#010D3# => romdata <= X"B00C7381";
    when 16#010D4# => romdata <= X"B9E00CFC";
    when 16#010D5# => romdata <= X"91397284";
    when 16#010D6# => romdata <= X"150CFDA3";
    when 16#010D7# => romdata <= X"390404FD";
    when 16#010D8# => romdata <= X"3D0D800B";
    when 16#010D9# => romdata <= X"81D6840C";
    when 16#010DA# => romdata <= X"765186CB";
    when 16#010DB# => romdata <= X"3FB00853";
    when 16#010DC# => romdata <= X"B008FF2E";
    when 16#010DD# => romdata <= X"883872B0";
    when 16#010DE# => romdata <= X"0C853D0D";
    when 16#010DF# => romdata <= X"0481D684";
    when 16#010E0# => romdata <= X"08547380";
    when 16#010E1# => romdata <= X"2EF03875";
    when 16#010E2# => romdata <= X"74710C52";
    when 16#010E3# => romdata <= X"72B00C85";
    when 16#010E4# => romdata <= X"3D0D04FB";
    when 16#010E5# => romdata <= X"3D0D7770";
    when 16#010E6# => romdata <= X"5256C23F";
    when 16#010E7# => romdata <= X"81B9EC0B";
    when 16#010E8# => romdata <= X"88050884";
    when 16#010E9# => romdata <= X"1108FC06";
    when 16#010EA# => romdata <= X"707B319F";
    when 16#010EB# => romdata <= X"EF05E080";
    when 16#010EC# => romdata <= X"06E08005";
    when 16#010ED# => romdata <= X"565653A0";
    when 16#010EE# => romdata <= X"80742494";
    when 16#010EF# => romdata <= X"38805275";
    when 16#010F0# => romdata <= X"51FF9C3F";
    when 16#010F1# => romdata <= X"81B9F408";
    when 16#010F2# => romdata <= X"155372B0";
    when 16#010F3# => romdata <= X"082E8F38";
    when 16#010F4# => romdata <= X"7551FF8A";
    when 16#010F5# => romdata <= X"3F805372";
    when 16#010F6# => romdata <= X"B00C873D";
    when 16#010F7# => romdata <= X"0D047330";
    when 16#010F8# => romdata <= X"527551FE";
    when 16#010F9# => romdata <= X"FA3FB008";
    when 16#010FA# => romdata <= X"FF2EA838";
    when 16#010FB# => romdata <= X"81B9EC0B";
    when 16#010FC# => romdata <= X"88050875";
    when 16#010FD# => romdata <= X"75318107";
    when 16#010FE# => romdata <= X"84120C53";
    when 16#010FF# => romdata <= X"81B9B008";
    when 16#01100# => romdata <= X"743181B9";
    when 16#01101# => romdata <= X"B00C7551";
    when 16#01102# => romdata <= X"FED43F81";
    when 16#01103# => romdata <= X"0BB00C87";
    when 16#01104# => romdata <= X"3D0D0480";
    when 16#01105# => romdata <= X"527551FE";
    when 16#01106# => romdata <= X"C63F81B9";
    when 16#01107# => romdata <= X"EC0B8805";
    when 16#01108# => romdata <= X"08B00871";
    when 16#01109# => romdata <= X"3156538F";
    when 16#0110A# => romdata <= X"7525FFA4";
    when 16#0110B# => romdata <= X"38B00881";
    when 16#0110C# => romdata <= X"B9E00831";
    when 16#0110D# => romdata <= X"81B9B00C";
    when 16#0110E# => romdata <= X"74810784";
    when 16#0110F# => romdata <= X"140C7551";
    when 16#01110# => romdata <= X"FE9C3F80";
    when 16#01111# => romdata <= X"53FF9039";
    when 16#01112# => romdata <= X"F63D0D7C";
    when 16#01113# => romdata <= X"7E545B72";
    when 16#01114# => romdata <= X"802E8283";
    when 16#01115# => romdata <= X"387A51FE";
    when 16#01116# => romdata <= X"843FF813";
    when 16#01117# => romdata <= X"84110870";
    when 16#01118# => romdata <= X"FE067013";
    when 16#01119# => romdata <= X"841108FC";
    when 16#0111A# => romdata <= X"065D5859";
    when 16#0111B# => romdata <= X"545881B9";
    when 16#0111C# => romdata <= X"F408752E";
    when 16#0111D# => romdata <= X"82DE3878";
    when 16#0111E# => romdata <= X"84160C80";
    when 16#0111F# => romdata <= X"73810654";
    when 16#01120# => romdata <= X"5A727A2E";
    when 16#01121# => romdata <= X"81D53878";
    when 16#01122# => romdata <= X"15841108";
    when 16#01123# => romdata <= X"81065153";
    when 16#01124# => romdata <= X"72A03878";
    when 16#01125# => romdata <= X"17577981";
    when 16#01126# => romdata <= X"E6388815";
    when 16#01127# => romdata <= X"08537281";
    when 16#01128# => romdata <= X"B9F42E82";
    when 16#01129# => romdata <= X"F9388C15";
    when 16#0112A# => romdata <= X"08708C15";
    when 16#0112B# => romdata <= X"0C738812";
    when 16#0112C# => romdata <= X"0C567681";
    when 16#0112D# => romdata <= X"0784190C";
    when 16#0112E# => romdata <= X"76187771";
    when 16#0112F# => romdata <= X"0C537981";
    when 16#01130# => romdata <= X"913883FF";
    when 16#01131# => romdata <= X"772781C8";
    when 16#01132# => romdata <= X"3876892A";
    when 16#01133# => romdata <= X"77832A56";
    when 16#01134# => romdata <= X"5372802E";
    when 16#01135# => romdata <= X"BF387686";
    when 16#01136# => romdata <= X"2AB80555";
    when 16#01137# => romdata <= X"847327B4";
    when 16#01138# => romdata <= X"3880DB13";
    when 16#01139# => romdata <= X"55947327";
    when 16#0113A# => romdata <= X"AB38768C";
    when 16#0113B# => romdata <= X"2A80EE05";
    when 16#0113C# => romdata <= X"5580D473";
    when 16#0113D# => romdata <= X"279E3876";
    when 16#0113E# => romdata <= X"8F2A80F7";
    when 16#0113F# => romdata <= X"055582D4";
    when 16#01140# => romdata <= X"73279138";
    when 16#01141# => romdata <= X"76922A80";
    when 16#01142# => romdata <= X"FC05558A";
    when 16#01143# => romdata <= X"D4732784";
    when 16#01144# => romdata <= X"3880FE55";
    when 16#01145# => romdata <= X"74101010";
    when 16#01146# => romdata <= X"81B9EC05";
    when 16#01147# => romdata <= X"88110855";
    when 16#01148# => romdata <= X"5673762E";
    when 16#01149# => romdata <= X"82B33884";
    when 16#0114A# => romdata <= X"1408FC06";
    when 16#0114B# => romdata <= X"53767327";
    when 16#0114C# => romdata <= X"8D388814";
    when 16#0114D# => romdata <= X"08547376";
    when 16#0114E# => romdata <= X"2E098106";
    when 16#0114F# => romdata <= X"EA388C14";
    when 16#01150# => romdata <= X"08708C1A";
    when 16#01151# => romdata <= X"0C74881A";
    when 16#01152# => romdata <= X"0C788812";
    when 16#01153# => romdata <= X"0C56778C";
    when 16#01154# => romdata <= X"150C7A51";
    when 16#01155# => romdata <= X"FC883F8C";
    when 16#01156# => romdata <= X"3D0D0477";
    when 16#01157# => romdata <= X"08787131";
    when 16#01158# => romdata <= X"59770588";
    when 16#01159# => romdata <= X"19085457";
    when 16#0115A# => romdata <= X"7281B9F4";
    when 16#0115B# => romdata <= X"2E80E038";
    when 16#0115C# => romdata <= X"8C180870";
    when 16#0115D# => romdata <= X"8C150C73";
    when 16#0115E# => romdata <= X"88120C56";
    when 16#0115F# => romdata <= X"FE893988";
    when 16#01160# => romdata <= X"15088C16";
    when 16#01161# => romdata <= X"08708C13";
    when 16#01162# => romdata <= X"0C578817";
    when 16#01163# => romdata <= X"0CFEA339";
    when 16#01164# => romdata <= X"76832A70";
    when 16#01165# => romdata <= X"54558075";
    when 16#01166# => romdata <= X"24819838";
    when 16#01167# => romdata <= X"72822C81";
    when 16#01168# => romdata <= X"712B81B9";
    when 16#01169# => romdata <= X"F0080781";
    when 16#0116A# => romdata <= X"B9EC0B84";
    when 16#0116B# => romdata <= X"050C5374";
    when 16#0116C# => romdata <= X"10101081";
    when 16#0116D# => romdata <= X"B9EC0588";
    when 16#0116E# => romdata <= X"11085556";
    when 16#0116F# => romdata <= X"758C190C";
    when 16#01170# => romdata <= X"7388190C";
    when 16#01171# => romdata <= X"7788170C";
    when 16#01172# => romdata <= X"778C150C";
    when 16#01173# => romdata <= X"FF843981";
    when 16#01174# => romdata <= X"5AFDB439";
    when 16#01175# => romdata <= X"78177381";
    when 16#01176# => romdata <= X"06545772";
    when 16#01177# => romdata <= X"98387708";
    when 16#01178# => romdata <= X"78713159";
    when 16#01179# => romdata <= X"77058C19";
    when 16#0117A# => romdata <= X"08881A08";
    when 16#0117B# => romdata <= X"718C120C";
    when 16#0117C# => romdata <= X"88120C57";
    when 16#0117D# => romdata <= X"57768107";
    when 16#0117E# => romdata <= X"84190C77";
    when 16#0117F# => romdata <= X"81B9EC0B";
    when 16#01180# => romdata <= X"88050C81";
    when 16#01181# => romdata <= X"B9E80877";
    when 16#01182# => romdata <= X"26FEC738";
    when 16#01183# => romdata <= X"81B9E408";
    when 16#01184# => romdata <= X"527A51FA";
    when 16#01185# => romdata <= X"FE3F7A51";
    when 16#01186# => romdata <= X"FAC43FFE";
    when 16#01187# => romdata <= X"BA398178";
    when 16#01188# => romdata <= X"8C150C78";
    when 16#01189# => romdata <= X"88150C73";
    when 16#0118A# => romdata <= X"8C1A0C73";
    when 16#0118B# => romdata <= X"881A0C5A";
    when 16#0118C# => romdata <= X"FD803983";
    when 16#0118D# => romdata <= X"1570822C";
    when 16#0118E# => romdata <= X"81712B81";
    when 16#0118F# => romdata <= X"B9F00807";
    when 16#01190# => romdata <= X"81B9EC0B";
    when 16#01191# => romdata <= X"84050C51";
    when 16#01192# => romdata <= X"53741010";
    when 16#01193# => romdata <= X"1081B9EC";
    when 16#01194# => romdata <= X"05881108";
    when 16#01195# => romdata <= X"5556FEE4";
    when 16#01196# => romdata <= X"39745380";
    when 16#01197# => romdata <= X"7524A738";
    when 16#01198# => romdata <= X"72822C81";
    when 16#01199# => romdata <= X"712B81B9";
    when 16#0119A# => romdata <= X"F0080781";
    when 16#0119B# => romdata <= X"B9EC0B84";
    when 16#0119C# => romdata <= X"050C5375";
    when 16#0119D# => romdata <= X"8C190C73";
    when 16#0119E# => romdata <= X"88190C77";
    when 16#0119F# => romdata <= X"88170C77";
    when 16#011A0# => romdata <= X"8C150CFD";
    when 16#011A1# => romdata <= X"CD398315";
    when 16#011A2# => romdata <= X"70822C81";
    when 16#011A3# => romdata <= X"712B81B9";
    when 16#011A4# => romdata <= X"F0080781";
    when 16#011A5# => romdata <= X"B9EC0B84";
    when 16#011A6# => romdata <= X"050C5153";
    when 16#011A7# => romdata <= X"D639810B";
    when 16#011A8# => romdata <= X"B00C0480";
    when 16#011A9# => romdata <= X"3D0D7281";
    when 16#011AA# => romdata <= X"2E893880";
    when 16#011AB# => romdata <= X"0BB00C82";
    when 16#011AC# => romdata <= X"3D0D0473";
    when 16#011AD# => romdata <= X"51B23FFE";
    when 16#011AE# => romdata <= X"3D0D81D6";
    when 16#011AF# => romdata <= X"80085170";
    when 16#011B0# => romdata <= X"8A3881D6";
    when 16#011B1# => romdata <= X"887081D6";
    when 16#011B2# => romdata <= X"800C5170";
    when 16#011B3# => romdata <= X"75125252";
    when 16#011B4# => romdata <= X"FF537087";
    when 16#011B5# => romdata <= X"FB808026";
    when 16#011B6# => romdata <= X"88387081";
    when 16#011B7# => romdata <= X"D6800C71";
    when 16#011B8# => romdata <= X"5372B00C";
    when 16#011B9# => romdata <= X"843D0D04";
    when 16#011BA# => romdata <= X"00FF3900";
    when 16#011BB# => romdata <= X"00000000";
    when 16#011BC# => romdata <= X"00000000";
    when 16#011BD# => romdata <= X"00000000";
    when 16#011BE# => romdata <= X"00000000";
    when 16#011BF# => romdata <= X"00CAC5CA";
    when 16#011C0# => romdata <= X"C5C0C0C0";
    when 16#011C1# => romdata <= X"C0C0C0C0";
    when 16#011C2# => romdata <= X"C0C0C0CF";
    when 16#011C3# => romdata <= X"CFCFCF00";
    when 16#011C4# => romdata <= X"00000F0F";
    when 16#011C5# => romdata <= X"0F0F8F8F";
    when 16#011C6# => romdata <= X"CFCFCFCF";
    when 16#011C7# => romdata <= X"CFCF4F0F";
    when 16#011C8# => romdata <= X"0F0F0000";
    when 16#011C9# => romdata <= X"CFCFCFCF";
    when 16#011CA# => romdata <= X"0F0F0F0F";
    when 16#011CB# => romdata <= X"0F0F0F0F";
    when 16#011CC# => romdata <= X"0F0FFEFE";
    when 16#011CD# => romdata <= X"FEFC0000";
    when 16#011CE# => romdata <= X"CFCFCFCF";
    when 16#011CF# => romdata <= X"CFCFCFCF";
    when 16#011D0# => romdata <= X"CFCFCFCF";
    when 16#011D1# => romdata <= X"CFFFFF7E";
    when 16#011D2# => romdata <= X"7E000000";
    when 16#011D3# => romdata <= X"00000000";
    when 16#011D4# => romdata <= X"00000000";
    when 16#011D5# => romdata <= X"00000000";
    when 16#011D6# => romdata <= X"00003F3F";
    when 16#011D7# => romdata <= X"3F3F0101";
    when 16#011D8# => romdata <= X"01010101";
    when 16#011D9# => romdata <= X"01010101";
    when 16#011DA# => romdata <= X"3F3F3F3F";
    when 16#011DB# => romdata <= X"0000383C";
    when 16#011DC# => romdata <= X"3E3E3F3F";
    when 16#011DD# => romdata <= X"3F3B3B39";
    when 16#011DE# => romdata <= X"39383838";
    when 16#011DF# => romdata <= X"38383800";
    when 16#011E0# => romdata <= X"003F3F3F";
    when 16#011E1# => romdata <= X"3F383838";
    when 16#011E2# => romdata <= X"38383838";
    when 16#011E3# => romdata <= X"38383C3F";
    when 16#011E4# => romdata <= X"3F1F0F00";
    when 16#011E5# => romdata <= X"003F3F3F";
    when 16#011E6# => romdata <= X"3F030303";
    when 16#011E7# => romdata <= X"03030303";
    when 16#011E8# => romdata <= X"03033F3F";
    when 16#011E9# => romdata <= X"3F3E0000";
    when 16#011EA# => romdata <= X"00000000";
    when 16#011EB# => romdata <= X"00000000";
    when 16#011EC# => romdata <= X"00000000";
    when 16#011ED# => romdata <= X"00000000";
    when 16#011EE# => romdata <= X"00000000";
    when 16#011EF# => romdata <= X"00000000";
    when 16#011F0# => romdata <= X"00000000";
    when 16#011F1# => romdata <= X"00000000";
    when 16#011F2# => romdata <= X"00000000";
    when 16#011F3# => romdata <= X"00000000";
    when 16#011F4# => romdata <= X"00000000";
    when 16#011F5# => romdata <= X"00000000";
    when 16#011F6# => romdata <= X"00000000";
    when 16#011F7# => romdata <= X"00000000";
    when 16#011F8# => romdata <= X"00000000";
    when 16#011F9# => romdata <= X"00000000";
    when 16#011FA# => romdata <= X"00000000";
    when 16#011FB# => romdata <= X"00000000";
    when 16#011FC# => romdata <= X"00000000";
    when 16#011FD# => romdata <= X"00000000";
    when 16#011FE# => romdata <= X"00000000";
    when 16#011FF# => romdata <= X"00000000";
    when 16#01200# => romdata <= X"00000000";
    when 16#01201# => romdata <= X"00000000";
    when 16#01202# => romdata <= X"8080C0C0";
    when 16#01203# => romdata <= X"E0E06000";
    when 16#01204# => romdata <= X"00000000";
    when 16#01205# => romdata <= X"00000000";
    when 16#01206# => romdata <= X"00000000";
    when 16#01207# => romdata <= X"00000000";
    when 16#01208# => romdata <= X"00000000";
    when 16#01209# => romdata <= X"00000000";
    when 16#0120A# => romdata <= X"00000000";
    when 16#0120B# => romdata <= X"00000000";
    when 16#0120C# => romdata <= X"00000000";
    when 16#0120D# => romdata <= X"00000000";
    when 16#0120E# => romdata <= X"00000000";
    when 16#0120F# => romdata <= X"00000000";
    when 16#01210# => romdata <= X"00000000";
    when 16#01211# => romdata <= X"00000000";
    when 16#01212# => romdata <= X"00000000";
    when 16#01213# => romdata <= X"00000000";
    when 16#01214# => romdata <= X"00000000";
    when 16#01215# => romdata <= X"00000000";
    when 16#01216# => romdata <= X"00000000";
    when 16#01217# => romdata <= X"00000000";
    when 16#01218# => romdata <= X"806098EE";
    when 16#01219# => romdata <= X"77BBDDEC";
    when 16#0121A# => romdata <= X"EE6E0200";
    when 16#0121B# => romdata <= X"00000000";
    when 16#0121C# => romdata <= X"00E08080";
    when 16#0121D# => romdata <= X"E00000E0";
    when 16#0121E# => romdata <= X"A0A00000";
    when 16#0121F# => romdata <= X"E0000000";
    when 16#01220# => romdata <= X"00E0C000";
    when 16#01221# => romdata <= X"C0E00000";
    when 16#01222# => romdata <= X"E08080E0";
    when 16#01223# => romdata <= X"0000C020";
    when 16#01224# => romdata <= X"20C00000";
    when 16#01225# => romdata <= X"E0000000";
    when 16#01226# => romdata <= X"20E02000";
    when 16#01227# => romdata <= X"0020A060";
    when 16#01228# => romdata <= X"20000000";
    when 16#01229# => romdata <= X"00000000";
    when 16#0122A# => romdata <= X"00000000";
    when 16#0122B# => romdata <= X"00000000";
    when 16#0122C# => romdata <= X"00000000";
    when 16#0122D# => romdata <= X"00000000";
    when 16#0122E# => romdata <= X"00000000";
    when 16#0122F# => romdata <= X"00030007";
    when 16#01230# => romdata <= X"00070701";
    when 16#01231# => romdata <= X"00000000";
    when 16#01232# => romdata <= X"00000000";
    when 16#01233# => romdata <= X"00000300";
    when 16#01234# => romdata <= X"C0030000";
    when 16#01235# => romdata <= X"034242C0";
    when 16#01236# => romdata <= X"00C34242";
    when 16#01237# => romdata <= X"0000C380";
    when 16#01238# => romdata <= X"01C00340";
    when 16#01239# => romdata <= X"C04300C0";
    when 16#0123A# => romdata <= X"43408001";
    when 16#0123B# => romdata <= X"C20201C0";
    when 16#0123C# => romdata <= X"00C38202";
    when 16#0123D# => romdata <= X"80C00300";
    when 16#0123E# => romdata <= X"00C04342";
    when 16#0123F# => romdata <= X"8202C040";
    when 16#01240# => romdata <= X"40800000";
    when 16#01241# => romdata <= X"C0404000";
    when 16#01242# => romdata <= X"80404000";
    when 16#01243# => romdata <= X"00C04040";
    when 16#01244# => romdata <= X"8000C040";
    when 16#01245# => romdata <= X"4000C080";
    when 16#01246# => romdata <= X"00C00000";
    when 16#01247# => romdata <= X"00000000";
    when 16#01248# => romdata <= X"00000000";
    when 16#01249# => romdata <= X"00000000";
    when 16#0124A# => romdata <= X"00000000";
    when 16#0124B# => romdata <= X"00FF0000";
    when 16#0124C# => romdata <= X"0000C645";
    when 16#0124D# => romdata <= X"44800785";
    when 16#0124E# => romdata <= X"45408007";
    when 16#0124F# => romdata <= X"80424700";
    when 16#01250# => romdata <= X"80474000";
    when 16#01251# => romdata <= X"07C14344";
    when 16#01252# => romdata <= X"00C38404";
    when 16#01253# => romdata <= X"C30007C1";
    when 16#01254# => romdata <= X"42418700";
    when 16#01255# => romdata <= X"80404784";
    when 16#01256# => romdata <= X"04C34047";
    when 16#01257# => romdata <= X"8101C640";
    when 16#01258# => romdata <= X"40070505";
    when 16#01259# => romdata <= X"00040502";
    when 16#0125A# => romdata <= X"00000704";
    when 16#0125B# => romdata <= X"04030007";
    when 16#0125C# => romdata <= X"05050007";
    when 16#0125D# => romdata <= X"00020700";
    when 16#0125E# => romdata <= X"00000000";
    when 16#0125F# => romdata <= X"00000000";
    when 16#01260# => romdata <= X"00000000";
    when 16#01261# => romdata <= X"00000000";
    when 16#01262# => romdata <= X"0000FF00";
    when 16#01263# => romdata <= X"00000007";
    when 16#01264# => romdata <= X"01030500";
    when 16#01265# => romdata <= X"03040403";
    when 16#01266# => romdata <= X"00040502";
    when 16#01267# => romdata <= X"00040502";
    when 16#01268# => romdata <= X"00000705";
    when 16#01269# => romdata <= X"05000700";
    when 16#0126A# => romdata <= X"02070000";
    when 16#0126B# => romdata <= X"07040403";
    when 16#0126C# => romdata <= X"00030404";
    when 16#0126D# => romdata <= X"03000701";
    when 16#0126E# => romdata <= X"03050007";
    when 16#0126F# => romdata <= X"01010000";
    when 16#01270# => romdata <= X"00000000";
    when 16#01271# => romdata <= X"00000000";
    when 16#01272# => romdata <= X"00000000";
    when 16#01273# => romdata <= X"00000000";
    when 16#01274# => romdata <= X"00000000";
    when 16#01275# => romdata <= X"71756974";
    when 16#01276# => romdata <= X"00000000";
    when 16#01277# => romdata <= X"68656C70";
    when 16#01278# => romdata <= X"00000000";
    when 16#01279# => romdata <= X"73686F77";
    when 16#0127A# => romdata <= X"2042504D";
    when 16#0127B# => romdata <= X"20726567";
    when 16#0127C# => romdata <= X"69737465";
    when 16#0127D# => romdata <= X"72730000";
    when 16#0127E# => romdata <= X"62706D00";
    when 16#0127F# => romdata <= X"73686F77";
    when 16#01280# => romdata <= X"2F736574";
    when 16#01281# => romdata <= X"20646562";
    when 16#01282# => romdata <= X"75672072";
    when 16#01283# => romdata <= X"65676973";
    when 16#01284# => romdata <= X"74657273";
    when 16#01285# => romdata <= X"203C7365";
    when 16#01286# => romdata <= X"74206D6F";
    when 16#01287# => romdata <= X"64653E00";
    when 16#01288# => romdata <= X"64656275";
    when 16#01289# => romdata <= X"67000000";
    when 16#0128A# => romdata <= X"73797374";
    when 16#0128B# => romdata <= X"656D2072";
    when 16#0128C# => romdata <= X"65736574";
    when 16#0128D# => romdata <= X"00000000";
    when 16#0128E# => romdata <= X"72657365";
    when 16#0128F# => romdata <= X"74000000";
    when 16#01290# => romdata <= X"73686F77";
    when 16#01291# => romdata <= X"20646562";
    when 16#01292# => romdata <= X"75672062";
    when 16#01293# => romdata <= X"75666665";
    when 16#01294# => romdata <= X"72203C6C";
    when 16#01295# => romdata <= X"656E6774";
    when 16#01296# => romdata <= X"683E0000";
    when 16#01297# => romdata <= X"646F776E";
    when 16#01298# => romdata <= X"6C6F6164";
    when 16#01299# => romdata <= X"20646562";
    when 16#0129A# => romdata <= X"75672062";
    when 16#0129B# => romdata <= X"75666665";
    when 16#0129C# => romdata <= X"72202878";
    when 16#0129D# => romdata <= X"6D6F6465";
    when 16#0129E# => romdata <= X"6D290000";
    when 16#0129F# => romdata <= X"62726561";
    when 16#012A0# => romdata <= X"64000000";
    when 16#012A1# => romdata <= X"75706C6F";
    when 16#012A2# => romdata <= X"61642064";
    when 16#012A3# => romdata <= X"65627567";
    when 16#012A4# => romdata <= X"20627566";
    when 16#012A5# => romdata <= X"66657220";
    when 16#012A6# => romdata <= X"28786D6F";
    when 16#012A7# => romdata <= X"64656D29";
    when 16#012A8# => romdata <= X"00000000";
    when 16#012A9# => romdata <= X"62777269";
    when 16#012AA# => romdata <= X"74650000";
    when 16#012AB# => romdata <= X"636C6561";
    when 16#012AC# => romdata <= X"72206465";
    when 16#012AD# => romdata <= X"62756720";
    when 16#012AE# => romdata <= X"62756666";
    when 16#012AF# => romdata <= X"65720000";
    when 16#012B0# => romdata <= X"62636C65";
    when 16#012B1# => romdata <= X"61720000";
    when 16#012B2# => romdata <= X"73657475";
    when 16#012B3# => romdata <= X"70206368";
    when 16#012B4# => romdata <= X"616E6E65";
    when 16#012B5# => romdata <= X"6C207465";
    when 16#012B6# => romdata <= X"7374203C";
    when 16#012B7# => romdata <= X"70302E2E";
    when 16#012B8# => romdata <= X"353E0000";
    when 16#012B9# => romdata <= X"63687465";
    when 16#012BA# => romdata <= X"73740000";
    when 16#012BB# => romdata <= X"74657374";
    when 16#012BC# => romdata <= X"67656E65";
    when 16#012BD# => romdata <= X"7261746F";
    when 16#012BE# => romdata <= X"72203C73";
    when 16#012BF# => romdata <= X"63616C65";
    when 16#012C0# => romdata <= X"723E203C";
    when 16#012C1# => romdata <= X"72657374";
    when 16#012C2# => romdata <= X"6172743E";
    when 16#012C3# => romdata <= X"00000000";
    when 16#012C4# => romdata <= X"74657374";
    when 16#012C5# => romdata <= X"67656E00";
    when 16#012C6# => romdata <= X"3C6D7574";
    when 16#012C7# => romdata <= X"655F6E3E";
    when 16#012C8# => romdata <= X"203C7273";
    when 16#012C9# => romdata <= X"745F6E3E";
    when 16#012CA# => romdata <= X"203C6270";
    when 16#012CB# => romdata <= X"625F6E3E";
    when 16#012CC# => romdata <= X"203C6F73";
    when 16#012CD# => romdata <= X"72313E20";
    when 16#012CE# => romdata <= X"3C6F7372";
    when 16#012CF# => romdata <= X"323E0000";
    when 16#012D0# => romdata <= X"64616363";
    when 16#012D1# => romdata <= X"6F6E6600";
    when 16#012D2# => romdata <= X"636C6B20";
    when 16#012D3# => romdata <= X"3C73656C";
    when 16#012D4# => romdata <= X"6563743E";
    when 16#012D5# => romdata <= X"2030203D";
    when 16#012D6# => romdata <= X"20696E74";
    when 16#012D7# => romdata <= X"2C203120";
    when 16#012D8# => romdata <= X"3D206578";
    when 16#012D9# => romdata <= X"74000000";
    when 16#012DA# => romdata <= X"636C6B00";
    when 16#012DB# => romdata <= X"73686F77";
    when 16#012DC# => romdata <= X"20737973";
    when 16#012DD# => romdata <= X"74656D20";
    when 16#012DE# => romdata <= X"696E666F";
    when 16#012DF# => romdata <= X"203C7665";
    when 16#012E0# => romdata <= X"72626F73";
    when 16#012E1# => romdata <= X"653E0000";
    when 16#012E2# => romdata <= X"73797369";
    when 16#012E3# => romdata <= X"6E666F00";
    when 16#012E4# => romdata <= X"72756E6E";
    when 16#012E5# => romdata <= X"696E6720";
    when 16#012E6# => romdata <= X"6C696768";
    when 16#012E7# => romdata <= X"74000000";
    when 16#012E8# => romdata <= X"72756E00";
    when 16#012E9# => romdata <= X"72756E20";
    when 16#012EA# => romdata <= X"64697370";
    when 16#012EB# => romdata <= X"6C617920";
    when 16#012EC# => romdata <= X"74657374";
    when 16#012ED# => romdata <= X"2066756E";
    when 16#012EE# => romdata <= X"6374696F";
    when 16#012EF# => romdata <= X"6E000000";
    when 16#012F0# => romdata <= X"64697370";
    when 16#012F1# => romdata <= X"6C617900";
    when 16#012F2# => romdata <= X"73657420";
    when 16#012F3# => romdata <= X"6261636B";
    when 16#012F4# => romdata <= X"6C696768";
    when 16#012F5# => romdata <= X"74203C30";
    when 16#012F6# => romdata <= X"2E2E3331";
    when 16#012F7# => romdata <= X"3E000000";
    when 16#012F8# => romdata <= X"6261636B";
    when 16#012F9# => romdata <= X"00000000";
    when 16#012FA# => romdata <= X"73686F77";
    when 16#012FB# => romdata <= X"206C6F67";
    when 16#012FC# => romdata <= X"6F206F6E";
    when 16#012FD# => romdata <= X"20676C63";
    when 16#012FE# => romdata <= X"64000000";
    when 16#012FF# => romdata <= X"6C6F676F";
    when 16#01300# => romdata <= X"00000000";
    when 16#01301# => romdata <= X"63686563";
    when 16#01302# => romdata <= X"6B204932";
    when 16#01303# => romdata <= X"43206164";
    when 16#01304# => romdata <= X"64726573";
    when 16#01305# => romdata <= X"73000000";
    when 16#01306# => romdata <= X"69326300";
    when 16#01307# => romdata <= X"72656164";
    when 16#01308# => romdata <= X"20454550";
    when 16#01309# => romdata <= X"524F4D20";
    when 16#0130A# => romdata <= X"3C627573";
    when 16#0130B# => romdata <= X"3E203C69";
    when 16#0130C# => romdata <= X"32635F61";
    when 16#0130D# => romdata <= X"6464723E";
    when 16#0130E# => romdata <= X"203C6C65";
    when 16#0130F# => romdata <= X"6E677468";
    when 16#01310# => romdata <= X"3E000000";
    when 16#01311# => romdata <= X"65657072";
    when 16#01312# => romdata <= X"6F6D0000";
    when 16#01313# => romdata <= X"41444320";
    when 16#01314# => romdata <= X"72656769";
    when 16#01315# => romdata <= X"73746572";
    when 16#01316# => romdata <= X"20747261";
    when 16#01317# => romdata <= X"6E736665";
    when 16#01318# => romdata <= X"72203C76";
    when 16#01319# => romdata <= X"616C7565";
    when 16#0131A# => romdata <= X"3E000000";
    when 16#0131B# => romdata <= X"61747261";
    when 16#0131C# => romdata <= X"6E730000";
    when 16#0131D# => romdata <= X"696E6974";
    when 16#0131E# => romdata <= X"20414443";
    when 16#0131F# => romdata <= X"20726567";
    when 16#01320# => romdata <= X"69737465";
    when 16#01321# => romdata <= X"72730000";
    when 16#01322# => romdata <= X"61696E69";
    when 16#01323# => romdata <= X"74000000";
    when 16#01324# => romdata <= X"616C6961";
    when 16#01325# => romdata <= X"7320666F";
    when 16#01326# => romdata <= X"72207800";
    when 16#01327# => romdata <= X"6D656D00";
    when 16#01328# => romdata <= X"77726974";
    when 16#01329# => romdata <= X"6520776F";
    when 16#0132A# => romdata <= X"7264203C";
    when 16#0132B# => romdata <= X"61646472";
    when 16#0132C# => romdata <= X"3E203C6C";
    when 16#0132D# => romdata <= X"656E6774";
    when 16#0132E# => romdata <= X"683E203C";
    when 16#0132F# => romdata <= X"76616C75";
    when 16#01330# => romdata <= X"65287329";
    when 16#01331# => romdata <= X"3E000000";
    when 16#01332# => romdata <= X"776D656D";
    when 16#01333# => romdata <= X"00000000";
    when 16#01334# => romdata <= X"6558616D";
    when 16#01335# => romdata <= X"696E6520";
    when 16#01336# => romdata <= X"6D656D6F";
    when 16#01337# => romdata <= X"72790000";
    when 16#01338# => romdata <= X"636C6561";
    when 16#01339# => romdata <= X"72207363";
    when 16#0133A# => romdata <= X"7265656E";
    when 16#0133B# => romdata <= X"00000000";
    when 16#0133C# => romdata <= X"636C6561";
    when 16#0133D# => romdata <= X"72000000";
    when 16#0133E# => romdata <= X"0A307800";
    when 16#0133F# => romdata <= X"69326320";
    when 16#01340# => romdata <= X"464D430A";
    when 16#01341# => romdata <= X"00000000";
    when 16#01342# => romdata <= X"61646472";
    when 16#01343# => romdata <= X"6573733A";
    when 16#01344# => romdata <= X"20307800";
    when 16#01345# => romdata <= X"2020202D";
    when 16#01346# => romdata <= X"2D3E2020";
    when 16#01347# => romdata <= X"2041434B";
    when 16#01348# => romdata <= X"0A000000";
    when 16#01349# => romdata <= X"72656164";
    when 16#0134A# => romdata <= X"20646174";
    when 16#0134B# => romdata <= X"61202800";
    when 16#0134C# => romdata <= X"20627974";
    when 16#0134D# => romdata <= X"65732920";
    when 16#0134E# => romdata <= X"66726F6D";
    when 16#0134F# => romdata <= X"20493243";
    when 16#01350# => romdata <= X"2D616464";
    when 16#01351# => romdata <= X"72657373";
    when 16#01352# => romdata <= X"20307800";
    when 16#01353# => romdata <= X"0A0A0000";
    when 16#01354# => romdata <= X"6E6F6163";
    when 16#01355# => romdata <= X"6B200000";
    when 16#01356# => romdata <= X"6368726F";
    when 16#01357# => romdata <= X"6E74656C";
    when 16#01358# => romdata <= X"20726567";
    when 16#01359# => romdata <= X"20307800";
    when 16#0135A# => romdata <= X"3A203078";
    when 16#0135B# => romdata <= X"00000000";
    when 16#0135C# => romdata <= X"206E6163";
    when 16#0135D# => romdata <= X"6B000000";
    when 16#0135E# => romdata <= X"6572726F";
    when 16#0135F# => romdata <= X"7220286E";
    when 16#01360# => romdata <= X"61636B29";
    when 16#01361# => romdata <= X"0A000000";
    when 16#01362# => romdata <= X"6265616D";
    when 16#01363# => romdata <= X"20706F73";
    when 16#01364# => romdata <= X"6974696F";
    when 16#01365# => romdata <= X"6E206D6F";
    when 16#01366# => romdata <= X"6E69746F";
    when 16#01367# => romdata <= X"72207265";
    when 16#01368# => romdata <= X"67697374";
    when 16#01369# => romdata <= X"65727300";
    when 16#0136A# => romdata <= X"0A202020";
    when 16#0136B# => romdata <= X"20202020";
    when 16#0136C# => romdata <= X"20202020";
    when 16#0136D# => romdata <= X"20202020";
    when 16#0136E# => romdata <= X"20202020";
    when 16#0136F# => romdata <= X"20202020";
    when 16#01370# => romdata <= X"20636861";
    when 16#01371# => romdata <= X"6E6E656C";
    when 16#01372# => romdata <= X"20302020";
    when 16#01373# => romdata <= X"20636861";
    when 16#01374# => romdata <= X"6E6E656C";
    when 16#01375# => romdata <= X"20312020";
    when 16#01376# => romdata <= X"20636861";
    when 16#01377# => romdata <= X"6E6E656C";
    when 16#01378# => romdata <= X"20322020";
    when 16#01379# => romdata <= X"20636861";
    when 16#0137A# => romdata <= X"6E6E656C";
    when 16#0137B# => romdata <= X"20330000";
    when 16#0137C# => romdata <= X"0A202020";
    when 16#0137D# => romdata <= X"20202020";
    when 16#0137E# => romdata <= X"20202020";
    when 16#0137F# => romdata <= X"20202020";
    when 16#01380# => romdata <= X"20202020";
    when 16#01381# => romdata <= X"20202020";
    when 16#01382# => romdata <= X"202D2D2D";
    when 16#01383# => romdata <= X"2D20686F";
    when 16#01384# => romdata <= X"72697A6F";
    when 16#01385# => romdata <= X"6E74616C";
    when 16#01386# => romdata <= X"202D2D2D";
    when 16#01387# => romdata <= X"2D2D2020";
    when 16#01388# => romdata <= X"202D2D2D";
    when 16#01389# => romdata <= X"2D2D2D20";
    when 16#0138A# => romdata <= X"76657274";
    when 16#0138B# => romdata <= X"6963616C";
    when 16#0138C# => romdata <= X"202D2D2D";
    when 16#0138D# => romdata <= X"2D2D0000";
    when 16#0138E# => romdata <= X"0A736361";
    when 16#0138F# => romdata <= X"6C657220";
    when 16#01390# => romdata <= X"76616C75";
    when 16#01391# => romdata <= X"65732020";
    when 16#01392# => romdata <= X"20202020";
    when 16#01393# => romdata <= X"20202020";
    when 16#01394# => romdata <= X"20000000";
    when 16#01395# => romdata <= X"0A6E6F69";
    when 16#01396# => romdata <= X"73652063";
    when 16#01397# => romdata <= X"6F6D7065";
    when 16#01398# => romdata <= X"6E736174";
    when 16#01399# => romdata <= X"696F6E20";
    when 16#0139A# => romdata <= X"20202020";
    when 16#0139B# => romdata <= X"20000000";
    when 16#0139C# => romdata <= X"0A6D6561";
    when 16#0139D# => romdata <= X"73757265";
    when 16#0139E# => romdata <= X"6D656E74";
    when 16#0139F# => romdata <= X"20202020";
    when 16#013A0# => romdata <= X"20202020";
    when 16#013A1# => romdata <= X"20202020";
    when 16#013A2# => romdata <= X"20000000";
    when 16#013A3# => romdata <= X"0A73756D";
    when 16#013A4# => romdata <= X"20636861";
    when 16#013A5# => romdata <= X"6E6E656C";
    when 16#013A6# => romdata <= X"2020203A";
    when 16#013A7# => romdata <= X"20000000";
    when 16#013A8# => romdata <= X"0A706F73";
    when 16#013A9# => romdata <= X"6974696F";
    when 16#013AA# => romdata <= X"6E20636F";
    when 16#013AB# => romdata <= X"6D707574";
    when 16#013AC# => romdata <= X"6174696F";
    when 16#013AD# => romdata <= X"6E000000";
    when 16#013AE# => romdata <= X"0A202073";
    when 16#013AF# => romdata <= X"63616C65";
    when 16#013B0# => romdata <= X"72207661";
    when 16#013B1# => romdata <= X"6C756573";
    when 16#013B2# => romdata <= X"20202020";
    when 16#013B3# => romdata <= X"20202020";
    when 16#013B4# => romdata <= X"20000000";
    when 16#013B5# => romdata <= X"0A20206F";
    when 16#013B6# => romdata <= X"66667365";
    when 16#013B7# => romdata <= X"74202020";
    when 16#013B8# => romdata <= X"20202020";
    when 16#013B9# => romdata <= X"20202020";
    when 16#013BA# => romdata <= X"20202020";
    when 16#013BB# => romdata <= X"20000000";
    when 16#013BC# => romdata <= X"0A6F7574";
    when 16#013BD# => romdata <= X"70757420";
    when 16#013BE# => romdata <= X"73656C65";
    when 16#013BF# => romdata <= X"6374203A";
    when 16#013C0# => romdata <= X"20000000";
    when 16#013C1# => romdata <= X"6368616E";
    when 16#013C2# => romdata <= X"6E656C20";
    when 16#013C3# => romdata <= X"30000000";
    when 16#013C4# => romdata <= X"0A63616C";
    when 16#013C5# => romdata <= X"63207374";
    when 16#013C6# => romdata <= X"61746520";
    when 16#013C7# => romdata <= X"2020203A";
    when 16#013C8# => romdata <= X"20307800";
    when 16#013C9# => romdata <= X"0A202064";
    when 16#013CA# => romdata <= X"69766964";
    when 16#013CB# => romdata <= X"656E6420";
    when 16#013CC# => romdata <= X"63757474";
    when 16#013CD# => romdata <= X"65640000";
    when 16#013CE# => romdata <= X"0A20206E";
    when 16#013CF# => romdata <= X"6F697365";
    when 16#013D0# => romdata <= X"20636F6D";
    when 16#013D1# => romdata <= X"70656E73";
    when 16#013D2# => romdata <= X"6174696F";
    when 16#013D3# => romdata <= X"6E20746F";
    when 16#013D4# => romdata <= X"20626967";
    when 16#013D5# => romdata <= X"00000000";
    when 16#013D6# => romdata <= X"0A20206E";
    when 16#013D7# => romdata <= X"6F697365";
    when 16#013D8# => romdata <= X"2076616C";
    when 16#013D9# => romdata <= X"75652063";
    when 16#013DA# => romdata <= X"75747465";
    when 16#013DB# => romdata <= X"64000000";
    when 16#013DC# => romdata <= X"0A202073";
    when 16#013DD# => romdata <= X"756D2076";
    when 16#013DE# => romdata <= X"616C7565";
    when 16#013DF# => romdata <= X"20637574";
    when 16#013E0# => romdata <= X"74656400";
    when 16#013E1# => romdata <= X"76657274";
    when 16#013E2# => romdata <= X"6963616C";
    when 16#013E3# => romdata <= X"00000000";
    when 16#013E4# => romdata <= X"686F7269";
    when 16#013E5# => romdata <= X"7A6F6E74";
    when 16#013E6# => romdata <= X"616C0000";
    when 16#013E7# => romdata <= X"73756D00";
    when 16#013E8# => romdata <= X"6368616E";
    when 16#013E9# => romdata <= X"6E656C20";
    when 16#013EA# => romdata <= X"33000000";
    when 16#013EB# => romdata <= X"6368616E";
    when 16#013EC# => romdata <= X"6E656C20";
    when 16#013ED# => romdata <= X"32000000";
    when 16#013EE# => romdata <= X"6368616E";
    when 16#013EF# => romdata <= X"6E656C20";
    when 16#013F0# => romdata <= X"31000000";
    when 16#013F1# => romdata <= X"786D6F64";
    when 16#013F2# => romdata <= X"656D2074";
    when 16#013F3# => romdata <= X"72616E73";
    when 16#013F4# => romdata <= X"6D69742E";
    when 16#013F5# => romdata <= X"2E2E0A00";
    when 16#013F6# => romdata <= X"20627974";
    when 16#013F7# => romdata <= X"65732074";
    when 16#013F8# => romdata <= X"72616E73";
    when 16#013F9# => romdata <= X"6D697474";
    when 16#013FA# => romdata <= X"65640A00";
    when 16#013FB# => romdata <= X"63616E63";
    when 16#013FC# => romdata <= X"656C0A00";
    when 16#013FD# => romdata <= X"72657472";
    when 16#013FE# => romdata <= X"79206F75";
    when 16#013FF# => romdata <= X"740A0000";
    when 16#01400# => romdata <= X"786D6F64";
    when 16#01401# => romdata <= X"656D2072";
    when 16#01402# => romdata <= X"65636569";
    when 16#01403# => romdata <= X"76652E2E";
    when 16#01404# => romdata <= X"2E0A0000";
    when 16#01405# => romdata <= X"20627974";
    when 16#01406# => romdata <= X"65732072";
    when 16#01407# => romdata <= X"65636569";
    when 16#01408# => romdata <= X"7665640A";
    when 16#01409# => romdata <= X"00000000";
    when 16#0140A# => romdata <= X"72782062";
    when 16#0140B# => romdata <= X"75666665";
    when 16#0140C# => romdata <= X"72206675";
    when 16#0140D# => romdata <= X"6C6C0A00";
    when 16#0140E# => romdata <= X"74696D65";
    when 16#0140F# => romdata <= X"206F7574";
    when 16#01410# => romdata <= X"0A000000";
    when 16#01411# => romdata <= X"64656275";
    when 16#01412# => romdata <= X"67207265";
    when 16#01413# => romdata <= X"67697374";
    when 16#01414# => romdata <= X"65727300";
    when 16#01415# => romdata <= X"0A6D6F64";
    when 16#01416# => romdata <= X"65202020";
    when 16#01417# => romdata <= X"20202020";
    when 16#01418# => romdata <= X"203A2000";
    when 16#01419# => romdata <= X"0A616464";
    when 16#0141A# => romdata <= X"72657373";
    when 16#0141B# => romdata <= X"20302020";
    when 16#0141C# => romdata <= X"203A2030";
    when 16#0141D# => romdata <= X"78000000";
    when 16#0141E# => romdata <= X"0A616464";
    when 16#0141F# => romdata <= X"72657373";
    when 16#01420# => romdata <= X"20312020";
    when 16#01421# => romdata <= X"203A2030";
    when 16#01422# => romdata <= X"78000000";
    when 16#01423# => romdata <= X"0A627566";
    when 16#01424# => romdata <= X"66657220";
    when 16#01425# => romdata <= X"73697A65";
    when 16#01426# => romdata <= X"203A2000";
    when 16#01427# => romdata <= X"65787465";
    when 16#01428# => romdata <= X"726E616C";
    when 16#01429# => romdata <= X"20636C6F";
    when 16#0142A# => romdata <= X"636B2000";
    when 16#0142B# => romdata <= X"61637469";
    when 16#0142C# => romdata <= X"76650A00";
    when 16#0142D# => romdata <= X"4E4F5420";
    when 16#0142E# => romdata <= X"00000000";
    when 16#0142F# => romdata <= X"6265616D";
    when 16#01430# => romdata <= X"20706F73";
    when 16#01431# => romdata <= X"6974696F";
    when 16#01432# => romdata <= X"6E206D6F";
    when 16#01433# => romdata <= X"6E69746F";
    when 16#01434# => romdata <= X"72000000";
    when 16#01435# => romdata <= X"20286F6E";
    when 16#01436# => romdata <= X"2073696D";
    when 16#01437# => romdata <= X"290A0000";
    when 16#01438# => romdata <= X"0A636F6D";
    when 16#01439# => romdata <= X"70696C65";
    when 16#0143A# => romdata <= X"643A204A";
    when 16#0143B# => romdata <= X"756C2020";
    when 16#0143C# => romdata <= X"31203230";
    when 16#0143D# => romdata <= X"31312020";
    when 16#0143E# => romdata <= X"30393A30";
    when 16#0143F# => romdata <= X"353A3030";
    when 16#01440# => romdata <= X"00000000";
    when 16#01441# => romdata <= X"0A737973";
    when 16#01442# => romdata <= X"74656D20";
    when 16#01443# => romdata <= X"636C6F63";
    when 16#01444# => romdata <= X"6B3A2000";
    when 16#01445# => romdata <= X"204D487A";
    when 16#01446# => romdata <= X"0A000000";
    when 16#01447# => romdata <= X"44454255";
    when 16#01448# => romdata <= X"47204D4F";
    when 16#01449# => romdata <= X"44450000";
    when 16#0144A# => romdata <= X"204F4E0A";
    when 16#0144B# => romdata <= X"00000000";
    when 16#0144C# => romdata <= X"00000EF0";
    when 16#0144D# => romdata <= X"00000FDE";
    when 16#0144E# => romdata <= X"00000FD3";
    when 16#0144F# => romdata <= X"00000FC8";
    when 16#01450# => romdata <= X"00000FBD";
    when 16#01451# => romdata <= X"00000FB2";
    when 16#01452# => romdata <= X"00000FA7";
    when 16#01453# => romdata <= X"0187FC09";
    when 16#01454# => romdata <= X"026F0000";
    when 16#01455# => romdata <= X"0003FFF6";
    when 16#01456# => romdata <= X"00060000";
    when 16#01457# => romdata <= X"3E200000";
    when 16#01458# => romdata <= X"636F6D6D";
    when 16#01459# => romdata <= X"616E6420";
    when 16#0145A# => romdata <= X"6E6F7420";
    when 16#0145B# => romdata <= X"666F756E";
    when 16#0145C# => romdata <= X"642E0A00";
    when 16#0145D# => romdata <= X"73757070";
    when 16#0145E# => romdata <= X"6F727465";
    when 16#0145F# => romdata <= X"6420636F";
    when 16#01460# => romdata <= X"6D6D616E";
    when 16#01461# => romdata <= X"64733A0A";
    when 16#01462# => romdata <= X"0A000000";
    when 16#01463# => romdata <= X"202D2000";
    when 16#01464# => romdata <= X"76656E64";
    when 16#01465# => romdata <= X"6F723F20";
    when 16#01466# => romdata <= X"20000000";
    when 16#01467# => romdata <= X"67616973";
    when 16#01468# => romdata <= X"6C657220";
    when 16#01469# => romdata <= X"20000000";
    when 16#0146A# => romdata <= X"756E6B6E";
    when 16#0146B# => romdata <= X"6F776E20";
    when 16#0146C# => romdata <= X"64657669";
    when 16#0146D# => romdata <= X"63650000";
    when 16#0146E# => romdata <= X"485A4452";
    when 16#0146F# => romdata <= X"20202020";
    when 16#01470# => romdata <= X"20000000";
    when 16#01471# => romdata <= X"47656E65";
    when 16#01472# => romdata <= X"72616C20";
    when 16#01473# => romdata <= X"50757270";
    when 16#01474# => romdata <= X"6F736520";
    when 16#01475# => romdata <= X"492F4F20";
    when 16#01476# => romdata <= X"706F7274";
    when 16#01477# => romdata <= X"00000000";
    when 16#01478# => romdata <= X"56474120";
    when 16#01479# => romdata <= X"636F6E74";
    when 16#0147A# => romdata <= X"726F6C6C";
    when 16#0147B# => romdata <= X"65720000";
    when 16#0147C# => romdata <= X"4475616C";
    when 16#0147D# => romdata <= X"2D706F72";
    when 16#0147E# => romdata <= X"74204148";
    when 16#0147F# => romdata <= X"42205352";
    when 16#01480# => romdata <= X"414D206D";
    when 16#01481# => romdata <= X"6F64756C";
    when 16#01482# => romdata <= X"65000000";
    when 16#01483# => romdata <= X"64656275";
    when 16#01484# => romdata <= X"67206275";
    when 16#01485# => romdata <= X"66666572";
    when 16#01486# => romdata <= X"20636F6E";
    when 16#01487# => romdata <= X"74726F6C";
    when 16#01488# => romdata <= X"00000000";
    when 16#01489# => romdata <= X"74726967";
    when 16#0148A# => romdata <= X"67657220";
    when 16#0148B# => romdata <= X"67656E65";
    when 16#0148C# => romdata <= X"7261746F";
    when 16#0148D# => romdata <= X"72000000";
    when 16#0148E# => romdata <= X"64656275";
    when 16#0148F# => romdata <= X"6720636F";
    when 16#01490# => romdata <= X"6E736F6C";
    when 16#01491# => romdata <= X"65000000";
    when 16#01492# => romdata <= X"44434D20";
    when 16#01493# => romdata <= X"70686173";
    when 16#01494# => romdata <= X"65207368";
    when 16#01495# => romdata <= X"69667420";
    when 16#01496# => romdata <= X"636F6E74";
    when 16#01497# => romdata <= X"726F6C00";
    when 16#01498# => romdata <= X"5A505520";
    when 16#01499# => romdata <= X"4D656D6F";
    when 16#0149A# => romdata <= X"72792077";
    when 16#0149B# => romdata <= X"72617070";
    when 16#0149C# => romdata <= X"65720000";
    when 16#0149D# => romdata <= X"5A505520";
    when 16#0149E# => romdata <= X"41484220";
    when 16#0149F# => romdata <= X"57726170";
    when 16#014A0# => romdata <= X"70657200";
    when 16#014A1# => romdata <= X"4148422F";
    when 16#014A2# => romdata <= X"41504220";
    when 16#014A3# => romdata <= X"42726964";
    when 16#014A4# => romdata <= X"67650000";
    when 16#014A5# => romdata <= X"4D6F6475";
    when 16#014A6# => romdata <= X"6C617220";
    when 16#014A7# => romdata <= X"54696D65";
    when 16#014A8# => romdata <= X"7220556E";
    when 16#014A9# => romdata <= X"69740000";
    when 16#014AA# => romdata <= X"414D4241";
    when 16#014AB# => romdata <= X"20577261";
    when 16#014AC# => romdata <= X"70706572";
    when 16#014AD# => romdata <= X"20666F72";
    when 16#014AE# => romdata <= X"204F4320";
    when 16#014AF# => romdata <= X"4932432D";
    when 16#014B0# => romdata <= X"6D617374";
    when 16#014B1# => romdata <= X"65720000";
    when 16#014B2# => romdata <= X"47656E65";
    when 16#014B3# => romdata <= X"72696320";
    when 16#014B4# => romdata <= X"55415254";
    when 16#014B5# => romdata <= X"00000000";
    when 16#014B6# => romdata <= X"20206170";
    when 16#014B7# => romdata <= X"62736C76";
    when 16#014B8# => romdata <= X"00000000";
    when 16#014B9# => romdata <= X"76656E64";
    when 16#014BA# => romdata <= X"20307800";
    when 16#014BB# => romdata <= X"64657620";
    when 16#014BC# => romdata <= X"30780000";
    when 16#014BD# => romdata <= X"76657220";
    when 16#014BE# => romdata <= X"00000000";
    when 16#014BF# => romdata <= X"69727120";
    when 16#014C0# => romdata <= X"00000000";
    when 16#014C1# => romdata <= X"61646472";
    when 16#014C2# => romdata <= X"20307800";
    when 16#014C3# => romdata <= X"6168626D";
    when 16#014C4# => romdata <= X"73740000";
    when 16#014C5# => romdata <= X"61686273";
    when 16#014C6# => romdata <= X"6C760000";
    when 16#014C7# => romdata <= X"00002201";
    when 16#014C8# => romdata <= X"000022AC";
    when 16#014C9# => romdata <= X"000022A1";
    when 16#014CA# => romdata <= X"00002296";
    when 16#014CB# => romdata <= X"0000228B";
    when 16#014CC# => romdata <= X"00002280";
    when 16#014CD# => romdata <= X"00002275";
    when 16#014CE# => romdata <= X"0000226A";
    when 16#014CF# => romdata <= X"04580808";
    when 16#014D0# => romdata <= X"20FF0000";
    when 16#014D1# => romdata <= X"0000534C";
    when 16#014D2# => romdata <= X"0000542C";
    when 16#014D3# => romdata <= X"02010305";
    when 16#014D4# => romdata <= X"05070501";
    when 16#014D5# => romdata <= X"03030505";
    when 16#014D6# => romdata <= X"02030104";
    when 16#014D7# => romdata <= X"05050505";
    when 16#014D8# => romdata <= X"05050505";
    when 16#014D9# => romdata <= X"05050101";
    when 16#014DA# => romdata <= X"04050404";
    when 16#014DB# => romdata <= X"07050505";
    when 16#014DC# => romdata <= X"05050505";
    when 16#014DD# => romdata <= X"05030405";
    when 16#014DE# => romdata <= X"05050505";
    when 16#014DF# => romdata <= X"05050505";
    when 16#014E0# => romdata <= X"05050505";
    when 16#014E1# => romdata <= X"05050503";
    when 16#014E2# => romdata <= X"04030505";
    when 16#014E3# => romdata <= X"02050504";
    when 16#014E4# => romdata <= X"05050405";
    when 16#014E5# => romdata <= X"04010204";
    when 16#014E6# => romdata <= X"02050404";
    when 16#014E7# => romdata <= X"05050404";
    when 16#014E8# => romdata <= X"04040507";
    when 16#014E9# => romdata <= X"05040404";
    when 16#014EA# => romdata <= X"02040500";
    when 16#014EB# => romdata <= X"04050200";
    when 16#014EC# => romdata <= X"04080303";
    when 16#014ED# => romdata <= X"04090003";
    when 16#014EE# => romdata <= X"06000000";
    when 16#014EF# => romdata <= X"00020204";
    when 16#014F0# => romdata <= X"04040400";
    when 16#014F1# => romdata <= X"04060003";
    when 16#014F2# => romdata <= X"05000000";
    when 16#014F3# => romdata <= X"00000404";
    when 16#014F4# => romdata <= X"05050204";
    when 16#014F5# => romdata <= X"05060305";
    when 16#014F6# => romdata <= X"04030705";
    when 16#014F7# => romdata <= X"04050303";
    when 16#014F8# => romdata <= X"02040502";
    when 16#014F9# => romdata <= X"03020405";
    when 16#014FA# => romdata <= X"06060604";
    when 16#014FB# => romdata <= X"05050505";
    when 16#014FC# => romdata <= X"05050504";
    when 16#014FD# => romdata <= X"04040404";
    when 16#014FE# => romdata <= X"03030303";
    when 16#014FF# => romdata <= X"05050505";
    when 16#01500# => romdata <= X"05050505";
    when 16#01501# => romdata <= X"05040404";
    when 16#01502# => romdata <= X"04050404";
    when 16#01503# => romdata <= X"04040404";
    when 16#01504# => romdata <= X"04040503";
    when 16#01505# => romdata <= X"04040404";
    when 16#01506# => romdata <= X"02020303";
    when 16#01507# => romdata <= X"04040404";
    when 16#01508# => romdata <= X"04040405";
    when 16#01509# => romdata <= X"04040404";
    when 16#0150A# => romdata <= X"04030303";
    when 16#0150B# => romdata <= X"00005F07";
    when 16#0150C# => romdata <= X"0007741C";
    when 16#0150D# => romdata <= X"771C172E";
    when 16#0150E# => romdata <= X"6A3E2B3A";
    when 16#0150F# => romdata <= X"06493608";
    when 16#01510# => romdata <= X"36493036";
    when 16#01511# => romdata <= X"49597648";
    when 16#01512# => romdata <= X"073C4281";
    when 16#01513# => romdata <= X"81423C0A";
    when 16#01514# => romdata <= X"041F040A";
    when 16#01515# => romdata <= X"08083E08";
    when 16#01516# => romdata <= X"08806008";
    when 16#01517# => romdata <= X"080840C0";
    when 16#01518# => romdata <= X"300C033E";
    when 16#01519# => romdata <= X"4141413E";
    when 16#0151A# => romdata <= X"44427F40";
    when 16#0151B# => romdata <= X"40466151";
    when 16#0151C# => romdata <= X"49462241";
    when 16#0151D# => romdata <= X"49493618";
    when 16#0151E# => romdata <= X"14127F10";
    when 16#0151F# => romdata <= X"27454545";
    when 16#01520# => romdata <= X"393E4949";
    when 16#01521# => romdata <= X"49300101";
    when 16#01522# => romdata <= X"710D0336";
    when 16#01523# => romdata <= X"49494936";
    when 16#01524# => romdata <= X"06494929";
    when 16#01525# => romdata <= X"1E36D008";
    when 16#01526# => romdata <= X"14224114";
    when 16#01527# => romdata <= X"14141414";
    when 16#01528# => romdata <= X"41221408";
    when 16#01529# => romdata <= X"02510906";
    when 16#0152A# => romdata <= X"3C4299A5";
    when 16#0152B# => romdata <= X"BD421C7C";
    when 16#0152C# => romdata <= X"1211127C";
    when 16#0152D# => romdata <= X"7F494949";
    when 16#0152E# => romdata <= X"363E4141";
    when 16#0152F# => romdata <= X"41227F41";
    when 16#01530# => romdata <= X"41413E7F";
    when 16#01531# => romdata <= X"49494941";
    when 16#01532# => romdata <= X"7F090909";
    when 16#01533# => romdata <= X"013E4149";
    when 16#01534# => romdata <= X"497A7F08";
    when 16#01535# => romdata <= X"08087F41";
    when 16#01536# => romdata <= X"7F414041";
    when 16#01537# => romdata <= X"413F7F08";
    when 16#01538# => romdata <= X"1422417F";
    when 16#01539# => romdata <= X"40404040";
    when 16#0153A# => romdata <= X"7F060C06";
    when 16#0153B# => romdata <= X"7F7F0608";
    when 16#0153C# => romdata <= X"307F3E41";
    when 16#0153D# => romdata <= X"41413E7F";
    when 16#0153E# => romdata <= X"09090906";
    when 16#0153F# => romdata <= X"3E4161C1";
    when 16#01540# => romdata <= X"BE7F0919";
    when 16#01541# => romdata <= X"29462649";
    when 16#01542# => romdata <= X"49493201";
    when 16#01543# => romdata <= X"017F0101";
    when 16#01544# => romdata <= X"3F404040";
    when 16#01545# => romdata <= X"3F073840";
    when 16#01546# => romdata <= X"38071F60";
    when 16#01547# => romdata <= X"1F601F63";
    when 16#01548# => romdata <= X"14081463";
    when 16#01549# => romdata <= X"01067806";
    when 16#0154A# => romdata <= X"01615149";
    when 16#0154B# => romdata <= X"45437F41";
    when 16#0154C# => romdata <= X"41030C30";
    when 16#0154D# => romdata <= X"C041417F";
    when 16#0154E# => romdata <= X"04020102";
    when 16#0154F# => romdata <= X"04808080";
    when 16#01550# => romdata <= X"80800102";
    when 16#01551# => romdata <= X"20545454";
    when 16#01552# => romdata <= X"787F4444";
    when 16#01553# => romdata <= X"44383844";
    when 16#01554# => romdata <= X"44443844";
    when 16#01555# => romdata <= X"44447F38";
    when 16#01556# => romdata <= X"54545458";
    when 16#01557# => romdata <= X"087E0901";
    when 16#01558# => romdata <= X"18A4A4A4";
    when 16#01559# => romdata <= X"787F0404";
    when 16#0155A# => romdata <= X"787D807D";
    when 16#0155B# => romdata <= X"7F102844";
    when 16#0155C# => romdata <= X"3F407C04";
    when 16#0155D# => romdata <= X"7804787C";
    when 16#0155E# => romdata <= X"04047838";
    when 16#0155F# => romdata <= X"444438FC";
    when 16#01560# => romdata <= X"24242418";
    when 16#01561# => romdata <= X"18242424";
    when 16#01562# => romdata <= X"FC7C0804";
    when 16#01563# => romdata <= X"04485454";
    when 16#01564# => romdata <= X"24043F44";
    when 16#01565# => romdata <= X"403C4040";
    when 16#01566# => romdata <= X"7C1C2040";
    when 16#01567# => romdata <= X"201C1C60";
    when 16#01568# => romdata <= X"601C6060";
    when 16#01569# => romdata <= X"1C442810";
    when 16#0156A# => romdata <= X"28449CA0";
    when 16#0156B# => romdata <= X"601C6454";
    when 16#0156C# => romdata <= X"544C187E";
    when 16#0156D# => romdata <= X"8181FFFF";
    when 16#0156E# => romdata <= X"81817E18";
    when 16#0156F# => romdata <= X"18040810";
    when 16#01570# => romdata <= X"0C143E55";
    when 16#01571# => romdata <= X"55FF8181";
    when 16#01572# => romdata <= X"81FF8060";
    when 16#01573# => romdata <= X"80608060";
    when 16#01574# => romdata <= X"60600060";
    when 16#01575# => romdata <= X"60006060";
    when 16#01576# => romdata <= X"047F0414";
    when 16#01577# => romdata <= X"7F140201";
    when 16#01578# => romdata <= X"01024629";
    when 16#01579# => romdata <= X"1608344A";
    when 16#0157A# => romdata <= X"31483000";
    when 16#0157B# => romdata <= X"18243E41";
    when 16#0157C# => romdata <= X"227F4941";
    when 16#0157D# => romdata <= X"03040403";
    when 16#0157E# => romdata <= X"03040304";
    when 16#0157F# => romdata <= X"04030403";
    when 16#01580# => romdata <= X"183C3C18";
    when 16#01581# => romdata <= X"08080808";
    when 16#01582# => romdata <= X"03010203";
    when 16#01583# => romdata <= X"020E020E";
    when 16#01584# => romdata <= X"060E0048";
    when 16#01585# => romdata <= X"30384438";
    when 16#01586# => romdata <= X"54483844";
    when 16#01587# => romdata <= X"FE44487E";
    when 16#01588# => romdata <= X"49014438";
    when 16#01589# => romdata <= X"28384403";
    when 16#0158A# => romdata <= X"147C1403";
    when 16#0158B# => romdata <= X"E7E74E55";
    when 16#0158C# => romdata <= X"55390101";
    when 16#0158D# => romdata <= X"0001011C";
    when 16#0158E# => romdata <= X"2A555522";
    when 16#0158F# => romdata <= X"1C1D151E";
    when 16#01590# => romdata <= X"18240018";
    when 16#01591# => romdata <= X"24080808";
    when 16#01592# => romdata <= X"18080808";
    when 16#01593# => romdata <= X"3C42BD95";
    when 16#01594# => romdata <= X"A9423C01";
    when 16#01595# => romdata <= X"01010101";
    when 16#01596# => romdata <= X"06090906";
    when 16#01597# => romdata <= X"44445F44";
    when 16#01598# => romdata <= X"44191512";
    when 16#01599# => romdata <= X"15150A02";
    when 16#0159A# => romdata <= X"01FC2020";
    when 16#0159B# => romdata <= X"1C0E7F01";
    when 16#0159C# => romdata <= X"7F011818";
    when 16#0159D# => romdata <= X"00804002";
    when 16#0159E# => romdata <= X"1F060909";
    when 16#0159F# => romdata <= X"06241800";
    when 16#015A0# => romdata <= X"2418824F";
    when 16#015A1# => romdata <= X"304C62F1";
    when 16#015A2# => romdata <= X"824F300C";
    when 16#015A3# => romdata <= X"D2B1955F";
    when 16#015A4# => romdata <= X"304C62F1";
    when 16#015A5# => romdata <= X"30484520";
    when 16#015A6# => romdata <= X"60392E38";
    when 16#015A7# => romdata <= X"6060382E";
    when 16#015A8# => romdata <= X"3960701D";
    when 16#015A9# => romdata <= X"131D7072";
    when 16#015AA# => romdata <= X"1D121E71";
    when 16#015AB# => romdata <= X"701D121D";
    when 16#015AC# => romdata <= X"70603B25";
    when 16#015AD# => romdata <= X"3B607E11";
    when 16#015AE# => romdata <= X"7F49411E";
    when 16#015AF# => romdata <= X"2161927C";
    when 16#015B0# => romdata <= X"5556447C";
    when 16#015B1# => romdata <= X"5655447C";
    when 16#015B2# => romdata <= X"5655467D";
    when 16#015B3# => romdata <= X"54544545";
    when 16#015B4# => romdata <= X"7E44447E";
    when 16#015B5# => romdata <= X"45467D46";
    when 16#015B6# => romdata <= X"457C4508";
    when 16#015B7# => romdata <= X"7F49413E";
    when 16#015B8# => romdata <= X"7E091222";
    when 16#015B9# => romdata <= X"7D384546";
    when 16#015BA# => romdata <= X"44383844";
    when 16#015BB# => romdata <= X"46453838";
    when 16#015BC# => romdata <= X"46454638";
    when 16#015BD# => romdata <= X"3A454546";
    when 16#015BE# => romdata <= X"39384544";
    when 16#015BF# => romdata <= X"45382214";
    when 16#015C0# => romdata <= X"081422BC";
    when 16#015C1# => romdata <= X"625A463D";
    when 16#015C2# => romdata <= X"3C41423C";
    when 16#015C3# => romdata <= X"3C42413C";
    when 16#015C4# => romdata <= X"3C42413E";
    when 16#015C5# => romdata <= X"3D40403D";
    when 16#015C6# => romdata <= X"0608F209";
    when 16#015C7# => romdata <= X"067F2222";
    when 16#015C8# => romdata <= X"1CFE0989";
    when 16#015C9# => romdata <= X"76205556";
    when 16#015CA# => romdata <= X"78205655";
    when 16#015CB# => romdata <= X"78225555";
    when 16#015CC# => romdata <= X"7A235556";
    when 16#015CD# => romdata <= X"7B205554";
    when 16#015CE# => romdata <= X"79275557";
    when 16#015CF# => romdata <= X"78205438";
    when 16#015D0# => romdata <= X"54483844";
    when 16#015D1# => romdata <= X"C4385556";
    when 16#015D2# => romdata <= X"58385655";
    when 16#015D3# => romdata <= X"583A5555";
    when 16#015D4# => romdata <= X"5A395454";
    when 16#015D5# => romdata <= X"59017A7A";
    when 16#015D6# => romdata <= X"01027902";
    when 16#015D7# => romdata <= X"02780260";
    when 16#015D8# => romdata <= X"91927C7B";
    when 16#015D9# => romdata <= X"090A7338";
    when 16#015DA# => romdata <= X"45463838";
    when 16#015DB# => romdata <= X"4645383A";
    when 16#015DC# => romdata <= X"45453A3B";
    when 16#015DD# => romdata <= X"45463B39";
    when 16#015DE# => romdata <= X"44443908";
    when 16#015DF# => romdata <= X"082A0808";
    when 16#015E0# => romdata <= X"B8644C3A";
    when 16#015E1# => romdata <= X"3C41427C";
    when 16#015E2# => romdata <= X"3C42417C";
    when 16#015E3# => romdata <= X"3A41417A";
    when 16#015E4# => romdata <= X"3D40407D";
    when 16#015E5# => romdata <= X"986219FF";
    when 16#015E6# => romdata <= X"423C9A60";
    when 16#015E7# => romdata <= X"1A000000";
    when 16#015E8# => romdata <= X"30622020";
    when 16#015E9# => romdata <= X"20202020";
    when 16#015EA# => romdata <= X"20202020";
    when 16#015EB# => romdata <= X"20202020";
    when 16#015EC# => romdata <= X"20202020";
    when 16#015ED# => romdata <= X"20202020";
    when 16#015EE# => romdata <= X"20202020";
    when 16#015EF# => romdata <= X"20202020";
    when 16#015F0# => romdata <= X"20200000";
    when 16#015F1# => romdata <= X"20202020";
    when 16#015F2# => romdata <= X"20202020";
    when 16#015F3# => romdata <= X"00000000";
    when 16#015F4# => romdata <= X"00202020";
    when 16#015F5# => romdata <= X"20202020";
    when 16#015F6# => romdata <= X"20202828";
    when 16#015F7# => romdata <= X"28282820";
    when 16#015F8# => romdata <= X"20202020";
    when 16#015F9# => romdata <= X"20202020";
    when 16#015FA# => romdata <= X"20202020";
    when 16#015FB# => romdata <= X"20202020";
    when 16#015FC# => romdata <= X"20881010";
    when 16#015FD# => romdata <= X"10101010";
    when 16#015FE# => romdata <= X"10101010";
    when 16#015FF# => romdata <= X"10101010";
    when 16#01600# => romdata <= X"10040404";
    when 16#01601# => romdata <= X"04040404";
    when 16#01602# => romdata <= X"04040410";
    when 16#01603# => romdata <= X"10101010";
    when 16#01604# => romdata <= X"10104141";
    when 16#01605# => romdata <= X"41414141";
    when 16#01606# => romdata <= X"01010101";
    when 16#01607# => romdata <= X"01010101";
    when 16#01608# => romdata <= X"01010101";
    when 16#01609# => romdata <= X"01010101";
    when 16#0160A# => romdata <= X"01010101";
    when 16#0160B# => romdata <= X"10101010";
    when 16#0160C# => romdata <= X"10104242";
    when 16#0160D# => romdata <= X"42424242";
    when 16#0160E# => romdata <= X"02020202";
    when 16#0160F# => romdata <= X"02020202";
    when 16#01610# => romdata <= X"02020202";
    when 16#01611# => romdata <= X"02020202";
    when 16#01612# => romdata <= X"02020202";
    when 16#01613# => romdata <= X"10101010";
    when 16#01614# => romdata <= X"20000000";
    when 16#01615# => romdata <= X"00000000";
    when 16#01616# => romdata <= X"00000000";
    when 16#01617# => romdata <= X"00000000";
    when 16#01618# => romdata <= X"00000000";
    when 16#01619# => romdata <= X"00000000";
    when 16#0161A# => romdata <= X"00000000";
    when 16#0161B# => romdata <= X"00000000";
    when 16#0161C# => romdata <= X"00000000";
    when 16#0161D# => romdata <= X"00000000";
    when 16#0161E# => romdata <= X"00000000";
    when 16#0161F# => romdata <= X"00000000";
    when 16#01620# => romdata <= X"00000000";
    when 16#01621# => romdata <= X"00000000";
    when 16#01622# => romdata <= X"00000000";
    when 16#01623# => romdata <= X"00000000";
    when 16#01624# => romdata <= X"00000000";
    when 16#01625# => romdata <= X"00000000";
    when 16#01626# => romdata <= X"00000000";
    when 16#01627# => romdata <= X"00000000";
    when 16#01628# => romdata <= X"00000000";
    when 16#01629# => romdata <= X"00000000";
    when 16#0162A# => romdata <= X"00000000";
    when 16#0162B# => romdata <= X"00000000";
    when 16#0162C# => romdata <= X"00000000";
    when 16#0162D# => romdata <= X"00000000";
    when 16#0162E# => romdata <= X"00000000";
    when 16#0162F# => romdata <= X"00000000";
    when 16#01630# => romdata <= X"00000000";
    when 16#01631# => romdata <= X"00000000";
    when 16#01632# => romdata <= X"00000000";
    when 16#01633# => romdata <= X"00000000";
    when 16#01634# => romdata <= X"00000000";
    when 16#01635# => romdata <= X"43000000";
    when 16#01636# => romdata <= X"00000000";
    when 16#01637# => romdata <= X"80000C00";
    when 16#01638# => romdata <= X"80000B00";
    when 16#01639# => romdata <= X"80000800";
    when 16#0163A# => romdata <= X"00000000";
    when 16#0163B# => romdata <= X"FF000000";
    when 16#0163C# => romdata <= X"00000000";
    when 16#0163D# => romdata <= X"00000000";
    when 16#0163E# => romdata <= X"00FFFFFF";
    when 16#0163F# => romdata <= X"FF00FFFF";
    when 16#01640# => romdata <= X"FFFF00FF";
    when 16#01641# => romdata <= X"FFFFFF00";
    when 16#01642# => romdata <= X"00000000";
    when 16#01643# => romdata <= X"00000000";
    when 16#01644# => romdata <= X"80000A00";
    when 16#01645# => romdata <= X"80000700";
    when 16#01646# => romdata <= X"80000600";
    when 16#01647# => romdata <= X"80000400";
    when 16#01648# => romdata <= X"80000200";
    when 16#01649# => romdata <= X"80000100";
    when 16#0164A# => romdata <= X"80000004";
    when 16#0164B# => romdata <= X"80000000";
    when 16#0164C# => romdata <= X"00005934";
    when 16#0164D# => romdata <= X"00000000";
    when 16#0164E# => romdata <= X"00005B9C";
    when 16#0164F# => romdata <= X"00005BF8";
    when 16#01650# => romdata <= X"00005C54";
    when 16#01651# => romdata <= X"00000000";
    when 16#01652# => romdata <= X"00000000";
    when 16#01653# => romdata <= X"00000000";
    when 16#01654# => romdata <= X"00000000";
    when 16#01655# => romdata <= X"00000000";
    when 16#01656# => romdata <= X"00000000";
    when 16#01657# => romdata <= X"00000000";
    when 16#01658# => romdata <= X"00000000";
    when 16#01659# => romdata <= X"00000000";
    when 16#0165A# => romdata <= X"000058D4";
    when 16#0165B# => romdata <= X"00000000";
    when 16#0165C# => romdata <= X"00000000";
    when 16#0165D# => romdata <= X"00000000";
    when 16#0165E# => romdata <= X"00000000";
    when 16#0165F# => romdata <= X"00000000";
    when 16#01660# => romdata <= X"00000000";
    when 16#01661# => romdata <= X"00000000";
    when 16#01662# => romdata <= X"00000000";
    when 16#01663# => romdata <= X"00000000";
    when 16#01664# => romdata <= X"00000000";
    when 16#01665# => romdata <= X"00000000";
    when 16#01666# => romdata <= X"00000000";
    when 16#01667# => romdata <= X"00000000";
    when 16#01668# => romdata <= X"00000000";
    when 16#01669# => romdata <= X"00000000";
    when 16#0166A# => romdata <= X"00000000";
    when 16#0166B# => romdata <= X"00000000";
    when 16#0166C# => romdata <= X"00000000";
    when 16#0166D# => romdata <= X"00000000";
    when 16#0166E# => romdata <= X"00000000";
    when 16#0166F# => romdata <= X"00000000";
    when 16#01670# => romdata <= X"00000000";
    when 16#01671# => romdata <= X"00000000";
    when 16#01672# => romdata <= X"00000000";
    when 16#01673# => romdata <= X"00000000";
    when 16#01674# => romdata <= X"00000000";
    when 16#01675# => romdata <= X"00000000";
    when 16#01676# => romdata <= X"00000000";
    when 16#01677# => romdata <= X"00000001";
    when 16#01678# => romdata <= X"330EABCD";
    when 16#01679# => romdata <= X"1234E66D";
    when 16#0167A# => romdata <= X"DEEC0005";
    when 16#0167B# => romdata <= X"000B0000";
    when 16#0167C# => romdata <= X"00000000";
    when 16#0167D# => romdata <= X"00000000";
    when 16#0167E# => romdata <= X"00000000";
    when 16#0167F# => romdata <= X"00000000";
    when 16#01680# => romdata <= X"00000000";
    when 16#01681# => romdata <= X"00000000";
    when 16#01682# => romdata <= X"00000000";
    when 16#01683# => romdata <= X"00000000";
    when 16#01684# => romdata <= X"00000000";
    when 16#01685# => romdata <= X"00000000";
    when 16#01686# => romdata <= X"00000000";
    when 16#01687# => romdata <= X"00000000";
    when 16#01688# => romdata <= X"00000000";
    when 16#01689# => romdata <= X"00000000";
    when 16#0168A# => romdata <= X"00000000";
    when 16#0168B# => romdata <= X"00000000";
    when 16#0168C# => romdata <= X"00000000";
    when 16#0168D# => romdata <= X"00000000";
    when 16#0168E# => romdata <= X"00000000";
    when 16#0168F# => romdata <= X"00000000";
    when 16#01690# => romdata <= X"00000000";
    when 16#01691# => romdata <= X"00000000";
    when 16#01692# => romdata <= X"00000000";
    when 16#01693# => romdata <= X"00000000";
    when 16#01694# => romdata <= X"00000000";
    when 16#01695# => romdata <= X"00000000";
    when 16#01696# => romdata <= X"00000000";
    when 16#01697# => romdata <= X"00000000";
    when 16#01698# => romdata <= X"00000000";
    when 16#01699# => romdata <= X"00000000";
    when 16#0169A# => romdata <= X"00000000";
    when 16#0169B# => romdata <= X"00000000";
    when 16#0169C# => romdata <= X"00000000";
    when 16#0169D# => romdata <= X"00000000";
    when 16#0169E# => romdata <= X"00000000";
    when 16#0169F# => romdata <= X"00000000";
    when 16#016A0# => romdata <= X"00000000";
    when 16#016A1# => romdata <= X"00000000";
    when 16#016A2# => romdata <= X"00000000";
    when 16#016A3# => romdata <= X"00000000";
    when 16#016A4# => romdata <= X"00000000";
    when 16#016A5# => romdata <= X"00000000";
    when 16#016A6# => romdata <= X"00000000";
    when 16#016A7# => romdata <= X"00000000";
    when 16#016A8# => romdata <= X"00000000";
    when 16#016A9# => romdata <= X"00000000";
    when 16#016AA# => romdata <= X"00000000";
    when 16#016AB# => romdata <= X"00000000";
    when 16#016AC# => romdata <= X"00000000";
    when 16#016AD# => romdata <= X"00000000";
    when 16#016AE# => romdata <= X"00000000";
    when 16#016AF# => romdata <= X"00000000";
    when 16#016B0# => romdata <= X"00000000";
    when 16#016B1# => romdata <= X"00000000";
    when 16#016B2# => romdata <= X"00000000";
    when 16#016B3# => romdata <= X"00000000";
    when 16#016B4# => romdata <= X"00000000";
    when 16#016B5# => romdata <= X"00000000";
    when 16#016B6# => romdata <= X"00000000";
    when 16#016B7# => romdata <= X"00000000";
    when 16#016B8# => romdata <= X"00000000";
    when 16#016B9# => romdata <= X"00000000";
    when 16#016BA# => romdata <= X"00000000";
    when 16#016BB# => romdata <= X"00000000";
    when 16#016BC# => romdata <= X"00000000";
    when 16#016BD# => romdata <= X"00000000";
    when 16#016BE# => romdata <= X"00000000";
    when 16#016BF# => romdata <= X"00000000";
    when 16#016C0# => romdata <= X"00000000";
    when 16#016C1# => romdata <= X"00000000";
    when 16#016C2# => romdata <= X"00000000";
    when 16#016C3# => romdata <= X"00000000";
    when 16#016C4# => romdata <= X"00000000";
    when 16#016C5# => romdata <= X"00000000";
    when 16#016C6# => romdata <= X"00000000";
    when 16#016C7# => romdata <= X"00000000";
    when 16#016C8# => romdata <= X"00000000";
    when 16#016C9# => romdata <= X"00000000";
    when 16#016CA# => romdata <= X"00000000";
    when 16#016CB# => romdata <= X"00000000";
    when 16#016CC# => romdata <= X"00000000";
    when 16#016CD# => romdata <= X"00000000";
    when 16#016CE# => romdata <= X"00000000";
    when 16#016CF# => romdata <= X"00000000";
    when 16#016D0# => romdata <= X"00000000";
    when 16#016D1# => romdata <= X"00000000";
    when 16#016D2# => romdata <= X"00000000";
    when 16#016D3# => romdata <= X"00000000";
    when 16#016D4# => romdata <= X"00000000";
    when 16#016D5# => romdata <= X"00000000";
    when 16#016D6# => romdata <= X"00000000";
    when 16#016D7# => romdata <= X"00000000";
    when 16#016D8# => romdata <= X"00000000";
    when 16#016D9# => romdata <= X"00000000";
    when 16#016DA# => romdata <= X"00000000";
    when 16#016DB# => romdata <= X"00000000";
    when 16#016DC# => romdata <= X"00000000";
    when 16#016DD# => romdata <= X"00000000";
    when 16#016DE# => romdata <= X"00000000";
    when 16#016DF# => romdata <= X"00000000";
    when 16#016E0# => romdata <= X"00000000";
    when 16#016E1# => romdata <= X"00000000";
    when 16#016E2# => romdata <= X"00000000";
    when 16#016E3# => romdata <= X"00000000";
    when 16#016E4# => romdata <= X"00000000";
    when 16#016E5# => romdata <= X"00000000";
    when 16#016E6# => romdata <= X"00000000";
    when 16#016E7# => romdata <= X"00000000";
    when 16#016E8# => romdata <= X"00000000";
    when 16#016E9# => romdata <= X"00000000";
    when 16#016EA# => romdata <= X"00000000";
    when 16#016EB# => romdata <= X"00000000";
    when 16#016EC# => romdata <= X"00000000";
    when 16#016ED# => romdata <= X"00000000";
    when 16#016EE# => romdata <= X"00000000";
    when 16#016EF# => romdata <= X"00000000";
    when 16#016F0# => romdata <= X"00000000";
    when 16#016F1# => romdata <= X"00000000";
    when 16#016F2# => romdata <= X"00000000";
    when 16#016F3# => romdata <= X"00000000";
    when 16#016F4# => romdata <= X"00000000";
    when 16#016F5# => romdata <= X"00000000";
    when 16#016F6# => romdata <= X"00000000";
    when 16#016F7# => romdata <= X"00000000";
    when 16#016F8# => romdata <= X"00000000";
    when 16#016F9# => romdata <= X"00000000";
    when 16#016FA# => romdata <= X"00000000";
    when 16#016FB# => romdata <= X"00000000";
    when 16#016FC# => romdata <= X"00000000";
    when 16#016FD# => romdata <= X"00000000";
    when 16#016FE# => romdata <= X"00000000";
    when 16#016FF# => romdata <= X"00000000";
    when 16#01700# => romdata <= X"00000000";
    when 16#01701# => romdata <= X"00000000";
    when 16#01702# => romdata <= X"00000000";
    when 16#01703# => romdata <= X"00000000";
    when 16#01704# => romdata <= X"00000000";
    when 16#01705# => romdata <= X"00000000";
    when 16#01706# => romdata <= X"00000000";
    when 16#01707# => romdata <= X"00000000";
    when 16#01708# => romdata <= X"00000000";
    when 16#01709# => romdata <= X"00000000";
    when 16#0170A# => romdata <= X"00000000";
    when 16#0170B# => romdata <= X"00000000";
    when 16#0170C# => romdata <= X"00000000";
    when 16#0170D# => romdata <= X"00000000";
    when 16#0170E# => romdata <= X"00000000";
    when 16#0170F# => romdata <= X"00000000";
    when 16#01710# => romdata <= X"00000000";
    when 16#01711# => romdata <= X"00000000";
    when 16#01712# => romdata <= X"00000000";
    when 16#01713# => romdata <= X"00000000";
    when 16#01714# => romdata <= X"00000000";
    when 16#01715# => romdata <= X"00000000";
    when 16#01716# => romdata <= X"00000000";
    when 16#01717# => romdata <= X"00000000";
    when 16#01718# => romdata <= X"00000000";
    when 16#01719# => romdata <= X"00000000";
    when 16#0171A# => romdata <= X"00000000";
    when 16#0171B# => romdata <= X"00000000";
    when 16#0171C# => romdata <= X"00000000";
    when 16#0171D# => romdata <= X"00000000";
    when 16#0171E# => romdata <= X"00000000";
    when 16#0171F# => romdata <= X"00000000";
    when 16#01720# => romdata <= X"00000000";
    when 16#01721# => romdata <= X"00000000";
    when 16#01722# => romdata <= X"00000000";
    when 16#01723# => romdata <= X"00000000";
    when 16#01724# => romdata <= X"00000000";
    when 16#01725# => romdata <= X"00000000";
    when 16#01726# => romdata <= X"00000000";
    when 16#01727# => romdata <= X"00000000";
    when 16#01728# => romdata <= X"00000000";
    when 16#01729# => romdata <= X"00000000";
    when 16#0172A# => romdata <= X"00000000";
    when 16#0172B# => romdata <= X"00000000";
    when 16#0172C# => romdata <= X"00000000";
    when 16#0172D# => romdata <= X"00000000";
    when 16#0172E# => romdata <= X"00000000";
    when 16#0172F# => romdata <= X"00000000";
    when 16#01730# => romdata <= X"00000000";
    when 16#01731# => romdata <= X"00000000";
    when 16#01732# => romdata <= X"00000000";
    when 16#01733# => romdata <= X"00000000";
    when 16#01734# => romdata <= X"00000000";
    when 16#01735# => romdata <= X"00000000";
    when 16#01736# => romdata <= X"00000000";
    when 16#01737# => romdata <= X"00000000";
    when 16#01738# => romdata <= X"FFFFFFFF";
    when 16#01739# => romdata <= X"00000000";
    when 16#0173A# => romdata <= X"00020000";
    when 16#0173B# => romdata <= X"00000000";
    when 16#0173C# => romdata <= X"00000000";
    when 16#0173D# => romdata <= X"00005CEC";
    when 16#0173E# => romdata <= X"00005CEC";
    when 16#0173F# => romdata <= X"00005CF4";
    when 16#01740# => romdata <= X"00005CF4";
    when 16#01741# => romdata <= X"00005CFC";
    when 16#01742# => romdata <= X"00005CFC";
    when 16#01743# => romdata <= X"00005D04";
    when 16#01744# => romdata <= X"00005D04";
    when 16#01745# => romdata <= X"00005D0C";
    when 16#01746# => romdata <= X"00005D0C";
    when 16#01747# => romdata <= X"00005D14";
    when 16#01748# => romdata <= X"00005D14";
    when 16#01749# => romdata <= X"00005D1C";
    when 16#0174A# => romdata <= X"00005D1C";
    when 16#0174B# => romdata <= X"00005D24";
    when 16#0174C# => romdata <= X"00005D24";
    when 16#0174D# => romdata <= X"00005D2C";
    when 16#0174E# => romdata <= X"00005D2C";
    when 16#0174F# => romdata <= X"00005D34";
    when 16#01750# => romdata <= X"00005D34";
    when 16#01751# => romdata <= X"00005D3C";
    when 16#01752# => romdata <= X"00005D3C";
    when 16#01753# => romdata <= X"00005D44";
    when 16#01754# => romdata <= X"00005D44";
    when 16#01755# => romdata <= X"00005D4C";
    when 16#01756# => romdata <= X"00005D4C";
    when 16#01757# => romdata <= X"00005D54";
    when 16#01758# => romdata <= X"00005D54";
    when 16#01759# => romdata <= X"00005D5C";
    when 16#0175A# => romdata <= X"00005D5C";
    when 16#0175B# => romdata <= X"00005D64";
    when 16#0175C# => romdata <= X"00005D64";
    when 16#0175D# => romdata <= X"00005D6C";
    when 16#0175E# => romdata <= X"00005D6C";
    when 16#0175F# => romdata <= X"00005D74";
    when 16#01760# => romdata <= X"00005D74";
    when 16#01761# => romdata <= X"00005D7C";
    when 16#01762# => romdata <= X"00005D7C";
    when 16#01763# => romdata <= X"00005D84";
    when 16#01764# => romdata <= X"00005D84";
    when 16#01765# => romdata <= X"00005D8C";
    when 16#01766# => romdata <= X"00005D8C";
    when 16#01767# => romdata <= X"00005D94";
    when 16#01768# => romdata <= X"00005D94";
    when 16#01769# => romdata <= X"00005D9C";
    when 16#0176A# => romdata <= X"00005D9C";
    when 16#0176B# => romdata <= X"00005DA4";
    when 16#0176C# => romdata <= X"00005DA4";
    when 16#0176D# => romdata <= X"00005DAC";
    when 16#0176E# => romdata <= X"00005DAC";
    when 16#0176F# => romdata <= X"00005DB4";
    when 16#01770# => romdata <= X"00005DB4";
    when 16#01771# => romdata <= X"00005DBC";
    when 16#01772# => romdata <= X"00005DBC";
    when 16#01773# => romdata <= X"00005DC4";
    when 16#01774# => romdata <= X"00005DC4";
    when 16#01775# => romdata <= X"00005DCC";
    when 16#01776# => romdata <= X"00005DCC";
    when 16#01777# => romdata <= X"00005DD4";
    when 16#01778# => romdata <= X"00005DD4";
    when 16#01779# => romdata <= X"00005DDC";
    when 16#0177A# => romdata <= X"00005DDC";
    when 16#0177B# => romdata <= X"00005DE4";
    when 16#0177C# => romdata <= X"00005DE4";
    when 16#0177D# => romdata <= X"00005DEC";
    when 16#0177E# => romdata <= X"00005DEC";
    when 16#0177F# => romdata <= X"00005DF4";
    when 16#01780# => romdata <= X"00005DF4";
    when 16#01781# => romdata <= X"00005DFC";
    when 16#01782# => romdata <= X"00005DFC";
    when 16#01783# => romdata <= X"00005E04";
    when 16#01784# => romdata <= X"00005E04";
    when 16#01785# => romdata <= X"00005E0C";
    when 16#01786# => romdata <= X"00005E0C";
    when 16#01787# => romdata <= X"00005E14";
    when 16#01788# => romdata <= X"00005E14";
    when 16#01789# => romdata <= X"00005E1C";
    when 16#0178A# => romdata <= X"00005E1C";
    when 16#0178B# => romdata <= X"00005E24";
    when 16#0178C# => romdata <= X"00005E24";
    when 16#0178D# => romdata <= X"00005E2C";
    when 16#0178E# => romdata <= X"00005E2C";
    when 16#0178F# => romdata <= X"00005E34";
    when 16#01790# => romdata <= X"00005E34";
    when 16#01791# => romdata <= X"00005E3C";
    when 16#01792# => romdata <= X"00005E3C";
    when 16#01793# => romdata <= X"00005E44";
    when 16#01794# => romdata <= X"00005E44";
    when 16#01795# => romdata <= X"00005E4C";
    when 16#01796# => romdata <= X"00005E4C";
    when 16#01797# => romdata <= X"00005E54";
    when 16#01798# => romdata <= X"00005E54";
    when 16#01799# => romdata <= X"00005E5C";
    when 16#0179A# => romdata <= X"00005E5C";
    when 16#0179B# => romdata <= X"00005E64";
    when 16#0179C# => romdata <= X"00005E64";
    when 16#0179D# => romdata <= X"00005E6C";
    when 16#0179E# => romdata <= X"00005E6C";
    when 16#0179F# => romdata <= X"00005E74";
    when 16#017A0# => romdata <= X"00005E74";
    when 16#017A1# => romdata <= X"00005E7C";
    when 16#017A2# => romdata <= X"00005E7C";
    when 16#017A3# => romdata <= X"00005E84";
    when 16#017A4# => romdata <= X"00005E84";
    when 16#017A5# => romdata <= X"00005E8C";
    when 16#017A6# => romdata <= X"00005E8C";
    when 16#017A7# => romdata <= X"00005E94";
    when 16#017A8# => romdata <= X"00005E94";
    when 16#017A9# => romdata <= X"00005E9C";
    when 16#017AA# => romdata <= X"00005E9C";
    when 16#017AB# => romdata <= X"00005EA4";
    when 16#017AC# => romdata <= X"00005EA4";
    when 16#017AD# => romdata <= X"00005EAC";
    when 16#017AE# => romdata <= X"00005EAC";
    when 16#017AF# => romdata <= X"00005EB4";
    when 16#017B0# => romdata <= X"00005EB4";
    when 16#017B1# => romdata <= X"00005EBC";
    when 16#017B2# => romdata <= X"00005EBC";
    when 16#017B3# => romdata <= X"00005EC4";
    when 16#017B4# => romdata <= X"00005EC4";
    when 16#017B5# => romdata <= X"00005ECC";
    when 16#017B6# => romdata <= X"00005ECC";
    when 16#017B7# => romdata <= X"00005ED4";
    when 16#017B8# => romdata <= X"00005ED4";
    when 16#017B9# => romdata <= X"00005EDC";
    when 16#017BA# => romdata <= X"00005EDC";
    when 16#017BB# => romdata <= X"00005EE4";
    when 16#017BC# => romdata <= X"00005EE4";
    when 16#017BD# => romdata <= X"00005EEC";
    when 16#017BE# => romdata <= X"00005EEC";
    when 16#017BF# => romdata <= X"00005EF4";
    when 16#017C0# => romdata <= X"00005EF4";
    when 16#017C1# => romdata <= X"00005EFC";
    when 16#017C2# => romdata <= X"00005EFC";
    when 16#017C3# => romdata <= X"00005F04";
    when 16#017C4# => romdata <= X"00005F04";
    when 16#017C5# => romdata <= X"00005F0C";
    when 16#017C6# => romdata <= X"00005F0C";
    when 16#017C7# => romdata <= X"00005F14";
    when 16#017C8# => romdata <= X"00005F14";
    when 16#017C9# => romdata <= X"00005F1C";
    when 16#017CA# => romdata <= X"00005F1C";
    when 16#017CB# => romdata <= X"00005F24";
    when 16#017CC# => romdata <= X"00005F24";
    when 16#017CD# => romdata <= X"00005F2C";
    when 16#017CE# => romdata <= X"00005F2C";
    when 16#017CF# => romdata <= X"00005F34";
    when 16#017D0# => romdata <= X"00005F34";
    when 16#017D1# => romdata <= X"00005F3C";
    when 16#017D2# => romdata <= X"00005F3C";
    when 16#017D3# => romdata <= X"00005F44";
    when 16#017D4# => romdata <= X"00005F44";
    when 16#017D5# => romdata <= X"00005F4C";
    when 16#017D6# => romdata <= X"00005F4C";
    when 16#017D7# => romdata <= X"00005F54";
    when 16#017D8# => romdata <= X"00005F54";
    when 16#017D9# => romdata <= X"00005F5C";
    when 16#017DA# => romdata <= X"00005F5C";
    when 16#017DB# => romdata <= X"00005F64";
    when 16#017DC# => romdata <= X"00005F64";
    when 16#017DD# => romdata <= X"00005F6C";
    when 16#017DE# => romdata <= X"00005F6C";
    when 16#017DF# => romdata <= X"00005F74";
    when 16#017E0# => romdata <= X"00005F74";
    when 16#017E1# => romdata <= X"00005F7C";
    when 16#017E2# => romdata <= X"00005F7C";
    when 16#017E3# => romdata <= X"00005F84";
    when 16#017E4# => romdata <= X"00005F84";
    when 16#017E5# => romdata <= X"00005F8C";
    when 16#017E6# => romdata <= X"00005F8C";
    when 16#017E7# => romdata <= X"00005F94";
    when 16#017E8# => romdata <= X"00005F94";
    when 16#017E9# => romdata <= X"00005F9C";
    when 16#017EA# => romdata <= X"00005F9C";
    when 16#017EB# => romdata <= X"00005FA4";
    when 16#017EC# => romdata <= X"00005FA4";
    when 16#017ED# => romdata <= X"00005FAC";
    when 16#017EE# => romdata <= X"00005FAC";
    when 16#017EF# => romdata <= X"00005FB4";
    when 16#017F0# => romdata <= X"00005FB4";
    when 16#017F1# => romdata <= X"00005FBC";
    when 16#017F2# => romdata <= X"00005FBC";
    when 16#017F3# => romdata <= X"00005FC4";
    when 16#017F4# => romdata <= X"00005FC4";
    when 16#017F5# => romdata <= X"00005FCC";
    when 16#017F6# => romdata <= X"00005FCC";
    when 16#017F7# => romdata <= X"00005FD4";
    when 16#017F8# => romdata <= X"00005FD4";
    when 16#017F9# => romdata <= X"00005FDC";
    when 16#017FA# => romdata <= X"00005FDC";
    when 16#017FB# => romdata <= X"00005FE4";
    when 16#017FC# => romdata <= X"00005FE4";
    when 16#017FD# => romdata <= X"00005FEC";
    when 16#017FE# => romdata <= X"00005FEC";
    when 16#017FF# => romdata <= X"00005FF4";
    when 16#01800# => romdata <= X"00005FF4";
    when 16#01801# => romdata <= X"00005FFC";
    when 16#01802# => romdata <= X"00005FFC";
    when 16#01803# => romdata <= X"00006004";
    when 16#01804# => romdata <= X"00006004";
    when 16#01805# => romdata <= X"0000600C";
    when 16#01806# => romdata <= X"0000600C";
    when 16#01807# => romdata <= X"00006014";
    when 16#01808# => romdata <= X"00006014";
    when 16#01809# => romdata <= X"0000601C";
    when 16#0180A# => romdata <= X"0000601C";
    when 16#0180B# => romdata <= X"00006024";
    when 16#0180C# => romdata <= X"00006024";
    when 16#0180D# => romdata <= X"0000602C";
    when 16#0180E# => romdata <= X"0000602C";
    when 16#0180F# => romdata <= X"00006034";
    when 16#01810# => romdata <= X"00006034";
    when 16#01811# => romdata <= X"0000603C";
    when 16#01812# => romdata <= X"0000603C";
    when 16#01813# => romdata <= X"00006044";
    when 16#01814# => romdata <= X"00006044";
    when 16#01815# => romdata <= X"0000604C";
    when 16#01816# => romdata <= X"0000604C";
    when 16#01817# => romdata <= X"00006054";
    when 16#01818# => romdata <= X"00006054";
    when 16#01819# => romdata <= X"0000605C";
    when 16#0181A# => romdata <= X"0000605C";
    when 16#0181B# => romdata <= X"00006064";
    when 16#0181C# => romdata <= X"00006064";
    when 16#0181D# => romdata <= X"0000606C";
    when 16#0181E# => romdata <= X"0000606C";
    when 16#0181F# => romdata <= X"00006074";
    when 16#01820# => romdata <= X"00006074";
    when 16#01821# => romdata <= X"0000607C";
    when 16#01822# => romdata <= X"0000607C";
    when 16#01823# => romdata <= X"00006084";
    when 16#01824# => romdata <= X"00006084";
    when 16#01825# => romdata <= X"0000608C";
    when 16#01826# => romdata <= X"0000608C";
    when 16#01827# => romdata <= X"00006094";
    when 16#01828# => romdata <= X"00006094";
    when 16#01829# => romdata <= X"0000609C";
    when 16#0182A# => romdata <= X"0000609C";
    when 16#0182B# => romdata <= X"000060A4";
    when 16#0182C# => romdata <= X"000060A4";
    when 16#0182D# => romdata <= X"000060AC";
    when 16#0182E# => romdata <= X"000060AC";
    when 16#0182F# => romdata <= X"000060B4";
    when 16#01830# => romdata <= X"000060B4";
    when 16#01831# => romdata <= X"000060BC";
    when 16#01832# => romdata <= X"000060BC";
    when 16#01833# => romdata <= X"000060C4";
    when 16#01834# => romdata <= X"000060C4";
    when 16#01835# => romdata <= X"000060CC";
    when 16#01836# => romdata <= X"000060CC";
    when 16#01837# => romdata <= X"000060D4";
    when 16#01838# => romdata <= X"000060D4";
    when 16#01839# => romdata <= X"000060DC";
    when 16#0183A# => romdata <= X"000060DC";
    when 16#0183B# => romdata <= X"000060E4";
    when 16#0183C# => romdata <= X"000060E4";
    when 16#0183D# => romdata <= X"000060E4";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
