-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0bba9c0c",
     3 => x"3a0b0b0b",
     4 => x"abbd0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b8ac52d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bba",
   162 => x"88738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b90",
   171 => x"c12d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b91",
   179 => x"f32d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bba980c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81fb3fa5",
   257 => x"9e3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104ba",
   280 => x"9808802e",
   281 => x"a338ba9c",
   282 => x"08822ebd",
   283 => x"38838080",
   284 => x"0b0b0b80",
   285 => x"caa00c82",
   286 => x"a0800b80",
   287 => x"caa40c82",
   288 => x"90800b80",
   289 => x"caa80c04",
   290 => x"f8808080",
   291 => x"a40b0b0b",
   292 => x"80caa00c",
   293 => x"f8808082",
   294 => x"800b80ca",
   295 => x"a40cf880",
   296 => x"8084800b",
   297 => x"80caa80c",
   298 => x"0480c0a8",
   299 => x"808c0b0b",
   300 => x"0b80caa0",
   301 => x"0c80c0a8",
   302 => x"80940b80",
   303 => x"caa40c0b",
   304 => x"0b0badd0",
   305 => x"0b80caa8",
   306 => x"0c04ff3d",
   307 => x"0d80caac",
   308 => x"335170a4",
   309 => x"38baa408",
   310 => x"70085252",
   311 => x"70802e92",
   312 => x"388412ba",
   313 => x"a40c702d",
   314 => x"baa40870",
   315 => x"08525270",
   316 => x"f038810b",
   317 => x"80caac34",
   318 => x"833d0d04",
   319 => x"04803d0d",
   320 => x"0b0b80ca",
   321 => x"9c08802e",
   322 => x"8e380b0b",
   323 => x"0b0b800b",
   324 => x"802e0981",
   325 => x"06853882",
   326 => x"3d0d040b",
   327 => x"0b80ca9c",
   328 => x"510b0b0b",
   329 => x"f5da3f82",
   330 => x"3d0d0404",
   331 => x"ff3d0d02",
   332 => x"8f053370",
   333 => x"52528490",
   334 => x"3f715185",
   335 => x"823f7180",
   336 => x"0c833d0d",
   337 => x"04ff3d0d",
   338 => x"800b80ca",
   339 => x"b4085252",
   340 => x"70722e09",
   341 => x"81068338",
   342 => x"81527180",
   343 => x"cab40cba",
   344 => x"b8085281",
   345 => x"800b8c13",
   346 => x"0c833d0d",
   347 => x"04f73d0d",
   348 => x"bab00870",
   349 => x"08810a06",
   350 => x"80cab00c",
   351 => x"5383843f",
   352 => x"83b13f8d",
   353 => x"a95280ca",
   354 => x"b0088438",
   355 => x"8aac5271",
   356 => x"80cab80c",
   357 => x"84863fba",
   358 => x"a80853fa",
   359 => x"c98e868c",
   360 => x"730c7208",
   361 => x"70842a81",
   362 => x"06515473",
   363 => x"f538bab0",
   364 => x"08881108",
   365 => x"81ff0788",
   366 => x"120c7480",
   367 => x"cab40c94",
   368 => x"11088180",
   369 => x"0794120c",
   370 => x"8c110881",
   371 => x"80078c12",
   372 => x"0c53bab8",
   373 => x"08528180",
   374 => x"0b80c013",
   375 => x"0cb9b051",
   376 => x"81dc3f80",
   377 => x"cab00880",
   378 => x"2e819838",
   379 => x"b9b85181",
   380 => x"cd3fb0c8",
   381 => x"5181c73f",
   382 => x"f881c08e",
   383 => x"8053a00b",
   384 => x"bab00855",
   385 => x"5580cab0",
   386 => x"08802e80",
   387 => x"d2387281",
   388 => x"ff068415",
   389 => x"0c80cab4",
   390 => x"08527180",
   391 => x"2e9f3872",
   392 => x"9f2a7310",
   393 => x"07537480",
   394 => x"2e9f38ff",
   395 => x"157381ff",
   396 => x"0684160c",
   397 => x"80cab408",
   398 => x"535571e3",
   399 => x"38720a10",
   400 => x"0a739f2b",
   401 => x"075374e3",
   402 => x"3887f23f",
   403 => x"720a100a",
   404 => x"739f2b07",
   405 => x"5380fd51",
   406 => x"81873fba",
   407 => x"b0085472",
   408 => x"81ff0684",
   409 => x"150c80ca",
   410 => x"b4085473",
   411 => x"802edd38",
   412 => x"729f2a73",
   413 => x"10075380",
   414 => x"fd5180e5",
   415 => x"3fbab008",
   416 => x"54dd39b9",
   417 => x"c451b73f",
   418 => x"b9d451b2",
   419 => x"3fb0c851",
   420 => x"ad3ff881",
   421 => x"c08e8053",
   422 => x"a00bbab0",
   423 => x"08555580",
   424 => x"cab008fe",
   425 => x"e938ffb7",
   426 => x"39ff3d0d",
   427 => x"028f0533",
   428 => x"baac0852",
   429 => x"710c800b",
   430 => x"800c833d",
   431 => x"0d04fe3d",
   432 => x"0d747033",
   433 => x"53537180",
   434 => x"2e933881",
   435 => x"13725280",
   436 => x"cab80853",
   437 => x"53712d72",
   438 => x"335271ef",
   439 => x"38843d0d",
   440 => x"04fd3d0d",
   441 => x"babc0876",
   442 => x"b0ea2994",
   443 => x"120c5485",
   444 => x"0b98150c",
   445 => x"98140870",
   446 => x"81065153",
   447 => x"72f63885",
   448 => x"3d0d0480",
   449 => x"3d0dbabc",
   450 => x"0851870b",
   451 => x"84120cff",
   452 => x"0bb4120c",
   453 => x"a70bb812",
   454 => x"0c87e80b",
   455 => x"a4120ca7",
   456 => x"0ba8120c",
   457 => x"b0ea0b94",
   458 => x"120c870b",
   459 => x"98120c82",
   460 => x"3d0d0480",
   461 => x"3d0dbac0",
   462 => x"0851b60b",
   463 => x"8c120c83",
   464 => x"0b88120c",
   465 => x"823d0d04",
   466 => x"fe3d0d02",
   467 => x"93053353",
   468 => x"728a2e9d",
   469 => x"38bac008",
   470 => x"52841208",
   471 => x"70822a70",
   472 => x"81065151",
   473 => x"5170802e",
   474 => x"f0387272",
   475 => x"0c843d0d",
   476 => x"04bac008",
   477 => x"52841208",
   478 => x"70822a70",
   479 => x"81065151",
   480 => x"5170802e",
   481 => x"f0388d72",
   482 => x"0c841208",
   483 => x"70822a70",
   484 => x"81065151",
   485 => x"5170802e",
   486 => x"c038cf39",
   487 => x"803d0dba",
   488 => x"b4085180",
   489 => x"0b84120c",
   490 => x"83fe800b",
   491 => x"88120c80",
   492 => x"0b80cabc",
   493 => x"34800b80",
   494 => x"cac03482",
   495 => x"3d0d04fa",
   496 => x"3d0d02a3",
   497 => x"0533bab4",
   498 => x"0880cabc",
   499 => x"337081ff",
   500 => x"06701010",
   501 => x"1180cac0",
   502 => x"337081ff",
   503 => x"06729029",
   504 => x"1170882b",
   505 => x"7807770c",
   506 => x"535b5b55",
   507 => x"55595454",
   508 => x"738a2e98",
   509 => x"387480cf",
   510 => x"2e923873",
   511 => x"8c2ea438",
   512 => x"81165372",
   513 => x"80cac034",
   514 => x"883d0d04",
   515 => x"71a326a3",
   516 => x"38811752",
   517 => x"7180cabc",
   518 => x"34800b80",
   519 => x"cac03488",
   520 => x"3d0d0480",
   521 => x"5271882b",
   522 => x"730c8112",
   523 => x"52979072",
   524 => x"26f33880",
   525 => x"0b80cabc",
   526 => x"34800b80",
   527 => x"cac034df",
   528 => x"398c0802",
   529 => x"8c0cf93d",
   530 => x"0d800b8c",
   531 => x"08fc050c",
   532 => x"8c088805",
   533 => x"088025ab",
   534 => x"388c0888",
   535 => x"0508308c",
   536 => x"0888050c",
   537 => x"800b8c08",
   538 => x"f4050c8c",
   539 => x"08fc0508",
   540 => x"8838810b",
   541 => x"8c08f405",
   542 => x"0c8c08f4",
   543 => x"05088c08",
   544 => x"fc050c8c",
   545 => x"088c0508",
   546 => x"8025ab38",
   547 => x"8c088c05",
   548 => x"08308c08",
   549 => x"8c050c80",
   550 => x"0b8c08f0",
   551 => x"050c8c08",
   552 => x"fc050888",
   553 => x"38810b8c",
   554 => x"08f0050c",
   555 => x"8c08f005",
   556 => x"088c08fc",
   557 => x"050c8053",
   558 => x"8c088c05",
   559 => x"08528c08",
   560 => x"88050851",
   561 => x"81a73f80",
   562 => x"08708c08",
   563 => x"f8050c54",
   564 => x"8c08fc05",
   565 => x"08802e8c",
   566 => x"388c08f8",
   567 => x"0508308c",
   568 => x"08f8050c",
   569 => x"8c08f805",
   570 => x"0870800c",
   571 => x"54893d0d",
   572 => x"8c0c048c",
   573 => x"08028c0c",
   574 => x"fb3d0d80",
   575 => x"0b8c08fc",
   576 => x"050c8c08",
   577 => x"88050880",
   578 => x"2593388c",
   579 => x"08880508",
   580 => x"308c0888",
   581 => x"050c810b",
   582 => x"8c08fc05",
   583 => x"0c8c088c",
   584 => x"05088025",
   585 => x"8c388c08",
   586 => x"8c050830",
   587 => x"8c088c05",
   588 => x"0c81538c",
   589 => x"088c0508",
   590 => x"528c0888",
   591 => x"050851ad",
   592 => x"3f800870",
   593 => x"8c08f805",
   594 => x"0c548c08",
   595 => x"fc050880",
   596 => x"2e8c388c",
   597 => x"08f80508",
   598 => x"308c08f8",
   599 => x"050c8c08",
   600 => x"f8050870",
   601 => x"800c5487",
   602 => x"3d0d8c0c",
   603 => x"048c0802",
   604 => x"8c0cfd3d",
   605 => x"0d810b8c",
   606 => x"08fc050c",
   607 => x"800b8c08",
   608 => x"f8050c8c",
   609 => x"088c0508",
   610 => x"8c088805",
   611 => x"0827ac38",
   612 => x"8c08fc05",
   613 => x"08802ea3",
   614 => x"38800b8c",
   615 => x"088c0508",
   616 => x"2499388c",
   617 => x"088c0508",
   618 => x"108c088c",
   619 => x"050c8c08",
   620 => x"fc050810",
   621 => x"8c08fc05",
   622 => x"0cc9398c",
   623 => x"08fc0508",
   624 => x"802e80c9",
   625 => x"388c088c",
   626 => x"05088c08",
   627 => x"88050826",
   628 => x"a1388c08",
   629 => x"8805088c",
   630 => x"088c0508",
   631 => x"318c0888",
   632 => x"050c8c08",
   633 => x"f805088c",
   634 => x"08fc0508",
   635 => x"078c08f8",
   636 => x"050c8c08",
   637 => x"fc050881",
   638 => x"2a8c08fc",
   639 => x"050c8c08",
   640 => x"8c050881",
   641 => x"2a8c088c",
   642 => x"050cffaf",
   643 => x"398c0890",
   644 => x"0508802e",
   645 => x"8f388c08",
   646 => x"88050870",
   647 => x"8c08f405",
   648 => x"0c518d39",
   649 => x"8c08f805",
   650 => x"08708c08",
   651 => x"f4050c51",
   652 => x"8c08f405",
   653 => x"08800c85",
   654 => x"3d0d8c0c",
   655 => x"04803d0d",
   656 => x"865182fd",
   657 => x"3f815197",
   658 => x"b53ffd3d",
   659 => x"0d755384",
   660 => x"d8130880",
   661 => x"2e8a3880",
   662 => x"5372800c",
   663 => x"853d0d04",
   664 => x"81805272",
   665 => x"5183d43f",
   666 => x"800884d8",
   667 => x"140cff53",
   668 => x"8008802e",
   669 => x"e4388008",
   670 => x"549f5380",
   671 => x"74708405",
   672 => x"560cff13",
   673 => x"53807324",
   674 => x"ce388074",
   675 => x"70840556",
   676 => x"0cff1353",
   677 => x"728025e3",
   678 => x"38ffbc39",
   679 => x"fd3d0d75",
   680 => x"7755539f",
   681 => x"74278d38",
   682 => x"96730cff",
   683 => x"5271800c",
   684 => x"853d0d04",
   685 => x"84d81308",
   686 => x"5271802e",
   687 => x"93387310",
   688 => x"10127008",
   689 => x"79720c51",
   690 => x"5271800c",
   691 => x"853d0d04",
   692 => x"7251fef6",
   693 => x"3fff5280",
   694 => x"08d33884",
   695 => x"d8130874",
   696 => x"10101170",
   697 => x"087a720c",
   698 => x"515152dd",
   699 => x"39f93d0d",
   700 => x"797b5856",
   701 => x"769f2680",
   702 => x"e83884d8",
   703 => x"16085473",
   704 => x"802eaa38",
   705 => x"76101014",
   706 => x"70085555",
   707 => x"73802eba",
   708 => x"38805873",
   709 => x"812e8f38",
   710 => x"73ff2ea3",
   711 => x"3880750c",
   712 => x"7651732d",
   713 => x"80587780",
   714 => x"0c893d0d",
   715 => x"047551fe",
   716 => x"993fff58",
   717 => x"8008ef38",
   718 => x"84d81608",
   719 => x"54c63996",
   720 => x"760c810b",
   721 => x"800c893d",
   722 => x"0d047551",
   723 => x"81e93f76",
   724 => x"53800852",
   725 => x"755181a9",
   726 => x"3f800880",
   727 => x"0c893d0d",
   728 => x"0496760c",
   729 => x"ff0b800c",
   730 => x"893d0d04",
   731 => x"fc3d0d76",
   732 => x"785653ff",
   733 => x"54749f26",
   734 => x"b13884d8",
   735 => x"13085271",
   736 => x"802eae38",
   737 => x"74101012",
   738 => x"70085353",
   739 => x"81547180",
   740 => x"2e983882",
   741 => x"5471ff2e",
   742 => x"91388354",
   743 => x"71812e8a",
   744 => x"3880730c",
   745 => x"7451712d",
   746 => x"80547380",
   747 => x"0c863d0d",
   748 => x"047251fd",
   749 => x"953f8008",
   750 => x"f13884d8",
   751 => x"130852c4",
   752 => x"39ff3d0d",
   753 => x"7352bac4",
   754 => x"0851fea1",
   755 => x"3f833d0d",
   756 => x"04fe3d0d",
   757 => x"75537452",
   758 => x"bac40851",
   759 => x"fdbe3f84",
   760 => x"3d0d0480",
   761 => x"3d0dbac4",
   762 => x"0851fcde",
   763 => x"3f823d0d",
   764 => x"04ff3d0d",
   765 => x"7352bac4",
   766 => x"0851fef0",
   767 => x"3f833d0d",
   768 => x"04fc3d0d",
   769 => x"800b80ca",
   770 => x"cc0c7852",
   771 => x"775192e7",
   772 => x"3f800854",
   773 => x"8008ff2e",
   774 => x"88387380",
   775 => x"0c863d0d",
   776 => x"0480cacc",
   777 => x"08557480",
   778 => x"2ef03876",
   779 => x"75710c53",
   780 => x"73800c86",
   781 => x"3d0d0492",
   782 => x"b93f04f3",
   783 => x"3d0d7f61",
   784 => x"8b1170f8",
   785 => x"065c5555",
   786 => x"5e729626",
   787 => x"83389059",
   788 => x"80792474",
   789 => x"7a260753",
   790 => x"80547274",
   791 => x"2e098106",
   792 => x"80cb387d",
   793 => x"518bca3f",
   794 => x"7883f726",
   795 => x"80c63878",
   796 => x"832a7010",
   797 => x"101080c2",
   798 => x"80058c11",
   799 => x"0859595a",
   800 => x"76782e83",
   801 => x"b0388417",
   802 => x"08fc0656",
   803 => x"8c170888",
   804 => x"1808718c",
   805 => x"120c8812",
   806 => x"0c587517",
   807 => x"84110881",
   808 => x"0784120c",
   809 => x"537d518b",
   810 => x"893f8817",
   811 => x"5473800c",
   812 => x"8f3d0d04",
   813 => x"78892a79",
   814 => x"832a5b53",
   815 => x"72802ebf",
   816 => x"3878862a",
   817 => x"b8055a84",
   818 => x"7327b438",
   819 => x"80db135a",
   820 => x"947327ab",
   821 => x"38788c2a",
   822 => x"80ee055a",
   823 => x"80d47327",
   824 => x"9e38788f",
   825 => x"2a80f705",
   826 => x"5a82d473",
   827 => x"27913878",
   828 => x"922a80fc",
   829 => x"055a8ad4",
   830 => x"73278438",
   831 => x"80fe5a79",
   832 => x"10101080",
   833 => x"c280058c",
   834 => x"11085855",
   835 => x"76752ea3",
   836 => x"38841708",
   837 => x"fc06707a",
   838 => x"31555673",
   839 => x"8f2488d5",
   840 => x"38738025",
   841 => x"fee6388c",
   842 => x"17085776",
   843 => x"752e0981",
   844 => x"06df3881",
   845 => x"1a5a80c2",
   846 => x"90085776",
   847 => x"80c2882e",
   848 => x"82c03884",
   849 => x"1708fc06",
   850 => x"707a3155",
   851 => x"56738f24",
   852 => x"81f93880",
   853 => x"c2880b80",
   854 => x"c2940c80",
   855 => x"c2880b80",
   856 => x"c2900c73",
   857 => x"8025feb2",
   858 => x"3883ff76",
   859 => x"2783df38",
   860 => x"75892a76",
   861 => x"832a5553",
   862 => x"72802ebf",
   863 => x"3875862a",
   864 => x"b8055484",
   865 => x"7327b438",
   866 => x"80db1354",
   867 => x"947327ab",
   868 => x"38758c2a",
   869 => x"80ee0554",
   870 => x"80d47327",
   871 => x"9e38758f",
   872 => x"2a80f705",
   873 => x"5482d473",
   874 => x"27913875",
   875 => x"922a80fc",
   876 => x"05548ad4",
   877 => x"73278438",
   878 => x"80fe5473",
   879 => x"10101080",
   880 => x"c2800588",
   881 => x"11085658",
   882 => x"74782e86",
   883 => x"cf388415",
   884 => x"08fc0653",
   885 => x"7573278d",
   886 => x"38881508",
   887 => x"5574782e",
   888 => x"098106ea",
   889 => x"388c1508",
   890 => x"80c2800b",
   891 => x"84050871",
   892 => x"8c1a0c76",
   893 => x"881a0c78",
   894 => x"88130c78",
   895 => x"8c180c5d",
   896 => x"58795380",
   897 => x"7a2483e6",
   898 => x"3872822c",
   899 => x"81712b5c",
   900 => x"537a7c26",
   901 => x"8198387b",
   902 => x"7b065372",
   903 => x"82f13879",
   904 => x"fc068405",
   905 => x"5a7a1070",
   906 => x"7d06545b",
   907 => x"7282e038",
   908 => x"841a5af1",
   909 => x"3988178c",
   910 => x"11085858",
   911 => x"76782e09",
   912 => x"8106fcc2",
   913 => x"38821a5a",
   914 => x"fdec3978",
   915 => x"17798107",
   916 => x"84190c70",
   917 => x"80c2940c",
   918 => x"7080c290",
   919 => x"0c80c288",
   920 => x"0b8c120c",
   921 => x"8c110888",
   922 => x"120c7481",
   923 => x"0784120c",
   924 => x"74117571",
   925 => x"0c51537d",
   926 => x"5187b73f",
   927 => x"881754fc",
   928 => x"ac3980c2",
   929 => x"800b8405",
   930 => x"087a545c",
   931 => x"798025fe",
   932 => x"f83882da",
   933 => x"397a097c",
   934 => x"067080c2",
   935 => x"800b8405",
   936 => x"0c5c7a10",
   937 => x"5b7a7c26",
   938 => x"85387a85",
   939 => x"b83880c2",
   940 => x"800b8805",
   941 => x"08708412",
   942 => x"08fc0670",
   943 => x"7c317c72",
   944 => x"268f7225",
   945 => x"0757575c",
   946 => x"5d557280",
   947 => x"2e80db38",
   948 => x"797a1680",
   949 => x"c1f8081b",
   950 => x"90115a55",
   951 => x"575b80c1",
   952 => x"f408ff2e",
   953 => x"8838a08f",
   954 => x"13e08006",
   955 => x"5776527d",
   956 => x"5186c03f",
   957 => x"80085480",
   958 => x"08ff2e90",
   959 => x"38800876",
   960 => x"27829938",
   961 => x"7480c280",
   962 => x"2e829138",
   963 => x"80c2800b",
   964 => x"88050855",
   965 => x"841508fc",
   966 => x"06707a31",
   967 => x"7a72268f",
   968 => x"72250752",
   969 => x"55537283",
   970 => x"e6387479",
   971 => x"81078417",
   972 => x"0c791670",
   973 => x"80c2800b",
   974 => x"88050c75",
   975 => x"81078412",
   976 => x"0c547e52",
   977 => x"5785eb3f",
   978 => x"881754fa",
   979 => x"e0397583",
   980 => x"2a705454",
   981 => x"80742481",
   982 => x"9b387282",
   983 => x"2c81712b",
   984 => x"80c28408",
   985 => x"077080c2",
   986 => x"800b8405",
   987 => x"0c751010",
   988 => x"1080c280",
   989 => x"05881108",
   990 => x"585a5d53",
   991 => x"778c180c",
   992 => x"7488180c",
   993 => x"7688190c",
   994 => x"768c160c",
   995 => x"fcf33979",
   996 => x"7a101010",
   997 => x"80c28005",
   998 => x"7057595d",
   999 => x"8c150857",
  1000 => x"76752ea3",
  1001 => x"38841708",
  1002 => x"fc06707a",
  1003 => x"31555673",
  1004 => x"8f2483ca",
  1005 => x"38738025",
  1006 => x"8481388c",
  1007 => x"17085776",
  1008 => x"752e0981",
  1009 => x"06df3888",
  1010 => x"15811b70",
  1011 => x"8306555b",
  1012 => x"5572c938",
  1013 => x"7c830653",
  1014 => x"72802efd",
  1015 => x"b838ff1d",
  1016 => x"f819595d",
  1017 => x"88180878",
  1018 => x"2eea38fd",
  1019 => x"b539831a",
  1020 => x"53fc9639",
  1021 => x"83147082",
  1022 => x"2c81712b",
  1023 => x"80c28408",
  1024 => x"077080c2",
  1025 => x"800b8405",
  1026 => x"0c761010",
  1027 => x"1080c280",
  1028 => x"05881108",
  1029 => x"595b5e51",
  1030 => x"53fee139",
  1031 => x"80c1c408",
  1032 => x"17588008",
  1033 => x"762e818d",
  1034 => x"3880c1f4",
  1035 => x"08ff2e83",
  1036 => x"ec387376",
  1037 => x"311880c1",
  1038 => x"c40c7387",
  1039 => x"06705753",
  1040 => x"72802e88",
  1041 => x"38887331",
  1042 => x"70155556",
  1043 => x"76149fff",
  1044 => x"06a08071",
  1045 => x"31177054",
  1046 => x"7f535753",
  1047 => x"83d53f80",
  1048 => x"08538008",
  1049 => x"ff2e81a0",
  1050 => x"3880c1c4",
  1051 => x"08167080",
  1052 => x"c1c40c74",
  1053 => x"7580c280",
  1054 => x"0b88050c",
  1055 => x"74763118",
  1056 => x"70810751",
  1057 => x"5556587b",
  1058 => x"80c2802e",
  1059 => x"839c3879",
  1060 => x"8f2682cb",
  1061 => x"38810b84",
  1062 => x"150c8415",
  1063 => x"08fc0670",
  1064 => x"7a317a72",
  1065 => x"268f7225",
  1066 => x"07525553",
  1067 => x"72802efc",
  1068 => x"f93880db",
  1069 => x"3980089f",
  1070 => x"ff065372",
  1071 => x"feeb3877",
  1072 => x"80c1c40c",
  1073 => x"80c2800b",
  1074 => x"8805087b",
  1075 => x"18810784",
  1076 => x"120c5580",
  1077 => x"c1f00878",
  1078 => x"27863877",
  1079 => x"80c1f00c",
  1080 => x"80c1ec08",
  1081 => x"7827fcac",
  1082 => x"387780c1",
  1083 => x"ec0c8415",
  1084 => x"08fc0670",
  1085 => x"7a317a72",
  1086 => x"268f7225",
  1087 => x"07525553",
  1088 => x"72802efc",
  1089 => x"a5388839",
  1090 => x"80745456",
  1091 => x"fedb397d",
  1092 => x"51829f3f",
  1093 => x"800b800c",
  1094 => x"8f3d0d04",
  1095 => x"73538074",
  1096 => x"24a93872",
  1097 => x"822c8171",
  1098 => x"2b80c284",
  1099 => x"08077080",
  1100 => x"c2800b84",
  1101 => x"050c5d53",
  1102 => x"778c180c",
  1103 => x"7488180c",
  1104 => x"7688190c",
  1105 => x"768c160c",
  1106 => x"f9b73983",
  1107 => x"1470822c",
  1108 => x"81712b80",
  1109 => x"c2840807",
  1110 => x"7080c280",
  1111 => x"0b84050c",
  1112 => x"5e5153d4",
  1113 => x"397b7b06",
  1114 => x"5372fca3",
  1115 => x"38841a7b",
  1116 => x"105c5af1",
  1117 => x"39ff1a81",
  1118 => x"11515af7",
  1119 => x"b9397817",
  1120 => x"79810784",
  1121 => x"190c8c18",
  1122 => x"08881908",
  1123 => x"718c120c",
  1124 => x"88120c59",
  1125 => x"7080c294",
  1126 => x"0c7080c2",
  1127 => x"900c80c2",
  1128 => x"880b8c12",
  1129 => x"0c8c1108",
  1130 => x"88120c74",
  1131 => x"81078412",
  1132 => x"0c741175",
  1133 => x"710c5153",
  1134 => x"f9bd3975",
  1135 => x"17841108",
  1136 => x"81078412",
  1137 => x"0c538c17",
  1138 => x"08881808",
  1139 => x"718c120c",
  1140 => x"88120c58",
  1141 => x"7d5180da",
  1142 => x"3f881754",
  1143 => x"f5cf3972",
  1144 => x"84150cf4",
  1145 => x"1af80670",
  1146 => x"841e0881",
  1147 => x"0607841e",
  1148 => x"0c701d54",
  1149 => x"5b850b84",
  1150 => x"140c850b",
  1151 => x"88140c8f",
  1152 => x"7b27fdcf",
  1153 => x"38881c52",
  1154 => x"7d518290",
  1155 => x"3f80c280",
  1156 => x"0b880508",
  1157 => x"80c1c408",
  1158 => x"5955fdb7",
  1159 => x"397780c1",
  1160 => x"c40c7380",
  1161 => x"c1f40cfc",
  1162 => x"91397284",
  1163 => x"150cfda3",
  1164 => x"390404fd",
  1165 => x"3d0d800b",
  1166 => x"80cacc0c",
  1167 => x"765186cc",
  1168 => x"3f800853",
  1169 => x"8008ff2e",
  1170 => x"88387280",
  1171 => x"0c853d0d",
  1172 => x"0480cacc",
  1173 => x"08547380",
  1174 => x"2ef03875",
  1175 => x"74710c52",
  1176 => x"72800c85",
  1177 => x"3d0d04fb",
  1178 => x"3d0d7770",
  1179 => x"5256c23f",
  1180 => x"80c2800b",
  1181 => x"88050884",
  1182 => x"1108fc06",
  1183 => x"707b319f",
  1184 => x"ef05e080",
  1185 => x"06e08005",
  1186 => x"565653a0",
  1187 => x"80742494",
  1188 => x"38805275",
  1189 => x"51ff9c3f",
  1190 => x"80c28808",
  1191 => x"15537280",
  1192 => x"082e8f38",
  1193 => x"7551ff8a",
  1194 => x"3f805372",
  1195 => x"800c873d",
  1196 => x"0d047330",
  1197 => x"527551fe",
  1198 => x"fa3f8008",
  1199 => x"ff2ea838",
  1200 => x"80c2800b",
  1201 => x"88050875",
  1202 => x"75318107",
  1203 => x"84120c53",
  1204 => x"80c1c408",
  1205 => x"743180c1",
  1206 => x"c40c7551",
  1207 => x"fed43f81",
  1208 => x"0b800c87",
  1209 => x"3d0d0480",
  1210 => x"527551fe",
  1211 => x"c63f80c2",
  1212 => x"800b8805",
  1213 => x"08800871",
  1214 => x"3156538f",
  1215 => x"7525ffa4",
  1216 => x"38800880",
  1217 => x"c1f40831",
  1218 => x"80c1c40c",
  1219 => x"74810784",
  1220 => x"140c7551",
  1221 => x"fe9c3f80",
  1222 => x"53ff9039",
  1223 => x"f63d0d7c",
  1224 => x"7e545b72",
  1225 => x"802e8283",
  1226 => x"387a51fe",
  1227 => x"843ff813",
  1228 => x"84110870",
  1229 => x"fe067013",
  1230 => x"841108fc",
  1231 => x"065d5859",
  1232 => x"545880c2",
  1233 => x"8808752e",
  1234 => x"82de3878",
  1235 => x"84160c80",
  1236 => x"73810654",
  1237 => x"5a727a2e",
  1238 => x"81d53878",
  1239 => x"15841108",
  1240 => x"81065153",
  1241 => x"72a03878",
  1242 => x"17577981",
  1243 => x"e6388815",
  1244 => x"08537280",
  1245 => x"c2882e82",
  1246 => x"f9388c15",
  1247 => x"08708c15",
  1248 => x"0c738812",
  1249 => x"0c567681",
  1250 => x"0784190c",
  1251 => x"76187771",
  1252 => x"0c537981",
  1253 => x"913883ff",
  1254 => x"772781c8",
  1255 => x"3876892a",
  1256 => x"77832a56",
  1257 => x"5372802e",
  1258 => x"bf387686",
  1259 => x"2ab80555",
  1260 => x"847327b4",
  1261 => x"3880db13",
  1262 => x"55947327",
  1263 => x"ab38768c",
  1264 => x"2a80ee05",
  1265 => x"5580d473",
  1266 => x"279e3876",
  1267 => x"8f2a80f7",
  1268 => x"055582d4",
  1269 => x"73279138",
  1270 => x"76922a80",
  1271 => x"fc05558a",
  1272 => x"d4732784",
  1273 => x"3880fe55",
  1274 => x"74101010",
  1275 => x"80c28005",
  1276 => x"88110855",
  1277 => x"5673762e",
  1278 => x"82b33884",
  1279 => x"1408fc06",
  1280 => x"53767327",
  1281 => x"8d388814",
  1282 => x"08547376",
  1283 => x"2e098106",
  1284 => x"ea388c14",
  1285 => x"08708c1a",
  1286 => x"0c74881a",
  1287 => x"0c788812",
  1288 => x"0c56778c",
  1289 => x"150c7a51",
  1290 => x"fc883f8c",
  1291 => x"3d0d0477",
  1292 => x"08787131",
  1293 => x"59770588",
  1294 => x"19085457",
  1295 => x"7280c288",
  1296 => x"2e80e038",
  1297 => x"8c180870",
  1298 => x"8c150c73",
  1299 => x"88120c56",
  1300 => x"fe893988",
  1301 => x"15088c16",
  1302 => x"08708c13",
  1303 => x"0c578817",
  1304 => x"0cfea339",
  1305 => x"76832a70",
  1306 => x"54558075",
  1307 => x"24819838",
  1308 => x"72822c81",
  1309 => x"712b80c2",
  1310 => x"84080780",
  1311 => x"c2800b84",
  1312 => x"050c5374",
  1313 => x"10101080",
  1314 => x"c2800588",
  1315 => x"11085556",
  1316 => x"758c190c",
  1317 => x"7388190c",
  1318 => x"7788170c",
  1319 => x"778c150c",
  1320 => x"ff843981",
  1321 => x"5afdb439",
  1322 => x"78177381",
  1323 => x"06545772",
  1324 => x"98387708",
  1325 => x"78713159",
  1326 => x"77058c19",
  1327 => x"08881a08",
  1328 => x"718c120c",
  1329 => x"88120c57",
  1330 => x"57768107",
  1331 => x"84190c77",
  1332 => x"80c2800b",
  1333 => x"88050c80",
  1334 => x"c1fc0877",
  1335 => x"26fec738",
  1336 => x"80c1f808",
  1337 => x"527a51fa",
  1338 => x"fe3f7a51",
  1339 => x"fac43ffe",
  1340 => x"ba398178",
  1341 => x"8c150c78",
  1342 => x"88150c73",
  1343 => x"8c1a0c73",
  1344 => x"881a0c5a",
  1345 => x"fd803983",
  1346 => x"1570822c",
  1347 => x"81712b80",
  1348 => x"c2840807",
  1349 => x"80c2800b",
  1350 => x"84050c51",
  1351 => x"53741010",
  1352 => x"1080c280",
  1353 => x"05881108",
  1354 => x"5556fee4",
  1355 => x"39745380",
  1356 => x"7524a738",
  1357 => x"72822c81",
  1358 => x"712b80c2",
  1359 => x"84080780",
  1360 => x"c2800b84",
  1361 => x"050c5375",
  1362 => x"8c190c73",
  1363 => x"88190c77",
  1364 => x"88170c77",
  1365 => x"8c150cfd",
  1366 => x"cd398315",
  1367 => x"70822c81",
  1368 => x"712b80c2",
  1369 => x"84080780",
  1370 => x"c2800b84",
  1371 => x"050c5153",
  1372 => x"d639810b",
  1373 => x"800c0480",
  1374 => x"3d0d7281",
  1375 => x"2e893880",
  1376 => x"0b800c82",
  1377 => x"3d0d0473",
  1378 => x"5180f33f",
  1379 => x"fe3d0d80",
  1380 => x"cac40851",
  1381 => x"708a3880",
  1382 => x"cad07080",
  1383 => x"cac40c51",
  1384 => x"70751252",
  1385 => x"52ff5370",
  1386 => x"87fb8080",
  1387 => x"26883870",
  1388 => x"80cac40c",
  1389 => x"71537280",
  1390 => x"0c843d0d",
  1391 => x"04fd3d0d",
  1392 => x"800bba9c",
  1393 => x"08545472",
  1394 => x"812e9a38",
  1395 => x"7380cac8",
  1396 => x"0cdd8c3f",
  1397 => x"dcaa3f80",
  1398 => x"ca885281",
  1399 => x"51df8e3f",
  1400 => x"8008519d",
  1401 => x"3f7280ca",
  1402 => x"c80cdcf3",
  1403 => x"3fdc913f",
  1404 => x"80ca8852",
  1405 => x"8151def5",
  1406 => x"3f800851",
  1407 => x"843f00ff",
  1408 => x"39f73d0d",
  1409 => x"7bbac408",
  1410 => x"82c81108",
  1411 => x"5a545a77",
  1412 => x"802e80d9",
  1413 => x"38818818",
  1414 => x"841908ff",
  1415 => x"0581712b",
  1416 => x"59555980",
  1417 => x"742480e9",
  1418 => x"38807424",
  1419 => x"b5387382",
  1420 => x"2b781188",
  1421 => x"05565681",
  1422 => x"80190877",
  1423 => x"06537280",
  1424 => x"2eb53878",
  1425 => x"16700853",
  1426 => x"53795174",
  1427 => x"0853722d",
  1428 => x"ff14fc17",
  1429 => x"fc177981",
  1430 => x"2c5a5757",
  1431 => x"54738025",
  1432 => x"d6387708",
  1433 => x"5877ffad",
  1434 => x"38bac408",
  1435 => x"53bc1308",
  1436 => x"a5387951",
  1437 => x"ff883f74",
  1438 => x"0853722d",
  1439 => x"ff14fc17",
  1440 => x"fc177981",
  1441 => x"2c5a5757",
  1442 => x"54738025",
  1443 => x"ffa938d2",
  1444 => x"398057ff",
  1445 => x"94397251",
  1446 => x"bc130853",
  1447 => x"722d7951",
  1448 => x"fedc3fff",
  1449 => x"3d0d80ca",
  1450 => x"900bfc05",
  1451 => x"70085252",
  1452 => x"70ff2e91",
  1453 => x"38702dfc",
  1454 => x"12700852",
  1455 => x"5270ff2e",
  1456 => x"098106f1",
  1457 => x"38833d0d",
  1458 => x"0404dbfe",
  1459 => x"3f040000",
  1460 => x"00000040",
  1461 => x"0a677265",
  1462 => x"74682072",
  1463 => x"65676973",
  1464 => x"74657273",
  1465 => x"3a000000",
  1466 => x"0a636f6e",
  1467 => x"74726f6c",
  1468 => x"3a202020",
  1469 => x"20202030",
  1470 => x"78000000",
  1471 => x"0a737461",
  1472 => x"7475733a",
  1473 => x"20202020",
  1474 => x"20202030",
  1475 => x"78000000",
  1476 => x"0a6d6163",
  1477 => x"5f6d7362",
  1478 => x"3a202020",
  1479 => x"20202030",
  1480 => x"78000000",
  1481 => x"0a6d6163",
  1482 => x"5f6c7362",
  1483 => x"3a202020",
  1484 => x"20202030",
  1485 => x"78000000",
  1486 => x"0a6d6469",
  1487 => x"6f5f636f",
  1488 => x"6e74726f",
  1489 => x"6c3a2030",
  1490 => x"78000000",
  1491 => x"0a74785f",
  1492 => x"706f696e",
  1493 => x"7465723a",
  1494 => x"20202030",
  1495 => x"78000000",
  1496 => x"0a72785f",
  1497 => x"706f696e",
  1498 => x"7465723a",
  1499 => x"20202030",
  1500 => x"78000000",
  1501 => x"0a656463",
  1502 => x"6c5f6970",
  1503 => x"3a202020",
  1504 => x"20202030",
  1505 => x"78000000",
  1506 => x"0a686173",
  1507 => x"685f6d73",
  1508 => x"623a2020",
  1509 => x"20202030",
  1510 => x"78000000",
  1511 => x"0a686173",
  1512 => x"685f6c73",
  1513 => x"623a2020",
  1514 => x"20202030",
  1515 => x"78000000",
  1516 => x"0a6d6469",
  1517 => x"6f207068",
  1518 => x"79207265",
  1519 => x"67697374",
  1520 => x"65727300",
  1521 => x"0a206d64",
  1522 => x"696f2070",
  1523 => x"68793a20",
  1524 => x"30780000",
  1525 => x"0a202072",
  1526 => x"65673a20",
  1527 => x"00000000",
  1528 => x"2d3e2030",
  1529 => x"78000000",
  1530 => x"67726574",
  1531 => x"682d3e63",
  1532 => x"6f6e7472",
  1533 => x"6f6c3a20",
  1534 => x"30780000",
  1535 => x"67726574",
  1536 => x"682d3e73",
  1537 => x"74617475",
  1538 => x"73203a20",
  1539 => x"30780000",
  1540 => x"64657363",
  1541 => x"722d3e63",
  1542 => x"6f6e7472",
  1543 => x"6f6c3a20",
  1544 => x"30780000",
  1545 => x"77726974",
  1546 => x"65206164",
  1547 => x"64726573",
  1548 => x"733a2030",
  1549 => x"78000000",
  1550 => x"20206c65",
  1551 => x"6e677468",
  1552 => x"3a203078",
  1553 => x"00000000",
  1554 => x"0a0a0000",
  1555 => x"72656164",
  1556 => x"20206164",
  1557 => x"64726573",
  1558 => x"733a2030",
  1559 => x"78000000",
  1560 => x"20206578",
  1561 => x"70656374",
  1562 => x"3a203078",
  1563 => x"00000000",
  1564 => x"2020676f",
  1565 => x"743a2030",
  1566 => x"78000000",
  1567 => x"20657272",
  1568 => x"6f720000",
  1569 => x"206f6b00",
  1570 => x"70686173",
  1571 => x"65207368",
  1572 => x"69667420",
  1573 => x"202d2020",
  1574 => x"76616c75",
  1575 => x"653a2000",
  1576 => x"20207374",
  1577 => x"61747573",
  1578 => x"3a203078",
  1579 => x"00000000",
  1580 => x"20202020",
  1581 => x"20000000",
  1582 => x"6f6b2020",
  1583 => x"00000000",
  1584 => x"0a307800",
  1585 => x"4641494c",
  1586 => x"00000000",
  1587 => x"44445220",
  1588 => x"6d656d6f",
  1589 => x"72792069",
  1590 => x"6e666f00",
  1591 => x"0a0a6175",
  1592 => x"746f2074",
  1593 => x"5f524552",
  1594 => x"45534820",
  1595 => x"3a000000",
  1596 => x"0a636c6f",
  1597 => x"636b2065",
  1598 => x"6e61626c",
  1599 => x"6520203a",
  1600 => x"30780000",
  1601 => x"0a696e69",
  1602 => x"74616c69",
  1603 => x"7a652020",
  1604 => x"2020203a",
  1605 => x"30780000",
  1606 => x"0a636f6c",
  1607 => x"756d6e20",
  1608 => x"73697a65",
  1609 => x"2020203a",
  1610 => x"00000000",
  1611 => x"0a62616e",
  1612 => x"6b73697a",
  1613 => x"65202020",
  1614 => x"2020203a",
  1615 => x"00000000",
  1616 => x"4d627974",
  1617 => x"65000000",
  1618 => x"0a745f52",
  1619 => x"43442020",
  1620 => x"20202020",
  1621 => x"2020203a",
  1622 => x"00000000",
  1623 => x"0a745f52",
  1624 => x"46432020",
  1625 => x"20202020",
  1626 => x"2020203a",
  1627 => x"00000000",
  1628 => x"0a745f52",
  1629 => x"50202020",
  1630 => x"20202020",
  1631 => x"2020203a",
  1632 => x"00000000",
  1633 => x"0a726566",
  1634 => x"72657368",
  1635 => x"20656e2e",
  1636 => x"2020203a",
  1637 => x"30780000",
  1638 => x"0a0a4444",
  1639 => x"52206672",
  1640 => x"65717565",
  1641 => x"6e637920",
  1642 => x"3a000000",
  1643 => x"0a444452",
  1644 => x"20646174",
  1645 => x"61207769",
  1646 => x"6474683a",
  1647 => x"00000000",
  1648 => x"0a6d6f62",
  1649 => x"696c6520",
  1650 => x"73757070",
  1651 => x"6f72743a",
  1652 => x"30780000",
  1653 => x"0a0a7374",
  1654 => x"61747573",
  1655 => x"20726561",
  1656 => x"64202020",
  1657 => x"3a307800",
  1658 => x"0a0a7365",
  1659 => x"6c662072",
  1660 => x"65667265",
  1661 => x"73682020",
  1662 => x"3a000000",
  1663 => x"20353132",
  1664 => x"00000000",
  1665 => x"34303639",
  1666 => x"00000000",
  1667 => x"312f3800",
  1668 => x"20617272",
  1669 => x"61790000",
  1670 => x"0a74656d",
  1671 => x"702d636f",
  1672 => x"6d702072",
  1673 => x"6566723a",
  1674 => x"00000000",
  1675 => x"c2b04300",
  1676 => x"0a647269",
  1677 => x"76652073",
  1678 => x"7472656e",
  1679 => x"6774683a",
  1680 => x"00000000",
  1681 => x"0a706f77",
  1682 => x"65722073",
  1683 => x"6176696e",
  1684 => x"6720203a",
  1685 => x"00000000",
  1686 => x"756e6b6e",
  1687 => x"6f776e00",
  1688 => x"0a745f58",
  1689 => x"50202020",
  1690 => x"20202020",
  1691 => x"2020203a",
  1692 => x"00000000",
  1693 => x"0a745f58",
  1694 => x"53522020",
  1695 => x"20202020",
  1696 => x"2020203a",
  1697 => x"00000000",
  1698 => x"0a745f43",
  1699 => x"4b452020",
  1700 => x"20202020",
  1701 => x"2020203a",
  1702 => x"00000000",
  1703 => x"0a434153",
  1704 => x"206c6174",
  1705 => x"656e6379",
  1706 => x"2020203a",
  1707 => x"00000000",
  1708 => x"0a6d6f62",
  1709 => x"696c6520",
  1710 => x"656e6162",
  1711 => x"6c65643a",
  1712 => x"30780000",
  1713 => x"0a0a7068",
  1714 => x"7920636f",
  1715 => x"6e666967",
  1716 => x"20302020",
  1717 => x"3a307800",
  1718 => x"0a0a7068",
  1719 => x"7920636f",
  1720 => x"6e666967",
  1721 => x"20312020",
  1722 => x"3a307800",
  1723 => x"31303234",
  1724 => x"00000000",
  1725 => x"32303438",
  1726 => x"00000000",
  1727 => x"66756c6c",
  1728 => x"00000000",
  1729 => x"37300000",
  1730 => x"64656570",
  1731 => x"20706f77",
  1732 => x"65722064",
  1733 => x"6f776e00",
  1734 => x"636c6f63",
  1735 => x"6b207374",
  1736 => x"6f700000",
  1737 => x"73656c66",
  1738 => x"20726566",
  1739 => x"72657368",
  1740 => x"00000000",
  1741 => x"706f7765",
  1742 => x"7220646f",
  1743 => x"776e0000",
  1744 => x"6e6f6e65",
  1745 => x"00000000",
  1746 => x"312f3200",
  1747 => x"312f3400",
  1748 => x"312f3100",
  1749 => x"332f3400",
  1750 => x"38350000",
  1751 => x"34350000",
  1752 => x"68616c66",
  1753 => x"00000000",
  1754 => x"31350000",
  1755 => x"61646472",
  1756 => x"6573733a",
  1757 => x"20307800",
  1758 => x"20646174",
  1759 => x"613a2030",
  1760 => x"78000000",
  1761 => x"0a0a4443",
  1762 => x"4d207068",
  1763 => x"61736520",
  1764 => x"73686966",
  1765 => x"74207465",
  1766 => x"7374696e",
  1767 => x"67000000",
  1768 => x"0a696e69",
  1769 => x"7469616c",
  1770 => x"3a200000",
  1771 => x"09000000",
  1772 => x"20202020",
  1773 => x"00000000",
  1774 => x"6c6f7720",
  1775 => x"666f756e",
  1776 => x"64000000",
  1777 => x"68696768",
  1778 => x"20666f75",
  1779 => x"6e640000",
  1780 => x"0a6c6f77",
  1781 => x"3a202020",
  1782 => x"20202020",
  1783 => x"20200000",
  1784 => x"0a686967",
  1785 => x"683a2020",
  1786 => x"20202020",
  1787 => x"20200000",
  1788 => x"0a646966",
  1789 => x"663a2020",
  1790 => x"20202020",
  1791 => x"20200000",
  1792 => x"0a6d696e",
  1793 => x"5f657272",
  1794 => x"3a202020",
  1795 => x"20200000",
  1796 => x"0a6d696e",
  1797 => x"5f657272",
  1798 => x"5f706f73",
  1799 => x"3a200000",
  1800 => x"676f206d",
  1801 => x"696e5f65",
  1802 => x"72726f72",
  1803 => x"00000000",
  1804 => x"0a66696e",
  1805 => x"616c3a20",
  1806 => x"20202020",
  1807 => x"20200000",
  1808 => x"6c6f7720",
  1809 => x"4e4f5420",
  1810 => x"666f756e",
  1811 => x"64000000",
  1812 => x"68696768",
  1813 => x"204e4f54",
  1814 => x"20666f75",
  1815 => x"6e640000",
  1816 => x"676f207a",
  1817 => x"65726f00",
  1818 => x"64617461",
  1819 => x"2076616c",
  1820 => x"69640000",
  1821 => x"6c6f7720",
  1822 => x"20666f75",
  1823 => x"6e640000",
  1824 => x"0a646966",
  1825 => x"662f323a",
  1826 => x"20202020",
  1827 => x"20200000",
  1828 => x"6c6f7720",
  1829 => x"204e4f54",
  1830 => x"20666f75",
  1831 => x"6e640000",
  1832 => x"64617461",
  1833 => x"204e4f54",
  1834 => x"2076616c",
  1835 => x"69640000",
  1836 => x"74657374",
  1837 => x"2e632000",
  1838 => x"286f6e20",
  1839 => x"73696d29",
  1840 => x"0a000000",
  1841 => x"286f6e20",
  1842 => x"68617264",
  1843 => x"77617265",
  1844 => x"290a0000",
  1845 => x"636f6d70",
  1846 => x"696c6564",
  1847 => x"3a204a61",
  1848 => x"6e203131",
  1849 => x"20323031",
  1850 => x"31202030",
  1851 => x"373a3438",
  1852 => x"3a33390a",
  1853 => x"00000000",
  1854 => x"43000000",
  1855 => x"64756d6d",
  1856 => x"792e6578",
  1857 => x"65000000",
  1858 => x"00ffffff",
  1859 => x"ff00ffff",
  1860 => x"ffff00ff",
  1861 => x"ffffff00",
  1862 => x"00000000",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00002518",
  1866 => x"fff00000",
  1867 => x"80000d00",
  1868 => x"80000800",
  1869 => x"80000600",
  1870 => x"80000300",
  1871 => x"80000200",
  1872 => x"80000100",
  1873 => x"00001d48",
  1874 => x"00000000",
  1875 => x"00001fb0",
  1876 => x"0000200c",
  1877 => x"00002068",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00000000",
  1887 => x"00001cf8",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000001",
  1917 => x"330eabcd",
  1918 => x"1234e66d",
  1919 => x"deec0005",
  1920 => x"000b0000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"00000000",
  1931 => x"00000000",
  1932 => x"00000000",
  1933 => x"00000000",
  1934 => x"00000000",
  1935 => x"00000000",
  1936 => x"00000000",
  1937 => x"00000000",
  1938 => x"00000000",
  1939 => x"00000000",
  1940 => x"00000000",
  1941 => x"00000000",
  1942 => x"00000000",
  1943 => x"00000000",
  1944 => x"00000000",
  1945 => x"00000000",
  1946 => x"00000000",
  1947 => x"00000000",
  1948 => x"00000000",
  1949 => x"00000000",
  1950 => x"00000000",
  1951 => x"00000000",
  1952 => x"00000000",
  1953 => x"00000000",
  1954 => x"00000000",
  1955 => x"00000000",
  1956 => x"00000000",
  1957 => x"00000000",
  1958 => x"00000000",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00000000",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00000000",
  1984 => x"00000000",
  1985 => x"00000000",
  1986 => x"00000000",
  1987 => x"00000000",
  1988 => x"00000000",
  1989 => x"00000000",
  1990 => x"00000000",
  1991 => x"00000000",
  1992 => x"00000000",
  1993 => x"00000000",
  1994 => x"00000000",
  1995 => x"00000000",
  1996 => x"00000000",
  1997 => x"00000000",
  1998 => x"00000000",
  1999 => x"00000000",
  2000 => x"00000000",
  2001 => x"00000000",
  2002 => x"00000000",
  2003 => x"00000000",
  2004 => x"00000000",
  2005 => x"00000000",
  2006 => x"00000000",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00000000",
  2010 => x"00000000",
  2011 => x"00000000",
  2012 => x"00000000",
  2013 => x"00000000",
  2014 => x"00000000",
  2015 => x"00000000",
  2016 => x"00000000",
  2017 => x"00000000",
  2018 => x"00000000",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00000000",
  2026 => x"00000000",
  2027 => x"00000000",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000000",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"00000000",
  2049 => x"00000000",
  2050 => x"00000000",
  2051 => x"00000000",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"ffffffff",
  2110 => x"00000000",
  2111 => x"00020000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00002100",
  2115 => x"00002100",
  2116 => x"00002108",
  2117 => x"00002108",
  2118 => x"00002110",
  2119 => x"00002110",
  2120 => x"00002118",
  2121 => x"00002118",
  2122 => x"00002120",
  2123 => x"00002120",
  2124 => x"00002128",
  2125 => x"00002128",
  2126 => x"00002130",
  2127 => x"00002130",
  2128 => x"00002138",
  2129 => x"00002138",
  2130 => x"00002140",
  2131 => x"00002140",
  2132 => x"00002148",
  2133 => x"00002148",
  2134 => x"00002150",
  2135 => x"00002150",
  2136 => x"00002158",
  2137 => x"00002158",
  2138 => x"00002160",
  2139 => x"00002160",
  2140 => x"00002168",
  2141 => x"00002168",
  2142 => x"00002170",
  2143 => x"00002170",
  2144 => x"00002178",
  2145 => x"00002178",
  2146 => x"00002180",
  2147 => x"00002180",
  2148 => x"00002188",
  2149 => x"00002188",
  2150 => x"00002190",
  2151 => x"00002190",
  2152 => x"00002198",
  2153 => x"00002198",
  2154 => x"000021a0",
  2155 => x"000021a0",
  2156 => x"000021a8",
  2157 => x"000021a8",
  2158 => x"000021b0",
  2159 => x"000021b0",
  2160 => x"000021b8",
  2161 => x"000021b8",
  2162 => x"000021c0",
  2163 => x"000021c0",
  2164 => x"000021c8",
  2165 => x"000021c8",
  2166 => x"000021d0",
  2167 => x"000021d0",
  2168 => x"000021d8",
  2169 => x"000021d8",
  2170 => x"000021e0",
  2171 => x"000021e0",
  2172 => x"000021e8",
  2173 => x"000021e8",
  2174 => x"000021f0",
  2175 => x"000021f0",
  2176 => x"000021f8",
  2177 => x"000021f8",
  2178 => x"00002200",
  2179 => x"00002200",
  2180 => x"00002208",
  2181 => x"00002208",
  2182 => x"00002210",
  2183 => x"00002210",
  2184 => x"00002218",
  2185 => x"00002218",
  2186 => x"00002220",
  2187 => x"00002220",
  2188 => x"00002228",
  2189 => x"00002228",
  2190 => x"00002230",
  2191 => x"00002230",
  2192 => x"00002238",
  2193 => x"00002238",
  2194 => x"00002240",
  2195 => x"00002240",
  2196 => x"00002248",
  2197 => x"00002248",
  2198 => x"00002250",
  2199 => x"00002250",
  2200 => x"00002258",
  2201 => x"00002258",
  2202 => x"00002260",
  2203 => x"00002260",
  2204 => x"00002268",
  2205 => x"00002268",
  2206 => x"00002270",
  2207 => x"00002270",
  2208 => x"00002278",
  2209 => x"00002278",
  2210 => x"00002280",
  2211 => x"00002280",
  2212 => x"00002288",
  2213 => x"00002288",
  2214 => x"00002290",
  2215 => x"00002290",
  2216 => x"00002298",
  2217 => x"00002298",
  2218 => x"000022a0",
  2219 => x"000022a0",
  2220 => x"000022a8",
  2221 => x"000022a8",
  2222 => x"000022b0",
  2223 => x"000022b0",
  2224 => x"000022b8",
  2225 => x"000022b8",
  2226 => x"000022c0",
  2227 => x"000022c0",
  2228 => x"000022c8",
  2229 => x"000022c8",
  2230 => x"000022d0",
  2231 => x"000022d0",
  2232 => x"000022d8",
  2233 => x"000022d8",
  2234 => x"000022e0",
  2235 => x"000022e0",
  2236 => x"000022e8",
  2237 => x"000022e8",
  2238 => x"000022f0",
  2239 => x"000022f0",
  2240 => x"000022f8",
  2241 => x"000022f8",
  2242 => x"00002300",
  2243 => x"00002300",
  2244 => x"00002308",
  2245 => x"00002308",
  2246 => x"00002310",
  2247 => x"00002310",
  2248 => x"00002318",
  2249 => x"00002318",
  2250 => x"00002320",
  2251 => x"00002320",
  2252 => x"00002328",
  2253 => x"00002328",
  2254 => x"00002330",
  2255 => x"00002330",
  2256 => x"00002338",
  2257 => x"00002338",
  2258 => x"00002340",
  2259 => x"00002340",
  2260 => x"00002348",
  2261 => x"00002348",
  2262 => x"00002350",
  2263 => x"00002350",
  2264 => x"00002358",
  2265 => x"00002358",
  2266 => x"00002360",
  2267 => x"00002360",
  2268 => x"00002368",
  2269 => x"00002368",
  2270 => x"00002370",
  2271 => x"00002370",
  2272 => x"00002378",
  2273 => x"00002378",
  2274 => x"00002380",
  2275 => x"00002380",
  2276 => x"00002388",
  2277 => x"00002388",
  2278 => x"00002390",
  2279 => x"00002390",
  2280 => x"00002398",
  2281 => x"00002398",
  2282 => x"000023a0",
  2283 => x"000023a0",
  2284 => x"000023a8",
  2285 => x"000023a8",
  2286 => x"000023b0",
  2287 => x"000023b0",
  2288 => x"000023b8",
  2289 => x"000023b8",
  2290 => x"000023c0",
  2291 => x"000023c0",
  2292 => x"000023c8",
  2293 => x"000023c8",
  2294 => x"000023d0",
  2295 => x"000023d0",
  2296 => x"000023d8",
  2297 => x"000023d8",
  2298 => x"000023e0",
  2299 => x"000023e0",
  2300 => x"000023e8",
  2301 => x"000023e8",
  2302 => x"000023f0",
  2303 => x"000023f0",
  2304 => x"000023f8",
  2305 => x"000023f8",
  2306 => x"00002400",
  2307 => x"00002400",
  2308 => x"00002408",
  2309 => x"00002408",
  2310 => x"00002410",
  2311 => x"00002410",
  2312 => x"00002418",
  2313 => x"00002418",
  2314 => x"00002420",
  2315 => x"00002420",
  2316 => x"00002428",
  2317 => x"00002428",
  2318 => x"00002430",
  2319 => x"00002430",
  2320 => x"00002438",
  2321 => x"00002438",
  2322 => x"00002440",
  2323 => x"00002440",
  2324 => x"00002448",
  2325 => x"00002448",
  2326 => x"00002450",
  2327 => x"00002450",
  2328 => x"00002458",
  2329 => x"00002458",
  2330 => x"00002460",
  2331 => x"00002460",
  2332 => x"00002468",
  2333 => x"00002468",
  2334 => x"00002470",
  2335 => x"00002470",
  2336 => x"00002478",
  2337 => x"00002478",
  2338 => x"00002480",
  2339 => x"00002480",
  2340 => x"00002488",
  2341 => x"00002488",
  2342 => x"00002490",
  2343 => x"00002490",
  2344 => x"00002498",
  2345 => x"00002498",
  2346 => x"000024a0",
  2347 => x"000024a0",
  2348 => x"000024a8",
  2349 => x"000024a8",
  2350 => x"000024b0",
  2351 => x"000024b0",
  2352 => x"000024b8",
  2353 => x"000024b8",
  2354 => x"000024c0",
  2355 => x"000024c0",
  2356 => x"000024c8",
  2357 => x"000024c8",
  2358 => x"000024d0",
  2359 => x"000024d0",
  2360 => x"000024d8",
  2361 => x"000024d8",
  2362 => x"000024e0",
  2363 => x"000024e0",
  2364 => x"000024e8",
  2365 => x"000024e8",
  2366 => x"000024f0",
  2367 => x"000024f0",
  2368 => x"000024f8",
  2369 => x"000024f8",
  2370 => x"00001cfc",
  2371 => x"ffffffff",
  2372 => x"00000000",
  2373 => x"ffffffff",
  2374 => x"00000000",
  2375 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
