library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


library zylin;
use zylin.zpu_config.all;
use zylin.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);


--shared variable ram : ram_type :=
signal ram : ram_type :=
(
0 => x"800b0b0b",
1 => x"0b0b8070",
2 => x"0b0b818a",
3 => x"dc0c3a0b",
4 => x"0b80dab4",
5 => x"04000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"80db972d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b0b2a",
20 => x"83ffff06",
21 => x"52810504",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b0b2b09",
29 => x"067383ff",
30 => x"ff0b0b0b",
31 => x"0b83a704",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53518105",
38 => x"04000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51810504",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53518105",
55 => x"04000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51810504",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"72ff0571",
65 => x"81050673",
66 => x"ff050972",
67 => x"74058005",
68 => x"06075350",
69 => x"50040000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b8c",
73 => x"f8040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535181",
82 => x"05040000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"81050400",
102 => x"00000000",
103 => x"00000000",
104 => x"71718105",
105 => x"53510406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515181",
111 => x"05040000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51810504",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53518105",
125 => x"04000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52810504",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"81050409",
139 => x"81058305",
140 => x"1010102b",
141 => x"0772fc06",
142 => x"0c515181",
143 => x"05040000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535181",
147 => x"05040000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"81050400",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b818a",
162 => x"88738306",
163 => x"10100508",
164 => x"067381ff",
165 => x"06738306",
166 => x"0b0b0b84",
167 => x"ab040000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0bb3",
171 => x"912d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c810551",
175 => x"04000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0bb4",
179 => x"8a2d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c810551",
183 => x"04000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547181",
188 => x"05067309",
189 => x"72740580",
190 => x"05060753",
191 => x"50500400",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"81050673",
197 => x"09727405",
198 => x"80050607",
199 => x"53505004",
200 => x"05800504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"818ad80c",
210 => x"51810504",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"72830610",
217 => x"10728306",
218 => x"0710100b",
219 => x"0b818a98",
220 => x"05080400",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"81050400",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"71710571",
249 => x"81055351",
250 => x"04000000",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"8db33f80",
257 => x"f39e3f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51810504",
267 => x"72fc0608",
268 => x"81ff0a06",
269 => x"72fc0670",
270 => x"5408fe80",
271 => x"0a060772",
272 => x"0c515181",
273 => x"050472fc",
274 => x"06080a10",
275 => x"10101010",
276 => x"1010100a",
277 => x"87fc8080",
278 => x"0672fc06",
279 => x"08f883ff",
280 => x"ff060772",
281 => x"fc060c51",
282 => x"51810504",
283 => x"72fc0608",
284 => x"0a101010",
285 => x"10101010",
286 => x"10101010",
287 => x"10101010",
288 => x"100a83fe",
289 => x"800672fc",
290 => x"0608fc81",
291 => x"ff060772",
292 => x"fc060c51",
293 => x"51810504",
294 => x"72fc0608",
295 => x"0a101010",
296 => x"10101010",
297 => x"10101010",
298 => x"10101010",
299 => x"10101010",
300 => x"10101010",
301 => x"100a81ff",
302 => x"0672fc06",
303 => x"08fe8006",
304 => x"0772fc06",
305 => x"0c515181",
306 => x"050472fc",
307 => x"06081010",
308 => x"10101010",
309 => x"101081ff",
310 => x"0a0672fc",
311 => x"0608fe80",
312 => x"0a060772",
313 => x"fc060c51",
314 => x"51810504",
315 => x"72fc0608",
316 => x"87fc8080",
317 => x"0672fc06",
318 => x"705408f8",
319 => x"83ffff06",
320 => x"07720c51",
321 => x"51810504",
322 => x"72fc0608",
323 => x"0a101010",
324 => x"10101010",
325 => x"100a83fe",
326 => x"800672fc",
327 => x"0608fc81",
328 => x"ff060772",
329 => x"fc060c51",
330 => x"51810504",
331 => x"72fc0608",
332 => x"0a101010",
333 => x"10101010",
334 => x"10101010",
335 => x"10101010",
336 => x"100a81ff",
337 => x"0672fc06",
338 => x"08fe8006",
339 => x"0772fc06",
340 => x"0c515181",
341 => x"050472fc",
342 => x"06081010",
343 => x"10101010",
344 => x"10101010",
345 => x"10101010",
346 => x"101081ff",
347 => x"0a0672fc",
348 => x"0608fe80",
349 => x"0a060772",
350 => x"fc060c51",
351 => x"51810504",
352 => x"72fc0608",
353 => x"10101010",
354 => x"10101010",
355 => x"87fc8080",
356 => x"0672fc06",
357 => x"08f883ff",
358 => x"ff060772",
359 => x"fc060c51",
360 => x"51810504",
361 => x"72fc0608",
362 => x"83fe8006",
363 => x"72fc0670",
364 => x"5408fc81",
365 => x"ff060772",
366 => x"0c515181",
367 => x"050472fc",
368 => x"06080a10",
369 => x"10101010",
370 => x"1010100a",
371 => x"81ff0672",
372 => x"fc0608fe",
373 => x"80060772",
374 => x"fc060c51",
375 => x"51810504",
376 => x"72fc0608",
377 => x"10101010",
378 => x"10101010",
379 => x"10101010",
380 => x"10101010",
381 => x"10101010",
382 => x"10101010",
383 => x"81ff0a06",
384 => x"72fc0608",
385 => x"fe800a06",
386 => x"0772fc06",
387 => x"0c515181",
388 => x"050472fc",
389 => x"06081010",
390 => x"10101010",
391 => x"10101010",
392 => x"10101010",
393 => x"101087fc",
394 => x"80800672",
395 => x"fc0608f8",
396 => x"83ffff06",
397 => x"0772fc06",
398 => x"0c515181",
399 => x"050472fc",
400 => x"06081010",
401 => x"10101010",
402 => x"101083fe",
403 => x"800672fc",
404 => x"0608fc81",
405 => x"ff060772",
406 => x"fc060c51",
407 => x"51810504",
408 => x"72fc0608",
409 => x"81ff0672",
410 => x"fc067054",
411 => x"08fe8006",
412 => x"07720c51",
413 => x"51810504",
414 => x"72728072",
415 => x"8106ff05",
416 => x"09720605",
417 => x"71105272",
418 => x"0a100a53",
419 => x"728106ff",
420 => x"05097206",
421 => x"05711052",
422 => x"720a100a",
423 => x"53728106",
424 => x"ff050972",
425 => x"06057110",
426 => x"52720a10",
427 => x"0a537281",
428 => x"06ff0509",
429 => x"72060571",
430 => x"1052720a",
431 => x"100a5372",
432 => x"8106ff05",
433 => x"09720605",
434 => x"71105272",
435 => x"0a100a53",
436 => x"728106ff",
437 => x"05097206",
438 => x"05711052",
439 => x"720a100a",
440 => x"53728106",
441 => x"ff050972",
442 => x"06057110",
443 => x"52720a10",
444 => x"0a537281",
445 => x"06ff0509",
446 => x"72060571",
447 => x"1052720a",
448 => x"100a5372",
449 => x"83a13772",
450 => x"8106ff05",
451 => x"09720605",
452 => x"71105272",
453 => x"0a100a53",
454 => x"728106ff",
455 => x"05097206",
456 => x"05711052",
457 => x"720a100a",
458 => x"53728106",
459 => x"ff050972",
460 => x"06057110",
461 => x"52720a10",
462 => x"0a537281",
463 => x"06ff0509",
464 => x"72060571",
465 => x"1052720a",
466 => x"100a5372",
467 => x"8106ff05",
468 => x"09720605",
469 => x"71105272",
470 => x"0a100a53",
471 => x"728106ff",
472 => x"05097206",
473 => x"05711052",
474 => x"720a100a",
475 => x"53728106",
476 => x"ff050972",
477 => x"06057110",
478 => x"52720a10",
479 => x"0a537281",
480 => x"06ff0509",
481 => x"72060571",
482 => x"1052720a",
483 => x"100a5372",
484 => x"82953772",
485 => x"8106ff05",
486 => x"09720605",
487 => x"71105272",
488 => x"0a100a53",
489 => x"728106ff",
490 => x"05097206",
491 => x"05711052",
492 => x"720a100a",
493 => x"53728106",
494 => x"ff050972",
495 => x"06057110",
496 => x"52720a10",
497 => x"0a537281",
498 => x"06ff0509",
499 => x"72060571",
500 => x"1052720a",
501 => x"100a5372",
502 => x"8106ff05",
503 => x"09720605",
504 => x"71105272",
505 => x"0a100a53",
506 => x"728106ff",
507 => x"05097206",
508 => x"05711052",
509 => x"720a100a",
510 => x"53728106",
511 => x"ff050972",
512 => x"06057110",
513 => x"52720a10",
514 => x"0a537281",
515 => x"06ff0509",
516 => x"72060571",
517 => x"1052720a",
518 => x"100a5372",
519 => x"81893772",
520 => x"8106ff05",
521 => x"09720605",
522 => x"71105272",
523 => x"0a100a53",
524 => x"728106ff",
525 => x"05097206",
526 => x"05711052",
527 => x"720a100a",
528 => x"53728106",
529 => x"ff050972",
530 => x"06057110",
531 => x"52720a10",
532 => x"0a537281",
533 => x"06ff0509",
534 => x"72060571",
535 => x"1052720a",
536 => x"100a5372",
537 => x"8106ff05",
538 => x"09720605",
539 => x"71105272",
540 => x"0a100a53",
541 => x"728106ff",
542 => x"05097206",
543 => x"05711052",
544 => x"720a100a",
545 => x"53728106",
546 => x"ff050972",
547 => x"06057110",
548 => x"52720a10",
549 => x"0a537281",
550 => x"06ff0509",
551 => x"72060571",
552 => x"1052720a",
553 => x"100a5351",
554 => x"51535181",
555 => x"05043c04",
556 => x"70700b0b",
557 => x"819acc08",
558 => x"52841208",
559 => x"70810651",
560 => x"51700970",
561 => x"81050906",
562 => x"0a098106",
563 => x"ff0509e9",
564 => x"0bf70506",
565 => x"84010505",
566 => x"04710881",
567 => x"ff06800c",
568 => x"50500470",
569 => x"700b0b81",
570 => x"9acc0852",
571 => x"84120870",
572 => x"0a100a70",
573 => x"81065151",
574 => x"51700970",
575 => x"81050906",
576 => x"0a098106",
577 => x"ff0509e4",
578 => x"0bf70506",
579 => x"84010505",
580 => x"0473720c",
581 => x"50500481",
582 => x"8ad80809",
583 => x"70810509",
584 => x"060a8106",
585 => x"ff0509b0",
586 => x"0bf70506",
587 => x"84010505",
588 => x"04838080",
589 => x"0b0b0b81",
590 => x"9acc0c82",
591 => x"a0800b0b",
592 => x"0b819ad0",
593 => x"0c829080",
594 => x"0b819ae0",
595 => x"0c0b0b81",
596 => x"9ad40b81",
597 => x"9ae40c04",
598 => x"f8808080",
599 => x"a40b0b0b",
600 => x"819acc0c",
601 => x"f8808082",
602 => x"800b0b0b",
603 => x"819ad00c",
604 => x"f8808084",
605 => x"800b819a",
606 => x"e00cf880",
607 => x"8080940b",
608 => x"819ae40c",
609 => x"f8808080",
610 => x"9c0b819a",
611 => x"dc0cf880",
612 => x"8080a00b",
613 => x"819ae80c",
614 => x"04f23d0d",
615 => x"600b0b81",
616 => x"9ad00856",
617 => x"5d82750c",
618 => x"8059805a",
619 => x"800b8f3d",
620 => x"71101017",
621 => x"70085957",
622 => x"5d5b8076",
623 => x"81ff067c",
624 => x"832b5658",
625 => x"5276537b",
626 => x"519ede3f",
627 => x"7d7f7a72",
628 => x"077c7207",
629 => x"71716081",
630 => x"05415f5d",
631 => x"5b595755",
632 => x"7a8724ff",
633 => x"050980ce",
634 => x"0bf70506",
635 => x"84010505",
636 => x"040b0b81",
637 => x"9ad0087b",
638 => x"10101170",
639 => x"08585155",
640 => x"807681ff",
641 => x"067c832b",
642 => x"56585276",
643 => x"537b519e",
644 => x"983f7d7f",
645 => x"7a72077c",
646 => x"72077171",
647 => x"60810541",
648 => x"5f5d5b59",
649 => x"5755877b",
650 => x"25ff0509",
651 => x"c40bf705",
652 => x"06840105",
653 => x"0504767d",
654 => x"0c77841e",
655 => x"0c7c800c",
656 => x"903d0d04",
657 => x"7070819a",
658 => x"d8335170",
659 => x"09708105",
660 => x"09060a09",
661 => x"8106ff05",
662 => x"0980d60b",
663 => x"f7050684",
664 => x"01050504",
665 => x"818ae408",
666 => x"70085252",
667 => x"70097081",
668 => x"0509060a",
669 => x"8106ff05",
670 => x"09b10bf7",
671 => x"05068401",
672 => x"05050484",
673 => x"12818ae4",
674 => x"0c702d81",
675 => x"8ae40870",
676 => x"08525270",
677 => x"09708105",
678 => x"09060a09",
679 => x"8106ff05",
680 => x"09e10bf7",
681 => x"05068401",
682 => x"05050481",
683 => x"0b819ad8",
684 => x"34505004",
685 => x"04700b0b",
686 => x"819ac808",
687 => x"09708105",
688 => x"09060a81",
689 => x"06ff0509",
690 => x"a50bf705",
691 => x"06840105",
692 => x"05040b0b",
693 => x"0b0b8009",
694 => x"70810509",
695 => x"060a0981",
696 => x"06ff0509",
697 => x"8b0bf705",
698 => x"06840105",
699 => x"05045004",
700 => x"0b0b819a",
701 => x"c8510b0b",
702 => x"0bea853f",
703 => x"50040470",
704 => x"70028f05",
705 => x"33527109",
706 => x"81058a05",
707 => x"09708105",
708 => x"09060a81",
709 => x"06ff0509",
710 => x"910bf705",
711 => x"06840105",
712 => x"05047151",
713 => x"fbbd3f50",
714 => x"50048d51",
715 => x"fbb53f71",
716 => x"51fbb03f",
717 => x"505004cd",
718 => x"3d0db63d",
719 => x"70708405",
720 => x"520895ff",
721 => x"5d56a63d",
722 => x"5f5d8075",
723 => x"70810557",
724 => x"33765c55",
725 => x"59730981",
726 => x"05790509",
727 => x"70810509",
728 => x"060a8106",
729 => x"ff050981",
730 => x"ad0bf705",
731 => x"06840105",
732 => x"05048f3d",
733 => x"5c730981",
734 => x"05a50509",
735 => x"70810509",
736 => x"060a0981",
737 => x"06ff0509",
738 => x"819c0bf7",
739 => x"05068401",
740 => x"05050479",
741 => x"7081055b",
742 => x"33547309",
743 => x"810580e4",
744 => x"05097081",
745 => x"0509060a",
746 => x"8106ff05",
747 => x"0982ee0b",
748 => x"f7050684",
749 => x"01050504",
750 => x"7380e424",
751 => x"ff050981",
752 => x"900bf705",
753 => x"06840105",
754 => x"05047309",
755 => x"810580e3",
756 => x"05097081",
757 => x"0509060a",
758 => x"8106ff05",
759 => x"09bf0bf7",
760 => x"05068401",
761 => x"05050480",
762 => x"52a5517a",
763 => x"2d805273",
764 => x"517a2d82",
765 => x"19597970",
766 => x"81055b33",
767 => x"54730970",
768 => x"81050906",
769 => x"0a098106",
770 => x"ff0509fe",
771 => x"e80bf705",
772 => x"06840105",
773 => x"05047880",
774 => x"0cb53d0d",
775 => x"047c841e",
776 => x"83123356",
777 => x"5e578052",
778 => x"73517a2d",
779 => x"81197a70",
780 => x"81055c33",
781 => x"55597309",
782 => x"70810509",
783 => x"060a0981",
784 => x"06ff0509",
785 => x"feaf0bf7",
786 => x"05068401",
787 => x"050504c6",
788 => x"39730981",
789 => x"0580f305",
790 => x"09708105",
791 => x"09060a09",
792 => x"8106ff05",
793 => x"09ff800b",
794 => x"f7050684",
795 => x"01050504",
796 => x"7c841e71",
797 => x"08595e56",
798 => x"80773356",
799 => x"56740981",
800 => x"05760509",
801 => x"70810509",
802 => x"060a8106",
803 => x"ff0509aa",
804 => x"0bf70506",
805 => x"84010505",
806 => x"04811670",
807 => x"1870335a",
808 => x"55567709",
809 => x"70810509",
810 => x"060a0981",
811 => x"06ff0509",
812 => x"e80bf705",
813 => x"06840105",
814 => x"0504ff16",
815 => x"55807625",
816 => x"ff0509fe",
817 => x"b10bf705",
818 => x"06840105",
819 => x"05047670",
820 => x"81055833",
821 => x"58805277",
822 => x"517a2d81",
823 => x"1975ff17",
824 => x"57575980",
825 => x"7625ff05",
826 => x"09fe8b0b",
827 => x"f7050684",
828 => x"01050504",
829 => x"76708105",
830 => x"58335880",
831 => x"5277517a",
832 => x"2d811975",
833 => x"ff175757",
834 => x"59758024",
835 => x"ff0509ff",
836 => x"bd0bf705",
837 => x"06840105",
838 => x"0504fdda",
839 => x"397c841e",
840 => x"71087071",
841 => x"9f2c5953",
842 => x"595e5680",
843 => x"7524ff05",
844 => x"0981f80b",
845 => x"f7050684",
846 => x"01050504",
847 => x"757e7d58",
848 => x"59558057",
849 => x"74098105",
850 => x"77050970",
851 => x"81050906",
852 => x"0a098106",
853 => x"ff050980",
854 => x"f40bf705",
855 => x"06840105",
856 => x"0504b07c",
857 => x"3402b905",
858 => x"567b0981",
859 => x"05760509",
860 => x"70810509",
861 => x"060a8106",
862 => x"ff0509b3",
863 => x"0bf70506",
864 => x"84010505",
865 => x"04ff1656",
866 => x"75787081",
867 => x"055a3b81",
868 => x"17577b09",
869 => x"81057605",
870 => x"09708105",
871 => x"09060a09",
872 => x"8106ff05",
873 => x"09df0bf7",
874 => x"05068401",
875 => x"05050480",
876 => x"7834767e",
877 => x"ff125758",
878 => x"56758024",
879 => x"ff0509fe",
880 => x"8d0bf705",
881 => x"06840105",
882 => x"0504fcaa",
883 => x"398a7536",
884 => x"0b0b80fb",
885 => x"fc055473",
886 => x"76708105",
887 => x"583b8a75",
888 => x"35557409",
889 => x"70810509",
890 => x"060a8106",
891 => x"ff0509fe",
892 => x"f80bf705",
893 => x"06840105",
894 => x"05048a75",
895 => x"360b0b80",
896 => x"fbfc0554",
897 => x"73767081",
898 => x"05583b8a",
899 => x"75355574",
900 => x"09708105",
901 => x"09060a09",
902 => x"8106ff05",
903 => x"09ffae0b",
904 => x"f7050684",
905 => x"01050504",
906 => x"febf3974",
907 => x"527653b5",
908 => x"3dffb805",
909 => x"5195c73f",
910 => x"a43d0856",
911 => x"fdfe3970",
912 => x"80c10b81",
913 => x"e9983480",
914 => x"0b81eaf0",
915 => x"0c70800c",
916 => x"50047070",
917 => x"800b81e9",
918 => x"98335252",
919 => x"70098105",
920 => x"80c10509",
921 => x"70810509",
922 => x"060a8106",
923 => x"ff0509a0",
924 => x"0bf70506",
925 => x"84010505",
926 => x"047181ea",
927 => x"f0080781",
928 => x"eaf00c80",
929 => x"c20b81e9",
930 => x"9c347080",
931 => x"0c505004",
932 => x"810b81ea",
933 => x"f0080781",
934 => x"eaf00c80",
935 => x"c20b81e9",
936 => x"9c347080",
937 => x"0c505004",
938 => x"70707070",
939 => x"7570088a",
940 => x"05535381",
941 => x"e9983351",
942 => x"70098105",
943 => x"80c10509",
944 => x"70810509",
945 => x"060a8106",
946 => x"ff0509a9",
947 => x"0bf70506",
948 => x"84010505",
949 => x"04730970",
950 => x"81050906",
951 => x"0a098106",
952 => x"ff0509cf",
953 => x"0bf70506",
954 => x"84010505",
955 => x"0470800c",
956 => x"50505050",
957 => x"04ff1270",
958 => x"81e99408",
959 => x"31740c80",
960 => x"0c505050",
961 => x"5004fc3d",
962 => x"0d81e9a0",
963 => x"08557409",
964 => x"70810509",
965 => x"060a8106",
966 => x"ff050994",
967 => x"0bf70506",
968 => x"84010505",
969 => x"04767508",
970 => x"710c81e9",
971 => x"a0085654",
972 => x"8c155381",
973 => x"e9940852",
974 => x"8a5190ac",
975 => x"3f73800c",
976 => x"863d0d04",
977 => x"fb3d0d77",
978 => x"70085656",
979 => x"b05381e9",
980 => x"a0085274",
981 => x"51acb53f",
982 => x"850b8c17",
983 => x"0c850b8c",
984 => x"160c7508",
985 => x"750c81e9",
986 => x"a0085473",
987 => x"09708105",
988 => x"09060a81",
989 => x"06ff0509",
990 => x"920bf705",
991 => x"06840105",
992 => x"05047308",
993 => x"750c81e9",
994 => x"a008548c",
995 => x"145381e9",
996 => x"9408528a",
997 => x"518fd13f",
998 => x"84150809",
999 => x"70810509",
1000 => x"060a0981",
1001 => x"06ff0509",
1002 => x"b50bf705",
1003 => x"06840105",
1004 => x"0504860b",
1005 => x"8c160c88",
1006 => x"15528816",
1007 => x"08518dd3",
1008 => x"3f81e9a0",
1009 => x"08700876",
1010 => x"0c548c15",
1011 => x"7054548a",
1012 => x"52730851",
1013 => x"8f923f73",
1014 => x"800c873d",
1015 => x"0d047508",
1016 => x"54b05373",
1017 => x"527551ab",
1018 => x"a33f7380",
1019 => x"0c873d0d",
1020 => x"04e13d0d",
1021 => x"b05196c2",
1022 => x"3f800881",
1023 => x"e9900cb0",
1024 => x"5196b73f",
1025 => x"800881e9",
1026 => x"a00c81e9",
1027 => x"90088008",
1028 => x"0c800b80",
1029 => x"0884050c",
1030 => x"820b8008",
1031 => x"88050ca8",
1032 => x"0b80088c",
1033 => x"050c9f53",
1034 => x"0b0b80fc",
1035 => x"88528008",
1036 => x"900551aa",
1037 => x"d73f993d",
1038 => x"5c9f530b",
1039 => x"0b80fca8",
1040 => x"527b51aa",
1041 => x"c73f8a0b",
1042 => x"81a7d80c",
1043 => x"0b0b8186",
1044 => x"cc51f5e3",
1045 => x"3f0b0b80",
1046 => x"fcc851f5",
1047 => x"da3f0b0b",
1048 => x"8186cc51",
1049 => x"f5d13f81",
1050 => x"8aec0809",
1051 => x"70810509",
1052 => x"060a8106",
1053 => x"ff05098a",
1054 => x"ef0bf705",
1055 => x"06840105",
1056 => x"05040b0b",
1057 => x"80fcf851",
1058 => x"f5ad3f0b",
1059 => x"0b8186cc",
1060 => x"51f5a43f",
1061 => x"818ae808",
1062 => x"520b0b80",
1063 => x"fda451f5",
1064 => x"963f8051",
1065 => x"80c5a13f",
1066 => x"8008819a",
1067 => x"f80c810b",
1068 => x"923d5c58",
1069 => x"800b818a",
1070 => x"e80825ff",
1071 => x"05098492",
1072 => x"0bf70506",
1073 => x"84010505",
1074 => x"048e3d5d",
1075 => x"80c10b81",
1076 => x"e9983481",
1077 => x"0b81eaf0",
1078 => x"0c80c20b",
1079 => x"81e99c34",
1080 => x"825e835a",
1081 => x"9f530b0b",
1082 => x"80fdd452",
1083 => x"7a51a99c",
1084 => x"3f815f80",
1085 => x"7b537c52",
1086 => x"558eba3f",
1087 => x"80080981",
1088 => x"05750509",
1089 => x"70810509",
1090 => x"060a0981",
1091 => x"06ff0509",
1092 => x"8b0bf705",
1093 => x"06840105",
1094 => x"05048155",
1095 => x"7481eaf0",
1096 => x"0c7d7057",
1097 => x"55748325",
1098 => x"ff0509b4",
1099 => x"0bf70506",
1100 => x"84010505",
1101 => x"04741010",
1102 => x"15fd0540",
1103 => x"a13dffbc",
1104 => x"05538352",
1105 => x"75518ca0",
1106 => x"3f811e70",
1107 => x"5f705755",
1108 => x"837524ff",
1109 => x"0509de0b",
1110 => x"f7050684",
1111 => x"01050504",
1112 => x"7f547453",
1113 => x"819afc52",
1114 => x"81e9a851",
1115 => x"8c863f81",
1116 => x"e9a00870",
1117 => x"085757b0",
1118 => x"53765275",
1119 => x"51a88d3f",
1120 => x"850b8c18",
1121 => x"0c850b8c",
1122 => x"170c7608",
1123 => x"760c81e9",
1124 => x"a0085574",
1125 => x"09708105",
1126 => x"09060a81",
1127 => x"06ff0509",
1128 => x"920bf705",
1129 => x"06840105",
1130 => x"05047408",
1131 => x"760c81e9",
1132 => x"a008558c",
1133 => x"155381e9",
1134 => x"9408528a",
1135 => x"518ba93f",
1136 => x"84160809",
1137 => x"70810509",
1138 => x"060a0981",
1139 => x"06ff0509",
1140 => x"889f0bf7",
1141 => x"05068401",
1142 => x"05050486",
1143 => x"0b8c170c",
1144 => x"88165288",
1145 => x"17085189",
1146 => x"aa3f81e9",
1147 => x"a0087008",
1148 => x"770c578c",
1149 => x"16705455",
1150 => x"8a527408",
1151 => x"518ae93f",
1152 => x"80c10b81",
1153 => x"e99c3356",
1154 => x"56757526",
1155 => x"ff050980",
1156 => x"cc0bf705",
1157 => x"06840105",
1158 => x"050480c3",
1159 => x"5275518b",
1160 => x"d33f8008",
1161 => x"0981057f",
1162 => x"05097081",
1163 => x"0509060a",
1164 => x"8106ff05",
1165 => x"0987f50b",
1166 => x"f7050684",
1167 => x"01050504",
1168 => x"81167081",
1169 => x"ff0681e9",
1170 => x"9c335257",
1171 => x"55747627",
1172 => x"ff0509c6",
1173 => x"0bf70506",
1174 => x"84010505",
1175 => x"04797e29",
1176 => x"60707235",
1177 => x"70417272",
1178 => x"31707011",
1179 => x"11111111",
1180 => x"11517231",
1181 => x"5e538a05",
1182 => x"81e99833",
1183 => x"81e99408",
1184 => x"5a525258",
1185 => x"55760981",
1186 => x"0580c105",
1187 => x"09708105",
1188 => x"09060a81",
1189 => x"06ff0509",
1190 => x"87c10bf7",
1191 => x"05068401",
1192 => x"05050478",
1193 => x"09708105",
1194 => x"09060a09",
1195 => x"8106ff05",
1196 => x"09d30bf7",
1197 => x"05068401",
1198 => x"05050481",
1199 => x"1858818a",
1200 => x"e8087825",
1201 => x"ff0509fc",
1202 => x"830bf705",
1203 => x"06840105",
1204 => x"05048051",
1205 => x"80c0f13f",
1206 => x"800881e9",
1207 => x"8c0c0b0b",
1208 => x"80fdf451",
1209 => x"f0d13f0b",
1210 => x"0b8186cc",
1211 => x"51f0c83f",
1212 => x"0b0b80fe",
1213 => x"8451f0bf",
1214 => x"3f0b0b81",
1215 => x"86cc51f0",
1216 => x"b63f81e9",
1217 => x"9408520b",
1218 => x"0b80febc",
1219 => x"51f0a83f",
1220 => x"85520b0b",
1221 => x"80fed851",
1222 => x"f09d3f81",
1223 => x"eaf00852",
1224 => x"0b0b80fe",
1225 => x"f451f08f",
1226 => x"3f81520b",
1227 => x"0b80fed8",
1228 => x"51f0843f",
1229 => x"81e99833",
1230 => x"520b0b80",
1231 => x"ff9051ef",
1232 => x"f63f80c1",
1233 => x"520b0b80",
1234 => x"ffac51ef",
1235 => x"ea3f81e9",
1236 => x"9c33520b",
1237 => x"0b80ffc8",
1238 => x"51efdc3f",
1239 => x"80c2520b",
1240 => x"0b80ffac",
1241 => x"51efd03f",
1242 => x"81e9c808",
1243 => x"520b0b80",
1244 => x"ffe451ef",
1245 => x"c23f8752",
1246 => x"0b0b80fe",
1247 => x"d851efb7",
1248 => x"3f81a7d8",
1249 => x"08520b0b",
1250 => x"81808051",
1251 => x"efa93f0b",
1252 => x"0b81809c",
1253 => x"51efa03f",
1254 => x"0b0b8180",
1255 => x"c851ef97",
1256 => x"3f81e9a0",
1257 => x"08700853",
1258 => x"560b0b81",
1259 => x"80d451ef",
1260 => x"863f0b0b",
1261 => x"8180f051",
1262 => x"eefd3f81",
1263 => x"e9a00884",
1264 => x"1108535d",
1265 => x"0b0b8181",
1266 => x"a451eeeb",
1267 => x"3f80520b",
1268 => x"0b80fed8",
1269 => x"51eee03f",
1270 => x"81e9a008",
1271 => x"88110853",
1272 => x"580b0b81",
1273 => x"81c051ee",
1274 => x"ce3f8252",
1275 => x"0b0b80fe",
1276 => x"d851eec3",
1277 => x"3f81e9a0",
1278 => x"088c1108",
1279 => x"53590b0b",
1280 => x"8181dc51",
1281 => x"eeb13f91",
1282 => x"520b0b80",
1283 => x"fed851ee",
1284 => x"a63f81e9",
1285 => x"a0089005",
1286 => x"520b0b81",
1287 => x"81f851ee",
1288 => x"963f0b0b",
1289 => x"81829451",
1290 => x"ee8d3f0b",
1291 => x"0b8182cc",
1292 => x"51ee843f",
1293 => x"81e99008",
1294 => x"70085357",
1295 => x"0b0b8180",
1296 => x"d451edf3",
1297 => x"3f0b0b81",
1298 => x"82e051ed",
1299 => x"ea3f81e9",
1300 => x"90088411",
1301 => x"0853550b",
1302 => x"0b8181a4",
1303 => x"51edd83f",
1304 => x"80520b0b",
1305 => x"80fed851",
1306 => x"edcd3f81",
1307 => x"e9900888",
1308 => x"11085356",
1309 => x"0b0b8181",
1310 => x"c051edbb",
1311 => x"3f81520b",
1312 => x"0b80fed8",
1313 => x"51edb03f",
1314 => x"81e99008",
1315 => x"8c110853",
1316 => x"5d0b0b81",
1317 => x"81dc51ed",
1318 => x"9e3f9252",
1319 => x"0b0b80fe",
1320 => x"d851ed93",
1321 => x"3f81e990",
1322 => x"08900552",
1323 => x"0b0b8181",
1324 => x"f851ed83",
1325 => x"3f0b0b81",
1326 => x"829451ec",
1327 => x"fa3f7d52",
1328 => x"0b0b8183",
1329 => x"a051ecef",
1330 => x"3f85520b",
1331 => x"0b80fed8",
1332 => x"51ece43f",
1333 => x"79520b0b",
1334 => x"8183bc51",
1335 => x"ecd93f8d",
1336 => x"520b0b80",
1337 => x"fed851ec",
1338 => x"ce3f7f52",
1339 => x"0b0b8183",
1340 => x"d851ecc3",
1341 => x"3f87520b",
1342 => x"0b80fed8",
1343 => x"51ecb83f",
1344 => x"7e520b0b",
1345 => x"8183f451",
1346 => x"ecad3f81",
1347 => x"520b0b80",
1348 => x"fed851ec",
1349 => x"a23f7b52",
1350 => x"0b0b8184",
1351 => x"9051ec97",
1352 => x"3f0b0b81",
1353 => x"84ac51ec",
1354 => x"8e3f7a52",
1355 => x"0b0b8184",
1356 => x"e451ec83",
1357 => x"3f0b0b81",
1358 => x"858051eb",
1359 => x"fa3f0b0b",
1360 => x"8186cc51",
1361 => x"ebf13f81",
1362 => x"e98c0881",
1363 => x"9af80831",
1364 => x"70819af4",
1365 => x"0c520b0b",
1366 => x"8185b851",
1367 => x"ebd93f81",
1368 => x"9af40856",
1369 => x"817625ff",
1370 => x"0509819d",
1371 => x"0bf70506",
1372 => x"84010505",
1373 => x"04818ae8",
1374 => x"087077bd",
1375 => x"84c0290b",
1376 => x"35819aec",
1377 => x"0c767135",
1378 => x"819af00c",
1379 => x"768ddd29",
1380 => x"7187e829",
1381 => x"0b3581e9",
1382 => x"a40c5b0b",
1383 => x"0b8185c8",
1384 => x"51eb943f",
1385 => x"819aec08",
1386 => x"520b0b81",
1387 => x"85f851eb",
1388 => x"863f0b0b",
1389 => x"81868051",
1390 => x"eafd3f81",
1391 => x"9af00852",
1392 => x"0b0b8185",
1393 => x"f851eaef",
1394 => x"3f81e9a4",
1395 => x"08520b0b",
1396 => x"8186b051",
1397 => x"eae13f0b",
1398 => x"0b8186cc",
1399 => x"51ead83f",
1400 => x"800b800c",
1401 => x"a13d0d04",
1402 => x"0b0b8186",
1403 => x"d051f598",
1404 => x"39760856",
1405 => x"b0537552",
1406 => x"76519f90",
1407 => x"3f80c10b",
1408 => x"81e99c33",
1409 => x"5656f881",
1410 => x"390b0b81",
1411 => x"878051ea",
1412 => x"a63f0b0b",
1413 => x"8187b851",
1414 => x"ea9d3f0b",
1415 => x"0b8186cc",
1416 => x"51ea943f",
1417 => x"800b800c",
1418 => x"a13d0d04",
1419 => x"a13dffb8",
1420 => x"05528051",
1421 => x"80dd3f9f",
1422 => x"530b0b81",
1423 => x"87d8527a",
1424 => x"519ec93f",
1425 => x"777881e9",
1426 => x"940c8117",
1427 => x"7081ff06",
1428 => x"81e99c33",
1429 => x"5258565a",
1430 => x"f7f339ff",
1431 => x"15707731",
1432 => x"7e0c5980",
1433 => x"0b811959",
1434 => x"59818ae8",
1435 => x"087825ff",
1436 => x"0509f4d8",
1437 => x"0bf70506",
1438 => x"84010505",
1439 => x"04f8d339",
1440 => x"70707382",
1441 => x"32703070",
1442 => x"72078025",
1443 => x"800c5252",
1444 => x"50500470",
1445 => x"70707476",
1446 => x"71535452",
1447 => x"71098105",
1448 => x"82050970",
1449 => x"81050906",
1450 => x"0a8106ff",
1451 => x"05098b0b",
1452 => x"f7050684",
1453 => x"01050504",
1454 => x"83517109",
1455 => x"81058105",
1456 => x"09708105",
1457 => x"09060a81",
1458 => x"06ff0509",
1459 => x"80dd0bf7",
1460 => x"05068401",
1461 => x"05050481",
1462 => x"7226ff05",
1463 => x"0980e10b",
1464 => x"f7050684",
1465 => x"01050504",
1466 => x"71098105",
1467 => x"82050970",
1468 => x"81050906",
1469 => x"0a8106ff",
1470 => x"050980e2",
1471 => x"0bf70506",
1472 => x"84010505",
1473 => x"04710981",
1474 => x"05840509",
1475 => x"70810509",
1476 => x"060a8106",
1477 => x"ff0509bc",
1478 => x"0bf70506",
1479 => x"84010505",
1480 => x"0470730c",
1481 => x"70800c50",
1482 => x"50500480",
1483 => x"e40b81e9",
1484 => x"940825ff",
1485 => x"0509930b",
1486 => x"f7050684",
1487 => x"01050504",
1488 => x"80730c70",
1489 => x"800c5050",
1490 => x"50048373",
1491 => x"0c70800c",
1492 => x"50505004",
1493 => x"82730c70",
1494 => x"800c5050",
1495 => x"50048173",
1496 => x"0c70800c",
1497 => x"50505004",
1498 => x"70747414",
1499 => x"8205710c",
1500 => x"800c5004",
1501 => x"f73d0d7b",
1502 => x"7d7f6185",
1503 => x"1270822b",
1504 => x"75117074",
1505 => x"71708405",
1506 => x"530c5a5a",
1507 => x"5d5b760c",
1508 => x"7980f818",
1509 => x"0c798612",
1510 => x"5257585a",
1511 => x"5a767624",
1512 => x"ff0509ac",
1513 => x"0bf70506",
1514 => x"84010505",
1515 => x"0476b329",
1516 => x"822b7911",
1517 => x"51537673",
1518 => x"70840555",
1519 => x"0c811454",
1520 => x"757425ff",
1521 => x"0509ef0b",
1522 => x"f7050684",
1523 => x"01050504",
1524 => x"7681cc29",
1525 => x"19fc1108",
1526 => x"8105fc12",
1527 => x"0c7a1970",
1528 => x"089fa013",
1529 => x"0c585685",
1530 => x"0b81e994",
1531 => x"0c75800c",
1532 => x"8b3d0d04",
1533 => x"70707002",
1534 => x"93053351",
1535 => x"80028405",
1536 => x"97053354",
1537 => x"52700981",
1538 => x"05730509",
1539 => x"70810509",
1540 => x"060a8106",
1541 => x"ff050990",
1542 => x"0bf70506",
1543 => x"84010505",
1544 => x"0471800c",
1545 => x"50505004",
1546 => x"7081e998",
1547 => x"34810b80",
1548 => x"0c505050",
1549 => x"04f83d0d",
1550 => x"7a7c5956",
1551 => x"820b8319",
1552 => x"55557416",
1553 => x"70337533",
1554 => x"5b515372",
1555 => x"09810579",
1556 => x"05097081",
1557 => x"0509060a",
1558 => x"8106ff05",
1559 => x"0981860b",
1560 => x"f7050684",
1561 => x"01050504",
1562 => x"80c10b81",
1563 => x"16811656",
1564 => x"56578275",
1565 => x"25ff0509",
1566 => x"c90bf705",
1567 => x"06840105",
1568 => x"0504ffa9",
1569 => x"177081ff",
1570 => x"06555973",
1571 => x"8226ff05",
1572 => x"098b0bf7",
1573 => x"05068401",
1574 => x"05050487",
1575 => x"55815376",
1576 => x"09810580",
1577 => x"d2050970",
1578 => x"81050906",
1579 => x"0a8106ff",
1580 => x"0509ab0b",
1581 => x"f7050684",
1582 => x"01050504",
1583 => x"77527551",
1584 => x"9cb43f80",
1585 => x"53728008",
1586 => x"25ff0509",
1587 => x"910bf705",
1588 => x"06840105",
1589 => x"05048715",
1590 => x"81e9940c",
1591 => x"81537280",
1592 => x"0c8a3d0d",
1593 => x"047281e9",
1594 => x"98348275",
1595 => x"25ff0509",
1596 => x"fed00bf7",
1597 => x"05068401",
1598 => x"050504ff",
1599 => x"8539f93d",
1600 => x"0d797b7d",
1601 => x"54587259",
1602 => x"77307970",
1603 => x"30707207",
1604 => x"9f2a7371",
1605 => x"315a5259",
1606 => x"77795673",
1607 => x"0c537384",
1608 => x"130c5480",
1609 => x"0c893d0d",
1610 => x"04f93d0d",
1611 => x"797b7d7f",
1612 => x"56545254",
1613 => x"72097081",
1614 => x"0509060a",
1615 => x"8106ff05",
1616 => x"09b30bf7",
1617 => x"05068401",
1618 => x"05050470",
1619 => x"577158a0",
1620 => x"73315280",
1621 => x"7225ff05",
1622 => x"09a90bf7",
1623 => x"05068401",
1624 => x"05050477",
1625 => x"70742b57",
1626 => x"70732a78",
1627 => x"752b0756",
1628 => x"51747653",
1629 => x"5170740c",
1630 => x"7184150c",
1631 => x"73800c89",
1632 => x"3d0d0480",
1633 => x"56777230",
1634 => x"0b2b5574",
1635 => x"765351e5",
1636 => x"39fb3d0d",
1637 => x"77795555",
1638 => x"80567575",
1639 => x"24ff0509",
1640 => x"80d00bf7",
1641 => x"05068401",
1642 => x"05050480",
1643 => x"7424ff05",
1644 => x"09b70bf7",
1645 => x"05068401",
1646 => x"05050480",
1647 => x"53735274",
1648 => x"51819c3f",
1649 => x"80085475",
1650 => x"09708105",
1651 => x"09060a81",
1652 => x"06ff0509",
1653 => x"8d0bf705",
1654 => x"06840105",
1655 => x"05048008",
1656 => x"30547380",
1657 => x"0c873d0d",
1658 => x"04733076",
1659 => x"81325754",
1660 => x"ca397430",
1661 => x"55815673",
1662 => x"8025ff05",
1663 => x"09ffbc0b",
1664 => x"f7050684",
1665 => x"01050504",
1666 => x"e039fa3d",
1667 => x"0d787a57",
1668 => x"55805776",
1669 => x"7524ff05",
1670 => x"09be0bf7",
1671 => x"05068401",
1672 => x"05050475",
1673 => x"9f2c5481",
1674 => x"53757432",
1675 => x"74315274",
1676 => x"51ad3f80",
1677 => x"08547609",
1678 => x"70810509",
1679 => x"060a8106",
1680 => x"ff05098d",
1681 => x"0bf70506",
1682 => x"84010505",
1683 => x"04800830",
1684 => x"5473800c",
1685 => x"883d0d04",
1686 => x"74305581",
1687 => x"57c539fc",
1688 => x"3d0d7678",
1689 => x"53548153",
1690 => x"80747326",
1691 => x"52557209",
1692 => x"70810509",
1693 => x"060a8106",
1694 => x"ff050980",
1695 => x"d50bf705",
1696 => x"06840105",
1697 => x"05047009",
1698 => x"70810509",
1699 => x"060a8106",
1700 => x"ff050980",
1701 => x"ea0bf705",
1702 => x"06840105",
1703 => x"05048072",
1704 => x"24ff0509",
1705 => x"80d90bf7",
1706 => x"05068401",
1707 => x"05050471",
1708 => x"10731075",
1709 => x"72265354",
1710 => x"52720970",
1711 => x"81050906",
1712 => x"0a098106",
1713 => x"ff0509ff",
1714 => x"bd0bf705",
1715 => x"06840105",
1716 => x"05047351",
1717 => x"78097081",
1718 => x"0509060a",
1719 => x"098106ff",
1720 => x"05098b0b",
1721 => x"f7050684",
1722 => x"01050504",
1723 => x"74517080",
1724 => x"0c863d0d",
1725 => x"04720a10",
1726 => x"0a720a10",
1727 => x"0a535372",
1728 => x"09708105",
1729 => x"09060a81",
1730 => x"06ff0509",
1731 => x"c50bf705",
1732 => x"06840105",
1733 => x"05047174",
1734 => x"26ff0509",
1735 => x"d80bf705",
1736 => x"06840105",
1737 => x"05047372",
1738 => x"31757407",
1739 => x"740a100a",
1740 => x"740a100a",
1741 => x"55555654",
1742 => x"c6397070",
1743 => x"73528193",
1744 => x"b4085193",
1745 => x"3f505004",
1746 => x"70707352",
1747 => x"8193b408",
1748 => x"519bc43f",
1749 => x"505004f4",
1750 => x"3d0d7e60",
1751 => x"8b1170f8",
1752 => x"065b5555",
1753 => x"5d729626",
1754 => x"ff05098b",
1755 => x"0bf70506",
1756 => x"84010505",
1757 => x"04905880",
1758 => x"78247479",
1759 => x"26075580",
1760 => x"54740981",
1761 => x"05740509",
1762 => x"70810509",
1763 => x"060a0981",
1764 => x"06ff0509",
1765 => x"80f40bf7",
1766 => x"05068401",
1767 => x"0505047c",
1768 => x"5195f13f",
1769 => x"7783f726",
1770 => x"ff050980",
1771 => x"e40bf705",
1772 => x"06840105",
1773 => x"05047783",
1774 => x"2a701010",
1775 => x"10818bac",
1776 => x"058c1108",
1777 => x"58585475",
1778 => x"09810577",
1779 => x"05097081",
1780 => x"0509060a",
1781 => x"8106ff05",
1782 => x"0983b60b",
1783 => x"f7050684",
1784 => x"01050504",
1785 => x"841608fc",
1786 => x"068c1708",
1787 => x"88180871",
1788 => x"8c120c88",
1789 => x"120c5b76",
1790 => x"05841108",
1791 => x"81078412",
1792 => x"0c537c51",
1793 => x"958f3f88",
1794 => x"16547380",
1795 => x"0c8e3d0d",
1796 => x"0477892a",
1797 => x"78832a58",
1798 => x"54730970",
1799 => x"81050906",
1800 => x"0a8106ff",
1801 => x"05098180",
1802 => x"0bf70506",
1803 => x"84010505",
1804 => x"0477862a",
1805 => x"b8055784",
1806 => x"7427ff05",
1807 => x"0980e90b",
1808 => x"f7050684",
1809 => x"01050504",
1810 => x"80db1457",
1811 => x"947427ff",
1812 => x"050980d4",
1813 => x"0bf70506",
1814 => x"84010505",
1815 => x"04778c2a",
1816 => x"80ee0557",
1817 => x"80d47427",
1818 => x"ff0509bc",
1819 => x"0bf70506",
1820 => x"84010505",
1821 => x"04778f2a",
1822 => x"80f70557",
1823 => x"82d47427",
1824 => x"ff0509a4",
1825 => x"0bf70506",
1826 => x"84010505",
1827 => x"0477922a",
1828 => x"80fc0557",
1829 => x"8ad47427",
1830 => x"ff05098c",
1831 => x"0bf70506",
1832 => x"84010505",
1833 => x"0480fe57",
1834 => x"76101010",
1835 => x"818bac05",
1836 => x"8c110856",
1837 => x"53740981",
1838 => x"05730509",
1839 => x"70810509",
1840 => x"060a8106",
1841 => x"ff050980",
1842 => x"d70bf705",
1843 => x"06840105",
1844 => x"05048415",
1845 => x"08fc0670",
1846 => x"79315556",
1847 => x"738f24ff",
1848 => x"05098fb7",
1849 => x"0bf70506",
1850 => x"84010505",
1851 => x"04738025",
1852 => x"ff05098f",
1853 => x"ae0bf705",
1854 => x"06840105",
1855 => x"05048c15",
1856 => x"08557409",
1857 => x"81057305",
1858 => x"09708105",
1859 => x"09060a09",
1860 => x"8106ff05",
1861 => x"09ffbb0b",
1862 => x"f7050684",
1863 => x"01050504",
1864 => x"81175981",
1865 => x"8bbc0856",
1866 => x"75098105",
1867 => x"818bb405",
1868 => x"09708105",
1869 => x"09060a81",
1870 => x"06ff0509",
1871 => x"84ce0bf7",
1872 => x"05068401",
1873 => x"05050484",
1874 => x"1608fc06",
1875 => x"70793155",
1876 => x"55738f24",
1877 => x"ff050980",
1878 => x"e30bf705",
1879 => x"06840105",
1880 => x"0504818b",
1881 => x"b40b818b",
1882 => x"c00c818b",
1883 => x"b40b818b",
1884 => x"bc0c8074",
1885 => x"24ff0509",
1886 => x"80f80bf7",
1887 => x"05068401",
1888 => x"05050474",
1889 => x"16841108",
1890 => x"81078412",
1891 => x"0c53fcf2",
1892 => x"3988168c",
1893 => x"11085759",
1894 => x"75098105",
1895 => x"79050970",
1896 => x"81050906",
1897 => x"0a098106",
1898 => x"ff0509fc",
1899 => x"b70bf705",
1900 => x"06840105",
1901 => x"05048214",
1902 => x"59fee839",
1903 => x"77167881",
1904 => x"0784180c",
1905 => x"70818bc0",
1906 => x"0c70818b",
1907 => x"bc0c818b",
1908 => x"b40b8c12",
1909 => x"0c8c1108",
1910 => x"88120c74",
1911 => x"81078412",
1912 => x"0c740574",
1913 => x"710c5b7c",
1914 => x"5191aa3f",
1915 => x"881654fc",
1916 => x"993983ff",
1917 => x"7527ff05",
1918 => x"0985ff0b",
1919 => x"f7050684",
1920 => x"01050504",
1921 => x"74892a75",
1922 => x"832a5454",
1923 => x"73097081",
1924 => x"0509060a",
1925 => x"8106ff05",
1926 => x"0981800b",
1927 => x"f7050684",
1928 => x"01050504",
1929 => x"74862ab8",
1930 => x"05538474",
1931 => x"27ff0509",
1932 => x"80e90bf7",
1933 => x"05068401",
1934 => x"05050480",
1935 => x"db145394",
1936 => x"7427ff05",
1937 => x"0980d40b",
1938 => x"f7050684",
1939 => x"01050504",
1940 => x"748c2a80",
1941 => x"ee055380",
1942 => x"d47427ff",
1943 => x"0509bc0b",
1944 => x"f7050684",
1945 => x"01050504",
1946 => x"748f2a80",
1947 => x"f7055382",
1948 => x"d47427ff",
1949 => x"0509a40b",
1950 => x"f7050684",
1951 => x"01050504",
1952 => x"74922a80",
1953 => x"fc05538a",
1954 => x"d47427ff",
1955 => x"05098c0b",
1956 => x"f7050684",
1957 => x"01050504",
1958 => x"80fe5372",
1959 => x"10101081",
1960 => x"8bac0588",
1961 => x"11085557",
1962 => x"73098105",
1963 => x"77050970",
1964 => x"81050906",
1965 => x"0a8106ff",
1966 => x"05098aec",
1967 => x"0bf70506",
1968 => x"84010505",
1969 => x"04841408",
1970 => x"fc065b74",
1971 => x"7b27ff05",
1972 => x"09aa0bf7",
1973 => x"05068401",
1974 => x"05050488",
1975 => x"14085473",
1976 => x"09810577",
1977 => x"05097081",
1978 => x"0509060a",
1979 => x"098106ff",
1980 => x"0509d20b",
1981 => x"f7050684",
1982 => x"01050504",
1983 => x"8c140881",
1984 => x"8bac0b84",
1985 => x"0508718c",
1986 => x"190c7588",
1987 => x"190c7788",
1988 => x"130c5c57",
1989 => x"758c150c",
1990 => x"78538079",
1991 => x"24ff0509",
1992 => x"86860bf7",
1993 => x"05068401",
1994 => x"05050472",
1995 => x"822c8171",
1996 => x"2b565674",
1997 => x"7b26ff05",
1998 => x"0981a80b",
1999 => x"f7050684",
2000 => x"01050504",
2001 => x"7a750657",
2002 => x"76097081",
2003 => x"0509060a",
2004 => x"098106ff",
2005 => x"050983ee",
2006 => x"0bf70506",
2007 => x"84010505",
2008 => x"0478fc06",
2009 => x"84055974",
2010 => x"10707c06",
2011 => x"55557309",
2012 => x"70810509",
2013 => x"060a0981",
2014 => x"06ff0509",
2015 => x"83c80bf7",
2016 => x"05068401",
2017 => x"05050484",
2018 => x"1959dc39",
2019 => x"818bac0b",
2020 => x"84050879",
2021 => x"545b7880",
2022 => x"25ff0509",
2023 => x"ff8d0bf7",
2024 => x"05068401",
2025 => x"05050484",
2026 => x"ff397409",
2027 => x"7b067081",
2028 => x"8bac0b84",
2029 => x"050c5b74",
2030 => x"1055747b",
2031 => x"26ff0509",
2032 => x"a20bf705",
2033 => x"06840105",
2034 => x"05047409",
2035 => x"70810509",
2036 => x"060a0981",
2037 => x"06ff0509",
2038 => x"899c0bf7",
2039 => x"05068401",
2040 => x"05050481",
2041 => x"8bac0b88",
2042 => x"05087084",
2043 => x"1208fc06",
2044 => x"707b317b",
2045 => x"72268f72",
2046 => x"25075d57",
2047 => x"5c5c5578",
2048 => x"09708105",
2049 => x"09060a81",
2050 => x"06ff0509",
2051 => x"81c60bf7",
2052 => x"05068401",
2053 => x"05050479",
2054 => x"15818ba4",
2055 => x"08199011",
2056 => x"59545681",
2057 => x"8ba00809",
2058 => x"8105ff05",
2059 => x"09708105",
2060 => x"09060a81",
2061 => x"06ff0509",
2062 => x"900bf705",
2063 => x"06840105",
2064 => x"0504a08f",
2065 => x"13e08006",
2066 => x"5776527c",
2067 => x"518cc73f",
2068 => x"80085480",
2069 => x"08098105",
2070 => x"ff050970",
2071 => x"81050906",
2072 => x"0a8106ff",
2073 => x"0509ba0b",
2074 => x"f7050684",
2075 => x"01050504",
2076 => x"80087627",
2077 => x"ff050983",
2078 => x"e90bf705",
2079 => x"06840105",
2080 => x"05047409",
2081 => x"8105818b",
2082 => x"ac050970",
2083 => x"81050906",
2084 => x"0a8106ff",
2085 => x"050983ca",
2086 => x"0bf70506",
2087 => x"84010505",
2088 => x"04818bac",
2089 => x"0b880508",
2090 => x"55841508",
2091 => x"fc067079",
2092 => x"31797226",
2093 => x"8f722507",
2094 => x"5d555a7a",
2095 => x"09708105",
2096 => x"09060a09",
2097 => x"8106ff05",
2098 => x"0986d00b",
2099 => x"f7050684",
2100 => x"01050504",
2101 => x"77810784",
2102 => x"160c7715",
2103 => x"70818bac",
2104 => x"0b88050c",
2105 => x"74810784",
2106 => x"120c567c",
2107 => x"518ba63f",
2108 => x"88155473",
2109 => x"800c8e3d",
2110 => x"0d047483",
2111 => x"2a705454",
2112 => x"807424ff",
2113 => x"050982a6",
2114 => x"0bf70506",
2115 => x"84010505",
2116 => x"0472822c",
2117 => x"81712b81",
2118 => x"8bb00807",
2119 => x"70818bac",
2120 => x"0b84050c",
2121 => x"75101010",
2122 => x"818bac05",
2123 => x"88110871",
2124 => x"8c1b0c70",
2125 => x"881b0c79",
2126 => x"88130c57",
2127 => x"555c5575",
2128 => x"8c150cfb",
2129 => x"d3397879",
2130 => x"10101081",
2131 => x"8bac0570",
2132 => x"565b5c8c",
2133 => x"14085675",
2134 => x"09810574",
2135 => x"05097081",
2136 => x"0509060a",
2137 => x"8106ff05",
2138 => x"0980d70b",
2139 => x"f7050684",
2140 => x"01050504",
2141 => x"841608fc",
2142 => x"06707931",
2143 => x"5853768f",
2144 => x"24ff0509",
2145 => x"86c10bf7",
2146 => x"05068401",
2147 => x"05050476",
2148 => x"8025ff05",
2149 => x"0986f40b",
2150 => x"f7050684",
2151 => x"01050504",
2152 => x"8c160856",
2153 => x"75098105",
2154 => x"74050970",
2155 => x"81050906",
2156 => x"0a098106",
2157 => x"ff0509ff",
2158 => x"bb0bf705",
2159 => x"06840105",
2160 => x"05048814",
2161 => x"811a7083",
2162 => x"06555a54",
2163 => x"72097081",
2164 => x"0509060a",
2165 => x"098106ff",
2166 => x"0509fef7",
2167 => x"0bf70506",
2168 => x"84010505",
2169 => x"047b8306",
2170 => x"56750970",
2171 => x"81050906",
2172 => x"0a8106ff",
2173 => x"0509fbb2",
2174 => x"0bf70506",
2175 => x"84010505",
2176 => x"04ff1cf8",
2177 => x"1b5b5c88",
2178 => x"1a080981",
2179 => x"057a0509",
2180 => x"70810509",
2181 => x"060a8106",
2182 => x"ff0509c9",
2183 => x"0bf70506",
2184 => x"84010505",
2185 => x"04fb9039",
2186 => x"831953f9",
2187 => x"fe398314",
2188 => x"70822c81",
2189 => x"712b818b",
2190 => x"b0080770",
2191 => x"818bac0b",
2192 => x"84050c76",
2193 => x"10101081",
2194 => x"8bac0588",
2195 => x"1108718c",
2196 => x"1c0c7088",
2197 => x"1c0c7a88",
2198 => x"130c5853",
2199 => x"5d5653fd",
2200 => x"de39818a",
2201 => x"f0081759",
2202 => x"80080981",
2203 => x"05760509",
2204 => x"70810509",
2205 => x"060a8106",
2206 => x"ff050982",
2207 => x"870bf705",
2208 => x"06840105",
2209 => x"0504818b",
2210 => x"a0080981",
2211 => x"05ff0509",
2212 => x"70810509",
2213 => x"060a8106",
2214 => x"ff050985",
2215 => x"db0bf705",
2216 => x"06840105",
2217 => x"05047376",
2218 => x"3119818a",
2219 => x"f00c7387",
2220 => x"06705653",
2221 => x"72097081",
2222 => x"0509060a",
2223 => x"8106ff05",
2224 => x"09900bf7",
2225 => x"05068401",
2226 => x"05050488",
2227 => x"73317015",
2228 => x"55557614",
2229 => x"9fff06a0",
2230 => x"80713116",
2231 => x"70547e53",
2232 => x"515387b2",
2233 => x"3f800856",
2234 => x"80080981",
2235 => x"05ff0509",
2236 => x"70810509",
2237 => x"060a8106",
2238 => x"ff050982",
2239 => x"970bf705",
2240 => x"06840105",
2241 => x"0504818a",
2242 => x"f0081370",
2243 => x"818af00c",
2244 => x"7475818b",
2245 => x"ac0b8805",
2246 => x"0c777631",
2247 => x"15810755",
2248 => x"56597a09",
2249 => x"8105818b",
2250 => x"ac050970",
2251 => x"81050906",
2252 => x"0a8106ff",
2253 => x"050984cd",
2254 => x"0bf70506",
2255 => x"84010505",
2256 => x"04798f26",
2257 => x"ff050983",
2258 => x"e60bf705",
2259 => x"06840105",
2260 => x"0504810b",
2261 => x"84150c84",
2262 => x"1508fc06",
2263 => x"70793179",
2264 => x"72268f72",
2265 => x"25075d55",
2266 => x"5a7a0970",
2267 => x"81050906",
2268 => x"0a8106ff",
2269 => x"0509fadc",
2270 => x"0bf70506",
2271 => x"84010505",
2272 => x"04819839",
2273 => x"80089fff",
2274 => x"06557409",
2275 => x"70810509",
2276 => x"060a0981",
2277 => x"06ff0509",
2278 => x"fdec0bf7",
2279 => x"05068401",
2280 => x"05050478",
2281 => x"818af00c",
2282 => x"818bac0b",
2283 => x"8805087a",
2284 => x"18810784",
2285 => x"120c5581",
2286 => x"8b9c0879",
2287 => x"27ff0509",
2288 => x"8e0bf705",
2289 => x"06840105",
2290 => x"05047881",
2291 => x"8b9c0c81",
2292 => x"8b980879",
2293 => x"27ff0509",
2294 => x"f9cf0bf7",
2295 => x"05068401",
2296 => x"05050478",
2297 => x"818b980c",
2298 => x"841508fc",
2299 => x"06707931",
2300 => x"7972268f",
2301 => x"7225075d",
2302 => x"555a7a09",
2303 => x"70810509",
2304 => x"060a8106",
2305 => x"ff0509f9",
2306 => x"cb0bf705",
2307 => x"06840105",
2308 => x"05048839",
2309 => x"80745753",
2310 => x"fdec397c",
2311 => x"5184f63f",
2312 => x"800b800c",
2313 => x"8e3d0d04",
2314 => x"807324ff",
2315 => x"0509ad0b",
2316 => x"f7050684",
2317 => x"01050504",
2318 => x"72822c81",
2319 => x"712b818b",
2320 => x"b0080770",
2321 => x"818bac0b",
2322 => x"84050c5c",
2323 => x"5a768c17",
2324 => x"0c738817",
2325 => x"0c758818",
2326 => x"0cf5b939",
2327 => x"83137082",
2328 => x"2c81712b",
2329 => x"818bb008",
2330 => x"0770818b",
2331 => x"ac0b8405",
2332 => x"0c5d5b53",
2333 => x"d8397a75",
2334 => x"065c7b09",
2335 => x"70810509",
2336 => x"060a0981",
2337 => x"06ff0509",
2338 => x"f9bc0bf7",
2339 => x"05068401",
2340 => x"05050484",
2341 => x"19751056",
2342 => x"59dc39ff",
2343 => x"17810559",
2344 => x"f181398c",
2345 => x"15088816",
2346 => x"08718c12",
2347 => x"0c88120c",
2348 => x"59751584",
2349 => x"11088107",
2350 => x"84120c58",
2351 => x"7c5183d5",
2352 => x"3f881554",
2353 => x"f8ad3977",
2354 => x"16788107",
2355 => x"84180c8c",
2356 => x"17088818",
2357 => x"08718c12",
2358 => x"0c88120c",
2359 => x"5c70818b",
2360 => x"c00c7081",
2361 => x"8bbc0c81",
2362 => x"8bb40b8c",
2363 => x"120c8c11",
2364 => x"0888120c",
2365 => x"77810784",
2366 => x"120c7705",
2367 => x"77710c55",
2368 => x"7c518391",
2369 => x"3f881654",
2370 => x"ee803972",
2371 => x"16841108",
2372 => x"81078412",
2373 => x"0c588c16",
2374 => x"08881708",
2375 => x"718c120c",
2376 => x"88120c57",
2377 => x"7c5182ed",
2378 => x"3f881654",
2379 => x"eddc3972",
2380 => x"84150cf4",
2381 => x"1af80670",
2382 => x"841d0881",
2383 => x"0607841d",
2384 => x"0c701c55",
2385 => x"56850b84",
2386 => x"150c850b",
2387 => x"88150c8f",
2388 => x"7627ff05",
2389 => x"09fce00b",
2390 => x"f7050684",
2391 => x"01050504",
2392 => x"881b527c",
2393 => x"5187b03f",
2394 => x"818bac0b",
2395 => x"88050881",
2396 => x"8af0085a",
2397 => x"55fcc039",
2398 => x"78818af0",
2399 => x"0c73818b",
2400 => x"a00cfaaa",
2401 => x"39728415",
2402 => x"0cfcac39",
2403 => x"fb3d0d77",
2404 => x"707a7c58",
2405 => x"5553568f",
2406 => x"7527ff05",
2407 => x"0981a40b",
2408 => x"f7050684",
2409 => x"01050504",
2410 => x"72760783",
2411 => x"06517009",
2412 => x"70810509",
2413 => x"060a0981",
2414 => x"06ff0509",
2415 => x"81850bf7",
2416 => x"05068401",
2417 => x"05050475",
2418 => x"73525470",
2419 => x"70840552",
2420 => x"08747084",
2421 => x"05560c73",
2422 => x"71708405",
2423 => x"53087170",
2424 => x"8405530c",
2425 => x"71708405",
2426 => x"53087170",
2427 => x"8405530c",
2428 => x"71708405",
2429 => x"53087170",
2430 => x"8405530c",
2431 => x"f0165654",
2432 => x"748f26ff",
2433 => x"0509c40b",
2434 => x"f7050684",
2435 => x"01050504",
2436 => x"837527ff",
2437 => x"0509a80b",
2438 => x"f7050684",
2439 => x"01050504",
2440 => x"70708405",
2441 => x"52087470",
2442 => x"8405560c",
2443 => x"fc155574",
2444 => x"8326ff05",
2445 => x"09ea0bf7",
2446 => x"05068401",
2447 => x"05050473",
2448 => x"715452ff",
2449 => x"15517009",
2450 => x"8105ff05",
2451 => x"09708105",
2452 => x"09060a81",
2453 => x"06ff0509",
2454 => x"b40bf705",
2455 => x"06840105",
2456 => x"05047270",
2457 => x"81055472",
2458 => x"70810554",
2459 => x"3bff1151",
2460 => x"70098105",
2461 => x"ff050970",
2462 => x"81050906",
2463 => x"0a098106",
2464 => x"ff0509de",
2465 => x"0bf70506",
2466 => x"84010505",
2467 => x"0475800c",
2468 => x"873d0d04",
2469 => x"04047070",
2470 => x"7070800b",
2471 => x"81eaf40c",
2472 => x"76518cc1",
2473 => x"3f800853",
2474 => x"80080981",
2475 => x"05ff0509",
2476 => x"70810509",
2477 => x"060a8106",
2478 => x"ff050991",
2479 => x"0bf70506",
2480 => x"84010505",
2481 => x"0472800c",
2482 => x"50505050",
2483 => x"0481eaf4",
2484 => x"08547309",
2485 => x"70810509",
2486 => x"060a8106",
2487 => x"ff0509e5",
2488 => x"0bf70506",
2489 => x"84010505",
2490 => x"04757471",
2491 => x"0c527280",
2492 => x"0c505050",
2493 => x"5004fb3d",
2494 => x"0d777970",
2495 => x"72078306",
2496 => x"53545270",
2497 => x"09708105",
2498 => x"09060a09",
2499 => x"8106ff05",
2500 => x"09b20bf7",
2501 => x"05068401",
2502 => x"05050471",
2503 => x"73730854",
2504 => x"56547109",
2505 => x"81057308",
2506 => x"05097081",
2507 => x"0509060a",
2508 => x"8106ff05",
2509 => x"0981890b",
2510 => x"f7050684",
2511 => x"01050504",
2512 => x"73755452",
2513 => x"71337081",
2514 => x"ff065254",
2515 => x"70097081",
2516 => x"0509060a",
2517 => x"8106ff05",
2518 => x"0980cf0b",
2519 => x"f7050684",
2520 => x"01050504",
2521 => x"72335570",
2522 => x"09810575",
2523 => x"05097081",
2524 => x"0509060a",
2525 => x"098106ff",
2526 => x"0509b20b",
2527 => x"f7050684",
2528 => x"01050504",
2529 => x"81128114",
2530 => x"71337081",
2531 => x"ff065456",
2532 => x"54527009",
2533 => x"70810509",
2534 => x"060a0981",
2535 => x"06ff0509",
2536 => x"c30bf705",
2537 => x"06840105",
2538 => x"05047233",
2539 => x"557381ff",
2540 => x"067581ff",
2541 => x"06717131",
2542 => x"800c5552",
2543 => x"873d0d04",
2544 => x"7109f7fb",
2545 => x"fdff1306",
2546 => x"f8848281",
2547 => x"80065271",
2548 => x"09708105",
2549 => x"09060a09",
2550 => x"8106ff05",
2551 => x"09b70bf7",
2552 => x"05068401",
2553 => x"05050484",
2554 => x"14841671",
2555 => x"08545654",
2556 => x"71098105",
2557 => x"75080509",
2558 => x"70810509",
2559 => x"060a8106",
2560 => x"ff0509ff",
2561 => x"bb0bf705",
2562 => x"06840105",
2563 => x"05047375",
2564 => x"5452feb0",
2565 => x"39800b80",
2566 => x"0c873d0d",
2567 => x"04fb3d0d",
2568 => x"77705256",
2569 => x"fcee3f81",
2570 => x"8bac0b88",
2571 => x"05088411",
2572 => x"08fc0670",
2573 => x"7b319fef",
2574 => x"05e08006",
2575 => x"e0800552",
2576 => x"5555a080",
2577 => x"7524ff05",
2578 => x"09b30bf7",
2579 => x"05068401",
2580 => x"05050480",
2581 => x"527551fc",
2582 => x"bd3f818b",
2583 => x"b4081453",
2584 => x"72098105",
2585 => x"80080509",
2586 => x"70810509",
2587 => x"060a8106",
2588 => x"ff050997",
2589 => x"0bf70506",
2590 => x"84010505",
2591 => x"047551fc",
2592 => x"943f8053",
2593 => x"72800c87",
2594 => x"3d0d0474",
2595 => x"30527551",
2596 => x"fc843f80",
2597 => x"08098105",
2598 => x"ff050970",
2599 => x"81050906",
2600 => x"0a8106ff",
2601 => x"0509b00b",
2602 => x"f7050684",
2603 => x"01050504",
2604 => x"818bac0b",
2605 => x"88050874",
2606 => x"76318107",
2607 => x"84120c53",
2608 => x"818af008",
2609 => x"7531818a",
2610 => x"f00c7551",
2611 => x"fbc73f81",
2612 => x"0b800c87",
2613 => x"3d0d0480",
2614 => x"527551fb",
2615 => x"b93f818b",
2616 => x"ac0b8805",
2617 => x"08800871",
2618 => x"3154548f",
2619 => x"7325ff05",
2620 => x"09ff8a0b",
2621 => x"f7050684",
2622 => x"01050504",
2623 => x"8008818b",
2624 => x"a0083181",
2625 => x"8af00c72",
2626 => x"81078415",
2627 => x"0c7551fb",
2628 => x"843f8053",
2629 => x"feee39f7",
2630 => x"3d0d7b7d",
2631 => x"545a7209",
2632 => x"70810509",
2633 => x"060a8106",
2634 => x"ff050984",
2635 => x"9e0bf705",
2636 => x"06840105",
2637 => x"05047951",
2638 => x"fada3ff8",
2639 => x"13841108",
2640 => x"70fe0670",
2641 => x"13841108",
2642 => x"fc065c57",
2643 => x"58545781",
2644 => x"8bb40809",
2645 => x"81057405",
2646 => x"09708105",
2647 => x"09060a81",
2648 => x"06ff0509",
2649 => x"85840bf7",
2650 => x"05068401",
2651 => x"05050477",
2652 => x"84150c80",
2653 => x"73810656",
2654 => x"59740981",
2655 => x"05790509",
2656 => x"70810509",
2657 => x"060a8106",
2658 => x"ff050983",
2659 => x"c20bf705",
2660 => x"06840105",
2661 => x"05047714",
2662 => x"84110881",
2663 => x"06565374",
2664 => x"09708105",
2665 => x"09060a09",
2666 => x"8106ff05",
2667 => x"0980d40b",
2668 => x"f7050684",
2669 => x"01050504",
2670 => x"77165678",
2671 => x"09708105",
2672 => x"09060a09",
2673 => x"8106ff05",
2674 => x"0983bf0b",
2675 => x"f7050684",
2676 => x"01050504",
2677 => x"88140855",
2678 => x"74098105",
2679 => x"818bb405",
2680 => x"09708105",
2681 => x"09060a81",
2682 => x"06ff0509",
2683 => x"84e60bf7",
2684 => x"05068401",
2685 => x"0505048c",
2686 => x"1408708c",
2687 => x"170c7588",
2688 => x"120c5875",
2689 => x"81078418",
2690 => x"0c751776",
2691 => x"710c5478",
2692 => x"09708105",
2693 => x"09060a09",
2694 => x"8106ff05",
2695 => x"0982a70b",
2696 => x"f7050684",
2697 => x"01050504",
2698 => x"83ff7627",
2699 => x"ff050982",
2700 => x"ea0bf705",
2701 => x"06840105",
2702 => x"05047589",
2703 => x"2a76832a",
2704 => x"54547309",
2705 => x"70810509",
2706 => x"060a8106",
2707 => x"ff050981",
2708 => x"800bf705",
2709 => x"06840105",
2710 => x"05047586",
2711 => x"2ab80553",
2712 => x"847427ff",
2713 => x"050980e9",
2714 => x"0bf70506",
2715 => x"84010505",
2716 => x"0480db14",
2717 => x"53947427",
2718 => x"ff050980",
2719 => x"d40bf705",
2720 => x"06840105",
2721 => x"0504758c",
2722 => x"2a80ee05",
2723 => x"5380d474",
2724 => x"27ff0509",
2725 => x"bc0bf705",
2726 => x"06840105",
2727 => x"0504758f",
2728 => x"2a80f705",
2729 => x"5382d474",
2730 => x"27ff0509",
2731 => x"a40bf705",
2732 => x"06840105",
2733 => x"05047592",
2734 => x"2a80fc05",
2735 => x"538ad474",
2736 => x"27ff0509",
2737 => x"8c0bf705",
2738 => x"06840105",
2739 => x"050480fe",
2740 => x"53721010",
2741 => x"10818bac",
2742 => x"05881108",
2743 => x"55557309",
2744 => x"81057505",
2745 => x"09708105",
2746 => x"09060a81",
2747 => x"06ff0509",
2748 => x"83a90bf7",
2749 => x"05068401",
2750 => x"05050484",
2751 => x"1408fc06",
2752 => x"59757927",
2753 => x"ff0509aa",
2754 => x"0bf70506",
2755 => x"84010505",
2756 => x"04881408",
2757 => x"54730981",
2758 => x"05750509",
2759 => x"70810509",
2760 => x"060a0981",
2761 => x"06ff0509",
2762 => x"d20bf705",
2763 => x"06840105",
2764 => x"05048c14",
2765 => x"08708c19",
2766 => x"0c748819",
2767 => x"0c778812",
2768 => x"0c55768c",
2769 => x"150c7951",
2770 => x"f6cb3f8b",
2771 => x"3d0d0476",
2772 => x"08777131",
2773 => x"58760588",
2774 => x"18085656",
2775 => x"74098105",
2776 => x"818bb405",
2777 => x"09708105",
2778 => x"09060a81",
2779 => x"06ff0509",
2780 => x"80f30bf7",
2781 => x"05068401",
2782 => x"0505048c",
2783 => x"1708708c",
2784 => x"170c7588",
2785 => x"120c53fc",
2786 => x"8d398814",
2787 => x"088c1508",
2788 => x"708c130c",
2789 => x"5988190c",
2790 => x"fce93975",
2791 => x"832a7054",
2792 => x"54807424",
2793 => x"ff050981",
2794 => x"c00bf705",
2795 => x"06840105",
2796 => x"05047282",
2797 => x"2c81712b",
2798 => x"818bb008",
2799 => x"07818bac",
2800 => x"0b84050c",
2801 => x"74101010",
2802 => x"818bac05",
2803 => x"88110871",
2804 => x"8c1b0c70",
2805 => x"881b0c79",
2806 => x"88130c56",
2807 => x"5a55768c",
2808 => x"150cfee2",
2809 => x"398159fb",
2810 => x"ad397716",
2811 => x"73810654",
2812 => x"55720970",
2813 => x"81050906",
2814 => x"0a098106",
2815 => x"ff0509a0",
2816 => x"0bf70506",
2817 => x"84010505",
2818 => x"04760877",
2819 => x"71315875",
2820 => x"058c1808",
2821 => x"88190871",
2822 => x"8c120c88",
2823 => x"120c5555",
2824 => x"74810784",
2825 => x"180c7681",
2826 => x"8bac0b88",
2827 => x"050c818b",
2828 => x"a8087526",
2829 => x"ff0509fe",
2830 => x"8d0bf705",
2831 => x"06840105",
2832 => x"0504818b",
2833 => x"a4085279",
2834 => x"51f7d23f",
2835 => x"7951f4c5",
2836 => x"3ffdf839",
2837 => x"81778c17",
2838 => x"0c778817",
2839 => x"0c758c19",
2840 => x"0c758819",
2841 => x"0c59fb9b",
2842 => x"39831470",
2843 => x"822c8171",
2844 => x"2b818bb0",
2845 => x"0807818b",
2846 => x"ac0b8405",
2847 => x"0c751010",
2848 => x"10818bac",
2849 => x"05881108",
2850 => x"718c1c0c",
2851 => x"70881c0c",
2852 => x"7a88130c",
2853 => x"575b5653",
2854 => x"fec43980",
2855 => x"7324ff05",
2856 => x"09ab0bf7",
2857 => x"05068401",
2858 => x"05050472",
2859 => x"822c8171",
2860 => x"2b818bb0",
2861 => x"0807818b",
2862 => x"ac0b8405",
2863 => x"0c58748c",
2864 => x"180c7388",
2865 => x"180c7688",
2866 => x"160cfcf6",
2867 => x"39831370",
2868 => x"822c8171",
2869 => x"2b818bb0",
2870 => x"0807818b",
2871 => x"ac0b8405",
2872 => x"0c5953da",
2873 => x"39707070",
2874 => x"81eaf808",
2875 => x"51700970",
2876 => x"81050906",
2877 => x"0a098106",
2878 => x"ff050992",
2879 => x"0bf70506",
2880 => x"84010505",
2881 => x"0481eb80",
2882 => x"7081eaf8",
2883 => x"0c517411",
2884 => x"52ff5371",
2885 => x"87fb8080",
2886 => x"26ff0509",
2887 => x"900bf705",
2888 => x"06840105",
2889 => x"05047181",
2890 => x"eaf80c70",
2891 => x"5372800c",
2892 => x"50505004",
2893 => x"70707070",
2894 => x"800b818a",
2895 => x"dc085454",
2896 => x"72098105",
2897 => x"81050970",
2898 => x"81050906",
2899 => x"0a8106ff",
2900 => x"0509a50b",
2901 => x"f7050684",
2902 => x"01050504",
2903 => x"7381eafc",
2904 => x"0cffb7b3",
2905 => x"3fffad98",
2906 => x"3f819ab4",
2907 => x"528151c5",
2908 => x"803f8008",
2909 => x"518cbe3f",
2910 => x"7281eafc",
2911 => x"0cffb797",
2912 => x"3fffacfc",
2913 => x"3f819ab4",
2914 => x"528151c4",
2915 => x"e43f8008",
2916 => x"518ca23f",
2917 => x"00ff3900",
2918 => x"ff39f53d",
2919 => x"0d7e6081",
2920 => x"eafc0870",
2921 => x"5b585b5b",
2922 => x"75097081",
2923 => x"0509060a",
2924 => x"098106ff",
2925 => x"050980fb",
2926 => x"0bf70506",
2927 => x"84010505",
2928 => x"04777a25",
2929 => x"ff050980",
2930 => x"cc0bf705",
2931 => x"06840105",
2932 => x"0504771b",
2933 => x"70337081",
2934 => x"ff065858",
2935 => x"59750981",
2936 => x"058a0509",
2937 => x"70810509",
2938 => x"060a8106",
2939 => x"ff0509ac",
2940 => x"0bf70506",
2941 => x"84010505",
2942 => x"047681ff",
2943 => x"0651ffb5",
2944 => x"e23f8118",
2945 => x"58797824",
2946 => x"ff0509c6",
2947 => x"0bf70506",
2948 => x"84010505",
2949 => x"0479800c",
2950 => x"8d3d0d04",
2951 => x"8d51ffb5",
2952 => x"c23f7833",
2953 => x"7081ff06",
2954 => x"5257ffb5",
2955 => x"b63f8118",
2956 => x"58d33979",
2957 => x"557a547d",
2958 => x"5385528d",
2959 => x"3dfc0551",
2960 => x"ffb4eb3f",
2961 => x"8008568a",
2962 => x"e53f7b80",
2963 => x"080c7580",
2964 => x"0c8d3d0d",
2965 => x"04f63d0d",
2966 => x"7d7f81ea",
2967 => x"fc08705a",
2968 => x"585a5a75",
2969 => x"09708105",
2970 => x"09060a09",
2971 => x"8106ff05",
2972 => x"0981930b",
2973 => x"f7050684",
2974 => x"01050504",
2975 => x"767925ff",
2976 => x"050980f4",
2977 => x"0bf70506",
2978 => x"84010505",
2979 => x"04761a58",
2980 => x"ffb49d3f",
2981 => x"80087834",
2982 => x"800b8008",
2983 => x"81ff0657",
2984 => x"58750981",
2985 => x"058a0509",
2986 => x"70810509",
2987 => x"060a8106",
2988 => x"ff050980",
2989 => x"cc0bf705",
2990 => x"06840105",
2991 => x"0504758d",
2992 => x"32703070",
2993 => x"80257a07",
2994 => x"51515675",
2995 => x"09708105",
2996 => x"09060a09",
2997 => x"8106ff05",
2998 => x"0980cd0b",
2999 => x"f7050684",
3000 => x"01050504",
3001 => x"81175778",
3002 => x"7724ff05",
3003 => x"09ff9e0b",
3004 => x"f7050684",
3005 => x"01050504",
3006 => x"76567580",
3007 => x"0c8c3d0d",
3008 => x"048158ff",
3009 => x"b9397855",
3010 => x"79547c53",
3011 => x"84528c3d",
3012 => x"fc0551ff",
3013 => x"b3983f80",
3014 => x"08568992",
3015 => x"3f7a8008",
3016 => x"0c75800c",
3017 => x"8c3d0d04",
3018 => x"811756ce",
3019 => x"39f93d0d",
3020 => x"795781ea",
3021 => x"fc080970",
3022 => x"81050906",
3023 => x"0a8106ff",
3024 => x"0509b50b",
3025 => x"f7050684",
3026 => x"01050504",
3027 => x"76518d88",
3028 => x"3f7b567a",
3029 => x"55800881",
3030 => x"05547653",
3031 => x"8252893d",
3032 => x"fc0551ff",
3033 => x"b2c83f80",
3034 => x"085788c2",
3035 => x"3f778008",
3036 => x"0c76800c",
3037 => x"893d0d04",
3038 => x"88b43f85",
3039 => x"0b80080c",
3040 => x"ff0b800c",
3041 => x"893d0d04",
3042 => x"fb3d0d81",
3043 => x"eafc0870",
3044 => x"56547309",
3045 => x"70810509",
3046 => x"060a0981",
3047 => x"06ff0509",
3048 => x"900bf705",
3049 => x"06840105",
3050 => x"05047480",
3051 => x"0c873d0d",
3052 => x"04775383",
3053 => x"52873dfc",
3054 => x"0551ffb1",
3055 => x"f13f8008",
3056 => x"5487eb3f",
3057 => x"7580080c",
3058 => x"73800c87",
3059 => x"3d0d04ff",
3060 => x"0b800c04",
3061 => x"fb3d0d77",
3062 => x"5581eafc",
3063 => x"08097081",
3064 => x"0509060a",
3065 => x"8106ff05",
3066 => x"09b10bf7",
3067 => x"05068401",
3068 => x"05050474",
3069 => x"518be13f",
3070 => x"80088105",
3071 => x"54745387",
3072 => x"52873dfc",
3073 => x"0551ffb1",
3074 => x"a53f8008",
3075 => x"55879f3f",
3076 => x"7580080c",
3077 => x"74800c87",
3078 => x"3d0d0487",
3079 => x"913f850b",
3080 => x"80080cff",
3081 => x"0b800c87",
3082 => x"3d0d04fa",
3083 => x"3d0d81ea",
3084 => x"fc080970",
3085 => x"81050906",
3086 => x"0a8106ff",
3087 => x"0509ab0b",
3088 => x"f7050684",
3089 => x"01050504",
3090 => x"7a557954",
3091 => x"78538652",
3092 => x"883dfc05",
3093 => x"51ffb0d6",
3094 => x"3f800856",
3095 => x"86d03f76",
3096 => x"80080c75",
3097 => x"800c883d",
3098 => x"0d0486c2",
3099 => x"3f9d0b80",
3100 => x"080cff0b",
3101 => x"800c883d",
3102 => x"0d04f73d",
3103 => x"0d7b7d5b",
3104 => x"59bc5380",
3105 => x"52795188",
3106 => x"cd3f8070",
3107 => x"56579856",
3108 => x"74197033",
3109 => x"70782b79",
3110 => x"078118f8",
3111 => x"1a5a5859",
3112 => x"55588475",
3113 => x"24ff0509",
3114 => x"e70bf705",
3115 => x"06840105",
3116 => x"0504767a",
3117 => x"23841958",
3118 => x"80705657",
3119 => x"98567418",
3120 => x"70337078",
3121 => x"2b790781",
3122 => x"18f81a5a",
3123 => x"58595154",
3124 => x"847524ff",
3125 => x"0509e70b",
3126 => x"f7050684",
3127 => x"01050504",
3128 => x"76821b23",
3129 => x"88195880",
3130 => x"70565798",
3131 => x"56741870",
3132 => x"3370782b",
3133 => x"79078118",
3134 => x"f81a5a58",
3135 => x"59515484",
3136 => x"7524ff05",
3137 => x"09e70bf7",
3138 => x"05068401",
3139 => x"05050476",
3140 => x"841b0c8c",
3141 => x"19588070",
3142 => x"56579856",
3143 => x"74187033",
3144 => x"70782b79",
3145 => x"078118f8",
3146 => x"1a5a5859",
3147 => x"51548475",
3148 => x"24ff0509",
3149 => x"e70bf705",
3150 => x"06840105",
3151 => x"05047688",
3152 => x"1b239019",
3153 => x"58807056",
3154 => x"57985674",
3155 => x"18703370",
3156 => x"782b7907",
3157 => x"8118f81a",
3158 => x"5a585951",
3159 => x"54847524",
3160 => x"ff0509e7",
3161 => x"0bf70506",
3162 => x"84010505",
3163 => x"04768a1b",
3164 => x"23941958",
3165 => x"80705657",
3166 => x"98567418",
3167 => x"70337078",
3168 => x"2b790781",
3169 => x"18f81a5a",
3170 => x"58595154",
3171 => x"847524ff",
3172 => x"0509e70b",
3173 => x"f7050684",
3174 => x"01050504",
3175 => x"768c1b23",
3176 => x"98195880",
3177 => x"70565798",
3178 => x"56741870",
3179 => x"3370782b",
3180 => x"79078118",
3181 => x"f81a5a58",
3182 => x"59515484",
3183 => x"7524ff05",
3184 => x"09e70bf7",
3185 => x"05068401",
3186 => x"05050476",
3187 => x"8e1b239c",
3188 => x"19588070",
3189 => x"5657b856",
3190 => x"74187033",
3191 => x"70782b79",
3192 => x"078118f8",
3193 => x"1a5a5859",
3194 => x"5a548875",
3195 => x"24ff0509",
3196 => x"e70bf705",
3197 => x"06840105",
3198 => x"05047690",
3199 => x"1b0c8b3d",
3200 => x"0d04e93d",
3201 => x"0d6a81ea",
3202 => x"fc085757",
3203 => x"75097081",
3204 => x"0509060a",
3205 => x"098106ff",
3206 => x"05099b0b",
3207 => x"f7050684",
3208 => x"01050504",
3209 => x"80c0800b",
3210 => x"84180c75",
3211 => x"ac180c75",
3212 => x"800c993d",
3213 => x"0d04893d",
3214 => x"70556a54",
3215 => x"558a5299",
3216 => x"3dffbc05",
3217 => x"51fface6",
3218 => x"3f800877",
3219 => x"53755256",
3220 => x"fca83f82",
3221 => x"d93f7780",
3222 => x"080c7580",
3223 => x"0c993d0d",
3224 => x"04e93d0d",
3225 => x"695781ea",
3226 => x"fc080970",
3227 => x"81050906",
3228 => x"0a8106ff",
3229 => x"0509be0b",
3230 => x"f7050684",
3231 => x"01050504",
3232 => x"765186d4",
3233 => x"3f893d70",
3234 => x"56800881",
3235 => x"05557754",
3236 => x"568f5299",
3237 => x"3dffbc05",
3238 => x"51ffac92",
3239 => x"3f80086b",
3240 => x"53765257",
3241 => x"fbd43f82",
3242 => x"853f7780",
3243 => x"080c7680",
3244 => x"0c993d0d",
3245 => x"0481f73f",
3246 => x"850b8008",
3247 => x"0cff0b80",
3248 => x"0c993d0d",
3249 => x"04fc3d0d",
3250 => x"815481ea",
3251 => x"fc080970",
3252 => x"81050906",
3253 => x"0a098106",
3254 => x"ff050990",
3255 => x"0bf70506",
3256 => x"84010505",
3257 => x"0473800c",
3258 => x"863d0d04",
3259 => x"765397b9",
3260 => x"52863dfc",
3261 => x"0551ffab",
3262 => x"b53f8008",
3263 => x"5481af3f",
3264 => x"7480080c",
3265 => x"73800c86",
3266 => x"3d0d04f4",
3267 => x"3d0d7e81",
3268 => x"9ae00870",
3269 => x"0881ff06",
3270 => x"913df805",
3271 => x"54515959",
3272 => x"ffacf63f",
3273 => x"77578054",
3274 => x"76557b7d",
3275 => x"58527653",
3276 => x"8e3df005",
3277 => x"5186e23f",
3278 => x"797b5879",
3279 => x"0c76841a",
3280 => x"0c78800c",
3281 => x"8e3d0d04",
3282 => x"f43d0d7e",
3283 => x"819ae008",
3284 => x"70087081",
3285 => x"ff06923d",
3286 => x"f8055551",
3287 => x"5a5759ff",
3288 => x"acb73f77",
3289 => x"57800b8b",
3290 => x"3d595476",
3291 => x"557b7d58",
3292 => x"52765377",
3293 => x"5186a23f",
3294 => x"8056bd84",
3295 => x"c0765555",
3296 => x"797b5852",
3297 => x"76537751",
3298 => x"868f3f7a",
3299 => x"57780970",
3300 => x"81050906",
3301 => x"0a8106ff",
3302 => x"05098c0b",
3303 => x"f7050684",
3304 => x"01050504",
3305 => x"76790c76",
3306 => x"800c8e3d",
3307 => x"0d048193",
3308 => x"b408800c",
3309 => x"04f73d0d",
3310 => x"7b8193b4",
3311 => x"0882c811",
3312 => x"085a545a",
3313 => x"77097081",
3314 => x"0509060a",
3315 => x"8106ff05",
3316 => x"0981ac0b",
3317 => x"f7050684",
3318 => x"01050504",
3319 => x"81881884",
3320 => x"1908ff05",
3321 => x"81712b59",
3322 => x"55598074",
3323 => x"24ff0509",
3324 => x"81d20bf7",
3325 => x"05068401",
3326 => x"05050480",
3327 => x"7424ff05",
3328 => x"0980db0b",
3329 => x"f7050684",
3330 => x"01050504",
3331 => x"73822b78",
3332 => x"11880556",
3333 => x"56818019",
3334 => x"08770653",
3335 => x"72097081",
3336 => x"0509060a",
3337 => x"8106ff05",
3338 => x"0980f30b",
3339 => x"f7050684",
3340 => x"01050504",
3341 => x"78167008",
3342 => x"53537951",
3343 => x"74085372",
3344 => x"2dff14fc",
3345 => x"17fc1779",
3346 => x"812c5a57",
3347 => x"57547380",
3348 => x"25ff0509",
3349 => x"c00bf705",
3350 => x"06840105",
3351 => x"05047708",
3352 => x"58770970",
3353 => x"81050906",
3354 => x"0a098106",
3355 => x"ff0509fe",
3356 => x"eb0bf705",
3357 => x"06840105",
3358 => x"05048193",
3359 => x"b40853bc",
3360 => x"13080970",
3361 => x"81050906",
3362 => x"0a098106",
3363 => x"ff0509b9",
3364 => x"0bf70506",
3365 => x"84010505",
3366 => x"047951f1",
3367 => x"f73f7408",
3368 => x"53722dff",
3369 => x"14fc17fc",
3370 => x"1779812c",
3371 => x"5a575754",
3372 => x"738025ff",
3373 => x"0509fedd",
3374 => x"0bf70506",
3375 => x"84010505",
3376 => x"04ff9b39",
3377 => x"8057feb3",
3378 => x"397251bc",
3379 => x"13085473",
3380 => x"2d7951f1",
3381 => x"bf3ffb3d",
3382 => x"0d777a71",
3383 => x"028c05a3",
3384 => x"05335854",
3385 => x"54568373",
3386 => x"27ff0509",
3387 => x"819d0bf7",
3388 => x"05068401",
3389 => x"05050475",
3390 => x"83065170",
3391 => x"09708105",
3392 => x"09060a09",
3393 => x"8106ff05",
3394 => x"0981800b",
3395 => x"f7050684",
3396 => x"01050504",
3397 => x"74882b75",
3398 => x"07707190",
3399 => x"2b075551",
3400 => x"8f7327ff",
3401 => x"0509ba0b",
3402 => x"f7050684",
3403 => x"01050504",
3404 => x"73727084",
3405 => x"05540c71",
3406 => x"74717084",
3407 => x"05530c74",
3408 => x"71708405",
3409 => x"530c7471",
3410 => x"70840553",
3411 => x"0cf01454",
3412 => x"52728f26",
3413 => x"ff0509d8",
3414 => x"0bf70506",
3415 => x"84010505",
3416 => x"04837327",
3417 => x"ff0509a3",
3418 => x"0bf70506",
3419 => x"84010505",
3420 => x"04737270",
3421 => x"8405540c",
3422 => x"fc135372",
3423 => x"8326ff05",
3424 => x"09ef0bf7",
3425 => x"05068401",
3426 => x"050504ff",
3427 => x"13517009",
3428 => x"8105ff05",
3429 => x"09708105",
3430 => x"09060a81",
3431 => x"06ff0509",
3432 => x"b00bf705",
3433 => x"06840105",
3434 => x"05047472",
3435 => x"70810554",
3436 => x"34ff1151",
3437 => x"70098105",
3438 => x"ff050970",
3439 => x"81050906",
3440 => x"0a098106",
3441 => x"ff0509e2",
3442 => x"0bf70506",
3443 => x"84010505",
3444 => x"0475800c",
3445 => x"873d0d04",
3446 => x"70707070",
3447 => x"75707183",
3448 => x"06535552",
3449 => x"70097081",
3450 => x"0509060a",
3451 => x"098106ff",
3452 => x"050980e3",
3453 => x"0bf70506",
3454 => x"84010505",
3455 => x"04717008",
3456 => x"7009f7fb",
3457 => x"fdff1206",
3458 => x"f8848281",
3459 => x"80065452",
3460 => x"53710970",
3461 => x"81050906",
3462 => x"0a098106",
3463 => x"ff0509b5",
3464 => x"0bf70506",
3465 => x"84010505",
3466 => x"04841370",
3467 => x"087009f7",
3468 => x"fbfdff12",
3469 => x"06f88482",
3470 => x"81800654",
3471 => x"52537109",
3472 => x"70810509",
3473 => x"060a8106",
3474 => x"ff0509dd",
3475 => x"0bf70506",
3476 => x"84010505",
3477 => x"04725271",
3478 => x"33537209",
3479 => x"70810509",
3480 => x"060a8106",
3481 => x"ff0509a7",
3482 => x"0bf70506",
3483 => x"84010505",
3484 => x"04811270",
3485 => x"33545272",
3486 => x"09708105",
3487 => x"09060a09",
3488 => x"8106ff05",
3489 => x"09eb0bf7",
3490 => x"05068401",
3491 => x"05050471",
3492 => x"7431800c",
3493 => x"50505050",
3494 => x"04e43d0d",
3495 => x"6ea13d08",
3496 => x"a33d0859",
3497 => x"575f8076",
3498 => x"4d774ea3",
3499 => x"3d08a53d",
3500 => x"08574b75",
3501 => x"4c5e7d6c",
3502 => x"24ff0509",
3503 => x"8b860bf7",
3504 => x"05068401",
3505 => x"05050480",
3506 => x"6a24ff05",
3507 => x"098b9b0b",
3508 => x"f7050684",
3509 => x"01050504",
3510 => x"696b5856",
3511 => x"6b6d5d46",
3512 => x"7b477544",
3513 => x"76456464",
3514 => x"68685c5c",
3515 => x"56567409",
3516 => x"70810509",
3517 => x"060a0981",
3518 => x"06ff0509",
3519 => x"82ee0bf7",
3520 => x"05068401",
3521 => x"05050478",
3522 => x"7627ff05",
3523 => x"09848f0b",
3524 => x"f7050684",
3525 => x"01050504",
3526 => x"7581ff26",
3527 => x"832b5583",
3528 => x"ffff7627",
3529 => x"ff05099f",
3530 => x"0bf70506",
3531 => x"84010505",
3532 => x"049055fe",
3533 => x"800a7627",
3534 => x"ff05098b",
3535 => x"0bf70506",
3536 => x"84010505",
3537 => x"04985575",
3538 => x"752a8188",
3539 => x"88057033",
3540 => x"a0773171",
3541 => x"31575557",
3542 => x"74097081",
3543 => x"0509060a",
3544 => x"8106ff05",
3545 => x"099d0bf7",
3546 => x"05068401",
3547 => x"05050475",
3548 => x"752ba076",
3549 => x"317a772b",
3550 => x"7c722a07",
3551 => x"7c782b5d",
3552 => x"5b595675",
3553 => x"902a7683",
3554 => x"ffff0671",
3555 => x"547a5359",
3556 => x"578c803f",
3557 => x"80085b8b",
3558 => x"e93f8008",
3559 => x"80087929",
3560 => x"7c902b7c",
3561 => x"902a0756",
3562 => x"56597375",
3563 => x"27ff0509",
3564 => x"b20bf705",
3565 => x"06840105",
3566 => x"05048008",
3567 => x"ff057615",
3568 => x"55597574",
3569 => x"26ff0509",
3570 => x"9a0bf705",
3571 => x"06840105",
3572 => x"05047474",
3573 => x"26ff0509",
3574 => x"8b9f0bf7",
3575 => x"05068401",
3576 => x"05050476",
3577 => x"52737531",
3578 => x"518ba83f",
3579 => x"8008558b",
3580 => x"913f8008",
3581 => x"80087929",
3582 => x"7b83ffff",
3583 => x"0677902b",
3584 => x"07565957",
3585 => x"737827ff",
3586 => x"0509a90b",
3587 => x"f7050684",
3588 => x"01050504",
3589 => x"8008ff05",
3590 => x"76155557",
3591 => x"757426ff",
3592 => x"0509910b",
3593 => x"f7050684",
3594 => x"01050504",
3595 => x"77742677",
3596 => x"71315856",
3597 => x"78902b77",
3598 => x"0758805b",
3599 => x"7a407741",
3600 => x"7f615654",
3601 => x"7d097081",
3602 => x"0509060a",
3603 => x"098106ff",
3604 => x"050981ac",
3605 => x"0bf70506",
3606 => x"84010505",
3607 => x"04737f0c",
3608 => x"747f8405",
3609 => x"0c7e800c",
3610 => x"9e3d0d04",
3611 => x"80705c58",
3612 => x"747926ff",
3613 => x"0509c50b",
3614 => x"f7050684",
3615 => x"01050504",
3616 => x"7481ff26",
3617 => x"832b5774",
3618 => x"83ffff26",
3619 => x"ff050983",
3620 => x"e90bf705",
3621 => x"06840105",
3622 => x"05047477",
3623 => x"2a818888",
3624 => x"057033a0",
3625 => x"79317131",
3626 => x"595c5d76",
3627 => x"09708105",
3628 => x"09060a09",
3629 => x"8106ff05",
3630 => x"0983ff0b",
3631 => x"f7050684",
3632 => x"01050504",
3633 => x"76547479",
3634 => x"27ff0509",
3635 => x"8b0bf705",
3636 => x"06840105",
3637 => x"05048154",
3638 => x"79762774",
3639 => x"07598158",
3640 => x"78097081",
3641 => x"0509060a",
3642 => x"098106ff",
3643 => x"0509feca",
3644 => x"0bf70506",
3645 => x"84010505",
3646 => x"04765880",
3647 => x"5bfebd39",
3648 => x"73527453",
3649 => x"9e3de805",
3650 => x"51ffbff2",
3651 => x"3f676956",
3652 => x"7f0c747f",
3653 => x"84050c7e",
3654 => x"800c9e3d",
3655 => x"0d047509",
3656 => x"70810509",
3657 => x"060a8106",
3658 => x"ff050982",
3659 => x"c00bf705",
3660 => x"06840105",
3661 => x"05047581",
3662 => x"ff26832b",
3663 => x"5583ffff",
3664 => x"7627ff05",
3665 => x"099f0bf7",
3666 => x"05068401",
3667 => x"05050490",
3668 => x"55fe800a",
3669 => x"7627ff05",
3670 => x"098b0bf7",
3671 => x"05068401",
3672 => x"05050498",
3673 => x"5575752a",
3674 => x"81888805",
3675 => x"7033a077",
3676 => x"31713157",
3677 => x"5e547409",
3678 => x"70810509",
3679 => x"060a0981",
3680 => x"06ff0509",
3681 => x"86810bf7",
3682 => x"05068401",
3683 => x"05050478",
3684 => x"76315481",
3685 => x"76902a77",
3686 => x"83ffff06",
3687 => x"5f5d5b7b",
3688 => x"52735187",
3689 => x"ee3f8008",
3690 => x"5787d73f",
3691 => x"80088008",
3692 => x"7e297890",
3693 => x"2b7c902a",
3694 => x"07565659",
3695 => x"737527ff",
3696 => x"0509b20b",
3697 => x"f7050684",
3698 => x"01050504",
3699 => x"8008ff05",
3700 => x"76155559",
3701 => x"757426ff",
3702 => x"05099a0b",
3703 => x"f7050684",
3704 => x"01050504",
3705 => x"747426ff",
3706 => x"05098784",
3707 => x"0bf70506",
3708 => x"84010505",
3709 => x"047b5273",
3710 => x"75315187",
3711 => x"963f8008",
3712 => x"5586ff3f",
3713 => x"80088008",
3714 => x"7e297b83",
3715 => x"ffff0677",
3716 => x"902b0756",
3717 => x"59577378",
3718 => x"27ff0509",
3719 => x"a90bf705",
3720 => x"06840105",
3721 => x"05048008",
3722 => x"ff057615",
3723 => x"55577574",
3724 => x"26ff0509",
3725 => x"910bf705",
3726 => x"06840105",
3727 => x"05047774",
3728 => x"26777131",
3729 => x"585a7890",
3730 => x"2b77077b",
3731 => x"41417f61",
3732 => x"56547d09",
3733 => x"70810509",
3734 => x"060a8106",
3735 => x"ff0509fb",
3736 => x"fc0bf705",
3737 => x"06840105",
3738 => x"0504fd94",
3739 => x"39755281",
3740 => x"51868f3f",
3741 => x"800856fd",
3742 => x"bd399057",
3743 => x"fe800a75",
3744 => x"27ff0509",
3745 => x"fc940bf7",
3746 => x"05068401",
3747 => x"05050498",
3748 => x"75712a81",
3749 => x"88880570",
3750 => x"33a07331",
3751 => x"7131535d",
3752 => x"5e577609",
3753 => x"70810509",
3754 => x"060a8106",
3755 => x"ff0509fc",
3756 => x"930bf705",
3757 => x"06840105",
3758 => x"0504a077",
3759 => x"3175782b",
3760 => x"77722a07",
3761 => x"77792b7b",
3762 => x"7a2b7d74",
3763 => x"2a077d7b",
3764 => x"2b73902a",
3765 => x"7483ffff",
3766 => x"0671597f",
3767 => x"772a585e",
3768 => x"5c415f58",
3769 => x"5c5485ab",
3770 => x"3f800854",
3771 => x"85943f80",
3772 => x"08800879",
3773 => x"2975902b",
3774 => x"7e902a07",
3775 => x"56565973",
3776 => x"7527ff05",
3777 => x"09b70bf7",
3778 => x"05068401",
3779 => x"05050480",
3780 => x"08ff057b",
3781 => x"1555597a",
3782 => x"7426ff05",
3783 => x"099f0bf7",
3784 => x"05068401",
3785 => x"05050473",
3786 => x"7527ff05",
3787 => x"098f0bf7",
3788 => x"05068401",
3789 => x"050504ff",
3790 => x"197b1555",
3791 => x"59765273",
3792 => x"75315184",
3793 => x"ce3f8008",
3794 => x"5584b73f",
3795 => x"80088008",
3796 => x"79297d83",
3797 => x"ffff0677",
3798 => x"902b0756",
3799 => x"59577378",
3800 => x"27ff0509",
3801 => x"b70bf705",
3802 => x"06840105",
3803 => x"05048008",
3804 => x"ff057b15",
3805 => x"55577a74",
3806 => x"26ff0509",
3807 => x"9f0bf705",
3808 => x"06840105",
3809 => x"05047378",
3810 => x"27ff0509",
3811 => x"8f0bf705",
3812 => x"06840105",
3813 => x"0504ff17",
3814 => x"7b155557",
3815 => x"73783179",
3816 => x"902b7807",
3817 => x"7083ffff",
3818 => x"0671902a",
3819 => x"7983ffff",
3820 => x"067a902a",
3821 => x"73722973",
3822 => x"73297473",
3823 => x"29767429",
3824 => x"73902a05",
3825 => x"72055755",
3826 => x"435f5b58",
3827 => x"5a57595a",
3828 => x"747c27ff",
3829 => x"05098e0b",
3830 => x"f7050684",
3831 => x"01050504",
3832 => x"84808017",
3833 => x"5774902a",
3834 => x"177983ff",
3835 => x"ff067684",
3836 => x"80802905",
3837 => x"5757767a",
3838 => x"26ff0509",
3839 => x"bf0bf705",
3840 => x"06840105",
3841 => x"0504767a",
3842 => x"32703070",
3843 => x"72078025",
3844 => x"565a5b7c",
3845 => x"7627ff05",
3846 => x"09f89f0b",
3847 => x"f7050684",
3848 => x"01050504",
3849 => x"73097081",
3850 => x"0509060a",
3851 => x"8106ff05",
3852 => x"09f8870b",
3853 => x"f7050684",
3854 => x"01050504",
3855 => x"ff185880",
3856 => x"5bf7f939",
3857 => x"ff765377",
3858 => x"549f3de8",
3859 => x"05525eff",
3860 => x"b9ac3f67",
3861 => x"69574c75",
3862 => x"4d698025",
3863 => x"ff0509f4",
3864 => x"f70bf705",
3865 => x"06840105",
3866 => x"05047d09",
3867 => x"6a6c5c53",
3868 => x"7a549f3d",
3869 => x"e805525e",
3870 => x"ffb9833f",
3871 => x"6769714c",
3872 => x"704d5856",
3873 => x"f4d639a0",
3874 => x"75317676",
3875 => x"2b7a772b",
3876 => x"7c732a07",
3877 => x"7c782b72",
3878 => x"902a7383",
3879 => x"ffff0671",
3880 => x"587e762a",
3881 => x"5742405d",
3882 => x"5d575881",
3883 => x"e63f8008",
3884 => x"5781cf3f",
3885 => x"80088008",
3886 => x"7e297890",
3887 => x"2b7d902a",
3888 => x"07565659",
3889 => x"737527ff",
3890 => x"0509b70b",
3891 => x"f7050684",
3892 => x"01050504",
3893 => x"8008ff05",
3894 => x"76155559",
3895 => x"757426ff",
3896 => x"05099f0b",
3897 => x"f7050684",
3898 => x"01050504",
3899 => x"737527ff",
3900 => x"05098f0b",
3901 => x"f7050684",
3902 => x"01050504",
3903 => x"ff197615",
3904 => x"55597b52",
3905 => x"73753151",
3906 => x"81893f80",
3907 => x"085580f2",
3908 => x"3f800880",
3909 => x"087e297c",
3910 => x"83ffff06",
3911 => x"7078902b",
3912 => x"07515658",
3913 => x"58737727",
3914 => x"ff0509b7",
3915 => x"0bf70506",
3916 => x"84010505",
3917 => x"048008ff",
3918 => x"05761555",
3919 => x"58757426",
3920 => x"ff05099f",
3921 => x"0bf70506",
3922 => x"84010505",
3923 => x"04737727",
3924 => x"ff05098f",
3925 => x"0bf70506",
3926 => x"84010505",
3927 => x"04ff1876",
3928 => x"15555878",
3929 => x"902b7807",
3930 => x"74783155",
3931 => x"5bf8b039",
3932 => x"ff197615",
3933 => x"5559f8fd",
3934 => x"39ff1976",
3935 => x"155559f4",
3936 => x"e2397070",
3937 => x"70805375",
3938 => x"527451ff",
3939 => x"b9d13f50",
3940 => x"50500470",
3941 => x"70708153",
3942 => x"75527451",
3943 => x"ffb9c03f",
3944 => x"50505004",
3945 => x"7070819a",
3946 => x"bc0bfc05",
3947 => x"70085252",
3948 => x"70098105",
3949 => x"ff050970",
3950 => x"81050906",
3951 => x"0a8106ff",
3952 => x"0509ae0b",
3953 => x"f7050684",
3954 => x"01050504",
3955 => x"702dfc12",
3956 => x"70085252",
3957 => x"70098105",
3958 => x"ff050970",
3959 => x"81050906",
3960 => x"0a098106",
3961 => x"ff0509e4",
3962 => x"0bf70506",
3963 => x"84010505",
3964 => x"04505004",
3965 => x"04ff98cc",
3966 => x"3f040000",
3967 => x"30313233",
3968 => x"34353637",
3969 => x"38390000",
3970 => x"44485259",
3971 => x"53544f4e",
3972 => x"45205052",
3973 => x"4f475241",
3974 => x"4d2c2053",
3975 => x"4f4d4520",
3976 => x"53545249",
3977 => x"4e470000",
3978 => x"44485259",
3979 => x"53544f4e",
3980 => x"45205052",
3981 => x"4f475241",
3982 => x"4d2c2031",
3983 => x"27535420",
3984 => x"53545249",
3985 => x"4e470000",
3986 => x"44687279",
3987 => x"73746f6e",
3988 => x"65204265",
3989 => x"6e63686d",
3990 => x"61726b2c",
3991 => x"20566572",
3992 => x"73696f6e",
3993 => x"20322e31",
3994 => x"20284c61",
3995 => x"6e677561",
3996 => x"67653a20",
3997 => x"43290a00",
3998 => x"50726f67",
3999 => x"72616d20",
4000 => x"636f6d70",
4001 => x"696c6564",
4002 => x"20776974",
4003 => x"68202772",
4004 => x"65676973",
4005 => x"74657227",
4006 => x"20617474",
4007 => x"72696275",
4008 => x"74650a00",
4009 => x"45786563",
4010 => x"7574696f",
4011 => x"6e207374",
4012 => x"61727473",
4013 => x"2c202564",
4014 => x"2072756e",
4015 => x"73207468",
4016 => x"726f7567",
4017 => x"68204468",
4018 => x"72797374",
4019 => x"6f6e650a",
4020 => x"00000000",
4021 => x"44485259",
4022 => x"53544f4e",
4023 => x"45205052",
4024 => x"4f475241",
4025 => x"4d2c2032",
4026 => x"274e4420",
4027 => x"53545249",
4028 => x"4e470000",
4029 => x"45786563",
4030 => x"7574696f",
4031 => x"6e20656e",
4032 => x"64730a00",
4033 => x"46696e61",
4034 => x"6c207661",
4035 => x"6c756573",
4036 => x"206f6620",
4037 => x"74686520",
4038 => x"76617269",
4039 => x"61626c65",
4040 => x"73207573",
4041 => x"65642069",
4042 => x"6e207468",
4043 => x"65206265",
4044 => x"6e63686d",
4045 => x"61726b3a",
4046 => x"0a000000",
4047 => x"496e745f",
4048 => x"476c6f62",
4049 => x"3a202020",
4050 => x"20202020",
4051 => x"20202020",
4052 => x"2025640a",
4053 => x"00000000",
4054 => x"20202020",
4055 => x"20202020",
4056 => x"73686f75",
4057 => x"6c642062",
4058 => x"653a2020",
4059 => x"2025640a",
4060 => x"00000000",
4061 => x"426f6f6c",
4062 => x"5f476c6f",
4063 => x"623a2020",
4064 => x"20202020",
4065 => x"20202020",
4066 => x"2025640a",
4067 => x"00000000",
4068 => x"43685f31",
4069 => x"5f476c6f",
4070 => x"623a2020",
4071 => x"20202020",
4072 => x"20202020",
4073 => x"2025630a",
4074 => x"00000000",
4075 => x"20202020",
4076 => x"20202020",
4077 => x"73686f75",
4078 => x"6c642062",
4079 => x"653a2020",
4080 => x"2025630a",
4081 => x"00000000",
4082 => x"43685f32",
4083 => x"5f476c6f",
4084 => x"623a2020",
4085 => x"20202020",
4086 => x"20202020",
4087 => x"2025630a",
4088 => x"00000000",
4089 => x"4172725f",
4090 => x"315f476c",
4091 => x"6f625b38",
4092 => x"5d3a2020",
4093 => x"20202020",
4094 => x"2025640a",
4095 => x"00000000",
4096 => x"4172725f",
4097 => x"325f476c",
4098 => x"6f625b38",
4099 => x"5d5b375d",
4100 => x"3a202020",
4101 => x"2025640a",
4102 => x"00000000",
4103 => x"20202020",
4104 => x"20202020",
4105 => x"73686f75",
4106 => x"6c642062",
4107 => x"653a2020",
4108 => x"204e756d",
4109 => x"6265725f",
4110 => x"4f665f52",
4111 => x"756e7320",
4112 => x"2b203130",
4113 => x"0a000000",
4114 => x"5074725f",
4115 => x"476c6f62",
4116 => x"2d3e0a00",
4117 => x"20205074",
4118 => x"725f436f",
4119 => x"6d703a20",
4120 => x"20202020",
4121 => x"20202020",
4122 => x"2025640a",
4123 => x"00000000",
4124 => x"20202020",
4125 => x"20202020",
4126 => x"73686f75",
4127 => x"6c642062",
4128 => x"653a2020",
4129 => x"2028696d",
4130 => x"706c656d",
4131 => x"656e7461",
4132 => x"74696f6e",
4133 => x"2d646570",
4134 => x"656e6465",
4135 => x"6e74290a",
4136 => x"00000000",
4137 => x"20204469",
4138 => x"7363723a",
4139 => x"20202020",
4140 => x"20202020",
4141 => x"20202020",
4142 => x"2025640a",
4143 => x"00000000",
4144 => x"2020456e",
4145 => x"756d5f43",
4146 => x"6f6d703a",
4147 => x"20202020",
4148 => x"20202020",
4149 => x"2025640a",
4150 => x"00000000",
4151 => x"2020496e",
4152 => x"745f436f",
4153 => x"6d703a20",
4154 => x"20202020",
4155 => x"20202020",
4156 => x"2025640a",
4157 => x"00000000",
4158 => x"20205374",
4159 => x"725f436f",
4160 => x"6d703a20",
4161 => x"20202020",
4162 => x"20202020",
4163 => x"2025730a",
4164 => x"00000000",
4165 => x"20202020",
4166 => x"20202020",
4167 => x"73686f75",
4168 => x"6c642062",
4169 => x"653a2020",
4170 => x"20444852",
4171 => x"5953544f",
4172 => x"4e452050",
4173 => x"524f4752",
4174 => x"414d2c20",
4175 => x"534f4d45",
4176 => x"20535452",
4177 => x"494e470a",
4178 => x"00000000",
4179 => x"4e657874",
4180 => x"5f507472",
4181 => x"5f476c6f",
4182 => x"622d3e0a",
4183 => x"00000000",
4184 => x"20202020",
4185 => x"20202020",
4186 => x"73686f75",
4187 => x"6c642062",
4188 => x"653a2020",
4189 => x"2028696d",
4190 => x"706c656d",
4191 => x"656e7461",
4192 => x"74696f6e",
4193 => x"2d646570",
4194 => x"656e6465",
4195 => x"6e74292c",
4196 => x"2073616d",
4197 => x"65206173",
4198 => x"2061626f",
4199 => x"76650a00",
4200 => x"496e745f",
4201 => x"315f4c6f",
4202 => x"633a2020",
4203 => x"20202020",
4204 => x"20202020",
4205 => x"2025640a",
4206 => x"00000000",
4207 => x"496e745f",
4208 => x"325f4c6f",
4209 => x"633a2020",
4210 => x"20202020",
4211 => x"20202020",
4212 => x"2025640a",
4213 => x"00000000",
4214 => x"496e745f",
4215 => x"335f4c6f",
4216 => x"633a2020",
4217 => x"20202020",
4218 => x"20202020",
4219 => x"2025640a",
4220 => x"00000000",
4221 => x"456e756d",
4222 => x"5f4c6f63",
4223 => x"3a202020",
4224 => x"20202020",
4225 => x"20202020",
4226 => x"2025640a",
4227 => x"00000000",
4228 => x"5374725f",
4229 => x"315f4c6f",
4230 => x"633a2020",
4231 => x"20202020",
4232 => x"20202020",
4233 => x"2025730a",
4234 => x"00000000",
4235 => x"20202020",
4236 => x"20202020",
4237 => x"73686f75",
4238 => x"6c642062",
4239 => x"653a2020",
4240 => x"20444852",
4241 => x"5953544f",
4242 => x"4e452050",
4243 => x"524f4752",
4244 => x"414d2c20",
4245 => x"31275354",
4246 => x"20535452",
4247 => x"494e470a",
4248 => x"00000000",
4249 => x"5374725f",
4250 => x"325f4c6f",
4251 => x"633a2020",
4252 => x"20202020",
4253 => x"20202020",
4254 => x"2025730a",
4255 => x"00000000",
4256 => x"20202020",
4257 => x"20202020",
4258 => x"73686f75",
4259 => x"6c642062",
4260 => x"653a2020",
4261 => x"20444852",
4262 => x"5953544f",
4263 => x"4e452050",
4264 => x"524f4752",
4265 => x"414d2c20",
4266 => x"32274e44",
4267 => x"20535452",
4268 => x"494e470a",
4269 => x"00000000",
4270 => x"55736572",
4271 => x"2074696d",
4272 => x"653a2025",
4273 => x"640a0000",
4274 => x"4d696372",
4275 => x"6f736563",
4276 => x"6f6e6473",
4277 => x"20666f72",
4278 => x"206f6e65",
4279 => x"2072756e",
4280 => x"20746872",
4281 => x"6f756768",
4282 => x"20446872",
4283 => x"7973746f",
4284 => x"6e653a20",
4285 => x"00000000",
4286 => x"2564200a",
4287 => x"00000000",
4288 => x"44687279",
4289 => x"73746f6e",
4290 => x"65732070",
4291 => x"65722053",
4292 => x"65636f6e",
4293 => x"643a2020",
4294 => x"20202020",
4295 => x"20202020",
4296 => x"20202020",
4297 => x"20202020",
4298 => x"20202020",
4299 => x"00000000",
4300 => x"56415820",
4301 => x"4d495053",
4302 => x"20726174",
4303 => x"696e6720",
4304 => x"2a203130",
4305 => x"3030203d",
4306 => x"20256420",
4307 => x"0a000000",
4308 => x"50726f67",
4309 => x"72616d20",
4310 => x"636f6d70",
4311 => x"696c6564",
4312 => x"20776974",
4313 => x"686f7574",
4314 => x"20277265",
4315 => x"67697374",
4316 => x"65722720",
4317 => x"61747472",
4318 => x"69627574",
4319 => x"650a0000",
4320 => x"4d656173",
4321 => x"75726564",
4322 => x"2074696d",
4323 => x"6520746f",
4324 => x"6f20736d",
4325 => x"616c6c20",
4326 => x"746f206f",
4327 => x"62746169",
4328 => x"6e206d65",
4329 => x"616e696e",
4330 => x"6766756c",
4331 => x"20726573",
4332 => x"756c7473",
4333 => x"0a000000",
4334 => x"506c6561",
4335 => x"73652069",
4336 => x"6e637265",
4337 => x"61736520",
4338 => x"6e756d62",
4339 => x"6572206f",
4340 => x"66207275",
4341 => x"6e730a00",
4342 => x"44485259",
4343 => x"53544f4e",
4344 => x"45205052",
4345 => x"4f475241",
4346 => x"4d2c2033",
4347 => x"27524420",
4348 => x"53545249",
4349 => x"4e470000",
4350 => x"43000000",
4351 => x"64756d6d",
4352 => x"792e6578",
4353 => x"65000000",
4354 => x"00010202",
4355 => x"03030303",
4356 => x"04040404",
4357 => x"04040404",
4358 => x"05050505",
4359 => x"05050505",
4360 => x"05050505",
4361 => x"05050505",
4362 => x"06060606",
4363 => x"06060606",
4364 => x"06060606",
4365 => x"06060606",
4366 => x"06060606",
4367 => x"06060606",
4368 => x"06060606",
4369 => x"06060606",
4370 => x"07070707",
4371 => x"07070707",
4372 => x"07070707",
4373 => x"07070707",
4374 => x"07070707",
4375 => x"07070707",
4376 => x"07070707",
4377 => x"07070707",
4378 => x"07070707",
4379 => x"07070707",
4380 => x"07070707",
4381 => x"07070707",
4382 => x"07070707",
4383 => x"07070707",
4384 => x"07070707",
4385 => x"07070707",
4386 => x"08080808",
4387 => x"08080808",
4388 => x"08080808",
4389 => x"08080808",
4390 => x"08080808",
4391 => x"08080808",
4392 => x"08080808",
4393 => x"08080808",
4394 => x"08080808",
4395 => x"08080808",
4396 => x"08080808",
4397 => x"08080808",
4398 => x"08080808",
4399 => x"08080808",
4400 => x"08080808",
4401 => x"08080808",
4402 => x"08080808",
4403 => x"08080808",
4404 => x"08080808",
4405 => x"08080808",
4406 => x"08080808",
4407 => x"08080808",
4408 => x"08080808",
4409 => x"08080808",
4410 => x"08080808",
4411 => x"08080808",
4412 => x"08080808",
4413 => x"08080808",
4414 => x"08080808",
4415 => x"08080808",
4416 => x"08080808",
4417 => x"08080808",
4418 => x"00ffffff",
4419 => x"ff00ffff",
4420 => x"ffff00ff",
4421 => x"ffffff00",
4422 => x"0000042c",
4423 => x"00000446",
4424 => x"0000046c",
4425 => x"00000498",
4426 => x"000004ca",
4427 => x"000004ec",
4428 => x"00000508",
4429 => x"0000052c",
4430 => x"00000556",
4431 => x"00000580",
4432 => x"000005a4",
4433 => x"000005be",
4434 => x"000005e0",
4435 => x"00000612",
4436 => x"0000063e",
4437 => x"00000660",
4438 => x"00000000",
4439 => x"00000000",
4440 => x"00000000",
4441 => x"00004d44",
4442 => x"0000c350",
4443 => x"00000000",
4444 => x"00000000",
4445 => x"00000000",
4446 => x"00000000",
4447 => x"00000000",
4448 => x"00000000",
4449 => x"00000000",
4450 => x"00000000",
4451 => x"00000000",
4452 => x"00000000",
4453 => x"00000000",
4454 => x"00000000",
4455 => x"00000000",
4456 => x"ffffffff",
4457 => x"00000000",
4458 => x"00020000",
4459 => x"00000000",
4460 => x"00000000",
4461 => x"000045ac",
4462 => x"000045ac",
4463 => x"000045b4",
4464 => x"000045b4",
4465 => x"000045bc",
4466 => x"000045bc",
4467 => x"000045c4",
4468 => x"000045c4",
4469 => x"000045cc",
4470 => x"000045cc",
4471 => x"000045d4",
4472 => x"000045d4",
4473 => x"000045dc",
4474 => x"000045dc",
4475 => x"000045e4",
4476 => x"000045e4",
4477 => x"000045ec",
4478 => x"000045ec",
4479 => x"000045f4",
4480 => x"000045f4",
4481 => x"000045fc",
4482 => x"000045fc",
4483 => x"00004604",
4484 => x"00004604",
4485 => x"0000460c",
4486 => x"0000460c",
4487 => x"00004614",
4488 => x"00004614",
4489 => x"0000461c",
4490 => x"0000461c",
4491 => x"00004624",
4492 => x"00004624",
4493 => x"0000462c",
4494 => x"0000462c",
4495 => x"00004634",
4496 => x"00004634",
4497 => x"0000463c",
4498 => x"0000463c",
4499 => x"00004644",
4500 => x"00004644",
4501 => x"0000464c",
4502 => x"0000464c",
4503 => x"00004654",
4504 => x"00004654",
4505 => x"0000465c",
4506 => x"0000465c",
4507 => x"00004664",
4508 => x"00004664",
4509 => x"0000466c",
4510 => x"0000466c",
4511 => x"00004674",
4512 => x"00004674",
4513 => x"0000467c",
4514 => x"0000467c",
4515 => x"00004684",
4516 => x"00004684",
4517 => x"0000468c",
4518 => x"0000468c",
4519 => x"00004694",
4520 => x"00004694",
4521 => x"0000469c",
4522 => x"0000469c",
4523 => x"000046a4",
4524 => x"000046a4",
4525 => x"000046ac",
4526 => x"000046ac",
4527 => x"000046b4",
4528 => x"000046b4",
4529 => x"000046bc",
4530 => x"000046bc",
4531 => x"000046c4",
4532 => x"000046c4",
4533 => x"000046cc",
4534 => x"000046cc",
4535 => x"000046d4",
4536 => x"000046d4",
4537 => x"000046dc",
4538 => x"000046dc",
4539 => x"000046e4",
4540 => x"000046e4",
4541 => x"000046ec",
4542 => x"000046ec",
4543 => x"000046f4",
4544 => x"000046f4",
4545 => x"000046fc",
4546 => x"000046fc",
4547 => x"00004704",
4548 => x"00004704",
4549 => x"0000470c",
4550 => x"0000470c",
4551 => x"00004714",
4552 => x"00004714",
4553 => x"0000471c",
4554 => x"0000471c",
4555 => x"00004724",
4556 => x"00004724",
4557 => x"0000472c",
4558 => x"0000472c",
4559 => x"00004734",
4560 => x"00004734",
4561 => x"0000473c",
4562 => x"0000473c",
4563 => x"00004744",
4564 => x"00004744",
4565 => x"0000474c",
4566 => x"0000474c",
4567 => x"00004754",
4568 => x"00004754",
4569 => x"0000475c",
4570 => x"0000475c",
4571 => x"00004764",
4572 => x"00004764",
4573 => x"0000476c",
4574 => x"0000476c",
4575 => x"00004774",
4576 => x"00004774",
4577 => x"0000477c",
4578 => x"0000477c",
4579 => x"00004784",
4580 => x"00004784",
4581 => x"0000478c",
4582 => x"0000478c",
4583 => x"00004794",
4584 => x"00004794",
4585 => x"0000479c",
4586 => x"0000479c",
4587 => x"000047a4",
4588 => x"000047a4",
4589 => x"000047ac",
4590 => x"000047ac",
4591 => x"000047b4",
4592 => x"000047b4",
4593 => x"000047bc",
4594 => x"000047bc",
4595 => x"000047c4",
4596 => x"000047c4",
4597 => x"000047cc",
4598 => x"000047cc",
4599 => x"000047d4",
4600 => x"000047d4",
4601 => x"000047dc",
4602 => x"000047dc",
4603 => x"000047e4",
4604 => x"000047e4",
4605 => x"000047ec",
4606 => x"000047ec",
4607 => x"000047f4",
4608 => x"000047f4",
4609 => x"000047fc",
4610 => x"000047fc",
4611 => x"00004804",
4612 => x"00004804",
4613 => x"0000480c",
4614 => x"0000480c",
4615 => x"00004814",
4616 => x"00004814",
4617 => x"0000481c",
4618 => x"0000481c",
4619 => x"00004824",
4620 => x"00004824",
4621 => x"0000482c",
4622 => x"0000482c",
4623 => x"00004834",
4624 => x"00004834",
4625 => x"0000483c",
4626 => x"0000483c",
4627 => x"00004844",
4628 => x"00004844",
4629 => x"0000484c",
4630 => x"0000484c",
4631 => x"00004854",
4632 => x"00004854",
4633 => x"0000485c",
4634 => x"0000485c",
4635 => x"00004864",
4636 => x"00004864",
4637 => x"0000486c",
4638 => x"0000486c",
4639 => x"00004874",
4640 => x"00004874",
4641 => x"0000487c",
4642 => x"0000487c",
4643 => x"00004884",
4644 => x"00004884",
4645 => x"0000488c",
4646 => x"0000488c",
4647 => x"00004894",
4648 => x"00004894",
4649 => x"0000489c",
4650 => x"0000489c",
4651 => x"000048a4",
4652 => x"000048a4",
4653 => x"000048ac",
4654 => x"000048ac",
4655 => x"000048b4",
4656 => x"000048b4",
4657 => x"000048bc",
4658 => x"000048bc",
4659 => x"000048c4",
4660 => x"000048c4",
4661 => x"000048cc",
4662 => x"000048cc",
4663 => x"000048d4",
4664 => x"000048d4",
4665 => x"000048dc",
4666 => x"000048dc",
4667 => x"000048e4",
4668 => x"000048e4",
4669 => x"000048ec",
4670 => x"000048ec",
4671 => x"000048f4",
4672 => x"000048f4",
4673 => x"000048fc",
4674 => x"000048fc",
4675 => x"00004904",
4676 => x"00004904",
4677 => x"0000490c",
4678 => x"0000490c",
4679 => x"00004914",
4680 => x"00004914",
4681 => x"0000491c",
4682 => x"0000491c",
4683 => x"00004924",
4684 => x"00004924",
4685 => x"0000492c",
4686 => x"0000492c",
4687 => x"00004934",
4688 => x"00004934",
4689 => x"0000493c",
4690 => x"0000493c",
4691 => x"00004944",
4692 => x"00004944",
4693 => x"0000494c",
4694 => x"0000494c",
4695 => x"00004954",
4696 => x"00004954",
4697 => x"0000495c",
4698 => x"0000495c",
4699 => x"00004964",
4700 => x"00004964",
4701 => x"0000496c",
4702 => x"0000496c",
4703 => x"00004974",
4704 => x"00004974",
4705 => x"0000497c",
4706 => x"0000497c",
4707 => x"00004984",
4708 => x"00004984",
4709 => x"0000498c",
4710 => x"0000498c",
4711 => x"00004994",
4712 => x"00004994",
4713 => x"0000499c",
4714 => x"0000499c",
4715 => x"000049a4",
4716 => x"000049a4",
4717 => x"000049b8",
4718 => x"00000000",
4719 => x"00004c20",
4720 => x"00004c7c",
4721 => x"00004cd8",
4722 => x"00000000",
4723 => x"00000000",
4724 => x"00000000",
4725 => x"00000000",
4726 => x"00000000",
4727 => x"00000000",
4728 => x"00000000",
4729 => x"00000000",
4730 => x"00000000",
4731 => x"000043f8",
4732 => x"00000000",
4733 => x"00000000",
4734 => x"00000000",
4735 => x"00000000",
4736 => x"00000000",
4737 => x"00000000",
4738 => x"00000000",
4739 => x"00000000",
4740 => x"00000000",
4741 => x"00000000",
4742 => x"00000000",
4743 => x"00000000",
4744 => x"00000000",
4745 => x"00000000",
4746 => x"00000000",
4747 => x"00000000",
4748 => x"00000000",
4749 => x"00000000",
4750 => x"00000000",
4751 => x"00000000",
4752 => x"00000000",
4753 => x"00000000",
4754 => x"00000000",
4755 => x"00000000",
4756 => x"00000000",
4757 => x"00000000",
4758 => x"00000000",
4759 => x"00000000",
4760 => x"00000001",
4761 => x"330eabcd",
4762 => x"1234e66d",
4763 => x"deec0005",
4764 => x"000b0000",
4765 => x"00000000",
4766 => x"00000000",
4767 => x"00000000",
4768 => x"00000000",
4769 => x"00000000",
4770 => x"00000000",
4771 => x"00000000",
4772 => x"00000000",
4773 => x"00000000",
4774 => x"00000000",
4775 => x"00000000",
4776 => x"00000000",
4777 => x"00000000",
4778 => x"00000000",
4779 => x"00000000",
4780 => x"00000000",
4781 => x"00000000",
4782 => x"00000000",
4783 => x"00000000",
4784 => x"00000000",
4785 => x"00000000",
4786 => x"00000000",
4787 => x"00000000",
4788 => x"00000000",
4789 => x"00000000",
4790 => x"00000000",
4791 => x"00000000",
4792 => x"00000000",
4793 => x"00000000",
4794 => x"00000000",
4795 => x"00000000",
4796 => x"00000000",
4797 => x"00000000",
4798 => x"00000000",
4799 => x"00000000",
4800 => x"00000000",
4801 => x"00000000",
4802 => x"00000000",
4803 => x"00000000",
4804 => x"00000000",
4805 => x"00000000",
4806 => x"00000000",
4807 => x"00000000",
4808 => x"00000000",
4809 => x"00000000",
4810 => x"00000000",
4811 => x"00000000",
4812 => x"00000000",
4813 => x"00000000",
4814 => x"00000000",
4815 => x"00000000",
4816 => x"00000000",
4817 => x"00000000",
4818 => x"00000000",
4819 => x"00000000",
4820 => x"00000000",
4821 => x"00000000",
4822 => x"00000000",
4823 => x"00000000",
4824 => x"00000000",
4825 => x"00000000",
4826 => x"00000000",
4827 => x"00000000",
4828 => x"00000000",
4829 => x"00000000",
4830 => x"00000000",
4831 => x"00000000",
4832 => x"00000000",
4833 => x"00000000",
4834 => x"00000000",
4835 => x"00000000",
4836 => x"00000000",
4837 => x"00000000",
4838 => x"00000000",
4839 => x"00000000",
4840 => x"00000000",
4841 => x"00000000",
4842 => x"00000000",
4843 => x"00000000",
4844 => x"00000000",
4845 => x"00000000",
4846 => x"00000000",
4847 => x"00000000",
4848 => x"00000000",
4849 => x"00000000",
4850 => x"00000000",
4851 => x"00000000",
4852 => x"00000000",
4853 => x"00000000",
4854 => x"00000000",
4855 => x"00000000",
4856 => x"00000000",
4857 => x"00000000",
4858 => x"00000000",
4859 => x"00000000",
4860 => x"00000000",
4861 => x"00000000",
4862 => x"00000000",
4863 => x"00000000",
4864 => x"00000000",
4865 => x"00000000",
4866 => x"00000000",
4867 => x"00000000",
4868 => x"00000000",
4869 => x"00000000",
4870 => x"00000000",
4871 => x"00000000",
4872 => x"00000000",
4873 => x"00000000",
4874 => x"00000000",
4875 => x"00000000",
4876 => x"00000000",
4877 => x"00000000",
4878 => x"00000000",
4879 => x"00000000",
4880 => x"00000000",
4881 => x"00000000",
4882 => x"00000000",
4883 => x"00000000",
4884 => x"00000000",
4885 => x"00000000",
4886 => x"00000000",
4887 => x"00000000",
4888 => x"00000000",
4889 => x"00000000",
4890 => x"00000000",
4891 => x"00000000",
4892 => x"00000000",
4893 => x"00000000",
4894 => x"00000000",
4895 => x"00000000",
4896 => x"00000000",
4897 => x"00000000",
4898 => x"00000000",
4899 => x"00000000",
4900 => x"00000000",
4901 => x"00000000",
4902 => x"00000000",
4903 => x"00000000",
4904 => x"00000000",
4905 => x"00000000",
4906 => x"00000000",
4907 => x"00000000",
4908 => x"00000000",
4909 => x"00000000",
4910 => x"00000000",
4911 => x"00000000",
4912 => x"00000000",
4913 => x"00000000",
4914 => x"00000000",
4915 => x"00000000",
4916 => x"00000000",
4917 => x"00000000",
4918 => x"00000000",
4919 => x"00000000",
4920 => x"00000000",
4921 => x"00000000",
4922 => x"00000000",
4923 => x"00000000",
4924 => x"00000000",
4925 => x"00000000",
4926 => x"00000000",
4927 => x"00000000",
4928 => x"00000000",
4929 => x"00000000",
4930 => x"00000000",
4931 => x"00000000",
4932 => x"00000000",
4933 => x"00000000",
4934 => x"00000000",
4935 => x"00000000",
4936 => x"00000000",
4937 => x"00000000",
4938 => x"00000000",
4939 => x"00000000",
4940 => x"00000000",
4941 => x"000043fc",
4942 => x"ffffffff",
4943 => x"00000000",
4944 => x"ffffffff",
4945 => x"00000000",
	others => x"00000000"
);

attribute syn_ramstyle : string;
attribute syn_ramstyle of ram : signal is "no_rw_check" ;

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') then
			ram(conv_integer(memAAddr)) <= memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(conv_integer(memAAddr));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(conv_integer(memBAddr)) <= memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(conv_integer(memBAddr));
		end if;
	end if;
end process;




end dualport_ram_arch;
