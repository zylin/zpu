-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80d1c40c",
     3 => x"3a0b0b80",
     4 => x"c9b30400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80c9fe2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80d1",
   162 => x"b0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8b",
   171 => x"932d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8c",
   179 => x"c52d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80d1c00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82c73f80",
   257 => x"c8c63f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"fe3d0d0b",
   281 => x"0b80e1ac",
   282 => x"08538413",
   283 => x"0870882a",
   284 => x"70810651",
   285 => x"52527080",
   286 => x"2ef03871",
   287 => x"81ff0680",
   288 => x"0c843d0d",
   289 => x"04ff3d0d",
   290 => x"0b0b80e1",
   291 => x"ac085271",
   292 => x"0870882a",
   293 => x"81327081",
   294 => x"06515151",
   295 => x"70f13873",
   296 => x"720c833d",
   297 => x"0d0480d1",
   298 => x"c008802e",
   299 => x"a43880d1",
   300 => x"c408822e",
   301 => x"bd388380",
   302 => x"800b0b0b",
   303 => x"80e1ac0c",
   304 => x"82a0800b",
   305 => x"80e1b00c",
   306 => x"8290800b",
   307 => x"80e1b40c",
   308 => x"04f88080",
   309 => x"80a40b0b",
   310 => x"0b80e1ac",
   311 => x"0cf88080",
   312 => x"82800b80",
   313 => x"e1b00cf8",
   314 => x"80808480",
   315 => x"0b80e1b4",
   316 => x"0c0480c0",
   317 => x"a8808c0b",
   318 => x"0b0b80e1",
   319 => x"ac0c80c0",
   320 => x"a880940b",
   321 => x"80e1b00c",
   322 => x"0b0b80d0",
   323 => x"f80b80e1",
   324 => x"b40c04ff",
   325 => x"3d0d80e1",
   326 => x"b8335170",
   327 => x"a73880d1",
   328 => x"cc087008",
   329 => x"52527080",
   330 => x"2e943884",
   331 => x"1280d1cc",
   332 => x"0c702d80",
   333 => x"d1cc0870",
   334 => x"08525270",
   335 => x"ee38810b",
   336 => x"80e1b834",
   337 => x"833d0d04",
   338 => x"04803d0d",
   339 => x"0b0b80e1",
   340 => x"a808802e",
   341 => x"8e380b0b",
   342 => x"0b0b800b",
   343 => x"802e0981",
   344 => x"06853882",
   345 => x"3d0d040b",
   346 => x"0b80e1a8",
   347 => x"510b0b0b",
   348 => x"f58e3f82",
   349 => x"3d0d0404",
   350 => x"ff3d0d80",
   351 => x"d0fc5185",
   352 => x"f43f80c0",
   353 => x"80a4b408",
   354 => x"5280d194",
   355 => x"5185e63f",
   356 => x"83fd3f8c",
   357 => x"08028c0c",
   358 => x"f93d0d80",
   359 => x"0b8c08fc",
   360 => x"050c8c08",
   361 => x"88050880",
   362 => x"25ab388c",
   363 => x"08880508",
   364 => x"308c0888",
   365 => x"050c800b",
   366 => x"8c08f405",
   367 => x"0c8c08fc",
   368 => x"05088838",
   369 => x"810b8c08",
   370 => x"f4050c8c",
   371 => x"08f40508",
   372 => x"8c08fc05",
   373 => x"0c8c088c",
   374 => x"05088025",
   375 => x"ab388c08",
   376 => x"8c050830",
   377 => x"8c088c05",
   378 => x"0c800b8c",
   379 => x"08f0050c",
   380 => x"8c08fc05",
   381 => x"08883881",
   382 => x"0b8c08f0",
   383 => x"050c8c08",
   384 => x"f005088c",
   385 => x"08fc050c",
   386 => x"80538c08",
   387 => x"8c050852",
   388 => x"8c088805",
   389 => x"085181a7",
   390 => x"3f800870",
   391 => x"8c08f805",
   392 => x"0c548c08",
   393 => x"fc050880",
   394 => x"2e8c388c",
   395 => x"08f80508",
   396 => x"308c08f8",
   397 => x"050c8c08",
   398 => x"f8050870",
   399 => x"800c5489",
   400 => x"3d0d8c0c",
   401 => x"048c0802",
   402 => x"8c0cfb3d",
   403 => x"0d800b8c",
   404 => x"08fc050c",
   405 => x"8c088805",
   406 => x"08802593",
   407 => x"388c0888",
   408 => x"0508308c",
   409 => x"0888050c",
   410 => x"810b8c08",
   411 => x"fc050c8c",
   412 => x"088c0508",
   413 => x"80258c38",
   414 => x"8c088c05",
   415 => x"08308c08",
   416 => x"8c050c81",
   417 => x"538c088c",
   418 => x"0508528c",
   419 => x"08880508",
   420 => x"51ad3f80",
   421 => x"08708c08",
   422 => x"f8050c54",
   423 => x"8c08fc05",
   424 => x"08802e8c",
   425 => x"388c08f8",
   426 => x"0508308c",
   427 => x"08f8050c",
   428 => x"8c08f805",
   429 => x"0870800c",
   430 => x"54873d0d",
   431 => x"8c0c048c",
   432 => x"08028c0c",
   433 => x"fd3d0d81",
   434 => x"0b8c08fc",
   435 => x"050c800b",
   436 => x"8c08f805",
   437 => x"0c8c088c",
   438 => x"05088c08",
   439 => x"88050827",
   440 => x"ac388c08",
   441 => x"fc050880",
   442 => x"2ea33880",
   443 => x"0b8c088c",
   444 => x"05082499",
   445 => x"388c088c",
   446 => x"0508108c",
   447 => x"088c050c",
   448 => x"8c08fc05",
   449 => x"08108c08",
   450 => x"fc050cc9",
   451 => x"398c08fc",
   452 => x"0508802e",
   453 => x"80c9388c",
   454 => x"088c0508",
   455 => x"8c088805",
   456 => x"0826a138",
   457 => x"8c088805",
   458 => x"088c088c",
   459 => x"0508318c",
   460 => x"0888050c",
   461 => x"8c08f805",
   462 => x"088c08fc",
   463 => x"0508078c",
   464 => x"08f8050c",
   465 => x"8c08fc05",
   466 => x"08812a8c",
   467 => x"08fc050c",
   468 => x"8c088c05",
   469 => x"08812a8c",
   470 => x"088c050c",
   471 => x"ffaf398c",
   472 => x"08900508",
   473 => x"802e8f38",
   474 => x"8c088805",
   475 => x"08708c08",
   476 => x"f4050c51",
   477 => x"8d398c08",
   478 => x"f8050870",
   479 => x"8c08f405",
   480 => x"0c518c08",
   481 => x"f4050880",
   482 => x"0c853d0d",
   483 => x"8c0c0480",
   484 => x"3d0d8651",
   485 => x"84e73f81",
   486 => x"51bae03f",
   487 => x"fc3d0d76",
   488 => x"70797b55",
   489 => x"5555558f",
   490 => x"72278c38",
   491 => x"72750783",
   492 => x"06517080",
   493 => x"2ea738ff",
   494 => x"125271ff",
   495 => x"2e983872",
   496 => x"70810554",
   497 => x"33747081",
   498 => x"055634ff",
   499 => x"125271ff",
   500 => x"2e098106",
   501 => x"ea387480",
   502 => x"0c863d0d",
   503 => x"04745172",
   504 => x"70840554",
   505 => x"08717084",
   506 => x"05530c72",
   507 => x"70840554",
   508 => x"08717084",
   509 => x"05530c72",
   510 => x"70840554",
   511 => x"08717084",
   512 => x"05530c72",
   513 => x"70840554",
   514 => x"08717084",
   515 => x"05530cf0",
   516 => x"1252718f",
   517 => x"26c93883",
   518 => x"72279538",
   519 => x"72708405",
   520 => x"54087170",
   521 => x"8405530c",
   522 => x"fc125271",
   523 => x"8326ed38",
   524 => x"7054ff83",
   525 => x"39f73d0d",
   526 => x"7c705253",
   527 => x"84bd3f72",
   528 => x"54800855",
   529 => x"80d19c56",
   530 => x"81578008",
   531 => x"81055a8b",
   532 => x"3de41159",
   533 => x"538259f4",
   534 => x"13527b88",
   535 => x"11085253",
   536 => x"84f83f80",
   537 => x"08307080",
   538 => x"08079f2c",
   539 => x"8a07800c",
   540 => x"538b3d0d",
   541 => x"04ff3d0d",
   542 => x"735280d1",
   543 => x"d00851ff",
   544 => x"b43f833d",
   545 => x"0d04fd3d",
   546 => x"0d755384",
   547 => x"d8130880",
   548 => x"2e8a3880",
   549 => x"5372800c",
   550 => x"853d0d04",
   551 => x"81805272",
   552 => x"518a9e3f",
   553 => x"800884d8",
   554 => x"140cff53",
   555 => x"8008802e",
   556 => x"e4388008",
   557 => x"549f5380",
   558 => x"74708405",
   559 => x"560cff13",
   560 => x"53807324",
   561 => x"ce388074",
   562 => x"70840556",
   563 => x"0cff1353",
   564 => x"728025e3",
   565 => x"38ffbc39",
   566 => x"fd3d0d75",
   567 => x"7755539f",
   568 => x"74278d38",
   569 => x"96730cff",
   570 => x"5271800c",
   571 => x"853d0d04",
   572 => x"84d81308",
   573 => x"5271802e",
   574 => x"93387310",
   575 => x"10127008",
   576 => x"79720c51",
   577 => x"5271800c",
   578 => x"853d0d04",
   579 => x"7251fef6",
   580 => x"3fff5280",
   581 => x"08d33884",
   582 => x"d8130874",
   583 => x"10101170",
   584 => x"087a720c",
   585 => x"515152dd",
   586 => x"39f93d0d",
   587 => x"797b5856",
   588 => x"769f2680",
   589 => x"e83884d8",
   590 => x"16085473",
   591 => x"802eaa38",
   592 => x"76101014",
   593 => x"70085555",
   594 => x"73802eba",
   595 => x"38805873",
   596 => x"812e8f38",
   597 => x"73ff2ea3",
   598 => x"3880750c",
   599 => x"7651732d",
   600 => x"80587780",
   601 => x"0c893d0d",
   602 => x"047551fe",
   603 => x"993fff58",
   604 => x"8008ef38",
   605 => x"84d81608",
   606 => x"54c63996",
   607 => x"760c810b",
   608 => x"800c893d",
   609 => x"0d047551",
   610 => x"81ed3f76",
   611 => x"53800852",
   612 => x"755181ad",
   613 => x"3f800880",
   614 => x"0c893d0d",
   615 => x"0496760c",
   616 => x"ff0b800c",
   617 => x"893d0d04",
   618 => x"fc3d0d76",
   619 => x"785653ff",
   620 => x"54749f26",
   621 => x"b13884d8",
   622 => x"13085271",
   623 => x"802eae38",
   624 => x"74101012",
   625 => x"70085353",
   626 => x"81547180",
   627 => x"2e983882",
   628 => x"5471ff2e",
   629 => x"91388354",
   630 => x"71812e8a",
   631 => x"3880730c",
   632 => x"7451712d",
   633 => x"80547380",
   634 => x"0c863d0d",
   635 => x"047251fd",
   636 => x"953f8008",
   637 => x"f13884d8",
   638 => x"130852c4",
   639 => x"39ff3d0d",
   640 => x"735280d1",
   641 => x"d00851fe",
   642 => x"a03f833d",
   643 => x"0d04fe3d",
   644 => x"0d755374",
   645 => x"5280d1d0",
   646 => x"0851fdbc",
   647 => x"3f843d0d",
   648 => x"04803d0d",
   649 => x"80d1d008",
   650 => x"51fcdb3f",
   651 => x"823d0d04",
   652 => x"ff3d0d73",
   653 => x"5280d1d0",
   654 => x"0851feec",
   655 => x"3f833d0d",
   656 => x"04fc3d0d",
   657 => x"800b80e1",
   658 => x"c40c7852",
   659 => x"7751b49d",
   660 => x"3f800854",
   661 => x"8008ff2e",
   662 => x"88387380",
   663 => x"0c863d0d",
   664 => x"0480e1c4",
   665 => x"08557480",
   666 => x"2ef03876",
   667 => x"75710c53",
   668 => x"73800c86",
   669 => x"3d0d04b3",
   670 => x"ef3f04fd",
   671 => x"3d0d7570",
   672 => x"71830653",
   673 => x"555270b8",
   674 => x"38717008",
   675 => x"7009f7fb",
   676 => x"fdff1206",
   677 => x"70f88482",
   678 => x"81800651",
   679 => x"51525370",
   680 => x"9d388413",
   681 => x"70087009",
   682 => x"f7fbfdff",
   683 => x"120670f8",
   684 => x"84828180",
   685 => x"06515152",
   686 => x"5370802e",
   687 => x"e5387252",
   688 => x"71335170",
   689 => x"802e8a38",
   690 => x"81127033",
   691 => x"525270f8",
   692 => x"38717431",
   693 => x"800c853d",
   694 => x"0d04f23d",
   695 => x"0d606288",
   696 => x"11087057",
   697 => x"575f5a74",
   698 => x"802e8190",
   699 => x"388c1a22",
   700 => x"70832a81",
   701 => x"32708106",
   702 => x"51555873",
   703 => x"8638901a",
   704 => x"08913879",
   705 => x"519ccd3f",
   706 => x"ff548008",
   707 => x"80ee388c",
   708 => x"1a22587d",
   709 => x"08578078",
   710 => x"83ffff06",
   711 => x"700a100a",
   712 => x"70810651",
   713 => x"56575573",
   714 => x"752e80d7",
   715 => x"38749038",
   716 => x"76088418",
   717 => x"08881959",
   718 => x"56597480",
   719 => x"2ef23874",
   720 => x"54888075",
   721 => x"27843888",
   722 => x"80547353",
   723 => x"78529c1a",
   724 => x"0851a41a",
   725 => x"0854732d",
   726 => x"800b8008",
   727 => x"2582e638",
   728 => x"80081975",
   729 => x"8008317f",
   730 => x"88050880",
   731 => x"08317061",
   732 => x"88050c56",
   733 => x"565973ff",
   734 => x"b4388054",
   735 => x"73800c90",
   736 => x"3d0d0475",
   737 => x"81327081",
   738 => x"06764151",
   739 => x"5473802e",
   740 => x"81c13874",
   741 => x"90387608",
   742 => x"84180888",
   743 => x"19595659",
   744 => x"74802ef2",
   745 => x"38881a08",
   746 => x"7883ffff",
   747 => x"0670892a",
   748 => x"70810651",
   749 => x"56595673",
   750 => x"802e82fa",
   751 => x"38757527",
   752 => x"8d387787",
   753 => x"2a708106",
   754 => x"51547382",
   755 => x"b5387476",
   756 => x"27833874",
   757 => x"56755378",
   758 => x"52790851",
   759 => x"90f83f88",
   760 => x"1a087631",
   761 => x"881b0c79",
   762 => x"08167a0c",
   763 => x"74567519",
   764 => x"7577317f",
   765 => x"88050878",
   766 => x"31706188",
   767 => x"050c5656",
   768 => x"5973802e",
   769 => x"fef4388c",
   770 => x"1a2258ff",
   771 => x"86397778",
   772 => x"5479537b",
   773 => x"525690be",
   774 => x"3f881a08",
   775 => x"7831881b",
   776 => x"0c790818",
   777 => x"7a0c7c76",
   778 => x"315d7c8e",
   779 => x"3879519c",
   780 => x"873f8008",
   781 => x"818f3880",
   782 => x"085f7519",
   783 => x"7577317f",
   784 => x"88050878",
   785 => x"31706188",
   786 => x"050c5656",
   787 => x"5973802e",
   788 => x"fea83874",
   789 => x"81833876",
   790 => x"08841808",
   791 => x"88195956",
   792 => x"5974802e",
   793 => x"f2387453",
   794 => x"8a527851",
   795 => x"8ec93f80",
   796 => x"08793181",
   797 => x"055d8008",
   798 => x"84388115",
   799 => x"5d815f7c",
   800 => x"58747d27",
   801 => x"83387458",
   802 => x"941a0888",
   803 => x"1b081157",
   804 => x"5c807a08",
   805 => x"5c54901a",
   806 => x"087b2783",
   807 => x"38815475",
   808 => x"78258438",
   809 => x"73ba387b",
   810 => x"7824fee2",
   811 => x"387b5378",
   812 => x"529c1a08",
   813 => x"51a41a08",
   814 => x"54732d80",
   815 => x"08568008",
   816 => x"8024fee2",
   817 => x"388c1a22",
   818 => x"80c00754",
   819 => x"738c1b23",
   820 => x"ff547380",
   821 => x"0c903d0d",
   822 => x"047effa3",
   823 => x"38ff8739",
   824 => x"75537852",
   825 => x"7a518eee",
   826 => x"3f790816",
   827 => x"7a0c7951",
   828 => x"9ac63f80",
   829 => x"08cf387c",
   830 => x"76315d7c",
   831 => x"febc38fe",
   832 => x"ac39901a",
   833 => x"087a0871",
   834 => x"31761170",
   835 => x"565a5752",
   836 => x"80d1d008",
   837 => x"5190843f",
   838 => x"8008802e",
   839 => x"ffa73880",
   840 => x"08901b0c",
   841 => x"8008167a",
   842 => x"0c77941b",
   843 => x"0c74881b",
   844 => x"0c7456fd",
   845 => x"99397908",
   846 => x"58901a08",
   847 => x"78278338",
   848 => x"81547575",
   849 => x"27843873",
   850 => x"b338941a",
   851 => x"08567575",
   852 => x"2680d338",
   853 => x"75537852",
   854 => x"9c1a0851",
   855 => x"a41a0854",
   856 => x"732d8008",
   857 => x"56800880",
   858 => x"24fd8338",
   859 => x"8c1a2280",
   860 => x"c0075473",
   861 => x"8c1b23ff",
   862 => x"54fed739",
   863 => x"75537852",
   864 => x"77518dd2",
   865 => x"3f790816",
   866 => x"7a0c7951",
   867 => x"99aa3f80",
   868 => x"08802efc",
   869 => x"d9388c1a",
   870 => x"2280c007",
   871 => x"54738c1b",
   872 => x"23ff54fe",
   873 => x"ad397475",
   874 => x"54795378",
   875 => x"52568da6",
   876 => x"3f881a08",
   877 => x"7531881b",
   878 => x"0c790815",
   879 => x"7a0cfcae",
   880 => x"39f33d0d",
   881 => x"7f618b11",
   882 => x"70f8065c",
   883 => x"55555e72",
   884 => x"96268338",
   885 => x"90598079",
   886 => x"24747a26",
   887 => x"07538054",
   888 => x"72742e09",
   889 => x"810680cb",
   890 => x"387d518e",
   891 => x"ac3f7883",
   892 => x"f72680c6",
   893 => x"3878832a",
   894 => x"70101010",
   895 => x"80d98c05",
   896 => x"8c110859",
   897 => x"595a7678",
   898 => x"2e83b038",
   899 => x"841708fc",
   900 => x"06568c17",
   901 => x"08881808",
   902 => x"718c120c",
   903 => x"88120c58",
   904 => x"75178411",
   905 => x"08810784",
   906 => x"120c537d",
   907 => x"518deb3f",
   908 => x"88175473",
   909 => x"800c8f3d",
   910 => x"0d047889",
   911 => x"2a79832a",
   912 => x"5b537280",
   913 => x"2ebf3878",
   914 => x"862ab805",
   915 => x"5a847327",
   916 => x"b43880db",
   917 => x"135a9473",
   918 => x"27ab3878",
   919 => x"8c2a80ee",
   920 => x"055a80d4",
   921 => x"73279e38",
   922 => x"788f2a80",
   923 => x"f7055a82",
   924 => x"d4732791",
   925 => x"3878922a",
   926 => x"80fc055a",
   927 => x"8ad47327",
   928 => x"843880fe",
   929 => x"5a791010",
   930 => x"1080d98c",
   931 => x"058c1108",
   932 => x"58557675",
   933 => x"2ea33884",
   934 => x"1708fc06",
   935 => x"707a3155",
   936 => x"56738f24",
   937 => x"88d53873",
   938 => x"8025fee6",
   939 => x"388c1708",
   940 => x"5776752e",
   941 => x"098106df",
   942 => x"38811a5a",
   943 => x"80d99c08",
   944 => x"577680d9",
   945 => x"942e82c0",
   946 => x"38841708",
   947 => x"fc06707a",
   948 => x"31555673",
   949 => x"8f2481f9",
   950 => x"3880d994",
   951 => x"0b80d9a0",
   952 => x"0c80d994",
   953 => x"0b80d99c",
   954 => x"0c738025",
   955 => x"feb23883",
   956 => x"ff762783",
   957 => x"df387589",
   958 => x"2a76832a",
   959 => x"55537280",
   960 => x"2ebf3875",
   961 => x"862ab805",
   962 => x"54847327",
   963 => x"b43880db",
   964 => x"13549473",
   965 => x"27ab3875",
   966 => x"8c2a80ee",
   967 => x"055480d4",
   968 => x"73279e38",
   969 => x"758f2a80",
   970 => x"f7055482",
   971 => x"d4732791",
   972 => x"3875922a",
   973 => x"80fc0554",
   974 => x"8ad47327",
   975 => x"843880fe",
   976 => x"54731010",
   977 => x"1080d98c",
   978 => x"05881108",
   979 => x"56587478",
   980 => x"2e86cf38",
   981 => x"841508fc",
   982 => x"06537573",
   983 => x"278d3888",
   984 => x"15085574",
   985 => x"782e0981",
   986 => x"06ea388c",
   987 => x"150880d9",
   988 => x"8c0b8405",
   989 => x"08718c1a",
   990 => x"0c76881a",
   991 => x"0c788813",
   992 => x"0c788c18",
   993 => x"0c5d5879",
   994 => x"53807a24",
   995 => x"83e63872",
   996 => x"822c8171",
   997 => x"2b5c537a",
   998 => x"7c268198",
   999 => x"387b7b06",
  1000 => x"537282f1",
  1001 => x"3879fc06",
  1002 => x"84055a7a",
  1003 => x"10707d06",
  1004 => x"545b7282",
  1005 => x"e038841a",
  1006 => x"5af13988",
  1007 => x"178c1108",
  1008 => x"58587678",
  1009 => x"2e098106",
  1010 => x"fcc23882",
  1011 => x"1a5afdec",
  1012 => x"39781779",
  1013 => x"81078419",
  1014 => x"0c7080d9",
  1015 => x"a00c7080",
  1016 => x"d99c0c80",
  1017 => x"d9940b8c",
  1018 => x"120c8c11",
  1019 => x"0888120c",
  1020 => x"74810784",
  1021 => x"120c7411",
  1022 => x"75710c51",
  1023 => x"537d518a",
  1024 => x"993f8817",
  1025 => x"54fcac39",
  1026 => x"80d98c0b",
  1027 => x"8405087a",
  1028 => x"545c7980",
  1029 => x"25fef838",
  1030 => x"82da397a",
  1031 => x"097c0670",
  1032 => x"80d98c0b",
  1033 => x"84050c5c",
  1034 => x"7a105b7a",
  1035 => x"7c268538",
  1036 => x"7a85b838",
  1037 => x"80d98c0b",
  1038 => x"88050870",
  1039 => x"841208fc",
  1040 => x"06707c31",
  1041 => x"7c72268f",
  1042 => x"72250757",
  1043 => x"575c5d55",
  1044 => x"72802e80",
  1045 => x"db38797a",
  1046 => x"1680d984",
  1047 => x"081b9011",
  1048 => x"5a55575b",
  1049 => x"80d98008",
  1050 => x"ff2e8838",
  1051 => x"a08f13e0",
  1052 => x"80065776",
  1053 => x"527d5191",
  1054 => x"a73f8008",
  1055 => x"548008ff",
  1056 => x"2e903880",
  1057 => x"08762782",
  1058 => x"99387480",
  1059 => x"d98c2e82",
  1060 => x"913880d9",
  1061 => x"8c0b8805",
  1062 => x"08558415",
  1063 => x"08fc0670",
  1064 => x"7a317a72",
  1065 => x"268f7225",
  1066 => x"07525553",
  1067 => x"7283e638",
  1068 => x"74798107",
  1069 => x"84170c79",
  1070 => x"167080d9",
  1071 => x"8c0b8805",
  1072 => x"0c758107",
  1073 => x"84120c54",
  1074 => x"7e525788",
  1075 => x"cd3f8817",
  1076 => x"54fae039",
  1077 => x"75832a70",
  1078 => x"54548074",
  1079 => x"24819b38",
  1080 => x"72822c81",
  1081 => x"712b80d9",
  1082 => x"90080770",
  1083 => x"80d98c0b",
  1084 => x"84050c75",
  1085 => x"10101080",
  1086 => x"d98c0588",
  1087 => x"1108585a",
  1088 => x"5d53778c",
  1089 => x"180c7488",
  1090 => x"180c7688",
  1091 => x"190c768c",
  1092 => x"160cfcf3",
  1093 => x"39797a10",
  1094 => x"101080d9",
  1095 => x"8c057057",
  1096 => x"595d8c15",
  1097 => x"08577675",
  1098 => x"2ea33884",
  1099 => x"1708fc06",
  1100 => x"707a3155",
  1101 => x"56738f24",
  1102 => x"83ca3873",
  1103 => x"80258481",
  1104 => x"388c1708",
  1105 => x"5776752e",
  1106 => x"098106df",
  1107 => x"38881581",
  1108 => x"1b708306",
  1109 => x"555b5572",
  1110 => x"c9387c83",
  1111 => x"06537280",
  1112 => x"2efdb838",
  1113 => x"ff1df819",
  1114 => x"595d8818",
  1115 => x"08782eea",
  1116 => x"38fdb539",
  1117 => x"831a53fc",
  1118 => x"96398314",
  1119 => x"70822c81",
  1120 => x"712b80d9",
  1121 => x"90080770",
  1122 => x"80d98c0b",
  1123 => x"84050c76",
  1124 => x"10101080",
  1125 => x"d98c0588",
  1126 => x"1108595b",
  1127 => x"5e5153fe",
  1128 => x"e13980d8",
  1129 => x"d0081758",
  1130 => x"8008762e",
  1131 => x"818d3880",
  1132 => x"d98008ff",
  1133 => x"2e83ec38",
  1134 => x"73763118",
  1135 => x"80d8d00c",
  1136 => x"73870670",
  1137 => x"57537280",
  1138 => x"2e883888",
  1139 => x"73317015",
  1140 => x"55567614",
  1141 => x"9fff06a0",
  1142 => x"80713117",
  1143 => x"70547f53",
  1144 => x"57538ebc",
  1145 => x"3f800853",
  1146 => x"8008ff2e",
  1147 => x"81a03880",
  1148 => x"d8d00816",
  1149 => x"7080d8d0",
  1150 => x"0c747580",
  1151 => x"d98c0b88",
  1152 => x"050c7476",
  1153 => x"31187081",
  1154 => x"07515556",
  1155 => x"587b80d9",
  1156 => x"8c2e839c",
  1157 => x"38798f26",
  1158 => x"82cb3881",
  1159 => x"0b84150c",
  1160 => x"841508fc",
  1161 => x"06707a31",
  1162 => x"7a72268f",
  1163 => x"72250752",
  1164 => x"55537280",
  1165 => x"2efcf938",
  1166 => x"80db3980",
  1167 => x"089fff06",
  1168 => x"5372feeb",
  1169 => x"387780d8",
  1170 => x"d00c80d9",
  1171 => x"8c0b8805",
  1172 => x"087b1881",
  1173 => x"0784120c",
  1174 => x"5580d8fc",
  1175 => x"08782786",
  1176 => x"387780d8",
  1177 => x"fc0c80d8",
  1178 => x"f8087827",
  1179 => x"fcac3877",
  1180 => x"80d8f80c",
  1181 => x"841508fc",
  1182 => x"06707a31",
  1183 => x"7a72268f",
  1184 => x"72250752",
  1185 => x"55537280",
  1186 => x"2efca538",
  1187 => x"88398074",
  1188 => x"5456fedb",
  1189 => x"397d5185",
  1190 => x"813f800b",
  1191 => x"800c8f3d",
  1192 => x"0d047353",
  1193 => x"807424a9",
  1194 => x"3872822c",
  1195 => x"81712b80",
  1196 => x"d9900807",
  1197 => x"7080d98c",
  1198 => x"0b84050c",
  1199 => x"5d53778c",
  1200 => x"180c7488",
  1201 => x"180c7688",
  1202 => x"190c768c",
  1203 => x"160cf9b7",
  1204 => x"39831470",
  1205 => x"822c8171",
  1206 => x"2b80d990",
  1207 => x"08077080",
  1208 => x"d98c0b84",
  1209 => x"050c5e51",
  1210 => x"53d4397b",
  1211 => x"7b065372",
  1212 => x"fca33884",
  1213 => x"1a7b105c",
  1214 => x"5af139ff",
  1215 => x"1a811151",
  1216 => x"5af7b939",
  1217 => x"78177981",
  1218 => x"0784190c",
  1219 => x"8c180888",
  1220 => x"1908718c",
  1221 => x"120c8812",
  1222 => x"0c597080",
  1223 => x"d9a00c70",
  1224 => x"80d99c0c",
  1225 => x"80d9940b",
  1226 => x"8c120c8c",
  1227 => x"11088812",
  1228 => x"0c748107",
  1229 => x"84120c74",
  1230 => x"1175710c",
  1231 => x"5153f9bd",
  1232 => x"39751784",
  1233 => x"11088107",
  1234 => x"84120c53",
  1235 => x"8c170888",
  1236 => x"1808718c",
  1237 => x"120c8812",
  1238 => x"0c587d51",
  1239 => x"83bc3f88",
  1240 => x"1754f5cf",
  1241 => x"39728415",
  1242 => x"0cf41af8",
  1243 => x"0670841e",
  1244 => x"08810607",
  1245 => x"841e0c70",
  1246 => x"1d545b85",
  1247 => x"0b84140c",
  1248 => x"850b8814",
  1249 => x"0c8f7b27",
  1250 => x"fdcf3888",
  1251 => x"1c527d51",
  1252 => x"93ee3f80",
  1253 => x"d98c0b88",
  1254 => x"050880d8",
  1255 => x"d0085955",
  1256 => x"fdb73977",
  1257 => x"80d8d00c",
  1258 => x"7380d980",
  1259 => x"0cfc9139",
  1260 => x"7284150c",
  1261 => x"fda339fa",
  1262 => x"3d0d7a79",
  1263 => x"028805a7",
  1264 => x"05335652",
  1265 => x"53837327",
  1266 => x"8a387083",
  1267 => x"06527180",
  1268 => x"2ea838ff",
  1269 => x"135372ff",
  1270 => x"2e973870",
  1271 => x"33527372",
  1272 => x"2e913881",
  1273 => x"11ff1454",
  1274 => x"5172ff2e",
  1275 => x"098106eb",
  1276 => x"38805170",
  1277 => x"800c883d",
  1278 => x"0d047072",
  1279 => x"57558351",
  1280 => x"75828029",
  1281 => x"14ff1252",
  1282 => x"56708025",
  1283 => x"f3388373",
  1284 => x"27bf3874",
  1285 => x"08763270",
  1286 => x"09f7fbfd",
  1287 => x"ff120670",
  1288 => x"f8848281",
  1289 => x"80065151",
  1290 => x"5170802e",
  1291 => x"99387451",
  1292 => x"80527033",
  1293 => x"5773772e",
  1294 => x"ffb93881",
  1295 => x"11811353",
  1296 => x"51837227",
  1297 => x"ed38fc13",
  1298 => x"84165653",
  1299 => x"728326c3",
  1300 => x"387451fe",
  1301 => x"fe39fa3d",
  1302 => x"0d787a7c",
  1303 => x"72727257",
  1304 => x"57575956",
  1305 => x"56747627",
  1306 => x"b2387615",
  1307 => x"51757127",
  1308 => x"aa387077",
  1309 => x"17ff1454",
  1310 => x"555371ff",
  1311 => x"2e9638ff",
  1312 => x"14ff1454",
  1313 => x"54723374",
  1314 => x"34ff1252",
  1315 => x"71ff2e09",
  1316 => x"8106ec38",
  1317 => x"75800c88",
  1318 => x"3d0d0476",
  1319 => x"8f269738",
  1320 => x"ff125271",
  1321 => x"ff2eed38",
  1322 => x"72708105",
  1323 => x"54337470",
  1324 => x"81055634",
  1325 => x"eb397476",
  1326 => x"07830651",
  1327 => x"70e23875",
  1328 => x"75545172",
  1329 => x"70840554",
  1330 => x"08717084",
  1331 => x"05530c72",
  1332 => x"70840554",
  1333 => x"08717084",
  1334 => x"05530c72",
  1335 => x"70840554",
  1336 => x"08717084",
  1337 => x"05530c72",
  1338 => x"70840554",
  1339 => x"08717084",
  1340 => x"05530cf0",
  1341 => x"1252718f",
  1342 => x"26c93883",
  1343 => x"72279538",
  1344 => x"72708405",
  1345 => x"54087170",
  1346 => x"8405530c",
  1347 => x"fc125271",
  1348 => x"8326ed38",
  1349 => x"7054ff88",
  1350 => x"390404ef",
  1351 => x"3d0d6365",
  1352 => x"67405d42",
  1353 => x"7b802e84",
  1354 => x"f9386151",
  1355 => x"ec3ff81c",
  1356 => x"70841208",
  1357 => x"70fc0670",
  1358 => x"628b0570",
  1359 => x"f8064159",
  1360 => x"455b5c41",
  1361 => x"57967427",
  1362 => x"82c33880",
  1363 => x"7b247e7c",
  1364 => x"26075980",
  1365 => x"5478742e",
  1366 => x"09810682",
  1367 => x"a938777b",
  1368 => x"2581fc38",
  1369 => x"771780d9",
  1370 => x"8c0b8805",
  1371 => x"085e567c",
  1372 => x"762e84bd",
  1373 => x"38841608",
  1374 => x"70fe0617",
  1375 => x"84110881",
  1376 => x"06515555",
  1377 => x"73828b38",
  1378 => x"74fc0659",
  1379 => x"7c762e84",
  1380 => x"dd387719",
  1381 => x"5f7e7b25",
  1382 => x"81fd3879",
  1383 => x"81065473",
  1384 => x"82bf3876",
  1385 => x"77083184",
  1386 => x"1108fc06",
  1387 => x"565a7580",
  1388 => x"2e91387c",
  1389 => x"762e84ea",
  1390 => x"38741918",
  1391 => x"59787b25",
  1392 => x"84893879",
  1393 => x"802e8299",
  1394 => x"38771556",
  1395 => x"7a762482",
  1396 => x"90388c1a",
  1397 => x"08881b08",
  1398 => x"718c120c",
  1399 => x"88120c55",
  1400 => x"79765957",
  1401 => x"881761fc",
  1402 => x"05575975",
  1403 => x"a42685ef",
  1404 => x"387b7955",
  1405 => x"55937627",
  1406 => x"80c9387b",
  1407 => x"7084055d",
  1408 => x"087c5679",
  1409 => x"0c747084",
  1410 => x"0556088c",
  1411 => x"180c9017",
  1412 => x"549b7627",
  1413 => x"ae387470",
  1414 => x"84055608",
  1415 => x"740c7470",
  1416 => x"84055608",
  1417 => x"94180c98",
  1418 => x"1754a376",
  1419 => x"27953874",
  1420 => x"70840556",
  1421 => x"08740c74",
  1422 => x"70840556",
  1423 => x"089c180c",
  1424 => x"a0175474",
  1425 => x"70840556",
  1426 => x"08747084",
  1427 => x"05560c74",
  1428 => x"70840556",
  1429 => x"08747084",
  1430 => x"05560c74",
  1431 => x"08740c77",
  1432 => x"7b315675",
  1433 => x"8f2680c9",
  1434 => x"38841708",
  1435 => x"81067807",
  1436 => x"84180c77",
  1437 => x"17841108",
  1438 => x"81078412",
  1439 => x"0c546151",
  1440 => x"fd983f88",
  1441 => x"17547380",
  1442 => x"0c933d0d",
  1443 => x"04905bfd",
  1444 => x"ba397856",
  1445 => x"fe85398c",
  1446 => x"16088817",
  1447 => x"08718c12",
  1448 => x"0c88120c",
  1449 => x"557e707c",
  1450 => x"3157588f",
  1451 => x"7627ffb9",
  1452 => x"387a1784",
  1453 => x"18088106",
  1454 => x"7c078419",
  1455 => x"0c768107",
  1456 => x"84120c76",
  1457 => x"11841108",
  1458 => x"81078412",
  1459 => x"0c558805",
  1460 => x"5261518d",
  1461 => x"ab3f6151",
  1462 => x"fcc03f88",
  1463 => x"1754ffa6",
  1464 => x"397d5261",
  1465 => x"51edda3f",
  1466 => x"80085980",
  1467 => x"08802e81",
  1468 => x"a3388008",
  1469 => x"f8056084",
  1470 => x"0508fe06",
  1471 => x"61055557",
  1472 => x"76742e83",
  1473 => x"e638fc18",
  1474 => x"5675a426",
  1475 => x"81aa387b",
  1476 => x"80085555",
  1477 => x"93762780",
  1478 => x"d8387470",
  1479 => x"84055608",
  1480 => x"80087084",
  1481 => x"05800c0c",
  1482 => x"80087570",
  1483 => x"84055708",
  1484 => x"71708405",
  1485 => x"530c549b",
  1486 => x"7627b638",
  1487 => x"74708405",
  1488 => x"56087470",
  1489 => x"8405560c",
  1490 => x"74708405",
  1491 => x"56087470",
  1492 => x"8405560c",
  1493 => x"a3762799",
  1494 => x"38747084",
  1495 => x"05560874",
  1496 => x"70840556",
  1497 => x"0c747084",
  1498 => x"05560874",
  1499 => x"70840556",
  1500 => x"0c747084",
  1501 => x"05560874",
  1502 => x"70840556",
  1503 => x"0c747084",
  1504 => x"05560874",
  1505 => x"70840556",
  1506 => x"0c740874",
  1507 => x"0c7b5261",
  1508 => x"518bed3f",
  1509 => x"6151fb82",
  1510 => x"3f785473",
  1511 => x"800c933d",
  1512 => x"0d047d52",
  1513 => x"6151ec99",
  1514 => x"3f800880",
  1515 => x"0c933d0d",
  1516 => x"04841608",
  1517 => x"55fbd139",
  1518 => x"75537b52",
  1519 => x"800851df",
  1520 => x"db3f7b52",
  1521 => x"61518bb8",
  1522 => x"3fca398c",
  1523 => x"16088817",
  1524 => x"08718c12",
  1525 => x"0c88120c",
  1526 => x"558c1a08",
  1527 => x"881b0871",
  1528 => x"8c120c88",
  1529 => x"120c5579",
  1530 => x"795957fb",
  1531 => x"f7397719",
  1532 => x"901c5555",
  1533 => x"737524fb",
  1534 => x"a2387a17",
  1535 => x"7080d98c",
  1536 => x"0b88050c",
  1537 => x"757c3181",
  1538 => x"0784120c",
  1539 => x"5d841708",
  1540 => x"81067b07",
  1541 => x"84180c61",
  1542 => x"51f9ff3f",
  1543 => x"881754fc",
  1544 => x"e5397419",
  1545 => x"18901c55",
  1546 => x"5d737d24",
  1547 => x"fb95388c",
  1548 => x"1a08881b",
  1549 => x"08718c12",
  1550 => x"0c88120c",
  1551 => x"55881a61",
  1552 => x"fc055759",
  1553 => x"75a42681",
  1554 => x"ae387b79",
  1555 => x"55559376",
  1556 => x"2780c938",
  1557 => x"7b708405",
  1558 => x"5d087c56",
  1559 => x"790c7470",
  1560 => x"84055608",
  1561 => x"8c1b0c90",
  1562 => x"1a549b76",
  1563 => x"27ae3874",
  1564 => x"70840556",
  1565 => x"08740c74",
  1566 => x"70840556",
  1567 => x"08941b0c",
  1568 => x"981a54a3",
  1569 => x"76279538",
  1570 => x"74708405",
  1571 => x"5608740c",
  1572 => x"74708405",
  1573 => x"56089c1b",
  1574 => x"0ca01a54",
  1575 => x"74708405",
  1576 => x"56087470",
  1577 => x"8405560c",
  1578 => x"74708405",
  1579 => x"56087470",
  1580 => x"8405560c",
  1581 => x"7408740c",
  1582 => x"7a1a7080",
  1583 => x"d98c0b88",
  1584 => x"050c7d7c",
  1585 => x"31810784",
  1586 => x"120c5484",
  1587 => x"1a088106",
  1588 => x"7b07841b",
  1589 => x"0c6151f8",
  1590 => x"c13f7854",
  1591 => x"fdbd3975",
  1592 => x"537b5278",
  1593 => x"51ddb53f",
  1594 => x"faf53984",
  1595 => x"1708fc06",
  1596 => x"18605858",
  1597 => x"fae93975",
  1598 => x"537b5278",
  1599 => x"51dd9d3f",
  1600 => x"7a1a7080",
  1601 => x"d98c0b88",
  1602 => x"050c7d7c",
  1603 => x"31810784",
  1604 => x"120c5484",
  1605 => x"1a088106",
  1606 => x"7b07841b",
  1607 => x"0cffb639",
  1608 => x"fd3d0d80",
  1609 => x"0b80e1c4",
  1610 => x"0c765196",
  1611 => x"d53f8008",
  1612 => x"538008ff",
  1613 => x"2e883872",
  1614 => x"800c853d",
  1615 => x"0d0480e1",
  1616 => x"c4085473",
  1617 => x"802ef038",
  1618 => x"7574710c",
  1619 => x"5272800c",
  1620 => x"853d0d04",
  1621 => x"fa3d0d78",
  1622 => x"80d1d008",
  1623 => x"5455b813",
  1624 => x"08802e81",
  1625 => x"b6388c15",
  1626 => x"227083ff",
  1627 => x"ff067083",
  1628 => x"2a813270",
  1629 => x"81065155",
  1630 => x"55567280",
  1631 => x"2e80dc38",
  1632 => x"73842a81",
  1633 => x"32810657",
  1634 => x"ff537680",
  1635 => x"f7387382",
  1636 => x"2a708106",
  1637 => x"51537280",
  1638 => x"2eb938b0",
  1639 => x"15085473",
  1640 => x"802e9c38",
  1641 => x"80c01553",
  1642 => x"73732e8f",
  1643 => x"38735280",
  1644 => x"d1d00851",
  1645 => x"87ca3f8c",
  1646 => x"15225676",
  1647 => x"b0160c75",
  1648 => x"db065372",
  1649 => x"8c162380",
  1650 => x"0b84160c",
  1651 => x"90150875",
  1652 => x"0c725675",
  1653 => x"88075372",
  1654 => x"8c162390",
  1655 => x"1508802e",
  1656 => x"80c1388c",
  1657 => x"15227081",
  1658 => x"06555373",
  1659 => x"9e38720a",
  1660 => x"100a7081",
  1661 => x"06515372",
  1662 => x"85389415",
  1663 => x"08547388",
  1664 => x"160c8053",
  1665 => x"72800c88",
  1666 => x"3d0d0480",
  1667 => x"0b88160c",
  1668 => x"94150830",
  1669 => x"98160c80",
  1670 => x"53ea3972",
  1671 => x"5182fb3f",
  1672 => x"fec43974",
  1673 => x"518ce83f",
  1674 => x"8c152270",
  1675 => x"81065553",
  1676 => x"73802eff",
  1677 => x"b938d439",
  1678 => x"f83d0d7a",
  1679 => x"5877802e",
  1680 => x"81993880",
  1681 => x"d1d00854",
  1682 => x"b8140880",
  1683 => x"2e80ed38",
  1684 => x"8c182270",
  1685 => x"902b7090",
  1686 => x"2c70832a",
  1687 => x"81328106",
  1688 => x"5c515754",
  1689 => x"7880cd38",
  1690 => x"90180857",
  1691 => x"76802e80",
  1692 => x"c3387708",
  1693 => x"77317779",
  1694 => x"0c768306",
  1695 => x"7a585555",
  1696 => x"73853894",
  1697 => x"18085675",
  1698 => x"88190c80",
  1699 => x"7525a538",
  1700 => x"74537652",
  1701 => x"9c180851",
  1702 => x"a4180854",
  1703 => x"732d800b",
  1704 => x"80082580",
  1705 => x"c9388008",
  1706 => x"17758008",
  1707 => x"31565774",
  1708 => x"8024dd38",
  1709 => x"800b800c",
  1710 => x"8a3d0d04",
  1711 => x"735181da",
  1712 => x"3f8c1822",
  1713 => x"70902b70",
  1714 => x"902c7083",
  1715 => x"2a813281",
  1716 => x"065c5157",
  1717 => x"5478dd38",
  1718 => x"ff8e39b4",
  1719 => x"b85280d1",
  1720 => x"d0085189",
  1721 => x"f13f8008",
  1722 => x"800c8a3d",
  1723 => x"0d048c18",
  1724 => x"2280c007",
  1725 => x"54738c19",
  1726 => x"23ff0b80",
  1727 => x"0c8a3d0d",
  1728 => x"04803d0d",
  1729 => x"72518071",
  1730 => x"0c800b84",
  1731 => x"120c800b",
  1732 => x"88120c02",
  1733 => x"8e05228c",
  1734 => x"12230292",
  1735 => x"05228e12",
  1736 => x"23800b90",
  1737 => x"120c800b",
  1738 => x"94120c80",
  1739 => x"0b98120c",
  1740 => x"709c120c",
  1741 => x"80c4a10b",
  1742 => x"a0120c80",
  1743 => x"c4ed0ba4",
  1744 => x"120c80c5",
  1745 => x"e90ba812",
  1746 => x"0c80c6ba",
  1747 => x"0bac120c",
  1748 => x"823d0d04",
  1749 => x"fa3d0d79",
  1750 => x"7080dc29",
  1751 => x"8c11547a",
  1752 => x"535657e4",
  1753 => x"dc3f8008",
  1754 => x"80085556",
  1755 => x"8008802e",
  1756 => x"a2388008",
  1757 => x"8c055480",
  1758 => x"0b80080c",
  1759 => x"76800884",
  1760 => x"050c7380",
  1761 => x"0888050c",
  1762 => x"74538052",
  1763 => x"73518c82",
  1764 => x"3f755473",
  1765 => x"800c883d",
  1766 => x"0d04fc3d",
  1767 => x"0d76b9ad",
  1768 => x"0bbc120c",
  1769 => x"55810bb8",
  1770 => x"160c800b",
  1771 => x"84dc160c",
  1772 => x"830b84e0",
  1773 => x"160c84e8",
  1774 => x"1584e416",
  1775 => x"0c745480",
  1776 => x"53845284",
  1777 => x"150851fe",
  1778 => x"b83f7454",
  1779 => x"81538952",
  1780 => x"88150851",
  1781 => x"feab3f74",
  1782 => x"5482538a",
  1783 => x"528c1508",
  1784 => x"51fe9e3f",
  1785 => x"863d0d04",
  1786 => x"f93d0d79",
  1787 => x"80d1d008",
  1788 => x"5457b813",
  1789 => x"08802e80",
  1790 => x"c83884dc",
  1791 => x"13568816",
  1792 => x"08841708",
  1793 => x"ff055555",
  1794 => x"8074249f",
  1795 => x"388c1522",
  1796 => x"70902b70",
  1797 => x"902c5154",
  1798 => x"5872802e",
  1799 => x"80ca3880",
  1800 => x"dc15ff15",
  1801 => x"55557380",
  1802 => x"25e33875",
  1803 => x"08537280",
  1804 => x"2e9f3872",
  1805 => x"56881608",
  1806 => x"841708ff",
  1807 => x"055555c8",
  1808 => x"397251fe",
  1809 => x"d53f80d1",
  1810 => x"d00884dc",
  1811 => x"0556ffae",
  1812 => x"39845276",
  1813 => x"51fdfd3f",
  1814 => x"8008760c",
  1815 => x"8008802e",
  1816 => x"80c03880",
  1817 => x"0856ce39",
  1818 => x"810b8c16",
  1819 => x"2372750c",
  1820 => x"7288160c",
  1821 => x"7284160c",
  1822 => x"7290160c",
  1823 => x"7294160c",
  1824 => x"7298160c",
  1825 => x"ff0b8e16",
  1826 => x"2372b016",
  1827 => x"0c72b416",
  1828 => x"0c7280c4",
  1829 => x"160c7280",
  1830 => x"c8160c74",
  1831 => x"800c893d",
  1832 => x"0d048c77",
  1833 => x"0c800b80",
  1834 => x"0c893d0d",
  1835 => x"04ff3d0d",
  1836 => x"b4b85273",
  1837 => x"51869f3f",
  1838 => x"833d0d04",
  1839 => x"803d0d80",
  1840 => x"d1d00851",
  1841 => x"e83f823d",
  1842 => x"0d04fb3d",
  1843 => x"0d777052",
  1844 => x"56f0c63f",
  1845 => x"80d98c0b",
  1846 => x"88050884",
  1847 => x"1108fc06",
  1848 => x"707b319f",
  1849 => x"ef05e080",
  1850 => x"06e08005",
  1851 => x"565653a0",
  1852 => x"80742494",
  1853 => x"38805275",
  1854 => x"51f8a53f",
  1855 => x"80d99408",
  1856 => x"15537280",
  1857 => x"082e8f38",
  1858 => x"7551f08e",
  1859 => x"3f805372",
  1860 => x"800c873d",
  1861 => x"0d047330",
  1862 => x"527551f8",
  1863 => x"833f8008",
  1864 => x"ff2ea838",
  1865 => x"80d98c0b",
  1866 => x"88050875",
  1867 => x"75318107",
  1868 => x"84120c53",
  1869 => x"80d8d008",
  1870 => x"743180d8",
  1871 => x"d00c7551",
  1872 => x"efd83f81",
  1873 => x"0b800c87",
  1874 => x"3d0d0480",
  1875 => x"527551f7",
  1876 => x"cf3f80d9",
  1877 => x"8c0b8805",
  1878 => x"08800871",
  1879 => x"3156538f",
  1880 => x"7525ffa4",
  1881 => x"38800880",
  1882 => x"d9800831",
  1883 => x"80d8d00c",
  1884 => x"74810784",
  1885 => x"140c7551",
  1886 => x"efa03f80",
  1887 => x"53ff9039",
  1888 => x"f63d0d7c",
  1889 => x"7e545b72",
  1890 => x"802e8283",
  1891 => x"387a51ef",
  1892 => x"883ff813",
  1893 => x"84110870",
  1894 => x"fe067013",
  1895 => x"841108fc",
  1896 => x"065d5859",
  1897 => x"545880d9",
  1898 => x"9408752e",
  1899 => x"82de3878",
  1900 => x"84160c80",
  1901 => x"73810654",
  1902 => x"5a727a2e",
  1903 => x"81d53878",
  1904 => x"15841108",
  1905 => x"81065153",
  1906 => x"72a03878",
  1907 => x"17577981",
  1908 => x"e6388815",
  1909 => x"08537280",
  1910 => x"d9942e82",
  1911 => x"f9388c15",
  1912 => x"08708c15",
  1913 => x"0c738812",
  1914 => x"0c567681",
  1915 => x"0784190c",
  1916 => x"76187771",
  1917 => x"0c537981",
  1918 => x"913883ff",
  1919 => x"772781c8",
  1920 => x"3876892a",
  1921 => x"77832a56",
  1922 => x"5372802e",
  1923 => x"bf387686",
  1924 => x"2ab80555",
  1925 => x"847327b4",
  1926 => x"3880db13",
  1927 => x"55947327",
  1928 => x"ab38768c",
  1929 => x"2a80ee05",
  1930 => x"5580d473",
  1931 => x"279e3876",
  1932 => x"8f2a80f7",
  1933 => x"055582d4",
  1934 => x"73279138",
  1935 => x"76922a80",
  1936 => x"fc05558a",
  1937 => x"d4732784",
  1938 => x"3880fe55",
  1939 => x"74101010",
  1940 => x"80d98c05",
  1941 => x"88110855",
  1942 => x"5673762e",
  1943 => x"82b33884",
  1944 => x"1408fc06",
  1945 => x"53767327",
  1946 => x"8d388814",
  1947 => x"08547376",
  1948 => x"2e098106",
  1949 => x"ea388c14",
  1950 => x"08708c1a",
  1951 => x"0c74881a",
  1952 => x"0c788812",
  1953 => x"0c56778c",
  1954 => x"150c7a51",
  1955 => x"ed8c3f8c",
  1956 => x"3d0d0477",
  1957 => x"08787131",
  1958 => x"59770588",
  1959 => x"19085457",
  1960 => x"7280d994",
  1961 => x"2e80e038",
  1962 => x"8c180870",
  1963 => x"8c150c73",
  1964 => x"88120c56",
  1965 => x"fe893988",
  1966 => x"15088c16",
  1967 => x"08708c13",
  1968 => x"0c578817",
  1969 => x"0cfea339",
  1970 => x"76832a70",
  1971 => x"54558075",
  1972 => x"24819838",
  1973 => x"72822c81",
  1974 => x"712b80d9",
  1975 => x"90080780",
  1976 => x"d98c0b84",
  1977 => x"050c5374",
  1978 => x"10101080",
  1979 => x"d98c0588",
  1980 => x"11085556",
  1981 => x"758c190c",
  1982 => x"7388190c",
  1983 => x"7788170c",
  1984 => x"778c150c",
  1985 => x"ff843981",
  1986 => x"5afdb439",
  1987 => x"78177381",
  1988 => x"06545772",
  1989 => x"98387708",
  1990 => x"78713159",
  1991 => x"77058c19",
  1992 => x"08881a08",
  1993 => x"718c120c",
  1994 => x"88120c57",
  1995 => x"57768107",
  1996 => x"84190c77",
  1997 => x"80d98c0b",
  1998 => x"88050c80",
  1999 => x"d9880877",
  2000 => x"26fec738",
  2001 => x"80d98408",
  2002 => x"527a51fa",
  2003 => x"fd3f7a51",
  2004 => x"ebc83ffe",
  2005 => x"ba398178",
  2006 => x"8c150c78",
  2007 => x"88150c73",
  2008 => x"8c1a0c73",
  2009 => x"881a0c5a",
  2010 => x"fd803983",
  2011 => x"1570822c",
  2012 => x"81712b80",
  2013 => x"d9900807",
  2014 => x"80d98c0b",
  2015 => x"84050c51",
  2016 => x"53741010",
  2017 => x"1080d98c",
  2018 => x"05881108",
  2019 => x"5556fee4",
  2020 => x"39745380",
  2021 => x"7524a738",
  2022 => x"72822c81",
  2023 => x"712b80d9",
  2024 => x"90080780",
  2025 => x"d98c0b84",
  2026 => x"050c5375",
  2027 => x"8c190c73",
  2028 => x"88190c77",
  2029 => x"88170c77",
  2030 => x"8c150cfd",
  2031 => x"cd398315",
  2032 => x"70822c81",
  2033 => x"712b80d9",
  2034 => x"90080780",
  2035 => x"d98c0b84",
  2036 => x"050c5153",
  2037 => x"d639f93d",
  2038 => x"0d797b58",
  2039 => x"53800b80",
  2040 => x"d1d00853",
  2041 => x"5672722e",
  2042 => x"80c03884",
  2043 => x"dc135574",
  2044 => x"762eb738",
  2045 => x"88150884",
  2046 => x"1608ff05",
  2047 => x"54548073",
  2048 => x"249d388c",
  2049 => x"14227090",
  2050 => x"2b70902c",
  2051 => x"51535871",
  2052 => x"80d83880",
  2053 => x"dc14ff14",
  2054 => x"54547280",
  2055 => x"25e53874",
  2056 => x"085574d0",
  2057 => x"3880d1d0",
  2058 => x"085284dc",
  2059 => x"12557480",
  2060 => x"2eb13888",
  2061 => x"15088416",
  2062 => x"08ff0554",
  2063 => x"54807324",
  2064 => x"9c388c14",
  2065 => x"2270902b",
  2066 => x"70902c51",
  2067 => x"535871ad",
  2068 => x"3880dc14",
  2069 => x"ff145454",
  2070 => x"728025e6",
  2071 => x"38740855",
  2072 => x"74d13875",
  2073 => x"800c893d",
  2074 => x"0d047351",
  2075 => x"762d7580",
  2076 => x"080780dc",
  2077 => x"15ff1555",
  2078 => x"5556ff9e",
  2079 => x"39735176",
  2080 => x"2d758008",
  2081 => x"0780dc15",
  2082 => x"ff155555",
  2083 => x"56ca39ea",
  2084 => x"3d0d688c",
  2085 => x"1122700a",
  2086 => x"100a8106",
  2087 => x"57585674",
  2088 => x"80e4388e",
  2089 => x"16227090",
  2090 => x"2b70902c",
  2091 => x"51555880",
  2092 => x"7424b138",
  2093 => x"983dc405",
  2094 => x"53735280",
  2095 => x"d1d00851",
  2096 => x"86803f80",
  2097 => x"0b800824",
  2098 => x"97387983",
  2099 => x"e0800654",
  2100 => x"7380c080",
  2101 => x"2e818f38",
  2102 => x"73828080",
  2103 => x"2e819138",
  2104 => x"8c162257",
  2105 => x"76908007",
  2106 => x"54738c17",
  2107 => x"23888052",
  2108 => x"80d1d008",
  2109 => x"51d9ca3f",
  2110 => x"80089d38",
  2111 => x"8c162282",
  2112 => x"0754738c",
  2113 => x"172380c3",
  2114 => x"1670770c",
  2115 => x"90170c81",
  2116 => x"0b94170c",
  2117 => x"983d0d04",
  2118 => x"80d1d008",
  2119 => x"b9ad0bbc",
  2120 => x"120c548c",
  2121 => x"16228180",
  2122 => x"0754738c",
  2123 => x"17238008",
  2124 => x"760c8008",
  2125 => x"90170c88",
  2126 => x"800b9417",
  2127 => x"0c74802e",
  2128 => x"d3388e16",
  2129 => x"2270902b",
  2130 => x"70902c53",
  2131 => x"55588ca1",
  2132 => x"3f800880",
  2133 => x"2effbd38",
  2134 => x"8c162281",
  2135 => x"0754738c",
  2136 => x"1723983d",
  2137 => x"0d04810b",
  2138 => x"8c172258",
  2139 => x"55fef539",
  2140 => x"a8160880",
  2141 => x"c5e92e09",
  2142 => x"8106fee4",
  2143 => x"388c1622",
  2144 => x"88800754",
  2145 => x"738c1723",
  2146 => x"88800b80",
  2147 => x"cc170cfe",
  2148 => x"dc39fc3d",
  2149 => x"0d767971",
  2150 => x"028c059f",
  2151 => x"05335755",
  2152 => x"53558372",
  2153 => x"278a3874",
  2154 => x"83065170",
  2155 => x"802ea238",
  2156 => x"ff125271",
  2157 => x"ff2e9338",
  2158 => x"73737081",
  2159 => x"055534ff",
  2160 => x"125271ff",
  2161 => x"2e098106",
  2162 => x"ef387480",
  2163 => x"0c863d0d",
  2164 => x"04747488",
  2165 => x"2b750770",
  2166 => x"71902b07",
  2167 => x"5154518f",
  2168 => x"7227a538",
  2169 => x"72717084",
  2170 => x"05530c72",
  2171 => x"71708405",
  2172 => x"530c7271",
  2173 => x"70840553",
  2174 => x"0c727170",
  2175 => x"8405530c",
  2176 => x"f0125271",
  2177 => x"8f26dd38",
  2178 => x"83722790",
  2179 => x"38727170",
  2180 => x"8405530c",
  2181 => x"fc125271",
  2182 => x"8326f238",
  2183 => x"7053ff90",
  2184 => x"39f93d0d",
  2185 => x"797c557b",
  2186 => x"548e1122",
  2187 => x"70902b70",
  2188 => x"902c5557",
  2189 => x"80d1d008",
  2190 => x"53585683",
  2191 => x"f33f8008",
  2192 => x"57800b80",
  2193 => x"08249338",
  2194 => x"80d01608",
  2195 => x"80080580",
  2196 => x"d0170c76",
  2197 => x"800c893d",
  2198 => x"0d048c16",
  2199 => x"2283dfff",
  2200 => x"0655748c",
  2201 => x"17237680",
  2202 => x"0c893d0d",
  2203 => x"04fa3d0d",
  2204 => x"788c1122",
  2205 => x"70882a70",
  2206 => x"81065157",
  2207 => x"585674a9",
  2208 => x"388c1622",
  2209 => x"83dfff06",
  2210 => x"55748c17",
  2211 => x"237a5479",
  2212 => x"538e1622",
  2213 => x"70902b70",
  2214 => x"902c5456",
  2215 => x"80d1d008",
  2216 => x"525681b2",
  2217 => x"3f883d0d",
  2218 => x"04825480",
  2219 => x"538e1622",
  2220 => x"70902b70",
  2221 => x"902c5456",
  2222 => x"80d1d008",
  2223 => x"525782b8",
  2224 => x"3f8c1622",
  2225 => x"83dfff06",
  2226 => x"55748c17",
  2227 => x"237a5479",
  2228 => x"538e1622",
  2229 => x"70902b70",
  2230 => x"902c5456",
  2231 => x"80d1d008",
  2232 => x"525680f2",
  2233 => x"3f883d0d",
  2234 => x"04f93d0d",
  2235 => x"797c557b",
  2236 => x"548e1122",
  2237 => x"70902b70",
  2238 => x"902c5557",
  2239 => x"80d1d008",
  2240 => x"53585681",
  2241 => x"f33f8008",
  2242 => x"578008ff",
  2243 => x"2e99388c",
  2244 => x"1622a080",
  2245 => x"0755748c",
  2246 => x"17238008",
  2247 => x"80d0170c",
  2248 => x"76800c89",
  2249 => x"3d0d048c",
  2250 => x"162283df",
  2251 => x"ff065574",
  2252 => x"8c172376",
  2253 => x"800c893d",
  2254 => x"0d04fe3d",
  2255 => x"0d748e11",
  2256 => x"2270902b",
  2257 => x"70902c55",
  2258 => x"51515380",
  2259 => x"d1d00851",
  2260 => x"bd3f843d",
  2261 => x"0d04fb3d",
  2262 => x"0d800b80",
  2263 => x"e1c40c7a",
  2264 => x"53795278",
  2265 => x"51839a3f",
  2266 => x"80085580",
  2267 => x"08ff2e88",
  2268 => x"3874800c",
  2269 => x"873d0d04",
  2270 => x"80e1c408",
  2271 => x"5675802e",
  2272 => x"f0387776",
  2273 => x"710c5474",
  2274 => x"800c873d",
  2275 => x"0d04fd3d",
  2276 => x"0d800b80",
  2277 => x"e1c40c76",
  2278 => x"5184ef3f",
  2279 => x"80085380",
  2280 => x"08ff2e88",
  2281 => x"3872800c",
  2282 => x"853d0d04",
  2283 => x"80e1c408",
  2284 => x"5473802e",
  2285 => x"f0387574",
  2286 => x"710c5272",
  2287 => x"800c853d",
  2288 => x"0d04fc3d",
  2289 => x"0d800b80",
  2290 => x"e1c40c78",
  2291 => x"52775186",
  2292 => x"d73f8008",
  2293 => x"548008ff",
  2294 => x"2e883873",
  2295 => x"800c863d",
  2296 => x"0d0480e1",
  2297 => x"c4085574",
  2298 => x"802ef038",
  2299 => x"7675710c",
  2300 => x"5373800c",
  2301 => x"863d0d04",
  2302 => x"fb3d0d80",
  2303 => x"0b80e1c4",
  2304 => x"0c7a5379",
  2305 => x"52785184",
  2306 => x"b33f8008",
  2307 => x"558008ff",
  2308 => x"2e883874",
  2309 => x"800c873d",
  2310 => x"0d0480e1",
  2311 => x"c4085675",
  2312 => x"802ef038",
  2313 => x"7776710c",
  2314 => x"5474800c",
  2315 => x"873d0d04",
  2316 => x"fb3d0d80",
  2317 => x"0b80e1c4",
  2318 => x"0c7a5379",
  2319 => x"52785182",
  2320 => x"b83f8008",
  2321 => x"558008ff",
  2322 => x"2e883874",
  2323 => x"800c873d",
  2324 => x"0d0480e1",
  2325 => x"c4085675",
  2326 => x"802ef038",
  2327 => x"7776710c",
  2328 => x"5474800c",
  2329 => x"873d0d04",
  2330 => x"810b800c",
  2331 => x"04803d0d",
  2332 => x"72812e89",
  2333 => x"38800b80",
  2334 => x"0c823d0d",
  2335 => x"04735180",
  2336 => x"fa3ffe3d",
  2337 => x"0d80e1bc",
  2338 => x"0851708a",
  2339 => x"3880e1c8",
  2340 => x"7080e1bc",
  2341 => x"0c517075",
  2342 => x"125252ff",
  2343 => x"537087fb",
  2344 => x"80802688",
  2345 => x"387080e1",
  2346 => x"bc0c7153",
  2347 => x"72800c84",
  2348 => x"3d0d04fd",
  2349 => x"3d0d800b",
  2350 => x"80d1c408",
  2351 => x"54547281",
  2352 => x"2e9d3873",
  2353 => x"80e1c00c",
  2354 => x"ffbfdb3f",
  2355 => x"ffbeb13f",
  2356 => x"80e19452",
  2357 => x"8151c1a0",
  2358 => x"3f800851",
  2359 => x"85ca3f72",
  2360 => x"80e1c00c",
  2361 => x"ffbfbf3f",
  2362 => x"ffbe953f",
  2363 => x"80e19452",
  2364 => x"8151c184",
  2365 => x"3f800851",
  2366 => x"85ae3f00",
  2367 => x"ff3900ff",
  2368 => x"39f53d0d",
  2369 => x"7e6080e1",
  2370 => x"c008705b",
  2371 => x"585b5b75",
  2372 => x"80c53877",
  2373 => x"7a25a238",
  2374 => x"771b7033",
  2375 => x"7081ff06",
  2376 => x"58585975",
  2377 => x"8a2e9938",
  2378 => x"7681ff06",
  2379 => x"51ffbed5",
  2380 => x"3f811858",
  2381 => x"797824e0",
  2382 => x"3879800c",
  2383 => x"8d3d0d04",
  2384 => x"8d51ffbe",
  2385 => x"c03f7833",
  2386 => x"7081ff06",
  2387 => x"5257ffbe",
  2388 => x"b43f8118",
  2389 => x"58de3979",
  2390 => x"557a547d",
  2391 => x"5385528d",
  2392 => x"3dfc0551",
  2393 => x"ffbddb3f",
  2394 => x"80085684",
  2395 => x"b43f7b80",
  2396 => x"080c7580",
  2397 => x"0c8d3d0d",
  2398 => x"04f63d0d",
  2399 => x"7d7f80e1",
  2400 => x"c008705b",
  2401 => x"585a5a75",
  2402 => x"80c43877",
  2403 => x"7925b638",
  2404 => x"ffbdcd3f",
  2405 => x"800881ff",
  2406 => x"06708d32",
  2407 => x"7030709f",
  2408 => x"2a515157",
  2409 => x"57768a2e",
  2410 => x"80c63875",
  2411 => x"802e80c0",
  2412 => x"38771a56",
  2413 => x"76763476",
  2414 => x"51ffbdc9",
  2415 => x"3f811858",
  2416 => x"787824cc",
  2417 => x"38775675",
  2418 => x"800c8c3d",
  2419 => x"0d047855",
  2420 => x"79547c53",
  2421 => x"84528c3d",
  2422 => x"fc0551ff",
  2423 => x"bce43f80",
  2424 => x"085683bd",
  2425 => x"3f7a8008",
  2426 => x"0c75800c",
  2427 => x"8c3d0d04",
  2428 => x"771a568a",
  2429 => x"76348118",
  2430 => x"588d51ff",
  2431 => x"bd873f8a",
  2432 => x"51ffbd81",
  2433 => x"3f7756ff",
  2434 => x"be39fb3d",
  2435 => x"0d80e1c0",
  2436 => x"08705654",
  2437 => x"73883874",
  2438 => x"800c873d",
  2439 => x"0d047753",
  2440 => x"8352873d",
  2441 => x"fc0551ff",
  2442 => x"bc983f80",
  2443 => x"085482f1",
  2444 => x"3f758008",
  2445 => x"0c73800c",
  2446 => x"873d0d04",
  2447 => x"fa3d0d80",
  2448 => x"e1c00880",
  2449 => x"2ea3387a",
  2450 => x"55795478",
  2451 => x"53865288",
  2452 => x"3dfc0551",
  2453 => x"ffbbeb3f",
  2454 => x"80085682",
  2455 => x"c43f7680",
  2456 => x"080c7580",
  2457 => x"0c883d0d",
  2458 => x"0482b63f",
  2459 => x"9d0b8008",
  2460 => x"0cff0b80",
  2461 => x"0c883d0d",
  2462 => x"04fb3d0d",
  2463 => x"77795656",
  2464 => x"80705454",
  2465 => x"7375259f",
  2466 => x"38741010",
  2467 => x"10f80552",
  2468 => x"72167033",
  2469 => x"70742b76",
  2470 => x"078116f8",
  2471 => x"16565656",
  2472 => x"51517473",
  2473 => x"24ea3873",
  2474 => x"800c873d",
  2475 => x"0d04fc3d",
  2476 => x"0d767855",
  2477 => x"55bc5380",
  2478 => x"527351f5",
  2479 => x"d53f8452",
  2480 => x"7451ffb5",
  2481 => x"3f800874",
  2482 => x"23845284",
  2483 => x"1551ffa9",
  2484 => x"3f800882",
  2485 => x"15238452",
  2486 => x"881551ff",
  2487 => x"9c3f8008",
  2488 => x"84150c84",
  2489 => x"528c1551",
  2490 => x"ff8f3f80",
  2491 => x"08881523",
  2492 => x"84529015",
  2493 => x"51ff823f",
  2494 => x"80088a15",
  2495 => x"23845294",
  2496 => x"1551fef5",
  2497 => x"3f80088c",
  2498 => x"15238452",
  2499 => x"981551fe",
  2500 => x"e83f8008",
  2501 => x"8e152388",
  2502 => x"529c1551",
  2503 => x"fedb3f80",
  2504 => x"0890150c",
  2505 => x"863d0d04",
  2506 => x"e93d0d6a",
  2507 => x"80e1c008",
  2508 => x"57577593",
  2509 => x"3880c080",
  2510 => x"0b84180c",
  2511 => x"75ac180c",
  2512 => x"75800c99",
  2513 => x"3d0d0489",
  2514 => x"3d70556a",
  2515 => x"54558a52",
  2516 => x"993dffbc",
  2517 => x"0551ffb9",
  2518 => x"e93f8008",
  2519 => x"77537552",
  2520 => x"56fecb3f",
  2521 => x"bc3f7780",
  2522 => x"080c7580",
  2523 => x"0c993d0d",
  2524 => x"04fc3d0d",
  2525 => x"815480e1",
  2526 => x"c0088838",
  2527 => x"73800c86",
  2528 => x"3d0d0476",
  2529 => x"5397b952",
  2530 => x"863dfc05",
  2531 => x"51ffb9b2",
  2532 => x"3f800854",
  2533 => x"8c3f7480",
  2534 => x"080c7380",
  2535 => x"0c863d0d",
  2536 => x"0480d1d0",
  2537 => x"08800c04",
  2538 => x"f73d0d7b",
  2539 => x"80d1d008",
  2540 => x"82c81108",
  2541 => x"5a545a77",
  2542 => x"802e80da",
  2543 => x"38818818",
  2544 => x"841908ff",
  2545 => x"0581712b",
  2546 => x"59555980",
  2547 => x"742480ea",
  2548 => x"38807424",
  2549 => x"b5387382",
  2550 => x"2b781188",
  2551 => x"05565681",
  2552 => x"80190877",
  2553 => x"06537280",
  2554 => x"2eb63878",
  2555 => x"16700853",
  2556 => x"53795174",
  2557 => x"0853722d",
  2558 => x"ff14fc17",
  2559 => x"fc177981",
  2560 => x"2c5a5757",
  2561 => x"54738025",
  2562 => x"d6387708",
  2563 => x"5877ffad",
  2564 => x"3880d1d0",
  2565 => x"0853bc13",
  2566 => x"08a53879",
  2567 => x"51f9dc3f",
  2568 => x"74085372",
  2569 => x"2dff14fc",
  2570 => x"17fc1779",
  2571 => x"812c5a57",
  2572 => x"57547380",
  2573 => x"25ffa838",
  2574 => x"d1398057",
  2575 => x"ff933972",
  2576 => x"51bc1308",
  2577 => x"53722d79",
  2578 => x"51f9b03f",
  2579 => x"ff3d0d80",
  2580 => x"e19c0bfc",
  2581 => x"05700852",
  2582 => x"5270ff2e",
  2583 => x"9138702d",
  2584 => x"fc127008",
  2585 => x"525270ff",
  2586 => x"2e098106",
  2587 => x"f138833d",
  2588 => x"0d0404ff",
  2589 => x"b99d3f04",
  2590 => x"00000040",
  2591 => x"72656164",
  2592 => x"2066726f",
  2593 => x"6d206164",
  2594 => x"72657373",
  2595 => x"20307831",
  2596 => x"32333400",
  2597 => x"656e642e",
  2598 => x"00000000",
  2599 => x"0a000000",
  2600 => x"43000000",
  2601 => x"64756d6d",
  2602 => x"792e6578",
  2603 => x"65000000",
  2604 => x"00ffffff",
  2605 => x"ff00ffff",
  2606 => x"ffff00ff",
  2607 => x"ffffff00",
  2608 => x"00000000",
  2609 => x"00000000",
  2610 => x"00000000",
  2611 => x"000030a4",
  2612 => x"000028d4",
  2613 => x"00000000",
  2614 => x"00002b3c",
  2615 => x"00002b98",
  2616 => x"00002bf4",
  2617 => x"00000000",
  2618 => x"00000000",
  2619 => x"00000000",
  2620 => x"00000000",
  2621 => x"00000000",
  2622 => x"00000000",
  2623 => x"00000000",
  2624 => x"00000000",
  2625 => x"00000000",
  2626 => x"000028a0",
  2627 => x"00000000",
  2628 => x"00000000",
  2629 => x"00000000",
  2630 => x"00000000",
  2631 => x"00000000",
  2632 => x"00000000",
  2633 => x"00000000",
  2634 => x"00000000",
  2635 => x"00000000",
  2636 => x"00000000",
  2637 => x"00000000",
  2638 => x"00000000",
  2639 => x"00000000",
  2640 => x"00000000",
  2641 => x"00000000",
  2642 => x"00000000",
  2643 => x"00000000",
  2644 => x"00000000",
  2645 => x"00000000",
  2646 => x"00000000",
  2647 => x"00000000",
  2648 => x"00000000",
  2649 => x"00000000",
  2650 => x"00000000",
  2651 => x"00000000",
  2652 => x"00000000",
  2653 => x"00000000",
  2654 => x"00000000",
  2655 => x"00000001",
  2656 => x"330eabcd",
  2657 => x"1234e66d",
  2658 => x"deec0005",
  2659 => x"000b0000",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000000",
  2683 => x"00000000",
  2684 => x"00000000",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000000",
  2712 => x"00000000",
  2713 => x"00000000",
  2714 => x"00000000",
  2715 => x"00000000",
  2716 => x"00000000",
  2717 => x"00000000",
  2718 => x"00000000",
  2719 => x"00000000",
  2720 => x"00000000",
  2721 => x"00000000",
  2722 => x"00000000",
  2723 => x"00000000",
  2724 => x"00000000",
  2725 => x"00000000",
  2726 => x"00000000",
  2727 => x"00000000",
  2728 => x"00000000",
  2729 => x"00000000",
  2730 => x"00000000",
  2731 => x"00000000",
  2732 => x"00000000",
  2733 => x"00000000",
  2734 => x"00000000",
  2735 => x"00000000",
  2736 => x"00000000",
  2737 => x"00000000",
  2738 => x"00000000",
  2739 => x"00000000",
  2740 => x"00000000",
  2741 => x"00000000",
  2742 => x"00000000",
  2743 => x"00000000",
  2744 => x"00000000",
  2745 => x"00000000",
  2746 => x"00000000",
  2747 => x"00000000",
  2748 => x"00000000",
  2749 => x"00000000",
  2750 => x"00000000",
  2751 => x"00000000",
  2752 => x"00000000",
  2753 => x"00000000",
  2754 => x"00000000",
  2755 => x"00000000",
  2756 => x"00000000",
  2757 => x"00000000",
  2758 => x"00000000",
  2759 => x"00000000",
  2760 => x"00000000",
  2761 => x"00000000",
  2762 => x"00000000",
  2763 => x"00000000",
  2764 => x"00000000",
  2765 => x"00000000",
  2766 => x"00000000",
  2767 => x"00000000",
  2768 => x"00000000",
  2769 => x"00000000",
  2770 => x"00000000",
  2771 => x"00000000",
  2772 => x"00000000",
  2773 => x"00000000",
  2774 => x"00000000",
  2775 => x"00000000",
  2776 => x"00000000",
  2777 => x"00000000",
  2778 => x"00000000",
  2779 => x"00000000",
  2780 => x"00000000",
  2781 => x"00000000",
  2782 => x"00000000",
  2783 => x"00000000",
  2784 => x"00000000",
  2785 => x"00000000",
  2786 => x"00000000",
  2787 => x"00000000",
  2788 => x"00000000",
  2789 => x"00000000",
  2790 => x"00000000",
  2791 => x"00000000",
  2792 => x"00000000",
  2793 => x"00000000",
  2794 => x"00000000",
  2795 => x"00000000",
  2796 => x"00000000",
  2797 => x"00000000",
  2798 => x"00000000",
  2799 => x"00000000",
  2800 => x"00000000",
  2801 => x"00000000",
  2802 => x"00000000",
  2803 => x"00000000",
  2804 => x"00000000",
  2805 => x"00000000",
  2806 => x"00000000",
  2807 => x"00000000",
  2808 => x"00000000",
  2809 => x"00000000",
  2810 => x"00000000",
  2811 => x"00000000",
  2812 => x"00000000",
  2813 => x"00000000",
  2814 => x"00000000",
  2815 => x"00000000",
  2816 => x"00000000",
  2817 => x"00000000",
  2818 => x"00000000",
  2819 => x"00000000",
  2820 => x"00000000",
  2821 => x"00000000",
  2822 => x"00000000",
  2823 => x"00000000",
  2824 => x"00000000",
  2825 => x"00000000",
  2826 => x"00000000",
  2827 => x"00000000",
  2828 => x"00000000",
  2829 => x"00000000",
  2830 => x"00000000",
  2831 => x"00000000",
  2832 => x"00000000",
  2833 => x"00000000",
  2834 => x"00000000",
  2835 => x"00000000",
  2836 => x"00000000",
  2837 => x"00000000",
  2838 => x"00000000",
  2839 => x"00000000",
  2840 => x"00000000",
  2841 => x"00000000",
  2842 => x"00000000",
  2843 => x"00000000",
  2844 => x"00000000",
  2845 => x"00000000",
  2846 => x"00000000",
  2847 => x"00000000",
  2848 => x"ffffffff",
  2849 => x"00000000",
  2850 => x"00020000",
  2851 => x"00000000",
  2852 => x"00000000",
  2853 => x"00002c8c",
  2854 => x"00002c8c",
  2855 => x"00002c94",
  2856 => x"00002c94",
  2857 => x"00002c9c",
  2858 => x"00002c9c",
  2859 => x"00002ca4",
  2860 => x"00002ca4",
  2861 => x"00002cac",
  2862 => x"00002cac",
  2863 => x"00002cb4",
  2864 => x"00002cb4",
  2865 => x"00002cbc",
  2866 => x"00002cbc",
  2867 => x"00002cc4",
  2868 => x"00002cc4",
  2869 => x"00002ccc",
  2870 => x"00002ccc",
  2871 => x"00002cd4",
  2872 => x"00002cd4",
  2873 => x"00002cdc",
  2874 => x"00002cdc",
  2875 => x"00002ce4",
  2876 => x"00002ce4",
  2877 => x"00002cec",
  2878 => x"00002cec",
  2879 => x"00002cf4",
  2880 => x"00002cf4",
  2881 => x"00002cfc",
  2882 => x"00002cfc",
  2883 => x"00002d04",
  2884 => x"00002d04",
  2885 => x"00002d0c",
  2886 => x"00002d0c",
  2887 => x"00002d14",
  2888 => x"00002d14",
  2889 => x"00002d1c",
  2890 => x"00002d1c",
  2891 => x"00002d24",
  2892 => x"00002d24",
  2893 => x"00002d2c",
  2894 => x"00002d2c",
  2895 => x"00002d34",
  2896 => x"00002d34",
  2897 => x"00002d3c",
  2898 => x"00002d3c",
  2899 => x"00002d44",
  2900 => x"00002d44",
  2901 => x"00002d4c",
  2902 => x"00002d4c",
  2903 => x"00002d54",
  2904 => x"00002d54",
  2905 => x"00002d5c",
  2906 => x"00002d5c",
  2907 => x"00002d64",
  2908 => x"00002d64",
  2909 => x"00002d6c",
  2910 => x"00002d6c",
  2911 => x"00002d74",
  2912 => x"00002d74",
  2913 => x"00002d7c",
  2914 => x"00002d7c",
  2915 => x"00002d84",
  2916 => x"00002d84",
  2917 => x"00002d8c",
  2918 => x"00002d8c",
  2919 => x"00002d94",
  2920 => x"00002d94",
  2921 => x"00002d9c",
  2922 => x"00002d9c",
  2923 => x"00002da4",
  2924 => x"00002da4",
  2925 => x"00002dac",
  2926 => x"00002dac",
  2927 => x"00002db4",
  2928 => x"00002db4",
  2929 => x"00002dbc",
  2930 => x"00002dbc",
  2931 => x"00002dc4",
  2932 => x"00002dc4",
  2933 => x"00002dcc",
  2934 => x"00002dcc",
  2935 => x"00002dd4",
  2936 => x"00002dd4",
  2937 => x"00002ddc",
  2938 => x"00002ddc",
  2939 => x"00002de4",
  2940 => x"00002de4",
  2941 => x"00002dec",
  2942 => x"00002dec",
  2943 => x"00002df4",
  2944 => x"00002df4",
  2945 => x"00002dfc",
  2946 => x"00002dfc",
  2947 => x"00002e04",
  2948 => x"00002e04",
  2949 => x"00002e0c",
  2950 => x"00002e0c",
  2951 => x"00002e14",
  2952 => x"00002e14",
  2953 => x"00002e1c",
  2954 => x"00002e1c",
  2955 => x"00002e24",
  2956 => x"00002e24",
  2957 => x"00002e2c",
  2958 => x"00002e2c",
  2959 => x"00002e34",
  2960 => x"00002e34",
  2961 => x"00002e3c",
  2962 => x"00002e3c",
  2963 => x"00002e44",
  2964 => x"00002e44",
  2965 => x"00002e4c",
  2966 => x"00002e4c",
  2967 => x"00002e54",
  2968 => x"00002e54",
  2969 => x"00002e5c",
  2970 => x"00002e5c",
  2971 => x"00002e64",
  2972 => x"00002e64",
  2973 => x"00002e6c",
  2974 => x"00002e6c",
  2975 => x"00002e74",
  2976 => x"00002e74",
  2977 => x"00002e7c",
  2978 => x"00002e7c",
  2979 => x"00002e84",
  2980 => x"00002e84",
  2981 => x"00002e8c",
  2982 => x"00002e8c",
  2983 => x"00002e94",
  2984 => x"00002e94",
  2985 => x"00002e9c",
  2986 => x"00002e9c",
  2987 => x"00002ea4",
  2988 => x"00002ea4",
  2989 => x"00002eac",
  2990 => x"00002eac",
  2991 => x"00002eb4",
  2992 => x"00002eb4",
  2993 => x"00002ebc",
  2994 => x"00002ebc",
  2995 => x"00002ec4",
  2996 => x"00002ec4",
  2997 => x"00002ecc",
  2998 => x"00002ecc",
  2999 => x"00002ed4",
  3000 => x"00002ed4",
  3001 => x"00002edc",
  3002 => x"00002edc",
  3003 => x"00002ee4",
  3004 => x"00002ee4",
  3005 => x"00002eec",
  3006 => x"00002eec",
  3007 => x"00002ef4",
  3008 => x"00002ef4",
  3009 => x"00002efc",
  3010 => x"00002efc",
  3011 => x"00002f04",
  3012 => x"00002f04",
  3013 => x"00002f0c",
  3014 => x"00002f0c",
  3015 => x"00002f14",
  3016 => x"00002f14",
  3017 => x"00002f1c",
  3018 => x"00002f1c",
  3019 => x"00002f24",
  3020 => x"00002f24",
  3021 => x"00002f2c",
  3022 => x"00002f2c",
  3023 => x"00002f34",
  3024 => x"00002f34",
  3025 => x"00002f3c",
  3026 => x"00002f3c",
  3027 => x"00002f44",
  3028 => x"00002f44",
  3029 => x"00002f4c",
  3030 => x"00002f4c",
  3031 => x"00002f54",
  3032 => x"00002f54",
  3033 => x"00002f5c",
  3034 => x"00002f5c",
  3035 => x"00002f64",
  3036 => x"00002f64",
  3037 => x"00002f6c",
  3038 => x"00002f6c",
  3039 => x"00002f74",
  3040 => x"00002f74",
  3041 => x"00002f7c",
  3042 => x"00002f7c",
  3043 => x"00002f84",
  3044 => x"00002f84",
  3045 => x"00002f8c",
  3046 => x"00002f8c",
  3047 => x"00002f94",
  3048 => x"00002f94",
  3049 => x"00002f9c",
  3050 => x"00002f9c",
  3051 => x"00002fa4",
  3052 => x"00002fa4",
  3053 => x"00002fac",
  3054 => x"00002fac",
  3055 => x"00002fb4",
  3056 => x"00002fb4",
  3057 => x"00002fbc",
  3058 => x"00002fbc",
  3059 => x"00002fc4",
  3060 => x"00002fc4",
  3061 => x"00002fcc",
  3062 => x"00002fcc",
  3063 => x"00002fd4",
  3064 => x"00002fd4",
  3065 => x"00002fdc",
  3066 => x"00002fdc",
  3067 => x"00002fe4",
  3068 => x"00002fe4",
  3069 => x"00002fec",
  3070 => x"00002fec",
  3071 => x"00002ff4",
  3072 => x"00002ff4",
  3073 => x"00002ffc",
  3074 => x"00002ffc",
  3075 => x"00003004",
  3076 => x"00003004",
  3077 => x"0000300c",
  3078 => x"0000300c",
  3079 => x"00003014",
  3080 => x"00003014",
  3081 => x"0000301c",
  3082 => x"0000301c",
  3083 => x"00003024",
  3084 => x"00003024",
  3085 => x"0000302c",
  3086 => x"0000302c",
  3087 => x"00003034",
  3088 => x"00003034",
  3089 => x"0000303c",
  3090 => x"0000303c",
  3091 => x"00003044",
  3092 => x"00003044",
  3093 => x"0000304c",
  3094 => x"0000304c",
  3095 => x"00003054",
  3096 => x"00003054",
  3097 => x"0000305c",
  3098 => x"0000305c",
  3099 => x"00003064",
  3100 => x"00003064",
  3101 => x"0000306c",
  3102 => x"0000306c",
  3103 => x"00003074",
  3104 => x"00003074",
  3105 => x"0000307c",
  3106 => x"0000307c",
  3107 => x"00003084",
  3108 => x"00003084",
  3109 => x"000028a4",
  3110 => x"ffffffff",
  3111 => x"00000000",
  3112 => x"ffffffff",
  3113 => x"00000000",
  3114 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
