-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b80f5",
     1 => x"e4040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b80f8",
     9 => x"cb040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b80f7",
    73 => x"fd040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b80f7e0",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b81ce",
   162 => x"d0738306",
   163 => x"10100508",
   164 => x"060b0b80",
   165 => x"f7e30400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b80f8",
   169 => x"b2040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b80f8",
   177 => x"99040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"81cee00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053370",
   258 => x"525280f5",
   259 => x"a63f7151",
   260 => x"80f6943f",
   261 => x"71b00c83",
   262 => x"3d0d04ff",
   263 => x"3d0d81ce",
   264 => x"bc08b811",
   265 => x"08535180",
   266 => x"0bb8120c",
   267 => x"71b00c83",
   268 => x"3d0d0480",
   269 => x"0b81f1f0",
   270 => x"34800bb0",
   271 => x"0c04fb3d",
   272 => x"0d815180",
   273 => x"c7ce3fb0",
   274 => x"08538251",
   275 => x"80c7c53f",
   276 => x"b00856b0",
   277 => x"08833890",
   278 => x"5672fc06",
   279 => x"5575812e",
   280 => x"80fb3880",
   281 => x"54737627",
   282 => x"ad387383",
   283 => x"06537280",
   284 => x"2eb23881",
   285 => x"c2c05180",
   286 => x"f0923f74",
   287 => x"70840556",
   288 => x"0852a051",
   289 => x"80f0a83f",
   290 => x"a05180ef",
   291 => x"e53f8114",
   292 => x"54757426",
   293 => x"d5388a51",
   294 => x"80efd73f",
   295 => x"800bb00c",
   296 => x"873d0d04",
   297 => x"81a7d051",
   298 => x"80efe13f",
   299 => x"7452a051",
   300 => x"80effc3f",
   301 => x"81b4bc51",
   302 => x"80efd13f",
   303 => x"81c2c051",
   304 => x"80efc93f",
   305 => x"74708405",
   306 => x"560852a0",
   307 => x"5180efdf",
   308 => x"3fa05180",
   309 => x"ef9c3f81",
   310 => x"1454ffb5",
   311 => x"3981c2c0",
   312 => x"5180efa8",
   313 => x"3f740852",
   314 => x"a05180ef",
   315 => x"c23f8a51",
   316 => x"80eeff3f",
   317 => x"800bb00c",
   318 => x"873d0d04",
   319 => x"fc3d0d81",
   320 => x"5180c690",
   321 => x"3fb00852",
   322 => x"825180c4",
   323 => x"d53fb008",
   324 => x"81ff0672",
   325 => x"56538354",
   326 => x"72802ea2",
   327 => x"38735180",
   328 => x"c5f23f81",
   329 => x"147081ff",
   330 => x"06ff1570",
   331 => x"81ff06b0",
   332 => x"08797084",
   333 => x"055b0c56",
   334 => x"52555272",
   335 => x"e03872b0",
   336 => x"0c863d0d",
   337 => x"04803d0d",
   338 => x"8c5180ee",
   339 => x"a53f800b",
   340 => x"b00c823d",
   341 => x"0d04fb3d",
   342 => x"0d800b81",
   343 => x"a7d45256",
   344 => x"80eea93f",
   345 => x"75557410",
   346 => x"81fe0653",
   347 => x"81d05281",
   348 => x"cee80851",
   349 => x"80d2d33f",
   350 => x"b008982b",
   351 => x"54807424",
   352 => x"a23881a7",
   353 => x"e05180ee",
   354 => x"833f7452",
   355 => x"885180ee",
   356 => x"9e3f81a7",
   357 => x"ec5180ed",
   358 => x"f33f8116",
   359 => x"7083ffff",
   360 => x"06575481",
   361 => x"157081ff",
   362 => x"0670982b",
   363 => x"52565473",
   364 => x"8025ffb2",
   365 => x"3875b00c",
   366 => x"873d0d04",
   367 => x"f33d0d7f",
   368 => x"02840580",
   369 => x"c3053302",
   370 => x"880580c6",
   371 => x"052281a7",
   372 => x"fc545b55",
   373 => x"5880edb4",
   374 => x"3f785180",
   375 => x"eef83f81",
   376 => x"a8885180",
   377 => x"eda63f73",
   378 => x"52885180",
   379 => x"edc13f81",
   380 => x"a8a45180",
   381 => x"ed963f80",
   382 => x"57767927",
   383 => x"81a13873",
   384 => x"108e3d5d",
   385 => x"5a7981ff",
   386 => x"06538190",
   387 => x"52775180",
   388 => x"d1b83f76",
   389 => x"882a5390",
   390 => x"52775180",
   391 => x"d1ac3f76",
   392 => x"81ff0653",
   393 => x"90527751",
   394 => x"80d19f3f",
   395 => x"811a7081",
   396 => x"ff065455",
   397 => x"81905277",
   398 => x"5180d18e",
   399 => x"3f805380",
   400 => x"e0527751",
   401 => x"80d1833f",
   402 => x"b008982b",
   403 => x"54807424",
   404 => x"8a388818",
   405 => x"087081ff",
   406 => x"065c567a",
   407 => x"81ff0681",
   408 => x"c2c05256",
   409 => x"80eca53f",
   410 => x"75528851",
   411 => x"80ecc03f",
   412 => x"81b29851",
   413 => x"80ec953f",
   414 => x"e0165480",
   415 => x"df7427b6",
   416 => x"38768706",
   417 => x"701d5755",
   418 => x"a0763474",
   419 => x"872eb938",
   420 => x"81177083",
   421 => x"ffff0658",
   422 => x"55787726",
   423 => x"fee73880",
   424 => x"e00b8c19",
   425 => x"0c8c1808",
   426 => x"70812a81",
   427 => x"06585a76",
   428 => x"f4388f3d",
   429 => x"0d047687",
   430 => x"06701d55",
   431 => x"55757434",
   432 => x"74872e09",
   433 => x"8106c938",
   434 => x"7b5180eb",
   435 => x"bf3f8a51",
   436 => x"80eb9f3f",
   437 => x"81177083",
   438 => x"ffff0658",
   439 => x"55787726",
   440 => x"fea338ff",
   441 => x"ba39fb3d",
   442 => x"0d815180",
   443 => x"c0f43fb0",
   444 => x"0881ff06",
   445 => x"54825180",
   446 => x"c29a3fb0",
   447 => x"0881ff06",
   448 => x"56835180",
   449 => x"c0dc3fb0",
   450 => x"0883ffff",
   451 => x"0655739c",
   452 => x"3881cee8",
   453 => x"08547484",
   454 => x"38818055",
   455 => x"74537552",
   456 => x"7351fd98",
   457 => x"3f74b00c",
   458 => x"873d0d04",
   459 => x"81ceec08",
   460 => x"54e439f8",
   461 => x"3d0d02aa",
   462 => x"052281ce",
   463 => x"c43381f7",
   464 => x"06585876",
   465 => x"81cec434",
   466 => x"81cee808",
   467 => x"5580c053",
   468 => x"81905274",
   469 => x"5180cef2",
   470 => x"3f745180",
   471 => x"cf9e3fb0",
   472 => x"0881ff06",
   473 => x"5473802e",
   474 => x"84903876",
   475 => x"5380d052",
   476 => x"745180ce",
   477 => x"d53f8059",
   478 => x"8f5781ce",
   479 => x"c43381fe",
   480 => x"06547381",
   481 => x"cec43481",
   482 => x"cee80874",
   483 => x"575580c0",
   484 => x"53819052",
   485 => x"745180ce",
   486 => x"b13f7451",
   487 => x"80cedd3f",
   488 => x"b00881ff",
   489 => x"06547380",
   490 => x"2e83c438",
   491 => x"755380d0",
   492 => x"52745180",
   493 => x"ce943f77",
   494 => x"772c8106",
   495 => x"5574802e",
   496 => x"83a23881",
   497 => x"cec43382",
   498 => x"07547381",
   499 => x"cec43481",
   500 => x"cee80874",
   501 => x"575580c0",
   502 => x"53819052",
   503 => x"745180cd",
   504 => x"e93f7451",
   505 => x"80ce953f",
   506 => x"b00881ff",
   507 => x"06547380",
   508 => x"2e82e638",
   509 => x"755380d0",
   510 => x"52745180",
   511 => x"cdcc3f81",
   512 => x"cee80855",
   513 => x"80c15381",
   514 => x"90527451",
   515 => x"80cdbb3f",
   516 => x"745180cd",
   517 => x"e73fb008",
   518 => x"81ff0656",
   519 => x"75802e82",
   520 => x"8c388053",
   521 => x"80e05274",
   522 => x"5180cd9e",
   523 => x"3f745180",
   524 => x"cdca3fb0",
   525 => x"0881ff06",
   526 => x"5473802e",
   527 => x"81ef3888",
   528 => x"15087090",
   529 => x"2b70902c",
   530 => x"56565673",
   531 => x"822a8106",
   532 => x"5473802e",
   533 => x"8d388177",
   534 => x"2b790770",
   535 => x"83ffff06",
   536 => x"5a5681ce",
   537 => x"c4338107",
   538 => x"547381ce",
   539 => x"c43481ce",
   540 => x"e8087457",
   541 => x"5580c053",
   542 => x"81905274",
   543 => x"5180ccca",
   544 => x"3f745180",
   545 => x"ccf63fb0",
   546 => x"0881ff06",
   547 => x"5473802e",
   548 => x"81a83875",
   549 => x"5380d052",
   550 => x"745180cc",
   551 => x"ad3f7681",
   552 => x"800a2981",
   553 => x"ff0a0570",
   554 => x"982c5856",
   555 => x"768025fd",
   556 => x"c93881ce",
   557 => x"c4338207",
   558 => x"577681ce",
   559 => x"c43481ce",
   560 => x"e8085580",
   561 => x"c0538190",
   562 => x"52745180",
   563 => x"cbfc3f74",
   564 => x"5180cca8",
   565 => x"3fb00881",
   566 => x"ff065877",
   567 => x"802e81b8",
   568 => x"38765380",
   569 => x"d0527451",
   570 => x"80cbdf3f",
   571 => x"81cec433",
   572 => x"88075776",
   573 => x"81cec434",
   574 => x"81cee808",
   575 => x"5580c053",
   576 => x"81905274",
   577 => x"5180cbc2",
   578 => x"3f745180",
   579 => x"cbee3fb0",
   580 => x"0881ff06",
   581 => x"5877802e",
   582 => x"80ef3876",
   583 => x"5380d052",
   584 => x"745180cb",
   585 => x"a53f78b0",
   586 => x"0c8a3d0d",
   587 => x"0481a8a8",
   588 => x"5180e6d8",
   589 => x"3fff54fe",
   590 => x"923981a8",
   591 => x"a85180e6",
   592 => x"cb3f7681",
   593 => x"800a2981",
   594 => x"ff0a0570",
   595 => x"982c5856",
   596 => x"768025fc",
   597 => x"a538feda",
   598 => x"3981a8a8",
   599 => x"5180e6ac",
   600 => x"3ffd9c39",
   601 => x"81cec433",
   602 => x"81fd0654",
   603 => x"fcdc3981",
   604 => x"a8a85180",
   605 => x"e6963ffc",
   606 => x"be3981a8",
   607 => x"a85180e6",
   608 => x"8b3f8059",
   609 => x"8f57fbf2",
   610 => x"3981a8a8",
   611 => x"5180e5fc",
   612 => x"3f78b00c",
   613 => x"8a3d0d04",
   614 => x"81a8a851",
   615 => x"80e5ed3f",
   616 => x"feca39ff",
   617 => x"3d0d8151",
   618 => x"bbb83fb0",
   619 => x"0881ff06",
   620 => x"52818051",
   621 => x"fafd3f82",
   622 => x"8051faf7",
   623 => x"3f848351",
   624 => x"faf13f86",
   625 => x"f151faeb",
   626 => x"3f71832b",
   627 => x"88830751",
   628 => x"fae13f71",
   629 => x"b00c833d",
   630 => x"0d04fe3d",
   631 => x"0d029305",
   632 => x"33028405",
   633 => x"97053354",
   634 => x"52717327",
   635 => x"9438a051",
   636 => x"80e4ff3f",
   637 => x"81127081",
   638 => x"ff065152",
   639 => x"727226ee",
   640 => x"38843d0d",
   641 => x"04fe3d0d",
   642 => x"74708106",
   643 => x"53537185",
   644 => x"d0387281",
   645 => x"2a708106",
   646 => x"51527185",
   647 => x"ac387282",
   648 => x"2a708106",
   649 => x"51527185",
   650 => x"88387283",
   651 => x"2a708106",
   652 => x"51527184",
   653 => x"e4387284",
   654 => x"2a708106",
   655 => x"51527184",
   656 => x"c0387285",
   657 => x"2a708106",
   658 => x"51527184",
   659 => x"9c387286",
   660 => x"2a708106",
   661 => x"51527183",
   662 => x"f8387287",
   663 => x"2a708106",
   664 => x"51527183",
   665 => x"d4387288",
   666 => x"2a708106",
   667 => x"51527183",
   668 => x"b0387289",
   669 => x"2a708106",
   670 => x"51527183",
   671 => x"8c38728a",
   672 => x"2a708106",
   673 => x"51527182",
   674 => x"e838728b",
   675 => x"2a708106",
   676 => x"51527182",
   677 => x"c438728c",
   678 => x"2a708106",
   679 => x"51527182",
   680 => x"a038728d",
   681 => x"2a708106",
   682 => x"51527181",
   683 => x"fc38728e",
   684 => x"2a708106",
   685 => x"51527181",
   686 => x"d838728f",
   687 => x"2a708106",
   688 => x"51527181",
   689 => x"b4387290",
   690 => x"2a708106",
   691 => x"51527181",
   692 => x"90387291",
   693 => x"2a708106",
   694 => x"51527180",
   695 => x"ec387292",
   696 => x"2a708106",
   697 => x"51527180",
   698 => x"c8387293",
   699 => x"2a708106",
   700 => x"515271a6",
   701 => x"3872942a",
   702 => x"70810651",
   703 => x"52718b38",
   704 => x"80732483",
   705 => x"f438843d",
   706 => x"0d0481a8",
   707 => x"e05180e2",
   708 => x"fb3f7280",
   709 => x"25f03883",
   710 => x"e03981a8",
   711 => x"fc5180e2",
   712 => x"eb3f7294",
   713 => x"2a708106",
   714 => x"51527180",
   715 => x"2ed238da",
   716 => x"3981a998",
   717 => x"5180e2d4",
   718 => x"3f72932a",
   719 => x"70810651",
   720 => x"5271802e",
   721 => x"ffaf38d2",
   722 => x"3981a9b4",
   723 => x"5180e2bc",
   724 => x"3f72922a",
   725 => x"70810651",
   726 => x"5271802e",
   727 => x"ff8c38d1",
   728 => x"3981a9d0",
   729 => x"5180e2a4",
   730 => x"3f72912a",
   731 => x"70810651",
   732 => x"5271802e",
   733 => x"fee838d1",
   734 => x"3981a9f0",
   735 => x"5180e28c",
   736 => x"3f72902a",
   737 => x"70810651",
   738 => x"5271802e",
   739 => x"fec438d1",
   740 => x"3981aa90",
   741 => x"5180e1f4",
   742 => x"3f728f2a",
   743 => x"70810651",
   744 => x"5271802e",
   745 => x"fea038d1",
   746 => x"3981aab0",
   747 => x"5180e1dc",
   748 => x"3f728e2a",
   749 => x"70810651",
   750 => x"5271802e",
   751 => x"fdfc38d1",
   752 => x"3981aad0",
   753 => x"5180e1c4",
   754 => x"3f728d2a",
   755 => x"70810651",
   756 => x"5271802e",
   757 => x"fdd838d1",
   758 => x"3981aae4",
   759 => x"5180e1ac",
   760 => x"3f728c2a",
   761 => x"70810651",
   762 => x"5271802e",
   763 => x"fdb438d1",
   764 => x"3981ab84",
   765 => x"5180e194",
   766 => x"3f728b2a",
   767 => x"70810651",
   768 => x"5271802e",
   769 => x"fd9038d1",
   770 => x"3981abac",
   771 => x"5180e0fc",
   772 => x"3f728a2a",
   773 => x"70810651",
   774 => x"5271802e",
   775 => x"fcec38d1",
   776 => x"3981abcc",
   777 => x"5180e0e4",
   778 => x"3f72892a",
   779 => x"70810651",
   780 => x"5271802e",
   781 => x"fcc838d1",
   782 => x"3981abec",
   783 => x"5180e0cc",
   784 => x"3f72882a",
   785 => x"70810651",
   786 => x"5271802e",
   787 => x"fca438d1",
   788 => x"3981ac94",
   789 => x"5180e0b4",
   790 => x"3f72872a",
   791 => x"70810651",
   792 => x"5271802e",
   793 => x"fc8038d1",
   794 => x"3981acb4",
   795 => x"5180e09c",
   796 => x"3f72862a",
   797 => x"70810651",
   798 => x"5271802e",
   799 => x"fbdc38d1",
   800 => x"3981acd4",
   801 => x"5180e084",
   802 => x"3f72852a",
   803 => x"70810651",
   804 => x"5271802e",
   805 => x"fbb838d1",
   806 => x"3981acfc",
   807 => x"5180dfec",
   808 => x"3f72842a",
   809 => x"70810651",
   810 => x"5271802e",
   811 => x"fb9438d1",
   812 => x"3981ad9c",
   813 => x"5180dfd4",
   814 => x"3f72832a",
   815 => x"70810651",
   816 => x"5271802e",
   817 => x"faf038d1",
   818 => x"3981adbc",
   819 => x"5180dfbc",
   820 => x"3f72822a",
   821 => x"70810651",
   822 => x"5271802e",
   823 => x"facc38d1",
   824 => x"3981ade4",
   825 => x"5180dfa4",
   826 => x"3f72812a",
   827 => x"70810651",
   828 => x"5271802e",
   829 => x"faa838d1",
   830 => x"3981ae84",
   831 => x"5180df8c",
   832 => x"3f843d0d",
   833 => x"04fd3d0d",
   834 => x"81ae9851",
   835 => x"80defd3f",
   836 => x"81cef408",
   837 => x"7008709e",
   838 => x"2a708106",
   839 => x"51525553",
   840 => x"81547283",
   841 => x"38725473",
   842 => x"802e88c4",
   843 => x"3881aeb4",
   844 => x"5180ded8",
   845 => x"3f81aebc",
   846 => x"5180ded0",
   847 => x"3f81cef4",
   848 => x"08841108",
   849 => x"709d2a81",
   850 => x"06515553",
   851 => x"73802e87",
   852 => x"b03881ae",
   853 => x"d85180de",
   854 => x"b33f81ae",
   855 => x"e45180de",
   856 => x"ab3f81ce",
   857 => x"bc0880d4",
   858 => x"11085254",
   859 => x"80dfe73f",
   860 => x"81af8051",
   861 => x"80de953f",
   862 => x"81cebc08",
   863 => x"80d01108",
   864 => x"525380df",
   865 => x"d13f8a51",
   866 => x"80dde73f",
   867 => x"81af9c51",
   868 => x"80ddf93f",
   869 => x"81afc051",
   870 => x"80ddf13f",
   871 => x"81b08851",
   872 => x"80dde93f",
   873 => x"81b0d051",
   874 => x"80dde13f",
   875 => x"81cebc08",
   876 => x"70085254",
   877 => x"80df9f3f",
   878 => x"b00881ff",
   879 => x"0653728c",
   880 => x"279438a0",
   881 => x"5180ddaa",
   882 => x"3f811370",
   883 => x"81ff0651",
   884 => x"538c7326",
   885 => x"ee3881ce",
   886 => x"bc088411",
   887 => x"08525480",
   888 => x"def43fb0",
   889 => x"0881ff06",
   890 => x"53728c27",
   891 => x"9438a051",
   892 => x"80dcff3f",
   893 => x"81137081",
   894 => x"ff065153",
   895 => x"8c7326ee",
   896 => x"3881cebc",
   897 => x"08881108",
   898 => x"525480de",
   899 => x"c93fb008",
   900 => x"81ff0653",
   901 => x"728c2794",
   902 => x"38a05180",
   903 => x"dcd43f81",
   904 => x"137081ff",
   905 => x"0651538c",
   906 => x"7326ee38",
   907 => x"81cebc08",
   908 => x"8c110852",
   909 => x"5480de9e",
   910 => x"3fb00881",
   911 => x"ff065372",
   912 => x"8c279438",
   913 => x"a05180dc",
   914 => x"a93f8113",
   915 => x"7081ff06",
   916 => x"51538c73",
   917 => x"26ee3881",
   918 => x"b0ec5180",
   919 => x"dcae3f81",
   920 => x"cebc0890",
   921 => x"11085254",
   922 => x"80ddeb3f",
   923 => x"b00881ff",
   924 => x"0653728c",
   925 => x"279438a0",
   926 => x"5180dbf6",
   927 => x"3f811370",
   928 => x"81ff0651",
   929 => x"538c7326",
   930 => x"ee3881ce",
   931 => x"bc089411",
   932 => x"08525480",
   933 => x"ddc03fb0",
   934 => x"0881ff06",
   935 => x"53728c27",
   936 => x"9438a051",
   937 => x"80dbcb3f",
   938 => x"81137081",
   939 => x"ff065153",
   940 => x"8c7326ee",
   941 => x"3881cebc",
   942 => x"08981108",
   943 => x"525480dd",
   944 => x"953fb008",
   945 => x"81ff0653",
   946 => x"728c2794",
   947 => x"38a05180",
   948 => x"dba03f81",
   949 => x"137081ff",
   950 => x"0651538c",
   951 => x"7326ee38",
   952 => x"81cebc08",
   953 => x"9c110852",
   954 => x"5480dcea",
   955 => x"3fb00881",
   956 => x"ff065372",
   957 => x"8c279438",
   958 => x"a05180da",
   959 => x"f53f8113",
   960 => x"7081ff06",
   961 => x"51538c73",
   962 => x"26ee3881",
   963 => x"b1885180",
   964 => x"dafa3f81",
   965 => x"cebc0854",
   966 => x"810bb015",
   967 => x"0cb01408",
   968 => x"53728025",
   969 => x"f838a014",
   970 => x"085180dc",
   971 => x"a93fb008",
   972 => x"81ff0653",
   973 => x"728c2794",
   974 => x"38a05180",
   975 => x"dab43f81",
   976 => x"137081ff",
   977 => x"0654548c",
   978 => x"7326ee38",
   979 => x"81cebc08",
   980 => x"a4110852",
   981 => x"5380dbfe",
   982 => x"3fb00881",
   983 => x"ff065372",
   984 => x"8c279438",
   985 => x"a05180da",
   986 => x"893f8113",
   987 => x"7081ff06",
   988 => x"54548c73",
   989 => x"26ee3881",
   990 => x"cebc08a8",
   991 => x"11085253",
   992 => x"80dbd33f",
   993 => x"b00881ff",
   994 => x"0653728c",
   995 => x"279438a0",
   996 => x"5180d9de",
   997 => x"3f811370",
   998 => x"81ff0654",
   999 => x"548c7326",
  1000 => x"ee3881ce",
  1001 => x"bc08ac11",
  1002 => x"08525380",
  1003 => x"dba83fb0",
  1004 => x"0881ff06",
  1005 => x"53728c27",
  1006 => x"9438a051",
  1007 => x"80d9b33f",
  1008 => x"81137081",
  1009 => x"ff065454",
  1010 => x"8c7326ee",
  1011 => x"3881b1a4",
  1012 => x"5180d9b8",
  1013 => x"3f81cebc",
  1014 => x"0880e011",
  1015 => x"08525380",
  1016 => x"daf43f81",
  1017 => x"b1b85180",
  1018 => x"d9a23f81",
  1019 => x"cebc08b0",
  1020 => x"1108fe0a",
  1021 => x"06525480",
  1022 => x"dadc3f81",
  1023 => x"cebc0854",
  1024 => x"800bb015",
  1025 => x"0c81b1cc",
  1026 => x"5180d980",
  1027 => x"3f81b1e4",
  1028 => x"5180d8f8",
  1029 => x"3f81cebc",
  1030 => x"0880c011",
  1031 => x"08525380",
  1032 => x"dab43fb0",
  1033 => x"0881ff06",
  1034 => x"53729827",
  1035 => x"9438a051",
  1036 => x"80d8bf3f",
  1037 => x"81137081",
  1038 => x"ff065454",
  1039 => x"987326ee",
  1040 => x"3881cebc",
  1041 => x"0880c811",
  1042 => x"08525380",
  1043 => x"da883fb0",
  1044 => x"0881ff06",
  1045 => x"53729827",
  1046 => x"9438a051",
  1047 => x"80d8933f",
  1048 => x"81137081",
  1049 => x"ff065454",
  1050 => x"987326ee",
  1051 => x"3881b280",
  1052 => x"5180d898",
  1053 => x"3f81cebc",
  1054 => x"0880c411",
  1055 => x"08525380",
  1056 => x"d9d43fb0",
  1057 => x"0881ff06",
  1058 => x"53729827",
  1059 => x"9438a051",
  1060 => x"80d7df3f",
  1061 => x"81137081",
  1062 => x"ff065454",
  1063 => x"987326ee",
  1064 => x"3881cebc",
  1065 => x"0880cc11",
  1066 => x"08525380",
  1067 => x"d9a83fb0",
  1068 => x"0881ff06",
  1069 => x"53729827",
  1070 => x"9438a051",
  1071 => x"80d7b33f",
  1072 => x"81137081",
  1073 => x"ff065454",
  1074 => x"987326ee",
  1075 => x"388a5180",
  1076 => x"d7a03f81",
  1077 => x"cebc08b4",
  1078 => x"110881b2",
  1079 => x"9c535153",
  1080 => x"80d7a93f",
  1081 => x"725180d8",
  1082 => x"ed3fa051",
  1083 => x"80d7833f",
  1084 => x"72862681",
  1085 => x"8e387210",
  1086 => x"1081bec0",
  1087 => x"05547308",
  1088 => x"0481b2b0",
  1089 => x"5180d784",
  1090 => x"3f81aee4",
  1091 => x"5180d6fc",
  1092 => x"3f81cebc",
  1093 => x"0880d411",
  1094 => x"08525480",
  1095 => x"d8b83f81",
  1096 => x"af805180",
  1097 => x"d6e63f81",
  1098 => x"cebc0880",
  1099 => x"d0110852",
  1100 => x"5380d8a2",
  1101 => x"3f8a5180",
  1102 => x"d6b83f81",
  1103 => x"af9c5180",
  1104 => x"d6ca3f81",
  1105 => x"afc05180",
  1106 => x"d6c23f81",
  1107 => x"b0885180",
  1108 => x"d6ba3f81",
  1109 => x"b0d05180",
  1110 => x"d6b23f81",
  1111 => x"cebc0870",
  1112 => x"08525480",
  1113 => x"d7f03fb0",
  1114 => x"0881ff06",
  1115 => x"53f8cf39",
  1116 => x"81b2b851",
  1117 => x"80d6953f",
  1118 => x"f7b33981",
  1119 => x"b2c05180",
  1120 => x"d68a3f81",
  1121 => x"cebc08b8",
  1122 => x"110881b2",
  1123 => x"cc535454",
  1124 => x"80d5f93f",
  1125 => x"7252a051",
  1126 => x"80d6943f",
  1127 => x"7251f0e5",
  1128 => x"3f8a5180",
  1129 => x"d5cc3f80",
  1130 => x"0bb00c85",
  1131 => x"3d0d0481",
  1132 => x"b2e05180",
  1133 => x"d5d63fcb",
  1134 => x"3981b2ec",
  1135 => x"5180d5cc",
  1136 => x"3fc13981",
  1137 => x"b2f85180",
  1138 => x"d5c23fff",
  1139 => x"b63981b2",
  1140 => x"fc5180d5",
  1141 => x"b73fffab",
  1142 => x"3981b388",
  1143 => x"5180d5ac",
  1144 => x"3fffa039",
  1145 => x"81b39451",
  1146 => x"80d5a13f",
  1147 => x"ff9539fe",
  1148 => x"3d0d8151",
  1149 => x"aaec3fb0",
  1150 => x"0881ff06",
  1151 => x"81cebc08",
  1152 => x"71b4120c",
  1153 => x"53b00c84",
  1154 => x"3d0d04fe",
  1155 => x"3d0d880a",
  1156 => x"53840a0b",
  1157 => x"81ceb808",
  1158 => x"8c110851",
  1159 => x"52528071",
  1160 => x"27953880",
  1161 => x"73708405",
  1162 => x"550c8072",
  1163 => x"70840554",
  1164 => x"0cff1151",
  1165 => x"70ed3880",
  1166 => x"0bb00c84",
  1167 => x"3d0d04fa",
  1168 => x"3d0d880a",
  1169 => x"57840a56",
  1170 => x"8151aa96",
  1171 => x"3fb00883",
  1172 => x"ffff0654",
  1173 => x"73833890",
  1174 => x"54805574",
  1175 => x"742781c2",
  1176 => x"38750870",
  1177 => x"902c5253",
  1178 => x"80d5eb3f",
  1179 => x"b00881ff",
  1180 => x"0652718a",
  1181 => x"279438a0",
  1182 => x"5180d3f6",
  1183 => x"3f811270",
  1184 => x"81ff0651",
  1185 => x"528a7226",
  1186 => x"ee387290",
  1187 => x"2b70902c",
  1188 => x"525280d5",
  1189 => x"c13fb008",
  1190 => x"81ff0652",
  1191 => x"718a2794",
  1192 => x"38a05180",
  1193 => x"d3cc3f81",
  1194 => x"127081ff",
  1195 => x"0653538a",
  1196 => x"7226ee38",
  1197 => x"76087090",
  1198 => x"2c525380",
  1199 => x"d5983fb0",
  1200 => x"0881ff06",
  1201 => x"52718a27",
  1202 => x"9438a051",
  1203 => x"80d3a33f",
  1204 => x"81127081",
  1205 => x"ff065152",
  1206 => x"8a7226ee",
  1207 => x"3872902b",
  1208 => x"70902c52",
  1209 => x"5280d4ee",
  1210 => x"3fb00881",
  1211 => x"ff065271",
  1212 => x"8a279438",
  1213 => x"a05180d2",
  1214 => x"f93f8112",
  1215 => x"7081ff06",
  1216 => x"53538a72",
  1217 => x"26ee388a",
  1218 => x"5180d2e6",
  1219 => x"3f841784",
  1220 => x"17811770",
  1221 => x"83ffff06",
  1222 => x"58545757",
  1223 => x"737526fe",
  1224 => x"c03873b0",
  1225 => x"0c883d0d",
  1226 => x"04fd3d0d",
  1227 => x"8151a8b2",
  1228 => x"3fb00881",
  1229 => x"ff065473",
  1230 => x"802ea438",
  1231 => x"73842690",
  1232 => x"3881ceb8",
  1233 => x"0874710c",
  1234 => x"5373b00c",
  1235 => x"853d0d04",
  1236 => x"81ceb808",
  1237 => x"5380730c",
  1238 => x"73b00c85",
  1239 => x"3d0d0481",
  1240 => x"b4a05180",
  1241 => x"d2a63f81",
  1242 => x"b4b05180",
  1243 => x"d29e3f81",
  1244 => x"ceb80870",
  1245 => x"08525380",
  1246 => x"d3dc3f81",
  1247 => x"b4c05180",
  1248 => x"d28a3f81",
  1249 => x"ceb80884",
  1250 => x"11085353",
  1251 => x"a05180d2",
  1252 => x"9e3f81b4",
  1253 => x"d45180d1",
  1254 => x"f33f81ce",
  1255 => x"b8088811",
  1256 => x"085353a0",
  1257 => x"5180d287",
  1258 => x"3f81b4e8",
  1259 => x"5180d1dc",
  1260 => x"3f81ceb8",
  1261 => x"088c1108",
  1262 => x"525380d3",
  1263 => x"993f8a51",
  1264 => x"80d1af3f",
  1265 => x"73b00c85",
  1266 => x"3d0d04bc",
  1267 => x"0802bc0c",
  1268 => x"f93d0d02",
  1269 => x"bc08fc05",
  1270 => x"0c880a0b",
  1271 => x"bc08f405",
  1272 => x"0cfc3d0d",
  1273 => x"823dbc08",
  1274 => x"f0050c81",
  1275 => x"51a6f33f",
  1276 => x"b00881ff",
  1277 => x"06bc08f8",
  1278 => x"050c8251",
  1279 => x"a6e43fb0",
  1280 => x"08bc08f0",
  1281 => x"05082383",
  1282 => x"51a6d73f",
  1283 => x"b008bc08",
  1284 => x"f0050882",
  1285 => x"05238451",
  1286 => x"a6c83fb0",
  1287 => x"08bc08f0",
  1288 => x"05088405",
  1289 => x"238551a6",
  1290 => x"b93fb008",
  1291 => x"bc08f005",
  1292 => x"08860523",
  1293 => x"8651a6aa",
  1294 => x"3fb008bc",
  1295 => x"08f00508",
  1296 => x"88052387",
  1297 => x"51a69b3f",
  1298 => x"b008bc08",
  1299 => x"f005088a",
  1300 => x"05238851",
  1301 => x"a68c3fb0",
  1302 => x"08bc08f0",
  1303 => x"05088c05",
  1304 => x"238951a5",
  1305 => x"fd3fb008",
  1306 => x"bc08f005",
  1307 => x"088e0523",
  1308 => x"800b81ce",
  1309 => x"b808708c",
  1310 => x"050851bc",
  1311 => x"08e4050c",
  1312 => x"bc08ec05",
  1313 => x"0cbc08ec",
  1314 => x"0508bc08",
  1315 => x"e4050827",
  1316 => x"818f38bc",
  1317 => x"08e40508",
  1318 => x"bc08e805",
  1319 => x"0cbc08f8",
  1320 => x"0508802e",
  1321 => x"81b638bc",
  1322 => x"08ec0508",
  1323 => x"10bc08f0",
  1324 => x"05080570",
  1325 => x"22bc08f4",
  1326 => x"05088205",
  1327 => x"2271902b",
  1328 => x"07bc08f4",
  1329 => x"05080cbc",
  1330 => x"08e4050c",
  1331 => x"bc08f805",
  1332 => x"0cbc08ec",
  1333 => x"05088105",
  1334 => x"7081ff06",
  1335 => x"bc08e405",
  1336 => x"0cbc08f8",
  1337 => x"050c860b",
  1338 => x"bc08ec05",
  1339 => x"08278838",
  1340 => x"800bbc08",
  1341 => x"e4050cbc",
  1342 => x"08e40508",
  1343 => x"bc08f405",
  1344 => x"088405bc",
  1345 => x"08e80508",
  1346 => x"ff05bc08",
  1347 => x"e8050cbc",
  1348 => x"08f4050c",
  1349 => x"bc08ec05",
  1350 => x"0cbc08e8",
  1351 => x"0508ff87",
  1352 => x"38bc08fc",
  1353 => x"05080d80",
  1354 => x"0bb00c89",
  1355 => x"3d0dbc0c",
  1356 => x"04bc08e4",
  1357 => x"0508bc08",
  1358 => x"f4050884",
  1359 => x"05bc08e8",
  1360 => x"0508ff05",
  1361 => x"bc08e805",
  1362 => x"0cbc08f4",
  1363 => x"050cbc08",
  1364 => x"ec050cbc",
  1365 => x"08e80508",
  1366 => x"802ec638",
  1367 => x"bc08ec05",
  1368 => x"0810bc08",
  1369 => x"f0050805",
  1370 => x"70227090",
  1371 => x"2bbc08f4",
  1372 => x"050808fc",
  1373 => x"80800671",
  1374 => x"902c07bc",
  1375 => x"08f40508",
  1376 => x"0c52bc08",
  1377 => x"e4050cbc",
  1378 => x"08f8050c",
  1379 => x"800bbc08",
  1380 => x"e4050cbc",
  1381 => x"08ec0508",
  1382 => x"8626ff95",
  1383 => x"38bc08ec",
  1384 => x"05088105",
  1385 => x"7081ff06",
  1386 => x"bc08f405",
  1387 => x"088405bc",
  1388 => x"08e80508",
  1389 => x"ff05bc08",
  1390 => x"e8050cbc",
  1391 => x"08f4050c",
  1392 => x"bc08ec05",
  1393 => x"0cbc08e4",
  1394 => x"050cbc08",
  1395 => x"e80508ff",
  1396 => x"8b38fecd",
  1397 => x"39fb3d0d",
  1398 => x"029f0533",
  1399 => x"79982b70",
  1400 => x"982c5154",
  1401 => x"55810a54",
  1402 => x"805672e8",
  1403 => x"25bd38e8",
  1404 => x"53751081",
  1405 => x"07738180",
  1406 => x"0a298180",
  1407 => x"0a057098",
  1408 => x"2c515456",
  1409 => x"807324e9",
  1410 => x"38807325",
  1411 => x"80c73873",
  1412 => x"812a810a",
  1413 => x"07738180",
  1414 => x"0a2981ff",
  1415 => x"0a057098",
  1416 => x"2c515454",
  1417 => x"728024e7",
  1418 => x"38ab3997",
  1419 => x"73259a38",
  1420 => x"9774812a",
  1421 => x"810a0771",
  1422 => x"81800a29",
  1423 => x"81ff0a05",
  1424 => x"70982c51",
  1425 => x"525553dc",
  1426 => x"39807324",
  1427 => x"ffa33872",
  1428 => x"8024ffbb",
  1429 => x"38745280",
  1430 => x"51b3af3f",
  1431 => x"7381ff06",
  1432 => x"51b4ad3f",
  1433 => x"74528151",
  1434 => x"b3a03f73",
  1435 => x"882a7081",
  1436 => x"ff065253",
  1437 => x"b49a3f74",
  1438 => x"528251b3",
  1439 => x"8d3f7390",
  1440 => x"2a7081ff",
  1441 => x"065253b4",
  1442 => x"873f7452",
  1443 => x"8351b2fa",
  1444 => x"3f73982a",
  1445 => x"51b3f93f",
  1446 => x"74528451",
  1447 => x"b2ec3f75",
  1448 => x"81ff0651",
  1449 => x"b3ea3f74",
  1450 => x"528551b2",
  1451 => x"dd3f7588",
  1452 => x"2a7081ff",
  1453 => x"065253b3",
  1454 => x"d73f7452",
  1455 => x"8651b2ca",
  1456 => x"3f75902a",
  1457 => x"7081ff06",
  1458 => x"5254b3c4",
  1459 => x"3f745287",
  1460 => x"51b2b73f",
  1461 => x"75982a51",
  1462 => x"b3b63f87",
  1463 => x"3d0d04f2",
  1464 => x"3d0d0280",
  1465 => x"c3053302",
  1466 => x"840580c7",
  1467 => x"05338180",
  1468 => x"0a712b98",
  1469 => x"2a81ceb8",
  1470 => x"088c1108",
  1471 => x"71084453",
  1472 => x"565c5557",
  1473 => x"80730c80",
  1474 => x"7071725c",
  1475 => x"5a5e5b80",
  1476 => x"56757a27",
  1477 => x"80d73881",
  1478 => x"772783ce",
  1479 => x"387783ff",
  1480 => x"ff068119",
  1481 => x"71101084",
  1482 => x"0a057930",
  1483 => x"7a823270",
  1484 => x"30728025",
  1485 => x"71802507",
  1486 => x"56585841",
  1487 => x"57595c7b",
  1488 => x"802e83d5",
  1489 => x"38821522",
  1490 => x"5372902b",
  1491 => x"70902c54",
  1492 => x"55727b25",
  1493 => x"8338725b",
  1494 => x"7c732583",
  1495 => x"38725d81",
  1496 => x"167081ff",
  1497 => x"06575e79",
  1498 => x"7626ffb1",
  1499 => x"38811970",
  1500 => x"81ff065a",
  1501 => x"5680e579",
  1502 => x"27ff9438",
  1503 => x"987d3590",
  1504 => x"2b70902c",
  1505 => x"7c309871",
  1506 => x"35902b70",
  1507 => x"902c5c5c",
  1508 => x"55565477",
  1509 => x"54777525",
  1510 => x"83387454",
  1511 => x"73902b70",
  1512 => x"902c5d55",
  1513 => x"7b54807c",
  1514 => x"2583d738",
  1515 => x"73902b70",
  1516 => x"902c5f56",
  1517 => x"80705d58",
  1518 => x"80705a56",
  1519 => x"757a2780",
  1520 => x"e4388177",
  1521 => x"27838c38",
  1522 => x"7783ffff",
  1523 => x"06811971",
  1524 => x"1010840a",
  1525 => x"0579307a",
  1526 => x"82327030",
  1527 => x"72802571",
  1528 => x"80250753",
  1529 => x"51575357",
  1530 => x"59547380",
  1531 => x"2e83a438",
  1532 => x"82152254",
  1533 => x"73902b70",
  1534 => x"902c719f",
  1535 => x"2c707232",
  1536 => x"7131799f",
  1537 => x"2c707b32",
  1538 => x"71315154",
  1539 => x"51565653",
  1540 => x"72742583",
  1541 => x"38745681",
  1542 => x"197081ff",
  1543 => x"065a5579",
  1544 => x"7926ffa4",
  1545 => x"387d7635",
  1546 => x"982b7098",
  1547 => x"2c53547b",
  1548 => x"51fba23f",
  1549 => x"811c7081",
  1550 => x"ff065d59",
  1551 => x"80e57c27",
  1552 => x"fef63881",
  1553 => x"ceb8087f",
  1554 => x"710c5880",
  1555 => x"5281c394",
  1556 => x"51b3ad3f",
  1557 => x"81f2d408",
  1558 => x"80f5c40b",
  1559 => x"81f2d40c",
  1560 => x"5f805280",
  1561 => x"51afa33f",
  1562 => x"81b4f851",
  1563 => x"80c89d3f",
  1564 => x"7c5180c9",
  1565 => x"e13f8052",
  1566 => x"8751af8e",
  1567 => x"3f81b580",
  1568 => x"5180c888",
  1569 => x"3f7a5180",
  1570 => x"c9cc3f80",
  1571 => x"d2528051",
  1572 => x"aef83f81",
  1573 => x"b5885180",
  1574 => x"c7f23f76",
  1575 => x"5180c9b6",
  1576 => x"3f80c052",
  1577 => x"8751aee2",
  1578 => x"3f81b590",
  1579 => x"5180c7dc",
  1580 => x"3f7980e6",
  1581 => x"295180c9",
  1582 => x"9d3f7e81",
  1583 => x"f2d40c90",
  1584 => x"3d0d0474",
  1585 => x"22537290",
  1586 => x"2b70902c",
  1587 => x"545c727b",
  1588 => x"25833872",
  1589 => x"5b7c7325",
  1590 => x"8338725d",
  1591 => x"81167081",
  1592 => x"ff06575e",
  1593 => x"757a27fd",
  1594 => x"84387783",
  1595 => x"ffff0681",
  1596 => x"19711010",
  1597 => x"880a0579",
  1598 => x"307a8232",
  1599 => x"70307280",
  1600 => x"25718025",
  1601 => x"07565840",
  1602 => x"41575954",
  1603 => x"73802eff",
  1604 => x"b2388215",
  1605 => x"2253ffae",
  1606 => x"39742253",
  1607 => x"fcab3974",
  1608 => x"22547390",
  1609 => x"2b70902c",
  1610 => x"719f2c70",
  1611 => x"72327131",
  1612 => x"799f2c70",
  1613 => x"7b327131",
  1614 => x"51545156",
  1615 => x"56537274",
  1616 => x"25833874",
  1617 => x"56811970",
  1618 => x"81ff065a",
  1619 => x"55787a27",
  1620 => x"fdd33877",
  1621 => x"83ffff06",
  1622 => x"81197110",
  1623 => x"10880a05",
  1624 => x"79307a82",
  1625 => x"32703072",
  1626 => x"80257180",
  1627 => x"25075351",
  1628 => x"57535759",
  1629 => x"5473802e",
  1630 => x"ffa53882",
  1631 => x"152254ff",
  1632 => x"a1398170",
  1633 => x"902b7090",
  1634 => x"2c405754",
  1635 => x"80705d58",
  1636 => x"fca63974",
  1637 => x"2254fcdc",
  1638 => x"39fa3d0d",
  1639 => x"8a5180c5",
  1640 => x"d13f97b9",
  1641 => x"3f9a8553",
  1642 => x"81b59852",
  1643 => x"81b5ac51",
  1644 => x"97be3fa3",
  1645 => x"ef5381b5",
  1646 => x"b05281b5",
  1647 => x"d85197b0",
  1648 => x"3fbbeb53",
  1649 => x"81b5e052",
  1650 => x"81b5f051",
  1651 => x"97a23fbb",
  1652 => x"d25381b5",
  1653 => x"f85281b6",
  1654 => x"94519794",
  1655 => x"3fa6a953",
  1656 => x"81b69c52",
  1657 => x"81b6c051",
  1658 => x"97863fbe",
  1659 => x"ae5381b6",
  1660 => x"c85281b6",
  1661 => x"e85196f8",
  1662 => x"3fbfcc53",
  1663 => x"81b6ec52",
  1664 => x"81b79051",
  1665 => x"96ea3fbc",
  1666 => x"825381b7",
  1667 => x"985281b2",
  1668 => x"b05196dc",
  1669 => x"3fbcc353",
  1670 => x"81b7bc52",
  1671 => x"81b7e451",
  1672 => x"96ce3fbd",
  1673 => x"eb5381b7",
  1674 => x"ec5281b8",
  1675 => x"8c5196c0",
  1676 => x"3f889b53",
  1677 => x"81b89452",
  1678 => x"81b8b051",
  1679 => x"96b23fa4",
  1680 => x"bf5381b8",
  1681 => x"b85281b8",
  1682 => x"845196a4",
  1683 => x"3fa48b53",
  1684 => x"81b8d452",
  1685 => x"81b8e851",
  1686 => x"96963fb9",
  1687 => x"905381b8",
  1688 => x"f05281b9",
  1689 => x"8c519688",
  1690 => x"3fb9b653",
  1691 => x"81b99452",
  1692 => x"81b9a851",
  1693 => x"95fa3fa7",
  1694 => x"cb5381b9",
  1695 => x"b05281b9",
  1696 => x"d45195ec",
  1697 => x"3f80c0aa",
  1698 => x"5381b9dc",
  1699 => x"5281b9ec",
  1700 => x"5195dd3f",
  1701 => x"80c2f553",
  1702 => x"81b9f052",
  1703 => x"81ba8c51",
  1704 => x"95ce3fbb",
  1705 => x"985381ba",
  1706 => x"945281ba",
  1707 => x"ac5195c0",
  1708 => x"3f80c2fd",
  1709 => x"5381bab4",
  1710 => x"5281bac8",
  1711 => x"5195b13f",
  1712 => x"8ad65381",
  1713 => x"bad05281",
  1714 => x"bae45195",
  1715 => x"a33f8de6",
  1716 => x"5381bae8",
  1717 => x"5281bb90",
  1718 => x"5195953f",
  1719 => x"bbb45381",
  1720 => x"bb985281",
  1721 => x"bbb85195",
  1722 => x"873f93a3",
  1723 => x"5381bbc0",
  1724 => x"5281bbd4",
  1725 => x"5194f93f",
  1726 => x"88be5381",
  1727 => x"bbdc5281",
  1728 => x"bbe85194",
  1729 => x"eb3f89fc",
  1730 => x"5381bbec",
  1731 => x"5281bc94",
  1732 => x"5194dd3f",
  1733 => x"88be5381",
  1734 => x"bc9c5281",
  1735 => x"b4d05194",
  1736 => x"cf3f8ac5",
  1737 => x"5381bcac",
  1738 => x"5281bcbc",
  1739 => x"5194c13f",
  1740 => x"88b35381",
  1741 => x"a7dc5281",
  1742 => x"a7c05194",
  1743 => x"b33f80d1",
  1744 => x"c65381a7",
  1745 => x"dc5281a7",
  1746 => x"c85194a4",
  1747 => x"3f9af73f",
  1748 => x"94ea3f81",
  1749 => x"0b81f1f0",
  1750 => x"3481ded0",
  1751 => x"337081ff",
  1752 => x"06555573",
  1753 => x"b23880c6",
  1754 => x"953fb008",
  1755 => x"903894da",
  1756 => x"3f81f1f0",
  1757 => x"335675e1",
  1758 => x"38883d0d",
  1759 => x"0480c691",
  1760 => x"3fb00881",
  1761 => x"ff065195",
  1762 => x"af3f94be",
  1763 => x"3f81f1f0",
  1764 => x"335675c5",
  1765 => x"38e33980",
  1766 => x"0b81ded0",
  1767 => x"349bc73f",
  1768 => x"81cef408",
  1769 => x"70087087",
  1770 => x"2a810652",
  1771 => x"57547380",
  1772 => x"2e8f3876",
  1773 => x"802e81c5",
  1774 => x"38ff1770",
  1775 => x"81ff0658",
  1776 => x"5475862a",
  1777 => x"81065574",
  1778 => x"802eaa38",
  1779 => x"7680f738",
  1780 => x"81960b81",
  1781 => x"cef40884",
  1782 => x"110870ef",
  1783 => x"ff0a06ae",
  1784 => x"800a0784",
  1785 => x"130c5784",
  1786 => x"110870be",
  1787 => x"800a0784",
  1788 => x"130c5755",
  1789 => x"5775852a",
  1790 => x"81065574",
  1791 => x"802e9638",
  1792 => x"76ba3881",
  1793 => x"960b81ce",
  1794 => x"bc08b811",
  1795 => x"08575557",
  1796 => x"800bb815",
  1797 => x"0c75842a",
  1798 => x"81065675",
  1799 => x"802efec6",
  1800 => x"3876802e",
  1801 => x"ac38ff17",
  1802 => x"7081ff06",
  1803 => x"585580c4",
  1804 => x"cd3fb008",
  1805 => x"802efeb6",
  1806 => x"38fec239",
  1807 => x"ff177081",
  1808 => x"ff065855",
  1809 => x"d039ff17",
  1810 => x"7081ff06",
  1811 => x"5854ffa5",
  1812 => x"3981960b",
  1813 => x"81cef408",
  1814 => x"84110884",
  1815 => x"0a078412",
  1816 => x"0c5657a8",
  1817 => x"c83f8052",
  1818 => x"81c39451",
  1819 => x"ab923f80",
  1820 => x"c48c3fb0",
  1821 => x"08802efd",
  1822 => x"f538fe81",
  1823 => x"39819676",
  1824 => x"822a8306",
  1825 => x"53768306",
  1826 => x"5257f4d3",
  1827 => x"3ffeb239",
  1828 => x"fe3d0d81",
  1829 => x"5195cb3f",
  1830 => x"b00881ff",
  1831 => x"06538251",
  1832 => x"95c03fb0",
  1833 => x"0881ff06",
  1834 => x"527251f4",
  1835 => x"b23f800b",
  1836 => x"b00c843d",
  1837 => x"0d04f93d",
  1838 => x"0d815195",
  1839 => x"a53fb008",
  1840 => x"81ff0681",
  1841 => x"bcc45257",
  1842 => x"bfc23f81",
  1843 => x"bcd851bf",
  1844 => x"bb3ff880",
  1845 => x"809a8054",
  1846 => x"80557370",
  1847 => x"84055508",
  1848 => x"74708405",
  1849 => x"56085456",
  1850 => x"72a03881",
  1851 => x"157081ff",
  1852 => x"06565687",
  1853 => x"7527e338",
  1854 => x"76812e80",
  1855 => x"d9388a51",
  1856 => x"bef03f76",
  1857 => x"b00c893d",
  1858 => x"0d048a51",
  1859 => x"bee43f72",
  1860 => x"5180c0c2",
  1861 => x"3fb00881",
  1862 => x"ff065372",
  1863 => x"8c279338",
  1864 => x"a051bece",
  1865 => x"3f811370",
  1866 => x"81ff0651",
  1867 => x"538c7326",
  1868 => x"ef3881bc",
  1869 => x"f051bed4",
  1870 => x"3f7552a0",
  1871 => x"51bef03f",
  1872 => x"7551d9c1",
  1873 => x"3f811570",
  1874 => x"81ff0656",
  1875 => x"56877527",
  1876 => x"ff8838ff",
  1877 => x"a339f880",
  1878 => x"809a8054",
  1879 => x"80538074",
  1880 => x"70840556",
  1881 => x"0c807470",
  1882 => x"8405560c",
  1883 => x"81137081",
  1884 => x"ff065455",
  1885 => x"728726ff",
  1886 => x"85388074",
  1887 => x"70840556",
  1888 => x"0c807470",
  1889 => x"8405560c",
  1890 => x"81137081",
  1891 => x"ff065455",
  1892 => x"877327ca",
  1893 => x"38fee739",
  1894 => x"fe3d0d81",
  1895 => x"5193c33f",
  1896 => x"b00881ff",
  1897 => x"0681ceb4",
  1898 => x"08718812",
  1899 => x"0c53b00c",
  1900 => x"843d0d04",
  1901 => x"803d0d81",
  1902 => x"5194d93f",
  1903 => x"b00883ff",
  1904 => x"ff0651d2",
  1905 => x"ee3fb008",
  1906 => x"83ffff06",
  1907 => x"b00c823d",
  1908 => x"0d04803d",
  1909 => x"0d815193",
  1910 => x"893fb008",
  1911 => x"81ff0651",
  1912 => x"9e863f80",
  1913 => x"0bb00c82",
  1914 => x"3d0d0480",
  1915 => x"3d0d81cf",
  1916 => x"800851f8",
  1917 => x"bb9586a1",
  1918 => x"710c810b",
  1919 => x"b00c823d",
  1920 => x"0d04fc3d",
  1921 => x"0d815192",
  1922 => x"d93fb008",
  1923 => x"81ff0654",
  1924 => x"825192ce",
  1925 => x"3fb00881",
  1926 => x"ff0681ce",
  1927 => x"f4088411",
  1928 => x"0870fe8f",
  1929 => x"0a067798",
  1930 => x"2b075154",
  1931 => x"56537280",
  1932 => x"2e863871",
  1933 => x"810a0752",
  1934 => x"7184160c",
  1935 => x"71b00c86",
  1936 => x"3d0d04fd",
  1937 => x"3d0d81ce",
  1938 => x"f4088411",
  1939 => x"08555381",
  1940 => x"51928f3f",
  1941 => x"b00881ff",
  1942 => x"0674dfff",
  1943 => x"ff065452",
  1944 => x"71802e87",
  1945 => x"3873a080",
  1946 => x"80075382",
  1947 => x"5191f33f",
  1948 => x"b00881ff",
  1949 => x"0673efff",
  1950 => x"0a065552",
  1951 => x"71802e87",
  1952 => x"38729080",
  1953 => x"0a075483",
  1954 => x"5191d73f",
  1955 => x"b00881ff",
  1956 => x"0674f7ff",
  1957 => x"0a065452",
  1958 => x"71802e87",
  1959 => x"38738880",
  1960 => x"0a075384",
  1961 => x"5191bb3f",
  1962 => x"b00881ff",
  1963 => x"0673fbff",
  1964 => x"0a065552",
  1965 => x"71802e87",
  1966 => x"38728480",
  1967 => x"0a075485",
  1968 => x"51919f3f",
  1969 => x"b00881ff",
  1970 => x"0674fdff",
  1971 => x"0a065452",
  1972 => x"71802e87",
  1973 => x"38738280",
  1974 => x"0a075381",
  1975 => x"cef40873",
  1976 => x"84120c54",
  1977 => x"72b00c85",
  1978 => x"3d0d04fa",
  1979 => x"3d0d880a",
  1980 => x"0b81ceb8",
  1981 => x"088c1108",
  1982 => x"59555681",
  1983 => x"5190e33f",
  1984 => x"b008902b",
  1985 => x"70902c56",
  1986 => x"53807727",
  1987 => x"99388077",
  1988 => x"54547383",
  1989 => x"ffff0676",
  1990 => x"70840558",
  1991 => x"0cff1375",
  1992 => x"15555372",
  1993 => x"ed38800b",
  1994 => x"b00c883d",
  1995 => x"0d04fc3d",
  1996 => x"0d81bcf8",
  1997 => x"51bad53f",
  1998 => x"81cef408",
  1999 => x"7008709e",
  2000 => x"2a708106",
  2001 => x"51545454",
  2002 => x"81537183",
  2003 => x"38715372",
  2004 => x"802e80d2",
  2005 => x"3881bd88",
  2006 => x"51bab13f",
  2007 => x"81519082",
  2008 => x"3fb00881",
  2009 => x"ff0681bc",
  2010 => x"f85255ba",
  2011 => x"9f3f7480",
  2012 => x"2eab3881",
  2013 => x"bd9051ba",
  2014 => x"933f81ce",
  2015 => x"f4088411",
  2016 => x"0870fd0a",
  2017 => x"06545454",
  2018 => x"74802e86",
  2019 => x"3872820a",
  2020 => x"07527184",
  2021 => x"150c71b0",
  2022 => x"0c863d0d",
  2023 => x"0481b2b8",
  2024 => x"51b9e93f",
  2025 => x"ce3981b2",
  2026 => x"b851b9e0",
  2027 => x"3f81bd88",
  2028 => x"51b9d93f",
  2029 => x"81518faa",
  2030 => x"3fb00881",
  2031 => x"ff0681bc",
  2032 => x"f85255b9",
  2033 => x"c73f74ff",
  2034 => x"aa38d239",
  2035 => x"fd3d0d81",
  2036 => x"518f8f3f",
  2037 => x"b00881ff",
  2038 => x"0681bd9c",
  2039 => x"5254b9ac",
  2040 => x"3f73a438",
  2041 => x"81b2b051",
  2042 => x"b9a23f81",
  2043 => x"cef40884",
  2044 => x"110870fb",
  2045 => x"0a068413",
  2046 => x"0c53538a",
  2047 => x"51b8f33f",
  2048 => x"73b00c85",
  2049 => x"3d0d0481",
  2050 => x"aed851b8",
  2051 => x"ff3f81ce",
  2052 => x"f4088411",
  2053 => x"0870840a",
  2054 => x"0784130c",
  2055 => x"53538a51",
  2056 => x"b8d03f73",
  2057 => x"b00c853d",
  2058 => x"0d04fd3d",
  2059 => x"0d81decc",
  2060 => x"0852f881",
  2061 => x"c08e800b",
  2062 => x"81cef408",
  2063 => x"55537180",
  2064 => x"2e80f738",
  2065 => x"7281ff06",
  2066 => x"84150c81",
  2067 => x"ceb03370",
  2068 => x"81ff0651",
  2069 => x"5271802e",
  2070 => x"80c23872",
  2071 => x"9f2a7310",
  2072 => x"075381de",
  2073 => x"d0337081",
  2074 => x"ff065152",
  2075 => x"71802ed4",
  2076 => x"38800b81",
  2077 => x"ded03491",
  2078 => x"ed3f81ce",
  2079 => x"c0335473",
  2080 => x"80e23881",
  2081 => x"cef40873",
  2082 => x"81ff0684",
  2083 => x"120c81ce",
  2084 => x"b0337081",
  2085 => x"ff065153",
  2086 => x"5471c038",
  2087 => x"72812a73",
  2088 => x"9f2b0753",
  2089 => x"ffbc3972",
  2090 => x"812a739f",
  2091 => x"2b075380",
  2092 => x"fd51baeb",
  2093 => x"3f81cef4",
  2094 => x"08547281",
  2095 => x"ff068415",
  2096 => x"0c81ceb0",
  2097 => x"337081ff",
  2098 => x"06535471",
  2099 => x"802ed838",
  2100 => x"729f2a73",
  2101 => x"10075380",
  2102 => x"fd51bac3",
  2103 => x"3f81cef4",
  2104 => x"0854d739",
  2105 => x"800bb00c",
  2106 => x"853d0d04",
  2107 => x"f73d0d85",
  2108 => x"3d549653",
  2109 => x"81bdb052",
  2110 => x"7351be85",
  2111 => x"3fa09f3f",
  2112 => x"81518cde",
  2113 => x"3f805280",
  2114 => x"519dff3f",
  2115 => x"73538052",
  2116 => x"81c39451",
  2117 => x"b2be3f80",
  2118 => x"5281519d",
  2119 => x"ed3f7353",
  2120 => x"825281c3",
  2121 => x"9451b2ac",
  2122 => x"3f805282",
  2123 => x"519ddb3f",
  2124 => x"73538152",
  2125 => x"81c39451",
  2126 => x"b29a3f80",
  2127 => x"5284519d",
  2128 => x"c93f7353",
  2129 => x"845281c3",
  2130 => x"9451b288",
  2131 => x"3f805285",
  2132 => x"519db73f",
  2133 => x"73539052",
  2134 => x"81c39451",
  2135 => x"b1f63f80",
  2136 => x"5286519d",
  2137 => x"a53f7353",
  2138 => x"835281c3",
  2139 => x"9451b1e4",
  2140 => x"3f8b3d0d",
  2141 => x"04fef53f",
  2142 => x"800bb00c",
  2143 => x"04fc3d0d",
  2144 => x"81a1d854",
  2145 => x"80558452",
  2146 => x"74519cfe",
  2147 => x"3f805373",
  2148 => x"70810555",
  2149 => x"33519df8",
  2150 => x"3f811370",
  2151 => x"81ff0651",
  2152 => x"5380dc73",
  2153 => x"27e93881",
  2154 => x"157081ff",
  2155 => x"06565387",
  2156 => x"7527d338",
  2157 => x"800bb00c",
  2158 => x"863d0d04",
  2159 => x"fd3d0d81",
  2160 => x"ceb03370",
  2161 => x"81ff0654",
  2162 => x"5472bf26",
  2163 => x"ac3881ce",
  2164 => x"b0337081",
  2165 => x"ff0681ce",
  2166 => x"b4085288",
  2167 => x"120c5480",
  2168 => x"e45280c3",
  2169 => x"bc518fde",
  2170 => x"3f81ceb0",
  2171 => x"33810553",
  2172 => x"7281ceb0",
  2173 => x"34853d0d",
  2174 => x"0480e452",
  2175 => x"80c49351",
  2176 => x"8fc43f81",
  2177 => x"ceb03381",
  2178 => x"05537281",
  2179 => x"ceb03485",
  2180 => x"3d0d04fd",
  2181 => x"3d0d81ce",
  2182 => x"b0337081",
  2183 => x"ff065454",
  2184 => x"72bf2680",
  2185 => x"c93881ce",
  2186 => x"b0337081",
  2187 => x"ff0681ce",
  2188 => x"b4085688",
  2189 => x"160c5381",
  2190 => x"ceb03370",
  2191 => x"81ff0655",
  2192 => x"5373bf2e",
  2193 => x"80d13880",
  2194 => x"e45280c4",
  2195 => x"93518ef6",
  2196 => x"3f81ceb0",
  2197 => x"33810553",
  2198 => x"7281ceb0",
  2199 => x"3481ceb0",
  2200 => x"3380ff06",
  2201 => x"537281ce",
  2202 => x"b034853d",
  2203 => x"0d0481ce",
  2204 => x"b0337081",
  2205 => x"ff0680ff",
  2206 => x"713181ce",
  2207 => x"b4085288",
  2208 => x"120c5553",
  2209 => x"81ceb033",
  2210 => x"7081ff06",
  2211 => x"555373bf",
  2212 => x"2e098106",
  2213 => x"ffb13880",
  2214 => x"ce905280",
  2215 => x"c493518e",
  2216 => x"a53f81ce",
  2217 => x"b0338105",
  2218 => x"537281ce",
  2219 => x"b03481ce",
  2220 => x"b03380ff",
  2221 => x"06537281",
  2222 => x"ceb03485",
  2223 => x"3d0d0481",
  2224 => x"0b81cec0",
  2225 => x"3404fe3d",
  2226 => x"0d81cef8",
  2227 => x"08981108",
  2228 => x"70842a70",
  2229 => x"81065153",
  2230 => x"53537080",
  2231 => x"2e8d3871",
  2232 => x"ef069814",
  2233 => x"0c810b81",
  2234 => x"ded03484",
  2235 => x"3d0d04fb",
  2236 => x"3d0d81ce",
  2237 => x"f4087008",
  2238 => x"810a0681",
  2239 => x"decc0c54",
  2240 => x"b6c03fb6",
  2241 => x"e33f8efb",
  2242 => x"3f81cef8",
  2243 => x"08981108",
  2244 => x"88079812",
  2245 => x"0c5481de",
  2246 => x"cc0880f8",
  2247 => x"dc555372",
  2248 => x"84388880",
  2249 => x"547381f2",
  2250 => x"d40c7280",
  2251 => x"2e849a38",
  2252 => x"81a8a451",
  2253 => x"b2d63f8c",
  2254 => x"51b2b73f",
  2255 => x"81bdb051",
  2256 => x"b2ca3f81",
  2257 => x"decc0880",
  2258 => x"2e81d238",
  2259 => x"81bdc851",
  2260 => x"b2ba3f81",
  2261 => x"decc0854",
  2262 => x"73802e82",
  2263 => x"bd3881ce",
  2264 => x"b8085481",
  2265 => x"740c81ce",
  2266 => x"f4088411",
  2267 => x"08705657",
  2268 => x"55805373",
  2269 => x"fe8f0a06",
  2270 => x"73982b07",
  2271 => x"7084170c",
  2272 => x"81147081",
  2273 => x"ff065154",
  2274 => x"548f7327",
  2275 => x"e6387584",
  2276 => x"160c81ce",
  2277 => x"bc085480",
  2278 => x"0bb8150c",
  2279 => x"825280c5",
  2280 => x"bf518ca2",
  2281 => x"3ff881c0",
  2282 => x"8e800b81",
  2283 => x"cef40856",
  2284 => x"5481decc",
  2285 => x"08802e81",
  2286 => x"b7387381",
  2287 => x"ff068416",
  2288 => x"0c81ceb0",
  2289 => x"337081ff",
  2290 => x"06545672",
  2291 => x"802e80c2",
  2292 => x"38739f2a",
  2293 => x"74100754",
  2294 => x"81ded033",
  2295 => x"7081ff06",
  2296 => x"57537580",
  2297 => x"2ed43880",
  2298 => x"0b81ded0",
  2299 => x"348af73f",
  2300 => x"81cec033",
  2301 => x"557482e2",
  2302 => x"3881cef4",
  2303 => x"087481ff",
  2304 => x"0684120c",
  2305 => x"81ceb033",
  2306 => x"7081ff06",
  2307 => x"55575572",
  2308 => x"c0387381",
  2309 => x"2a749f2b",
  2310 => x"0754ffbc",
  2311 => x"3981bdd4",
  2312 => x"51b0e93f",
  2313 => x"810a51b0",
  2314 => x"e33f81bd",
  2315 => x"e851b0dc",
  2316 => x"3f81be90",
  2317 => x"51b0d53f",
  2318 => x"b451b29a",
  2319 => x"3f81bea4",
  2320 => x"51b0c93f",
  2321 => x"81beac51",
  2322 => x"b0c23f81",
  2323 => x"beb851b0",
  2324 => x"bb3f81de",
  2325 => x"cc085473",
  2326 => x"fe8438be",
  2327 => x"3973812a",
  2328 => x"749f2b07",
  2329 => x"5480fd51",
  2330 => x"b3b53f81",
  2331 => x"cef40855",
  2332 => x"7381ff06",
  2333 => x"84160c81",
  2334 => x"ceb03370",
  2335 => x"81ff0656",
  2336 => x"5674802e",
  2337 => x"d838739f",
  2338 => x"2a741007",
  2339 => x"5480fd51",
  2340 => x"b38d3f81",
  2341 => x"cef40855",
  2342 => x"d73981ce",
  2343 => x"bc0874b4",
  2344 => x"120c5681",
  2345 => x"8051c58b",
  2346 => x"3f828051",
  2347 => x"c5853f84",
  2348 => x"8351c4ff",
  2349 => x"3f86f151",
  2350 => x"c4f93f88",
  2351 => x"8351c4f3",
  2352 => x"3f81cef4",
  2353 => x"08700870",
  2354 => x"9e2a7081",
  2355 => x"06515556",
  2356 => x"54815572",
  2357 => x"802e80fd",
  2358 => x"387481ff",
  2359 => x"06841508",
  2360 => x"70fd0a06",
  2361 => x"58565372",
  2362 => x"802e8638",
  2363 => x"74820a07",
  2364 => x"56758415",
  2365 => x"0c841408",
  2366 => x"be800a07",
  2367 => x"84150c84",
  2368 => x"1408840a",
  2369 => x"0784150c",
  2370 => x"81cebc08",
  2371 => x"55800bb8",
  2372 => x"160c81ce",
  2373 => x"b8085481",
  2374 => x"740c93c4",
  2375 => x"5280c2fd",
  2376 => x"5189a33f",
  2377 => x"87e85280",
  2378 => x"c3bc5189",
  2379 => x"993fe8e9",
  2380 => x"3f81ceb8",
  2381 => x"08548174",
  2382 => x"0c81cef4",
  2383 => x"08841108",
  2384 => x"70565755",
  2385 => x"8053fcab",
  2386 => x"39b3b83f",
  2387 => x"93c43f97",
  2388 => x"cd3ffbdc",
  2389 => x"397255ff",
  2390 => x"8039b598",
  2391 => x"3f800b81",
  2392 => x"f1e83480",
  2393 => x"0b81f1e4",
  2394 => x"34800b81",
  2395 => x"f1ec0c04",
  2396 => x"fc3d0d76",
  2397 => x"5281f1e4",
  2398 => x"33701010",
  2399 => x"10711005",
  2400 => x"81ded405",
  2401 => x"5254ba87",
  2402 => x"3f775281",
  2403 => x"f1e43370",
  2404 => x"90297131",
  2405 => x"70101081",
  2406 => x"e1940553",
  2407 => x"5555b9ef",
  2408 => x"3f81f1e4",
  2409 => x"33701010",
  2410 => x"81f09405",
  2411 => x"7a710c54",
  2412 => x"81055372",
  2413 => x"81f1e434",
  2414 => x"863d0d04",
  2415 => x"803d0d81",
  2416 => x"befc51ad",
  2417 => x"c73f823d",
  2418 => x"0d04fe3d",
  2419 => x"0d81f1ec",
  2420 => x"08537285",
  2421 => x"38843d0d",
  2422 => x"04722db0",
  2423 => x"0853800b",
  2424 => x"81f1ec0c",
  2425 => x"b0088c38",
  2426 => x"81befc51",
  2427 => x"ad9e3f84",
  2428 => x"3d0d0481",
  2429 => x"c2c051ad",
  2430 => x"933f7283",
  2431 => x"ffff26aa",
  2432 => x"3881ff73",
  2433 => x"27963872",
  2434 => x"529051ad",
  2435 => x"a23f8a51",
  2436 => x"ace03f81",
  2437 => x"befc51ac",
  2438 => x"f33fd439",
  2439 => x"72528851",
  2440 => x"ad8d3f8a",
  2441 => x"51accb3f",
  2442 => x"ea397252",
  2443 => x"a051acff",
  2444 => x"3f8a51ac",
  2445 => x"bd3fdc39",
  2446 => x"fa3d0d02",
  2447 => x"a3053356",
  2448 => x"758d2e80",
  2449 => x"f4387588",
  2450 => x"32703077",
  2451 => x"80ff3270",
  2452 => x"30728025",
  2453 => x"71802507",
  2454 => x"54515658",
  2455 => x"55749538",
  2456 => x"9f76278c",
  2457 => x"3881f1e8",
  2458 => x"335580ce",
  2459 => x"7527ae38",
  2460 => x"883d0d04",
  2461 => x"81f1e833",
  2462 => x"5675802e",
  2463 => x"f3388851",
  2464 => x"abf03fa0",
  2465 => x"51abeb3f",
  2466 => x"8851abe6",
  2467 => x"3f81f1e8",
  2468 => x"33ff0557",
  2469 => x"7681f1e8",
  2470 => x"34883d0d",
  2471 => x"047551ab",
  2472 => x"d13f81f1",
  2473 => x"e8338111",
  2474 => x"55577381",
  2475 => x"f1e83475",
  2476 => x"81f19418",
  2477 => x"34883d0d",
  2478 => x"048a51ab",
  2479 => x"b53f81f1",
  2480 => x"e8338111",
  2481 => x"56547481",
  2482 => x"f1e83480",
  2483 => x"0b81f194",
  2484 => x"15348056",
  2485 => x"800b81f1",
  2486 => x"94173356",
  2487 => x"5474a02e",
  2488 => x"83388154",
  2489 => x"74802e90",
  2490 => x"3873802e",
  2491 => x"8b388116",
  2492 => x"7081ff06",
  2493 => x"5757dd39",
  2494 => x"75802ebf",
  2495 => x"38800b81",
  2496 => x"f1e43355",
  2497 => x"55747427",
  2498 => x"ab387357",
  2499 => x"74101010",
  2500 => x"75100576",
  2501 => x"5481f194",
  2502 => x"5381ded4",
  2503 => x"0551b8bb",
  2504 => x"3fb00880",
  2505 => x"2ea63881",
  2506 => x"157081ff",
  2507 => x"06565476",
  2508 => x"7526d938",
  2509 => x"81bf8051",
  2510 => x"aad23f81",
  2511 => x"befc51aa",
  2512 => x"cb3f800b",
  2513 => x"81f1e834",
  2514 => x"883d0d04",
  2515 => x"74101081",
  2516 => x"f0940570",
  2517 => x"0881f1ec",
  2518 => x"0c56800b",
  2519 => x"81f1e834",
  2520 => x"e739f73d",
  2521 => x"0d02af05",
  2522 => x"3359800b",
  2523 => x"81f19433",
  2524 => x"81f19459",
  2525 => x"555673a0",
  2526 => x"2e098106",
  2527 => x"96388116",
  2528 => x"7081ff06",
  2529 => x"81f19411",
  2530 => x"70335359",
  2531 => x"575473a0",
  2532 => x"2eec3880",
  2533 => x"58777927",
  2534 => x"80ea3880",
  2535 => x"77335654",
  2536 => x"74742e83",
  2537 => x"38815474",
  2538 => x"a02e9a38",
  2539 => x"7380c538",
  2540 => x"74a02e91",
  2541 => x"38811870",
  2542 => x"81ff0659",
  2543 => x"55787826",
  2544 => x"da3880c0",
  2545 => x"39811670",
  2546 => x"81ff0681",
  2547 => x"f1941170",
  2548 => x"33575257",
  2549 => x"5773a02e",
  2550 => x"098106d9",
  2551 => x"38811670",
  2552 => x"81ff0681",
  2553 => x"f1941170",
  2554 => x"33575257",
  2555 => x"5773a02e",
  2556 => x"d438c239",
  2557 => x"81167081",
  2558 => x"ff0681f1",
  2559 => x"94115957",
  2560 => x"55ff9839",
  2561 => x"8a538b3d",
  2562 => x"fc055276",
  2563 => x"51bb913f",
  2564 => x"8b3d0d04",
  2565 => x"f73d0d02",
  2566 => x"af053359",
  2567 => x"800b81f1",
  2568 => x"943381f1",
  2569 => x"94595556",
  2570 => x"73a02e09",
  2571 => x"81069638",
  2572 => x"81167081",
  2573 => x"ff0681f1",
  2574 => x"94117033",
  2575 => x"53595754",
  2576 => x"73a02eec",
  2577 => x"38805877",
  2578 => x"792780ea",
  2579 => x"38807733",
  2580 => x"56547474",
  2581 => x"2e833881",
  2582 => x"5474a02e",
  2583 => x"9a387380",
  2584 => x"c53874a0",
  2585 => x"2e913881",
  2586 => x"187081ff",
  2587 => x"06595578",
  2588 => x"7826da38",
  2589 => x"80c03981",
  2590 => x"167081ff",
  2591 => x"0681f194",
  2592 => x"11703357",
  2593 => x"52575773",
  2594 => x"a02e0981",
  2595 => x"06d93881",
  2596 => x"167081ff",
  2597 => x"0681f194",
  2598 => x"11703357",
  2599 => x"52575773",
  2600 => x"a02ed438",
  2601 => x"c2398116",
  2602 => x"7081ff06",
  2603 => x"81f19411",
  2604 => x"595755ff",
  2605 => x"98399053",
  2606 => x"8b3dfc05",
  2607 => x"527651bc",
  2608 => x"fc3f8b3d",
  2609 => x"0d04fc3d",
  2610 => x"0d8a51a7",
  2611 => x"a53f81bf",
  2612 => x"9451a7b8",
  2613 => x"3f800b81",
  2614 => x"f1e43353",
  2615 => x"53727227",
  2616 => x"80f53872",
  2617 => x"10101073",
  2618 => x"100581de",
  2619 => x"d4057052",
  2620 => x"54a7993f",
  2621 => x"72842b70",
  2622 => x"7431822b",
  2623 => x"81e19411",
  2624 => x"33515355",
  2625 => x"71802eb7",
  2626 => x"387351b3",
  2627 => x"ef3fb008",
  2628 => x"81ff0652",
  2629 => x"71892693",
  2630 => x"38a051a6",
  2631 => x"d53f8112",
  2632 => x"7081ff06",
  2633 => x"53548972",
  2634 => x"27ef3881",
  2635 => x"bfac51a6",
  2636 => x"db3f7473",
  2637 => x"31822b81",
  2638 => x"e1940551",
  2639 => x"a6ce3f8a",
  2640 => x"51a6af3f",
  2641 => x"81137081",
  2642 => x"ff0681f1",
  2643 => x"e4335454",
  2644 => x"55717326",
  2645 => x"ff8d388a",
  2646 => x"51a6973f",
  2647 => x"81f1e433",
  2648 => x"b00c863d",
  2649 => x"0d04fe3d",
  2650 => x"0d81f2c4",
  2651 => x"22ff0551",
  2652 => x"7081f2c4",
  2653 => x"237083ff",
  2654 => x"ff065170",
  2655 => x"80c43881",
  2656 => x"f2c83351",
  2657 => x"7081ff2e",
  2658 => x"b9387010",
  2659 => x"101081f1",
  2660 => x"f4055271",
  2661 => x"3381f2c8",
  2662 => x"34fe7234",
  2663 => x"81f2c833",
  2664 => x"70101010",
  2665 => x"81f1f405",
  2666 => x"52538211",
  2667 => x"2281f2c4",
  2668 => x"23841208",
  2669 => x"53722d81",
  2670 => x"f2c42251",
  2671 => x"70802eff",
  2672 => x"be38843d",
  2673 => x"0d04f93d",
  2674 => x"0d02aa05",
  2675 => x"22568055",
  2676 => x"74101010",
  2677 => x"81f1f405",
  2678 => x"70335252",
  2679 => x"7081fe2e",
  2680 => x"99388115",
  2681 => x"7081ff06",
  2682 => x"5652748a",
  2683 => x"2e098106",
  2684 => x"df38810b",
  2685 => x"b00c893d",
  2686 => x"0d0481f2",
  2687 => x"c8337081",
  2688 => x"ff0681f2",
  2689 => x"c4225354",
  2690 => x"587281ff",
  2691 => x"2eb03872",
  2692 => x"832b5470",
  2693 => x"762780de",
  2694 => x"38757131",
  2695 => x"7083ffff",
  2696 => x"067481f1",
  2697 => x"f4173370",
  2698 => x"832b81f1",
  2699 => x"f6112256",
  2700 => x"58565257",
  2701 => x"577281ff",
  2702 => x"2e098106",
  2703 => x"d6387272",
  2704 => x"34758213",
  2705 => x"23798413",
  2706 => x"0c7781ff",
  2707 => x"06547373",
  2708 => x"2e963876",
  2709 => x"10101081",
  2710 => x"f1f40553",
  2711 => x"74733480",
  2712 => x"5170b00c",
  2713 => x"893d0d04",
  2714 => x"7481f2c8",
  2715 => x"347581f2",
  2716 => x"c4238051",
  2717 => x"ec397076",
  2718 => x"31517081",
  2719 => x"f1f61523",
  2720 => x"ffbc39ff",
  2721 => x"3d0d8a52",
  2722 => x"71101010",
  2723 => x"81f1ec05",
  2724 => x"51fe7134",
  2725 => x"ff127081",
  2726 => x"ff065351",
  2727 => x"71ea38ff",
  2728 => x"0b81f2c8",
  2729 => x"34833d0d",
  2730 => x"04fe3d0d",
  2731 => x"02930533",
  2732 => x"02840597",
  2733 => x"05335452",
  2734 => x"71812e92",
  2735 => x"387180d5",
  2736 => x"2ebb3881",
  2737 => x"bfb051a3",
  2738 => x"c33f843d",
  2739 => x"0d0481bf",
  2740 => x"bc51a3b8",
  2741 => x"3f72912e",
  2742 => x"81ef3872",
  2743 => x"9124b538",
  2744 => x"728c2e81",
  2745 => x"fa38728c",
  2746 => x"2480dc38",
  2747 => x"72862e81",
  2748 => x"cd3881bf",
  2749 => x"c851a394",
  2750 => x"3f843d0d",
  2751 => x"0481bfd8",
  2752 => x"51a3893f",
  2753 => x"728926ea",
  2754 => x"38721010",
  2755 => x"81c2ec05",
  2756 => x"52710804",
  2757 => x"72a82e81",
  2758 => x"bb3872a8",
  2759 => x"24943872",
  2760 => x"9a2e0981",
  2761 => x"06cc3881",
  2762 => x"bfe451a2",
  2763 => x"df3f843d",
  2764 => x"0d047280",
  2765 => x"e12e0981",
  2766 => x"06ffb738",
  2767 => x"81c08051",
  2768 => x"a2ca3f84",
  2769 => x"3d0d0472",
  2770 => x"8f2e0981",
  2771 => x"06ffa338",
  2772 => x"81c09051",
  2773 => x"a2b63f84",
  2774 => x"3d0d0481",
  2775 => x"c0ac51a2",
  2776 => x"ab3f843d",
  2777 => x"0d0481bd",
  2778 => x"b051a2a0",
  2779 => x"3f843d0d",
  2780 => x"0481c0c4",
  2781 => x"51a2953f",
  2782 => x"843d0d04",
  2783 => x"81c0d851",
  2784 => x"a28a3f84",
  2785 => x"3d0d0481",
  2786 => x"c0e851a1",
  2787 => x"ff3f843d",
  2788 => x"0d0481c0",
  2789 => x"fc51a1f4",
  2790 => x"3f843d0d",
  2791 => x"0481c198",
  2792 => x"51a1e93f",
  2793 => x"843d0d04",
  2794 => x"81c1b051",
  2795 => x"a1de3f84",
  2796 => x"3d0d0481",
  2797 => x"c1c451a1",
  2798 => x"d33f843d",
  2799 => x"0d0481c1",
  2800 => x"d451a1c8",
  2801 => x"3f843d0d",
  2802 => x"0481c1e4",
  2803 => x"51a1bd3f",
  2804 => x"843d0d04",
  2805 => x"81c1f851",
  2806 => x"a1b23f84",
  2807 => x"3d0d0481",
  2808 => x"c29851a1",
  2809 => x"a73f843d",
  2810 => x"0d04f73d",
  2811 => x"0d02b305",
  2812 => x"337c7008",
  2813 => x"c0808006",
  2814 => x"59545a80",
  2815 => x"5675832b",
  2816 => x"7707bfe0",
  2817 => x"80077070",
  2818 => x"84055208",
  2819 => x"71088c2a",
  2820 => x"bffe8006",
  2821 => x"79077198",
  2822 => x"2a728c2a",
  2823 => x"9fff0673",
  2824 => x"852a708f",
  2825 => x"06759f06",
  2826 => x"5651585d",
  2827 => x"58525558",
  2828 => x"748d3881",
  2829 => x"16568f76",
  2830 => x"27c3388b",
  2831 => x"3d0d0481",
  2832 => x"c2a851a0",
  2833 => x"c73f7551",
  2834 => x"a28c3f84",
  2835 => x"52b00851",
  2836 => x"ffbb873f",
  2837 => x"81c2b451",
  2838 => x"a0b23f74",
  2839 => x"528851a0",
  2840 => x"ce3f8452",
  2841 => x"b00851ff",
  2842 => x"baf03f81",
  2843 => x"c2bc51a0",
  2844 => x"9b3f7852",
  2845 => x"9051a0b7",
  2846 => x"3f8652b0",
  2847 => x"0851ffba",
  2848 => x"d93f81c2",
  2849 => x"c451a084",
  2850 => x"3f7251a1",
  2851 => x"c93f8452",
  2852 => x"b00851ff",
  2853 => x"bac43f81",
  2854 => x"c2cc519f",
  2855 => x"ef3f7351",
  2856 => x"a1b43f84",
  2857 => x"52b00851",
  2858 => x"ffbaaf3f",
  2859 => x"81c2d451",
  2860 => x"9fda3f77",
  2861 => x"52a0519f",
  2862 => x"f63f8a52",
  2863 => x"b00851ff",
  2864 => x"ba983f79",
  2865 => x"92388a51",
  2866 => x"9fa83f81",
  2867 => x"16568f76",
  2868 => x"27feaa38",
  2869 => x"fee53978",
  2870 => x"81ff0652",
  2871 => x"7451fbc9",
  2872 => x"3f8a519f",
  2873 => x"8d3fe439",
  2874 => x"f83d0d02",
  2875 => x"ab053359",
  2876 => x"80567585",
  2877 => x"2be09011",
  2878 => x"e0801208",
  2879 => x"70982a71",
  2880 => x"8c2a9fff",
  2881 => x"0672852a",
  2882 => x"708f0674",
  2883 => x"9f065551",
  2884 => x"585b5356",
  2885 => x"59557480",
  2886 => x"2e81a738",
  2887 => x"75bf2681",
  2888 => x"af3881c2",
  2889 => x"dc519ee4",
  2890 => x"3f7551a0",
  2891 => x"a93f8652",
  2892 => x"b00851ff",
  2893 => x"b9a43f81",
  2894 => x"c2b4519e",
  2895 => x"cf3f7452",
  2896 => x"88519eeb",
  2897 => x"3f8452b0",
  2898 => x"0851ffb9",
  2899 => x"8d3f81c2",
  2900 => x"bc519eb8",
  2901 => x"3f765290",
  2902 => x"519ed43f",
  2903 => x"8652b008",
  2904 => x"51ffb8f6",
  2905 => x"3f81c2c4",
  2906 => x"519ea13f",
  2907 => x"72519fe6",
  2908 => x"3f8452b0",
  2909 => x"0851ffb8",
  2910 => x"e13f81c2",
  2911 => x"cc519e8c",
  2912 => x"3f73519f",
  2913 => x"d13f8452",
  2914 => x"b00851ff",
  2915 => x"b8cc3f81",
  2916 => x"c2d4519d",
  2917 => x"f73f7708",
  2918 => x"c0808006",
  2919 => x"52a0519e",
  2920 => x"8e3f8a52",
  2921 => x"b00851ff",
  2922 => x"b8b03f78",
  2923 => x"81b2388a",
  2924 => x"519dbf3f",
  2925 => x"80537481",
  2926 => x"2e81df38",
  2927 => x"76862e81",
  2928 => x"bb388116",
  2929 => x"5680ff76",
  2930 => x"27fea738",
  2931 => x"8a3d0d04",
  2932 => x"81c2e451",
  2933 => x"9db63fc0",
  2934 => x"16519efa",
  2935 => x"3f8652b0",
  2936 => x"0851ffb7",
  2937 => x"f53f81c2",
  2938 => x"b4519da0",
  2939 => x"3f745288",
  2940 => x"519dbc3f",
  2941 => x"8452b008",
  2942 => x"51ffb7de",
  2943 => x"3f81c2bc",
  2944 => x"519d893f",
  2945 => x"76529051",
  2946 => x"9da53f86",
  2947 => x"52b00851",
  2948 => x"ffb7c73f",
  2949 => x"81c2c451",
  2950 => x"9cf23f72",
  2951 => x"519eb73f",
  2952 => x"8452b008",
  2953 => x"51ffb7b2",
  2954 => x"3f81c2cc",
  2955 => x"519cdd3f",
  2956 => x"73519ea2",
  2957 => x"3f8452b0",
  2958 => x"0851ffb7",
  2959 => x"9d3f81c2",
  2960 => x"d4519cc8",
  2961 => x"3f7708c0",
  2962 => x"80800652",
  2963 => x"a0519cdf",
  2964 => x"3f8a52b0",
  2965 => x"0851ffb7",
  2966 => x"813f7880",
  2967 => x"2efed038",
  2968 => x"7681ff06",
  2969 => x"527451f8",
  2970 => x"c03f8a51",
  2971 => x"9c843f80",
  2972 => x"5374812e",
  2973 => x"098106fe",
  2974 => x"c3389f39",
  2975 => x"72810657",
  2976 => x"76802efe",
  2977 => x"bd387852",
  2978 => x"7751fade",
  2979 => x"3f811656",
  2980 => x"80ff7627",
  2981 => x"fcdc38fe",
  2982 => x"b3397453",
  2983 => x"76862e09",
  2984 => x"8106fe9e",
  2985 => x"38d63980",
  2986 => x"3d0d81ce",
  2987 => x"ec085199",
  2988 => x"710c8180",
  2989 => x"0b84120c",
  2990 => x"81cee808",
  2991 => x"5199710c",
  2992 => x"81800b84",
  2993 => x"120c823d",
  2994 => x"0d04fe3d",
  2995 => x"0d740284",
  2996 => x"05970533",
  2997 => x"0288059b",
  2998 => x"05338813",
  2999 => x"0c8c120c",
  3000 => x"538c1308",
  3001 => x"70812a81",
  3002 => x"06515271",
  3003 => x"f4388c13",
  3004 => x"087081ff",
  3005 => x"06b00c51",
  3006 => x"843d0d04",
  3007 => x"803d0d72",
  3008 => x"8c110870",
  3009 => x"872a8132",
  3010 => x"8106b00c",
  3011 => x"5151823d",
  3012 => x"0d04fe3d",
  3013 => x"0dff903f",
  3014 => x"81ec5381",
  3015 => x"905281ce",
  3016 => x"ec0851ff",
  3017 => x"a53f9d53",
  3018 => x"905281ce",
  3019 => x"ec0851ff",
  3020 => x"993f80c5",
  3021 => x"5380d052",
  3022 => x"81ceec08",
  3023 => x"51ff8b3f",
  3024 => x"81ec5381",
  3025 => x"905281ce",
  3026 => x"ec0851fe",
  3027 => x"fd3fa153",
  3028 => x"905281ce",
  3029 => x"ec0851fe",
  3030 => x"f13f8953",
  3031 => x"80d05281",
  3032 => x"ceec0851",
  3033 => x"fee43f81",
  3034 => x"ec538190",
  3035 => x"5281ceec",
  3036 => x"0851fed6",
  3037 => x"3fb35390",
  3038 => x"5281ceec",
  3039 => x"0851feca",
  3040 => x"3f885380",
  3041 => x"d05281ce",
  3042 => x"ec0851fe",
  3043 => x"bd3f81ec",
  3044 => x"53819052",
  3045 => x"81ceec08",
  3046 => x"51feaf3f",
  3047 => x"b4539052",
  3048 => x"81ceec08",
  3049 => x"51fea33f",
  3050 => x"965380d0",
  3051 => x"5281ceec",
  3052 => x"0851fe96",
  3053 => x"3f81ec53",
  3054 => x"81905281",
  3055 => x"ceec0851",
  3056 => x"fe883fb6",
  3057 => x"53905281",
  3058 => x"ceec0851",
  3059 => x"fdfc3f80",
  3060 => x"e05380d0",
  3061 => x"5281ceec",
  3062 => x"0851fdee",
  3063 => x"3f81ec53",
  3064 => x"81905281",
  3065 => x"ceec0851",
  3066 => x"fde03f80",
  3067 => x"c9539052",
  3068 => x"81ceec08",
  3069 => x"51fdd33f",
  3070 => x"81c05380",
  3071 => x"d05281ce",
  3072 => x"ec0851fd",
  3073 => x"c53f843d",
  3074 => x"0d04fd3d",
  3075 => x"0d029705",
  3076 => x"33028405",
  3077 => x"9b053371",
  3078 => x"81b00781",
  3079 => x"bf065354",
  3080 => x"54f88080",
  3081 => x"98807171",
  3082 => x"0c73842a",
  3083 => x"9007710c",
  3084 => x"738f0671",
  3085 => x"0c527281",
  3086 => x"cec83473",
  3087 => x"81cecc34",
  3088 => x"853d0d04",
  3089 => x"fd3d0d02",
  3090 => x"97053381",
  3091 => x"cecc3354",
  3092 => x"73058706",
  3093 => x"0284059a",
  3094 => x"052281ce",
  3095 => x"c8335473",
  3096 => x"057081ff",
  3097 => x"067281b0",
  3098 => x"07545154",
  3099 => x"54f88080",
  3100 => x"98807171",
  3101 => x"0c73842a",
  3102 => x"9007710c",
  3103 => x"738f0671",
  3104 => x"0c527281",
  3105 => x"cec83473",
  3106 => x"81cecc34",
  3107 => x"853d0d04",
  3108 => x"ff3d0d02",
  3109 => x"8f0533f8",
  3110 => x"80809884",
  3111 => x"0c81cec8",
  3112 => x"33810551",
  3113 => x"7081cec8",
  3114 => x"34833d0d",
  3115 => x"04ff3d0d",
  3116 => x"80527181",
  3117 => x"b00781bf",
  3118 => x"06f88080",
  3119 => x"98800c90",
  3120 => x"0bf88080",
  3121 => x"98800c80",
  3122 => x"0bf88080",
  3123 => x"98800c80",
  3124 => x"51800bf8",
  3125 => x"80809884",
  3126 => x"0c811170",
  3127 => x"81ff0651",
  3128 => x"5180e571",
  3129 => x"27eb3881",
  3130 => x"127081ff",
  3131 => x"06535187",
  3132 => x"7227ffbe",
  3133 => x"3881b00b",
  3134 => x"f8808098",
  3135 => x"800c900b",
  3136 => x"f8808098",
  3137 => x"800c800b",
  3138 => x"f8808098",
  3139 => x"800c800b",
  3140 => x"81cec834",
  3141 => x"800b81ce",
  3142 => x"cc34833d",
  3143 => x"0d04ff3d",
  3144 => x"0d80c00b",
  3145 => x"f8808098",
  3146 => x"800c81a1",
  3147 => x"0bf88080",
  3148 => x"98800c81",
  3149 => x"c00bf880",
  3150 => x"8098800c",
  3151 => x"81a40bf8",
  3152 => x"80809880",
  3153 => x"0c81a60b",
  3154 => x"f8808098",
  3155 => x"800c81a2",
  3156 => x"0bf88080",
  3157 => x"98800caf",
  3158 => x"0bf88080",
  3159 => x"98800ca5",
  3160 => x"0bf88080",
  3161 => x"98800c81",
  3162 => x"810bf880",
  3163 => x"8098800c",
  3164 => x"9d0bf880",
  3165 => x"8098800c",
  3166 => x"81fa0bf8",
  3167 => x"80809880",
  3168 => x"0c800bf8",
  3169 => x"80809880",
  3170 => x"0c805271",
  3171 => x"81b00781",
  3172 => x"bf06f880",
  3173 => x"8098800c",
  3174 => x"900bf880",
  3175 => x"8098800c",
  3176 => x"800bf880",
  3177 => x"8098800c",
  3178 => x"8051800b",
  3179 => x"f8808098",
  3180 => x"840c8111",
  3181 => x"7081ff06",
  3182 => x"515180e5",
  3183 => x"7127eb38",
  3184 => x"81127081",
  3185 => x"ff065351",
  3186 => x"877227ff",
  3187 => x"be3881b0",
  3188 => x"0bf88080",
  3189 => x"98800c90",
  3190 => x"0bf88080",
  3191 => x"98800c80",
  3192 => x"0bf88080",
  3193 => x"98800c80",
  3194 => x"0b81cec8",
  3195 => x"34800b81",
  3196 => x"cecc3481",
  3197 => x"af0bf880",
  3198 => x"8098800c",
  3199 => x"833d0d04",
  3200 => x"803d0d02",
  3201 => x"8f053373",
  3202 => x"81f2cc0c",
  3203 => x"517081f2",
  3204 => x"d034823d",
  3205 => x"0d04ee3d",
  3206 => x"0d640284",
  3207 => x"0580d705",
  3208 => x"33028805",
  3209 => x"80db0533",
  3210 => x"59575980",
  3211 => x"76810677",
  3212 => x"812a8106",
  3213 => x"78832b81",
  3214 => x"80067982",
  3215 => x"2a810657",
  3216 => x"5e415f5d",
  3217 => x"81ff4272",
  3218 => x"7d2e0981",
  3219 => x"0683387c",
  3220 => x"42768a2e",
  3221 => x"83b93888",
  3222 => x"19085574",
  3223 => x"802e83a4",
  3224 => x"38851933",
  3225 => x"5aff5376",
  3226 => x"7a268e38",
  3227 => x"84193354",
  3228 => x"73772685",
  3229 => x"38767431",
  3230 => x"53741370",
  3231 => x"33545872",
  3232 => x"81ff0683",
  3233 => x"1a337098",
  3234 => x"2b81ff0a",
  3235 => x"119b2a81",
  3236 => x"055b4542",
  3237 => x"40815374",
  3238 => x"83387453",
  3239 => x"7281ff06",
  3240 => x"43807a81",
  3241 => x"ff06545c",
  3242 => x"ff547673",
  3243 => x"268b3884",
  3244 => x"19335376",
  3245 => x"732783f4",
  3246 => x"38737481",
  3247 => x"ff065553",
  3248 => x"805a7973",
  3249 => x"24ab3874",
  3250 => x"7a2e0981",
  3251 => x"0682e138",
  3252 => x"60982b81",
  3253 => x"ff0a119b",
  3254 => x"2a821b33",
  3255 => x"71712911",
  3256 => x"7081ff06",
  3257 => x"7871298c",
  3258 => x"1f080552",
  3259 => x"455d575d",
  3260 => x"537f6305",
  3261 => x"7081ff06",
  3262 => x"70612b70",
  3263 => x"81ff067b",
  3264 => x"622b7081",
  3265 => x"ff067b83",
  3266 => x"2a81065f",
  3267 => x"5358525e",
  3268 => x"42557880",
  3269 => x"2e8f3881",
  3270 => x"cec83361",
  3271 => x"05567580",
  3272 => x"e62483c5",
  3273 => x"387f7829",
  3274 => x"61304157",
  3275 => x"7c7e2c98",
  3276 => x"2b70982c",
  3277 => x"55557377",
  3278 => x"25818238",
  3279 => x"ff1c7d81",
  3280 => x"065a537c",
  3281 => x"732e83c4",
  3282 => x"387e86a6",
  3283 => x"386184eb",
  3284 => x"387d802e",
  3285 => x"82a43879",
  3286 => x"14703370",
  3287 => x"58545580",
  3288 => x"5578752e",
  3289 => x"85387284",
  3290 => x"2a567583",
  3291 => x"2a708106",
  3292 => x"51537280",
  3293 => x"2e843881",
  3294 => x"c0557582",
  3295 => x"2a708106",
  3296 => x"51537280",
  3297 => x"2e853874",
  3298 => x"b0075575",
  3299 => x"812a7081",
  3300 => x"06515372",
  3301 => x"802e8538",
  3302 => x"748c0755",
  3303 => x"75810653",
  3304 => x"72802e85",
  3305 => x"38748307",
  3306 => x"557451f9",
  3307 => x"e33f7714",
  3308 => x"982b7098",
  3309 => x"2c555676",
  3310 => x"7424ff9b",
  3311 => x"3862802e",
  3312 => x"953861ff",
  3313 => x"1d54547c",
  3314 => x"732e81fb",
  3315 => x"387351f9",
  3316 => x"bf3f7e81",
  3317 => x"ea387f52",
  3318 => x"8151f8e8",
  3319 => x"3f811d70",
  3320 => x"81ff065e",
  3321 => x"547b7d26",
  3322 => x"fec23860",
  3323 => x"527b3070",
  3324 => x"982b7098",
  3325 => x"2c53585b",
  3326 => x"f8ca3f60",
  3327 => x"5372b00c",
  3328 => x"943d0d04",
  3329 => x"82193385",
  3330 => x"1a335b53",
  3331 => x"fcf13981",
  3332 => x"cecc3353",
  3333 => x"72872681",
  3334 => x"9a388113",
  3335 => x"56805275",
  3336 => x"81ff0651",
  3337 => x"f7e43f80",
  3338 => x"5372b00c",
  3339 => x"943d0d04",
  3340 => x"73802eaf",
  3341 => x"38ff1470",
  3342 => x"81ff0655",
  3343 => x"5a7381ff",
  3344 => x"2ea13874",
  3345 => x"70810556",
  3346 => x"337c0570",
  3347 => x"83ffff06",
  3348 => x"ff167081",
  3349 => x"ff06575c",
  3350 => x"5d537381",
  3351 => x"ff2e0981",
  3352 => x"06e13860",
  3353 => x"982b81ff",
  3354 => x"0a119b2a",
  3355 => x"707e291e",
  3356 => x"8c1c0805",
  3357 => x"5c4255fc",
  3358 => x"f8397914",
  3359 => x"70335259",
  3360 => x"f88e3f77",
  3361 => x"14982b70",
  3362 => x"982c5556",
  3363 => x"737725fe",
  3364 => x"ac387914",
  3365 => x"70335259",
  3366 => x"f7f63f77",
  3367 => x"14982b70",
  3368 => x"982c5556",
  3369 => x"767424d2",
  3370 => x"38fe9239",
  3371 => x"76733154",
  3372 => x"fc873980",
  3373 => x"528051f6",
  3374 => x"d13f8053",
  3375 => x"feeb3973",
  3376 => x"51f7cd3f",
  3377 => x"fe903961",
  3378 => x"7b327081",
  3379 => x"ff065555",
  3380 => x"7d802efd",
  3381 => x"f8387a81",
  3382 => x"2a743270",
  3383 => x"5254f7b0",
  3384 => x"3f7e802e",
  3385 => x"fdf038d7",
  3386 => x"3981cecc",
  3387 => x"337c0553",
  3388 => x"80527281",
  3389 => x"ff0651f6",
  3390 => x"913f8053",
  3391 => x"76a02efd",
  3392 => x"fc387f78",
  3393 => x"29613041",
  3394 => x"57fca139",
  3395 => x"7e87ad38",
  3396 => x"6185eb38",
  3397 => x"7d802e80",
  3398 => x"ec387914",
  3399 => x"70337c07",
  3400 => x"70525456",
  3401 => x"80557875",
  3402 => x"2e853872",
  3403 => x"842a5675",
  3404 => x"832a7081",
  3405 => x"06515372",
  3406 => x"802e8438",
  3407 => x"81c05575",
  3408 => x"822a7081",
  3409 => x"06515372",
  3410 => x"802e8538",
  3411 => x"74b00755",
  3412 => x"75812a70",
  3413 => x"81065153",
  3414 => x"72802e85",
  3415 => x"38748c07",
  3416 => x"55758106",
  3417 => x"5372802e",
  3418 => x"85387483",
  3419 => x"07557451",
  3420 => x"f69e3f77",
  3421 => x"14982b70",
  3422 => x"982c5553",
  3423 => x"767424ff",
  3424 => x"9938fcb9",
  3425 => x"39791470",
  3426 => x"337c0752",
  3427 => x"56f6813f",
  3428 => x"7714982b",
  3429 => x"70982c55",
  3430 => x"59737725",
  3431 => x"fc9f3879",
  3432 => x"1470337c",
  3433 => x"075256f5",
  3434 => x"e73f7714",
  3435 => x"982b7098",
  3436 => x"2c555976",
  3437 => x"7424ce38",
  3438 => x"fc83397d",
  3439 => x"802e80f0",
  3440 => x"38791470",
  3441 => x"33705854",
  3442 => x"55805578",
  3443 => x"752e8538",
  3444 => x"72842a56",
  3445 => x"75832a70",
  3446 => x"81065153",
  3447 => x"72802e84",
  3448 => x"3881c055",
  3449 => x"75822a70",
  3450 => x"81065153",
  3451 => x"72802e85",
  3452 => x"3874b007",
  3453 => x"5575812a",
  3454 => x"70810651",
  3455 => x"5372802e",
  3456 => x"8538748c",
  3457 => x"07557581",
  3458 => x"06537280",
  3459 => x"2e853874",
  3460 => x"83075574",
  3461 => x"097081ff",
  3462 => x"065253f4",
  3463 => x"f33f7714",
  3464 => x"982b7098",
  3465 => x"2c555676",
  3466 => x"7424ff95",
  3467 => x"38fb8e39",
  3468 => x"79147033",
  3469 => x"70097081",
  3470 => x"ff065458",
  3471 => x"5455f4d0",
  3472 => x"3f771498",
  3473 => x"2b70982c",
  3474 => x"55597377",
  3475 => x"25faee38",
  3476 => x"79147033",
  3477 => x"70097081",
  3478 => x"ff065458",
  3479 => x"5455f4b0",
  3480 => x"3f771498",
  3481 => x"2b70982c",
  3482 => x"55597674",
  3483 => x"24c238fa",
  3484 => x"cc396180",
  3485 => x"2e81ce38",
  3486 => x"7d802e80",
  3487 => x"f7387914",
  3488 => x"70337058",
  3489 => x"54558055",
  3490 => x"78752e85",
  3491 => x"3872842a",
  3492 => x"5675832a",
  3493 => x"70810651",
  3494 => x"5372802e",
  3495 => x"843881c0",
  3496 => x"5575822a",
  3497 => x"70810651",
  3498 => x"5372802e",
  3499 => x"853874b0",
  3500 => x"07557581",
  3501 => x"2a708106",
  3502 => x"51537280",
  3503 => x"2e853874",
  3504 => x"8c075575",
  3505 => x"81065372",
  3506 => x"802e8538",
  3507 => x"74830755",
  3508 => x"74097081",
  3509 => x"ff067053",
  3510 => x"5753f3b4",
  3511 => x"3f7551f3",
  3512 => x"af3f7714",
  3513 => x"982b7098",
  3514 => x"2c555576",
  3515 => x"7424ff8e",
  3516 => x"38f9ca39",
  3517 => x"79147033",
  3518 => x"70097081",
  3519 => x"ff067055",
  3520 => x"59555659",
  3521 => x"f38a3f75",
  3522 => x"51f3853f",
  3523 => x"7714982b",
  3524 => x"70982c55",
  3525 => x"59737725",
  3526 => x"f9a33879",
  3527 => x"14703370",
  3528 => x"097081ff",
  3529 => x"06705559",
  3530 => x"555659f2",
  3531 => x"e33f7551",
  3532 => x"f2de3f77",
  3533 => x"14982b70",
  3534 => x"982c5559",
  3535 => x"767424ff",
  3536 => x"b338f8f9",
  3537 => x"397d802e",
  3538 => x"80f43879",
  3539 => x"14703370",
  3540 => x"58545580",
  3541 => x"5578752e",
  3542 => x"85387284",
  3543 => x"2a567583",
  3544 => x"2a708106",
  3545 => x"51537280",
  3546 => x"2e843881",
  3547 => x"c0557582",
  3548 => x"2a708106",
  3549 => x"51537280",
  3550 => x"2e853874",
  3551 => x"b0075575",
  3552 => x"812a7081",
  3553 => x"06515372",
  3554 => x"802e8538",
  3555 => x"748c0755",
  3556 => x"75810653",
  3557 => x"72802e85",
  3558 => x"38748307",
  3559 => x"557481ff",
  3560 => x"06705256",
  3561 => x"f1ea3f75",
  3562 => x"51f1e53f",
  3563 => x"7714982b",
  3564 => x"70982c55",
  3565 => x"55767424",
  3566 => x"ff9138f8",
  3567 => x"80397914",
  3568 => x"70337053",
  3569 => x"5753f1c8",
  3570 => x"3f7551f1",
  3571 => x"c33f7714",
  3572 => x"982b7098",
  3573 => x"2c555973",
  3574 => x"7725f7e1",
  3575 => x"38791470",
  3576 => x"33705357",
  3577 => x"53f1a93f",
  3578 => x"7551f1a4",
  3579 => x"3f771498",
  3580 => x"2b70982c",
  3581 => x"55597674",
  3582 => x"24c438f7",
  3583 => x"c0397d80",
  3584 => x"2e80f238",
  3585 => x"79147033",
  3586 => x"7c077052",
  3587 => x"54568055",
  3588 => x"78752e85",
  3589 => x"3872842a",
  3590 => x"5675832a",
  3591 => x"70810651",
  3592 => x"5372802e",
  3593 => x"843881c0",
  3594 => x"5575822a",
  3595 => x"70810651",
  3596 => x"5372802e",
  3597 => x"853874b0",
  3598 => x"07557581",
  3599 => x"2a708106",
  3600 => x"51537280",
  3601 => x"2e853874",
  3602 => x"8c075575",
  3603 => x"81065372",
  3604 => x"802e8538",
  3605 => x"74830755",
  3606 => x"74097081",
  3607 => x"ff065256",
  3608 => x"f0ae3f77",
  3609 => x"14982b70",
  3610 => x"982c5553",
  3611 => x"767424ff",
  3612 => x"9338f6c9",
  3613 => x"39791470",
  3614 => x"337c0770",
  3615 => x"097081ff",
  3616 => x"06545556",
  3617 => x"59f0893f",
  3618 => x"7714982b",
  3619 => x"70982c55",
  3620 => x"59737725",
  3621 => x"f6a73879",
  3622 => x"1470337c",
  3623 => x"07700970",
  3624 => x"81ff0654",
  3625 => x"555659ef",
  3626 => x"e73f7714",
  3627 => x"982b7098",
  3628 => x"2c555976",
  3629 => x"7424ffbd",
  3630 => x"38f68239",
  3631 => x"61802e81",
  3632 => x"d4387d80",
  3633 => x"2e80f938",
  3634 => x"79147033",
  3635 => x"7c077052",
  3636 => x"54568055",
  3637 => x"78752e85",
  3638 => x"3872842a",
  3639 => x"5675832a",
  3640 => x"70810651",
  3641 => x"5372802e",
  3642 => x"843881c0",
  3643 => x"5575822a",
  3644 => x"70810651",
  3645 => x"5372802e",
  3646 => x"853874b0",
  3647 => x"07557581",
  3648 => x"2a708106",
  3649 => x"51537280",
  3650 => x"2e853874",
  3651 => x"8c075575",
  3652 => x"81065372",
  3653 => x"802e8538",
  3654 => x"74830755",
  3655 => x"74097081",
  3656 => x"ff067053",
  3657 => x"5456eee8",
  3658 => x"3f7251ee",
  3659 => x"e33f7714",
  3660 => x"982b7098",
  3661 => x"2c555676",
  3662 => x"7424ff8c",
  3663 => x"38f4fe39",
  3664 => x"79147033",
  3665 => x"7c077009",
  3666 => x"7081ff06",
  3667 => x"70555357",
  3668 => x"5753eebc",
  3669 => x"3f7251ee",
  3670 => x"b73f7714",
  3671 => x"982b7098",
  3672 => x"2c555973",
  3673 => x"7725f4d5",
  3674 => x"38791470",
  3675 => x"337c0770",
  3676 => x"097081ff",
  3677 => x"06705553",
  3678 => x"575753ee",
  3679 => x"933f7251",
  3680 => x"ee8e3f77",
  3681 => x"14982b70",
  3682 => x"982c5559",
  3683 => x"767424ff",
  3684 => x"af38f4a9",
  3685 => x"397d802e",
  3686 => x"80f63879",
  3687 => x"1470337c",
  3688 => x"07705254",
  3689 => x"56805578",
  3690 => x"752e8538",
  3691 => x"72842a56",
  3692 => x"75832a70",
  3693 => x"81065153",
  3694 => x"72802e84",
  3695 => x"3881c055",
  3696 => x"75822a70",
  3697 => x"81065153",
  3698 => x"72802e85",
  3699 => x"3874b007",
  3700 => x"5575812a",
  3701 => x"70810651",
  3702 => x"5372802e",
  3703 => x"8538748c",
  3704 => x"07557581",
  3705 => x"06537280",
  3706 => x"2e853874",
  3707 => x"83075574",
  3708 => x"81ff0670",
  3709 => x"5256ed98",
  3710 => x"3f7551ed",
  3711 => x"933f7714",
  3712 => x"982b7098",
  3713 => x"2c555376",
  3714 => x"7424ff8f",
  3715 => x"38f3ae39",
  3716 => x"79147033",
  3717 => x"7c077053",
  3718 => x"5456ecf4",
  3719 => x"3f7251ec",
  3720 => x"ef3f7714",
  3721 => x"982b7098",
  3722 => x"2c555973",
  3723 => x"7725f38d",
  3724 => x"38791470",
  3725 => x"337c0770",
  3726 => x"535456ec",
  3727 => x"d33f7251",
  3728 => x"ecce3f77",
  3729 => x"14982b70",
  3730 => x"982c5559",
  3731 => x"767424c0",
  3732 => x"38f2ea39",
  3733 => x"f83d0d7a",
  3734 => x"7d028805",
  3735 => x"af05335a",
  3736 => x"55598074",
  3737 => x"70810556",
  3738 => x"33755856",
  3739 => x"5774772e",
  3740 => x"09810688",
  3741 => x"3876b00c",
  3742 => x"8a3d0d04",
  3743 => x"74537752",
  3744 => x"7851ef92",
  3745 => x"3fb00881",
  3746 => x"ff067705",
  3747 => x"7083ffff",
  3748 => x"06777081",
  3749 => x"05593352",
  3750 => x"58557480",
  3751 => x"2ed73874",
  3752 => x"53775278",
  3753 => x"51eeef3f",
  3754 => x"b00881ff",
  3755 => x"06770570",
  3756 => x"83ffff06",
  3757 => x"77708105",
  3758 => x"59335258",
  3759 => x"5574ffbc",
  3760 => x"38ffb239",
  3761 => x"fe3d0d02",
  3762 => x"93053353",
  3763 => x"81f2d033",
  3764 => x"5281f2cc",
  3765 => x"0851eebe",
  3766 => x"3fb00881",
  3767 => x"ff06b00c",
  3768 => x"843d0d04",
  3769 => x"d0893f04",
  3770 => x"fb3d0d77",
  3771 => x"79555580",
  3772 => x"56757524",
  3773 => x"ab388074",
  3774 => x"249d3880",
  3775 => x"53735274",
  3776 => x"5180e13f",
  3777 => x"b0085475",
  3778 => x"802e8538",
  3779 => x"b0083054",
  3780 => x"73b00c87",
  3781 => x"3d0d0473",
  3782 => x"30768132",
  3783 => x"5754dc39",
  3784 => x"74305581",
  3785 => x"56738025",
  3786 => x"d238ec39",
  3787 => x"fa3d0d78",
  3788 => x"7a575580",
  3789 => x"57767524",
  3790 => x"a438759f",
  3791 => x"2c548153",
  3792 => x"75743274",
  3793 => x"31527451",
  3794 => x"9b3fb008",
  3795 => x"5476802e",
  3796 => x"8538b008",
  3797 => x"305473b0",
  3798 => x"0c883d0d",
  3799 => x"04743055",
  3800 => x"8157d739",
  3801 => x"fc3d0d76",
  3802 => x"78535481",
  3803 => x"53807473",
  3804 => x"26525572",
  3805 => x"802e9838",
  3806 => x"70802ea9",
  3807 => x"38807224",
  3808 => x"a4387110",
  3809 => x"73107572",
  3810 => x"26535452",
  3811 => x"72ea3873",
  3812 => x"51788338",
  3813 => x"745170b0",
  3814 => x"0c863d0d",
  3815 => x"0472812a",
  3816 => x"72812a53",
  3817 => x"5372802e",
  3818 => x"e6387174",
  3819 => x"26ef3873",
  3820 => x"72317574",
  3821 => x"0774812a",
  3822 => x"74812a55",
  3823 => x"555654e5",
  3824 => x"39101010",
  3825 => x"10101010",
  3826 => x"10101010",
  3827 => x"10101010",
  3828 => x"10101010",
  3829 => x"10101010",
  3830 => x"10101010",
  3831 => x"10101010",
  3832 => x"53510473",
  3833 => x"81ff0673",
  3834 => x"83060981",
  3835 => x"05830510",
  3836 => x"10102b07",
  3837 => x"72fc060c",
  3838 => x"5151043c",
  3839 => x"04727280",
  3840 => x"728106ff",
  3841 => x"05097206",
  3842 => x"05711052",
  3843 => x"720a100a",
  3844 => x"5372ed38",
  3845 => x"51515351",
  3846 => x"04b008b4",
  3847 => x"08b80875",
  3848 => x"7580f6ac",
  3849 => x"2d5050b0",
  3850 => x"0856b80c",
  3851 => x"b40cb00c",
  3852 => x"5104b008",
  3853 => x"b408b808",
  3854 => x"757580f5",
  3855 => x"e82d5050",
  3856 => x"b00856b8",
  3857 => x"0cb40cb0",
  3858 => x"0c5104b0",
  3859 => x"08b408b8",
  3860 => x"0880c5c6",
  3861 => x"2db80cb4",
  3862 => x"0cb00c04",
  3863 => x"ff3d0d02",
  3864 => x"8f053381",
  3865 => x"cf840852",
  3866 => x"710c800b",
  3867 => x"b00c833d",
  3868 => x"0d04ff3d",
  3869 => x"0d028f05",
  3870 => x"335181f2",
  3871 => x"d4085271",
  3872 => x"2db00881",
  3873 => x"ff06b00c",
  3874 => x"833d0d04",
  3875 => x"fe3d0d74",
  3876 => x"70335353",
  3877 => x"71802e93",
  3878 => x"38811372",
  3879 => x"5281f2d4",
  3880 => x"08535371",
  3881 => x"2d723352",
  3882 => x"71ef3884",
  3883 => x"3d0d04f4",
  3884 => x"3d0d7f02",
  3885 => x"8405bb05",
  3886 => x"33555788",
  3887 => x"0b8c3d5b",
  3888 => x"59895381",
  3889 => x"cc9c5279",
  3890 => x"5186b63f",
  3891 => x"73792e80",
  3892 => x"ff387856",
  3893 => x"73902e80",
  3894 => x"ec3802a7",
  3895 => x"0558768f",
  3896 => x"06547389",
  3897 => x"2680c238",
  3898 => x"7518b015",
  3899 => x"55557375",
  3900 => x"3476842a",
  3901 => x"ff177081",
  3902 => x"ff065855",
  3903 => x"5775df38",
  3904 => x"781a5575",
  3905 => x"75347970",
  3906 => x"33555573",
  3907 => x"802e9338",
  3908 => x"81157452",
  3909 => x"81f2d408",
  3910 => x"5755752d",
  3911 => x"74335473",
  3912 => x"ef3878b0",
  3913 => x"0c8e3d0d",
  3914 => x"047518b7",
  3915 => x"15555573",
  3916 => x"75347684",
  3917 => x"2aff1770",
  3918 => x"81ff0658",
  3919 => x"555775ff",
  3920 => x"9d38ffbc",
  3921 => x"39847057",
  3922 => x"5902a705",
  3923 => x"58ff8f39",
  3924 => x"82705759",
  3925 => x"f439f13d",
  3926 => x"0d618d3d",
  3927 => x"705b5c5a",
  3928 => x"807a5657",
  3929 => x"767a2481",
  3930 => x"85387817",
  3931 => x"548a5274",
  3932 => x"5184dc3f",
  3933 => x"b008b005",
  3934 => x"53727434",
  3935 => x"8117578a",
  3936 => x"52745184",
  3937 => x"a53fb008",
  3938 => x"55b008de",
  3939 => x"38b00877",
  3940 => x"9f2a1870",
  3941 => x"812c5a56",
  3942 => x"56807825",
  3943 => x"9e387817",
  3944 => x"ff055575",
  3945 => x"19703355",
  3946 => x"53743373",
  3947 => x"34737534",
  3948 => x"8116ff16",
  3949 => x"56567776",
  3950 => x"24e93876",
  3951 => x"19588078",
  3952 => x"34807a24",
  3953 => x"177081ff",
  3954 => x"067c7033",
  3955 => x"56575556",
  3956 => x"72802e93",
  3957 => x"38811573",
  3958 => x"5281f2d4",
  3959 => x"08585576",
  3960 => x"2d743353",
  3961 => x"72ef3873",
  3962 => x"b00c913d",
  3963 => x"0d04ad7b",
  3964 => x"3402ad05",
  3965 => x"7a307119",
  3966 => x"5656598a",
  3967 => x"52745183",
  3968 => x"ce3fb008",
  3969 => x"b0055372",
  3970 => x"74348117",
  3971 => x"578a5274",
  3972 => x"5183973f",
  3973 => x"b00855b0",
  3974 => x"08fecf38",
  3975 => x"feef39fd",
  3976 => x"3d0d81ce",
  3977 => x"f80876b2",
  3978 => x"e4299412",
  3979 => x"0c54850b",
  3980 => x"98150c98",
  3981 => x"14087081",
  3982 => x"06515372",
  3983 => x"f638853d",
  3984 => x"0d04803d",
  3985 => x"0d81cef8",
  3986 => x"0851870b",
  3987 => x"84120cff",
  3988 => x"0ba4120c",
  3989 => x"a70ba812",
  3990 => x"0cb2e40b",
  3991 => x"94120c87",
  3992 => x"0b98120c",
  3993 => x"823d0d04",
  3994 => x"803d0d81",
  3995 => x"cefc0851",
  3996 => x"b80b8c12",
  3997 => x"0c830b88",
  3998 => x"120c823d",
  3999 => x"0d04803d",
  4000 => x"0d81cefc",
  4001 => x"08841108",
  4002 => x"8106b00c",
  4003 => x"51823d0d",
  4004 => x"04ff3d0d",
  4005 => x"81cefc08",
  4006 => x"52841208",
  4007 => x"70810651",
  4008 => x"5170802e",
  4009 => x"f4387108",
  4010 => x"7081ff06",
  4011 => x"b00c5183",
  4012 => x"3d0d04fe",
  4013 => x"3d0d0293",
  4014 => x"05335372",
  4015 => x"8a2e9c38",
  4016 => x"81cefc08",
  4017 => x"52841208",
  4018 => x"70892a70",
  4019 => x"81065151",
  4020 => x"5170f238",
  4021 => x"72720c84",
  4022 => x"3d0d0481",
  4023 => x"cefc0852",
  4024 => x"84120870",
  4025 => x"892a7081",
  4026 => x"06515151",
  4027 => x"70f2388d",
  4028 => x"720c8412",
  4029 => x"0870892a",
  4030 => x"70810651",
  4031 => x"515170c5",
  4032 => x"38d23980",
  4033 => x"3d0d81ce",
  4034 => x"f0085180",
  4035 => x"0b84120c",
  4036 => x"83fe800b",
  4037 => x"88120c80",
  4038 => x"0b81f2d8",
  4039 => x"34800b81",
  4040 => x"f2dc3482",
  4041 => x"3d0d04fa",
  4042 => x"3d0d02a3",
  4043 => x"053381ce",
  4044 => x"f00881f2",
  4045 => x"d8337081",
  4046 => x"ff067010",
  4047 => x"101181f2",
  4048 => x"dc337081",
  4049 => x"ff067290",
  4050 => x"29117088",
  4051 => x"2b780777",
  4052 => x"0c535b5b",
  4053 => x"55555954",
  4054 => x"54738a2e",
  4055 => x"98387480",
  4056 => x"cf2e9238",
  4057 => x"738c2ea4",
  4058 => x"38811653",
  4059 => x"7281f2dc",
  4060 => x"34883d0d",
  4061 => x"0471a326",
  4062 => x"a3388117",
  4063 => x"527181f2",
  4064 => x"d834800b",
  4065 => x"81f2dc34",
  4066 => x"883d0d04",
  4067 => x"80527188",
  4068 => x"2b730c81",
  4069 => x"12529790",
  4070 => x"7226f338",
  4071 => x"800b81f2",
  4072 => x"d834800b",
  4073 => x"81f2dc34",
  4074 => x"df39bc08",
  4075 => x"02bc0cfd",
  4076 => x"3d0d8053",
  4077 => x"bc088c05",
  4078 => x"0852bc08",
  4079 => x"88050851",
  4080 => x"f7a23fb0",
  4081 => x"0870b00c",
  4082 => x"54853d0d",
  4083 => x"bc0c04bc",
  4084 => x"0802bc0c",
  4085 => x"fd3d0d81",
  4086 => x"53bc088c",
  4087 => x"050852bc",
  4088 => x"08880508",
  4089 => x"51f6fd3f",
  4090 => x"b00870b0",
  4091 => x"0c54853d",
  4092 => x"0dbc0c04",
  4093 => x"803d0d86",
  4094 => x"5184963f",
  4095 => x"8151a1d3",
  4096 => x"3ffc3d0d",
  4097 => x"7670797b",
  4098 => x"55555555",
  4099 => x"8f72278c",
  4100 => x"38727507",
  4101 => x"83065170",
  4102 => x"802ea738",
  4103 => x"ff125271",
  4104 => x"ff2e9838",
  4105 => x"72708105",
  4106 => x"54337470",
  4107 => x"81055634",
  4108 => x"ff125271",
  4109 => x"ff2e0981",
  4110 => x"06ea3874",
  4111 => x"b00c863d",
  4112 => x"0d047451",
  4113 => x"72708405",
  4114 => x"54087170",
  4115 => x"8405530c",
  4116 => x"72708405",
  4117 => x"54087170",
  4118 => x"8405530c",
  4119 => x"72708405",
  4120 => x"54087170",
  4121 => x"8405530c",
  4122 => x"72708405",
  4123 => x"54087170",
  4124 => x"8405530c",
  4125 => x"f0125271",
  4126 => x"8f26c938",
  4127 => x"83722795",
  4128 => x"38727084",
  4129 => x"05540871",
  4130 => x"70840553",
  4131 => x"0cfc1252",
  4132 => x"718326ed",
  4133 => x"387054ff",
  4134 => x"8339fd3d",
  4135 => x"0d755384",
  4136 => x"d8130880",
  4137 => x"2e8a3880",
  4138 => x"5372b00c",
  4139 => x"853d0d04",
  4140 => x"81805272",
  4141 => x"518d9b3f",
  4142 => x"b00884d8",
  4143 => x"140cff53",
  4144 => x"b008802e",
  4145 => x"e438b008",
  4146 => x"549f5380",
  4147 => x"74708405",
  4148 => x"560cff13",
  4149 => x"53807324",
  4150 => x"ce388074",
  4151 => x"70840556",
  4152 => x"0cff1353",
  4153 => x"728025e3",
  4154 => x"38ffbc39",
  4155 => x"fd3d0d75",
  4156 => x"7755539f",
  4157 => x"74278d38",
  4158 => x"96730cff",
  4159 => x"5271b00c",
  4160 => x"853d0d04",
  4161 => x"84d81308",
  4162 => x"5271802e",
  4163 => x"93387310",
  4164 => x"10127008",
  4165 => x"79720c51",
  4166 => x"5271b00c",
  4167 => x"853d0d04",
  4168 => x"7251fef6",
  4169 => x"3fff52b0",
  4170 => x"08d33884",
  4171 => x"d8130874",
  4172 => x"10101170",
  4173 => x"087a720c",
  4174 => x"515152dd",
  4175 => x"39f93d0d",
  4176 => x"797b5856",
  4177 => x"769f2680",
  4178 => x"e83884d8",
  4179 => x"16085473",
  4180 => x"802eaa38",
  4181 => x"76101014",
  4182 => x"70085555",
  4183 => x"73802eba",
  4184 => x"38805873",
  4185 => x"812e8f38",
  4186 => x"73ff2ea3",
  4187 => x"3880750c",
  4188 => x"7651732d",
  4189 => x"805877b0",
  4190 => x"0c893d0d",
  4191 => x"047551fe",
  4192 => x"993fff58",
  4193 => x"b008ef38",
  4194 => x"84d81608",
  4195 => x"54c63996",
  4196 => x"760c810b",
  4197 => x"b00c893d",
  4198 => x"0d047551",
  4199 => x"81ed3f76",
  4200 => x"53b00852",
  4201 => x"755181ad",
  4202 => x"3fb008b0",
  4203 => x"0c893d0d",
  4204 => x"0496760c",
  4205 => x"ff0bb00c",
  4206 => x"893d0d04",
  4207 => x"fc3d0d76",
  4208 => x"785653ff",
  4209 => x"54749f26",
  4210 => x"b13884d8",
  4211 => x"13085271",
  4212 => x"802eae38",
  4213 => x"74101012",
  4214 => x"70085353",
  4215 => x"81547180",
  4216 => x"2e983882",
  4217 => x"5471ff2e",
  4218 => x"91388354",
  4219 => x"71812e8a",
  4220 => x"3880730c",
  4221 => x"7451712d",
  4222 => x"805473b0",
  4223 => x"0c863d0d",
  4224 => x"047251fd",
  4225 => x"953fb008",
  4226 => x"f13884d8",
  4227 => x"130852c4",
  4228 => x"39ff3d0d",
  4229 => x"735281cf",
  4230 => x"880851fe",
  4231 => x"a03f833d",
  4232 => x"0d04fe3d",
  4233 => x"0d755374",
  4234 => x"5281cf88",
  4235 => x"0851fdbc",
  4236 => x"3f843d0d",
  4237 => x"04803d0d",
  4238 => x"81cf8808",
  4239 => x"51fcdb3f",
  4240 => x"823d0d04",
  4241 => x"ff3d0d73",
  4242 => x"5281cf88",
  4243 => x"0851feec",
  4244 => x"3f833d0d",
  4245 => x"04fc3d0d",
  4246 => x"800b81f2",
  4247 => x"e40c7852",
  4248 => x"77519caa",
  4249 => x"3fb00854",
  4250 => x"b008ff2e",
  4251 => x"883873b0",
  4252 => x"0c863d0d",
  4253 => x"0481f2e4",
  4254 => x"08557480",
  4255 => x"2ef03876",
  4256 => x"75710c53",
  4257 => x"73b00c86",
  4258 => x"3d0d049b",
  4259 => x"fc3f04fc",
  4260 => x"3d0d7670",
  4261 => x"79707307",
  4262 => x"83065454",
  4263 => x"54557080",
  4264 => x"c3387170",
  4265 => x"08700970",
  4266 => x"f7fbfdff",
  4267 => x"130670f8",
  4268 => x"84828180",
  4269 => x"06515153",
  4270 => x"535470a6",
  4271 => x"38841472",
  4272 => x"74708405",
  4273 => x"560c7008",
  4274 => x"700970f7",
  4275 => x"fbfdff13",
  4276 => x"0670f884",
  4277 => x"82818006",
  4278 => x"51515353",
  4279 => x"5470802e",
  4280 => x"dc387352",
  4281 => x"71708105",
  4282 => x"53335170",
  4283 => x"73708105",
  4284 => x"553470f0",
  4285 => x"3874b00c",
  4286 => x"863d0d04",
  4287 => x"fd3d0d75",
  4288 => x"70718306",
  4289 => x"53555270",
  4290 => x"b8387170",
  4291 => x"087009f7",
  4292 => x"fbfdff12",
  4293 => x"0670f884",
  4294 => x"82818006",
  4295 => x"51515253",
  4296 => x"709d3884",
  4297 => x"13700870",
  4298 => x"09f7fbfd",
  4299 => x"ff120670",
  4300 => x"f8848281",
  4301 => x"80065151",
  4302 => x"52537080",
  4303 => x"2ee53872",
  4304 => x"52713351",
  4305 => x"70802e8a",
  4306 => x"38811270",
  4307 => x"33525270",
  4308 => x"f8387174",
  4309 => x"31b00c85",
  4310 => x"3d0d04fa",
  4311 => x"3d0d787a",
  4312 => x"7c705455",
  4313 => x"55527280",
  4314 => x"2e80d938",
  4315 => x"71740783",
  4316 => x"06517080",
  4317 => x"2e80d438",
  4318 => x"ff135372",
  4319 => x"ff2eb138",
  4320 => x"71337433",
  4321 => x"56517471",
  4322 => x"2e098106",
  4323 => x"a9387280",
  4324 => x"2e818738",
  4325 => x"7081ff06",
  4326 => x"5170802e",
  4327 => x"80fc3881",
  4328 => x"128115ff",
  4329 => x"15555552",
  4330 => x"72ff2e09",
  4331 => x"8106d138",
  4332 => x"71337433",
  4333 => x"56517081",
  4334 => x"ff067581",
  4335 => x"ff067171",
  4336 => x"31515252",
  4337 => x"70b00c88",
  4338 => x"3d0d0471",
  4339 => x"74575583",
  4340 => x"73278838",
  4341 => x"71087408",
  4342 => x"2e883874",
  4343 => x"765552ff",
  4344 => x"9739fc13",
  4345 => x"5372802e",
  4346 => x"b1387408",
  4347 => x"7009f7fb",
  4348 => x"fdff1206",
  4349 => x"70f88482",
  4350 => x"81800651",
  4351 => x"5151709a",
  4352 => x"38841584",
  4353 => x"17575583",
  4354 => x"7327d038",
  4355 => x"74087608",
  4356 => x"2ed03874",
  4357 => x"765552fe",
  4358 => x"df39800b",
  4359 => x"b00c883d",
  4360 => x"0d04f33d",
  4361 => x"0d606264",
  4362 => x"725a5a5e",
  4363 => x"5e805c76",
  4364 => x"70810558",
  4365 => x"3381cca9",
  4366 => x"11337083",
  4367 => x"2a708106",
  4368 => x"51555556",
  4369 => x"72e93875",
  4370 => x"ad2e8288",
  4371 => x"3875ab2e",
  4372 => x"82843877",
  4373 => x"30707907",
  4374 => x"80257990",
  4375 => x"32703070",
  4376 => x"72078025",
  4377 => x"73075357",
  4378 => x"57515372",
  4379 => x"802e8738",
  4380 => x"75b02e81",
  4381 => x"eb38778a",
  4382 => x"38885875",
  4383 => x"b02e8338",
  4384 => x"8a58810a",
  4385 => x"5a7b8438",
  4386 => x"fe0a5a77",
  4387 => x"527951f6",
  4388 => x"be3fb008",
  4389 => x"78537a52",
  4390 => x"5bf68f3f",
  4391 => x"b0085a80",
  4392 => x"7081cca9",
  4393 => x"18337082",
  4394 => x"2a708106",
  4395 => x"5156565a",
  4396 => x"5572802e",
  4397 => x"80c138d0",
  4398 => x"16567578",
  4399 => x"2580d738",
  4400 => x"80792475",
  4401 => x"7b260753",
  4402 => x"72933874",
  4403 => x"7a2e80eb",
  4404 => x"387a7625",
  4405 => x"80ed3872",
  4406 => x"802e80e7",
  4407 => x"38ff7770",
  4408 => x"81055933",
  4409 => x"575981cc",
  4410 => x"a9163370",
  4411 => x"822a7081",
  4412 => x"06515454",
  4413 => x"72c13873",
  4414 => x"83065372",
  4415 => x"802e9738",
  4416 => x"738106c9",
  4417 => x"17555372",
  4418 => x"8538ffa9",
  4419 => x"16547356",
  4420 => x"777624ff",
  4421 => x"ab388079",
  4422 => x"2480f038",
  4423 => x"7b802e84",
  4424 => x"38743055",
  4425 => x"7c802e8c",
  4426 => x"38ff1753",
  4427 => x"7883387d",
  4428 => x"53727d0c",
  4429 => x"74b00c8f",
  4430 => x"3d0d0481",
  4431 => x"53757b24",
  4432 => x"ff953881",
  4433 => x"75792917",
  4434 => x"78708105",
  4435 => x"5a335856",
  4436 => x"59ff9339",
  4437 => x"815c7670",
  4438 => x"81055833",
  4439 => x"56fdf439",
  4440 => x"80773354",
  4441 => x"547280f8",
  4442 => x"2eb23872",
  4443 => x"80d83270",
  4444 => x"30708025",
  4445 => x"76075151",
  4446 => x"5372802e",
  4447 => x"fdf83881",
  4448 => x"17338218",
  4449 => x"58569058",
  4450 => x"fdf83981",
  4451 => x"0a557b84",
  4452 => x"38fe0a55",
  4453 => x"7f53a273",
  4454 => x"0cff8939",
  4455 => x"8154cc39",
  4456 => x"fd3d0d77",
  4457 => x"54765375",
  4458 => x"5281cf88",
  4459 => x"0851fcf2",
  4460 => x"3f853d0d",
  4461 => x"04f33d0d",
  4462 => x"60626472",
  4463 => x"5a5a5d5d",
  4464 => x"805e7670",
  4465 => x"81055833",
  4466 => x"81cca911",
  4467 => x"3370832a",
  4468 => x"70810651",
  4469 => x"55555672",
  4470 => x"e93875ad",
  4471 => x"2e81ff38",
  4472 => x"75ab2e81",
  4473 => x"fb387730",
  4474 => x"70790780",
  4475 => x"25799032",
  4476 => x"70307072",
  4477 => x"07802573",
  4478 => x"07535757",
  4479 => x"51537280",
  4480 => x"2e873875",
  4481 => x"b02e81e2",
  4482 => x"38778a38",
  4483 => x"885875b0",
  4484 => x"2e83388a",
  4485 => x"587752ff",
  4486 => x"51f38f3f",
  4487 => x"b0087853",
  4488 => x"5aff51f3",
  4489 => x"aa3fb008",
  4490 => x"5b80705a",
  4491 => x"5581cca9",
  4492 => x"16337082",
  4493 => x"2a708106",
  4494 => x"51545472",
  4495 => x"802e80c1",
  4496 => x"38d01656",
  4497 => x"75782580",
  4498 => x"d7388079",
  4499 => x"24757b26",
  4500 => x"07537293",
  4501 => x"38747a2e",
  4502 => x"80eb387a",
  4503 => x"762580ed",
  4504 => x"3872802e",
  4505 => x"80e738ff",
  4506 => x"77708105",
  4507 => x"59335759",
  4508 => x"81cca916",
  4509 => x"3370822a",
  4510 => x"70810651",
  4511 => x"545472c1",
  4512 => x"38738306",
  4513 => x"5372802e",
  4514 => x"97387381",
  4515 => x"06c91755",
  4516 => x"53728538",
  4517 => x"ffa91654",
  4518 => x"73567776",
  4519 => x"24ffab38",
  4520 => x"80792481",
  4521 => x"89387d80",
  4522 => x"2e843874",
  4523 => x"30557b80",
  4524 => x"2e8c38ff",
  4525 => x"17537883",
  4526 => x"387c5372",
  4527 => x"7c0c74b0",
  4528 => x"0c8f3d0d",
  4529 => x"04815375",
  4530 => x"7b24ff95",
  4531 => x"38817579",
  4532 => x"29177870",
  4533 => x"81055a33",
  4534 => x"585659ff",
  4535 => x"9339815e",
  4536 => x"76708105",
  4537 => x"583356fd",
  4538 => x"fd398077",
  4539 => x"33545472",
  4540 => x"80f82e80",
  4541 => x"c3387280",
  4542 => x"d8327030",
  4543 => x"70802576",
  4544 => x"07515153",
  4545 => x"72802efe",
  4546 => x"80388117",
  4547 => x"33821858",
  4548 => x"56907053",
  4549 => x"58ff51f1",
  4550 => x"913fb008",
  4551 => x"78535aff",
  4552 => x"51f1ac3f",
  4553 => x"b0085b80",
  4554 => x"705a55fe",
  4555 => x"8039ff60",
  4556 => x"5455a273",
  4557 => x"0cfef739",
  4558 => x"8154ffba",
  4559 => x"39fd3d0d",
  4560 => x"77547653",
  4561 => x"755281cf",
  4562 => x"880851fc",
  4563 => x"e83f853d",
  4564 => x"0d04f33d",
  4565 => x"0d7f618b",
  4566 => x"1170f806",
  4567 => x"5c55555e",
  4568 => x"72962683",
  4569 => x"38905980",
  4570 => x"7924747a",
  4571 => x"26075380",
  4572 => x"5472742e",
  4573 => x"09810680",
  4574 => x"cb387d51",
  4575 => x"8bca3f78",
  4576 => x"83f72680",
  4577 => x"c6387883",
  4578 => x"2a701010",
  4579 => x"1081d6c4",
  4580 => x"058c1108",
  4581 => x"59595a76",
  4582 => x"782e83b0",
  4583 => x"38841708",
  4584 => x"fc06568c",
  4585 => x"17088818",
  4586 => x"08718c12",
  4587 => x"0c88120c",
  4588 => x"58751784",
  4589 => x"11088107",
  4590 => x"84120c53",
  4591 => x"7d518b89",
  4592 => x"3f881754",
  4593 => x"73b00c8f",
  4594 => x"3d0d0478",
  4595 => x"892a7983",
  4596 => x"2a5b5372",
  4597 => x"802ebf38",
  4598 => x"78862ab8",
  4599 => x"055a8473",
  4600 => x"27b43880",
  4601 => x"db135a94",
  4602 => x"7327ab38",
  4603 => x"788c2a80",
  4604 => x"ee055a80",
  4605 => x"d473279e",
  4606 => x"38788f2a",
  4607 => x"80f7055a",
  4608 => x"82d47327",
  4609 => x"91387892",
  4610 => x"2a80fc05",
  4611 => x"5a8ad473",
  4612 => x"27843880",
  4613 => x"fe5a7910",
  4614 => x"101081d6",
  4615 => x"c4058c11",
  4616 => x"08585576",
  4617 => x"752ea338",
  4618 => x"841708fc",
  4619 => x"06707a31",
  4620 => x"5556738f",
  4621 => x"2488d538",
  4622 => x"738025fe",
  4623 => x"e6388c17",
  4624 => x"08577675",
  4625 => x"2e098106",
  4626 => x"df38811a",
  4627 => x"5a81d6d4",
  4628 => x"08577681",
  4629 => x"d6cc2e82",
  4630 => x"c0388417",
  4631 => x"08fc0670",
  4632 => x"7a315556",
  4633 => x"738f2481",
  4634 => x"f93881d6",
  4635 => x"cc0b81d6",
  4636 => x"d80c81d6",
  4637 => x"cc0b81d6",
  4638 => x"d40c7380",
  4639 => x"25feb238",
  4640 => x"83ff7627",
  4641 => x"83df3875",
  4642 => x"892a7683",
  4643 => x"2a555372",
  4644 => x"802ebf38",
  4645 => x"75862ab8",
  4646 => x"05548473",
  4647 => x"27b43880",
  4648 => x"db135494",
  4649 => x"7327ab38",
  4650 => x"758c2a80",
  4651 => x"ee055480",
  4652 => x"d473279e",
  4653 => x"38758f2a",
  4654 => x"80f70554",
  4655 => x"82d47327",
  4656 => x"91387592",
  4657 => x"2a80fc05",
  4658 => x"548ad473",
  4659 => x"27843880",
  4660 => x"fe547310",
  4661 => x"101081d6",
  4662 => x"c4058811",
  4663 => x"08565874",
  4664 => x"782e86cf",
  4665 => x"38841508",
  4666 => x"fc065375",
  4667 => x"73278d38",
  4668 => x"88150855",
  4669 => x"74782e09",
  4670 => x"8106ea38",
  4671 => x"8c150881",
  4672 => x"d6c40b84",
  4673 => x"0508718c",
  4674 => x"1a0c7688",
  4675 => x"1a0c7888",
  4676 => x"130c788c",
  4677 => x"180c5d58",
  4678 => x"7953807a",
  4679 => x"2483e638",
  4680 => x"72822c81",
  4681 => x"712b5c53",
  4682 => x"7a7c2681",
  4683 => x"98387b7b",
  4684 => x"06537282",
  4685 => x"f13879fc",
  4686 => x"0684055a",
  4687 => x"7a10707d",
  4688 => x"06545b72",
  4689 => x"82e03884",
  4690 => x"1a5af139",
  4691 => x"88178c11",
  4692 => x"08585876",
  4693 => x"782e0981",
  4694 => x"06fcc238",
  4695 => x"821a5afd",
  4696 => x"ec397817",
  4697 => x"79810784",
  4698 => x"190c7081",
  4699 => x"d6d80c70",
  4700 => x"81d6d40c",
  4701 => x"81d6cc0b",
  4702 => x"8c120c8c",
  4703 => x"11088812",
  4704 => x"0c748107",
  4705 => x"84120c74",
  4706 => x"1175710c",
  4707 => x"51537d51",
  4708 => x"87b73f88",
  4709 => x"1754fcac",
  4710 => x"3981d6c4",
  4711 => x"0b840508",
  4712 => x"7a545c79",
  4713 => x"8025fef8",
  4714 => x"3882da39",
  4715 => x"7a097c06",
  4716 => x"7081d6c4",
  4717 => x"0b84050c",
  4718 => x"5c7a105b",
  4719 => x"7a7c2685",
  4720 => x"387a85b8",
  4721 => x"3881d6c4",
  4722 => x"0b880508",
  4723 => x"70841208",
  4724 => x"fc06707c",
  4725 => x"317c7226",
  4726 => x"8f722507",
  4727 => x"57575c5d",
  4728 => x"5572802e",
  4729 => x"80db3879",
  4730 => x"7a1681d6",
  4731 => x"bc081b90",
  4732 => x"115a5557",
  4733 => x"5b81d6b8",
  4734 => x"08ff2e88",
  4735 => x"38a08f13",
  4736 => x"e0800657",
  4737 => x"76527d51",
  4738 => x"86c03fb0",
  4739 => x"0854b008",
  4740 => x"ff2e9038",
  4741 => x"b0087627",
  4742 => x"82993874",
  4743 => x"81d6c42e",
  4744 => x"82913881",
  4745 => x"d6c40b88",
  4746 => x"05085584",
  4747 => x"1508fc06",
  4748 => x"707a317a",
  4749 => x"72268f72",
  4750 => x"25075255",
  4751 => x"537283e6",
  4752 => x"38747981",
  4753 => x"0784170c",
  4754 => x"79167081",
  4755 => x"d6c40b88",
  4756 => x"050c7581",
  4757 => x"0784120c",
  4758 => x"547e5257",
  4759 => x"85eb3f88",
  4760 => x"1754fae0",
  4761 => x"3975832a",
  4762 => x"70545480",
  4763 => x"7424819b",
  4764 => x"3872822c",
  4765 => x"81712b81",
  4766 => x"d6c80807",
  4767 => x"7081d6c4",
  4768 => x"0b84050c",
  4769 => x"75101010",
  4770 => x"81d6c405",
  4771 => x"88110858",
  4772 => x"5a5d5377",
  4773 => x"8c180c74",
  4774 => x"88180c76",
  4775 => x"88190c76",
  4776 => x"8c160cfc",
  4777 => x"f339797a",
  4778 => x"10101081",
  4779 => x"d6c40570",
  4780 => x"57595d8c",
  4781 => x"15085776",
  4782 => x"752ea338",
  4783 => x"841708fc",
  4784 => x"06707a31",
  4785 => x"5556738f",
  4786 => x"2483ca38",
  4787 => x"73802584",
  4788 => x"81388c17",
  4789 => x"08577675",
  4790 => x"2e098106",
  4791 => x"df388815",
  4792 => x"811b7083",
  4793 => x"06555b55",
  4794 => x"72c9387c",
  4795 => x"83065372",
  4796 => x"802efdb8",
  4797 => x"38ff1df8",
  4798 => x"19595d88",
  4799 => x"1808782e",
  4800 => x"ea38fdb5",
  4801 => x"39831a53",
  4802 => x"fc963983",
  4803 => x"1470822c",
  4804 => x"81712b81",
  4805 => x"d6c80807",
  4806 => x"7081d6c4",
  4807 => x"0b84050c",
  4808 => x"76101010",
  4809 => x"81d6c405",
  4810 => x"88110859",
  4811 => x"5b5e5153",
  4812 => x"fee13981",
  4813 => x"d6880817",
  4814 => x"58b00876",
  4815 => x"2e818d38",
  4816 => x"81d6b808",
  4817 => x"ff2e83ec",
  4818 => x"38737631",
  4819 => x"1881d688",
  4820 => x"0c738706",
  4821 => x"70575372",
  4822 => x"802e8838",
  4823 => x"88733170",
  4824 => x"15555676",
  4825 => x"149fff06",
  4826 => x"a0807131",
  4827 => x"1770547f",
  4828 => x"53575383",
  4829 => x"d53fb008",
  4830 => x"53b008ff",
  4831 => x"2e81a038",
  4832 => x"81d68808",
  4833 => x"167081d6",
  4834 => x"880c7475",
  4835 => x"81d6c40b",
  4836 => x"88050c74",
  4837 => x"76311870",
  4838 => x"81075155",
  4839 => x"56587b81",
  4840 => x"d6c42e83",
  4841 => x"9c38798f",
  4842 => x"2682cb38",
  4843 => x"810b8415",
  4844 => x"0c841508",
  4845 => x"fc06707a",
  4846 => x"317a7226",
  4847 => x"8f722507",
  4848 => x"52555372",
  4849 => x"802efcf9",
  4850 => x"3880db39",
  4851 => x"b0089fff",
  4852 => x"065372fe",
  4853 => x"eb387781",
  4854 => x"d6880c81",
  4855 => x"d6c40b88",
  4856 => x"05087b18",
  4857 => x"81078412",
  4858 => x"0c5581d6",
  4859 => x"b4087827",
  4860 => x"86387781",
  4861 => x"d6b40c81",
  4862 => x"d6b00878",
  4863 => x"27fcac38",
  4864 => x"7781d6b0",
  4865 => x"0c841508",
  4866 => x"fc06707a",
  4867 => x"317a7226",
  4868 => x"8f722507",
  4869 => x"52555372",
  4870 => x"802efca5",
  4871 => x"38883980",
  4872 => x"745456fe",
  4873 => x"db397d51",
  4874 => x"829f3f80",
  4875 => x"0bb00c8f",
  4876 => x"3d0d0473",
  4877 => x"53807424",
  4878 => x"a9387282",
  4879 => x"2c81712b",
  4880 => x"81d6c808",
  4881 => x"077081d6",
  4882 => x"c40b8405",
  4883 => x"0c5d5377",
  4884 => x"8c180c74",
  4885 => x"88180c76",
  4886 => x"88190c76",
  4887 => x"8c160cf9",
  4888 => x"b7398314",
  4889 => x"70822c81",
  4890 => x"712b81d6",
  4891 => x"c8080770",
  4892 => x"81d6c40b",
  4893 => x"84050c5e",
  4894 => x"5153d439",
  4895 => x"7b7b0653",
  4896 => x"72fca338",
  4897 => x"841a7b10",
  4898 => x"5c5af139",
  4899 => x"ff1a8111",
  4900 => x"515af7b9",
  4901 => x"39781779",
  4902 => x"81078419",
  4903 => x"0c8c1808",
  4904 => x"88190871",
  4905 => x"8c120c88",
  4906 => x"120c5970",
  4907 => x"81d6d80c",
  4908 => x"7081d6d4",
  4909 => x"0c81d6cc",
  4910 => x"0b8c120c",
  4911 => x"8c110888",
  4912 => x"120c7481",
  4913 => x"0784120c",
  4914 => x"74117571",
  4915 => x"0c5153f9",
  4916 => x"bd397517",
  4917 => x"84110881",
  4918 => x"0784120c",
  4919 => x"538c1708",
  4920 => x"88180871",
  4921 => x"8c120c88",
  4922 => x"120c587d",
  4923 => x"5180da3f",
  4924 => x"881754f5",
  4925 => x"cf397284",
  4926 => x"150cf41a",
  4927 => x"f8067084",
  4928 => x"1e088106",
  4929 => x"07841e0c",
  4930 => x"701d545b",
  4931 => x"850b8414",
  4932 => x"0c850b88",
  4933 => x"140c8f7b",
  4934 => x"27fdcf38",
  4935 => x"881c527d",
  4936 => x"5182903f",
  4937 => x"81d6c40b",
  4938 => x"88050881",
  4939 => x"d6880859",
  4940 => x"55fdb739",
  4941 => x"7781d688",
  4942 => x"0c7381d6",
  4943 => x"b80cfc91",
  4944 => x"39728415",
  4945 => x"0cfda339",
  4946 => x"0404fd3d",
  4947 => x"0d800b81",
  4948 => x"f2e40c76",
  4949 => x"5186cb3f",
  4950 => x"b00853b0",
  4951 => x"08ff2e88",
  4952 => x"3872b00c",
  4953 => x"853d0d04",
  4954 => x"81f2e408",
  4955 => x"5473802e",
  4956 => x"f0387574",
  4957 => x"710c5272",
  4958 => x"b00c853d",
  4959 => x"0d04fb3d",
  4960 => x"0d777052",
  4961 => x"56c23f81",
  4962 => x"d6c40b88",
  4963 => x"05088411",
  4964 => x"08fc0670",
  4965 => x"7b319fef",
  4966 => x"05e08006",
  4967 => x"e0800556",
  4968 => x"5653a080",
  4969 => x"74249438",
  4970 => x"80527551",
  4971 => x"ff9c3f81",
  4972 => x"d6cc0815",
  4973 => x"5372b008",
  4974 => x"2e8f3875",
  4975 => x"51ff8a3f",
  4976 => x"805372b0",
  4977 => x"0c873d0d",
  4978 => x"04733052",
  4979 => x"7551fefa",
  4980 => x"3fb008ff",
  4981 => x"2ea83881",
  4982 => x"d6c40b88",
  4983 => x"05087575",
  4984 => x"31810784",
  4985 => x"120c5381",
  4986 => x"d6880874",
  4987 => x"3181d688",
  4988 => x"0c7551fe",
  4989 => x"d43f810b",
  4990 => x"b00c873d",
  4991 => x"0d048052",
  4992 => x"7551fec6",
  4993 => x"3f81d6c4",
  4994 => x"0b880508",
  4995 => x"b0087131",
  4996 => x"56538f75",
  4997 => x"25ffa438",
  4998 => x"b00881d6",
  4999 => x"b8083181",
  5000 => x"d6880c74",
  5001 => x"81078414",
  5002 => x"0c7551fe",
  5003 => x"9c3f8053",
  5004 => x"ff9039f6",
  5005 => x"3d0d7c7e",
  5006 => x"545b7280",
  5007 => x"2e828338",
  5008 => x"7a51fe84",
  5009 => x"3ff81384",
  5010 => x"110870fe",
  5011 => x"06701384",
  5012 => x"1108fc06",
  5013 => x"5d585954",
  5014 => x"5881d6cc",
  5015 => x"08752e82",
  5016 => x"de387884",
  5017 => x"160c8073",
  5018 => x"8106545a",
  5019 => x"727a2e81",
  5020 => x"d5387815",
  5021 => x"84110881",
  5022 => x"06515372",
  5023 => x"a0387817",
  5024 => x"577981e6",
  5025 => x"38881508",
  5026 => x"537281d6",
  5027 => x"cc2e82f9",
  5028 => x"388c1508",
  5029 => x"708c150c",
  5030 => x"7388120c",
  5031 => x"56768107",
  5032 => x"84190c76",
  5033 => x"1877710c",
  5034 => x"53798191",
  5035 => x"3883ff77",
  5036 => x"2781c838",
  5037 => x"76892a77",
  5038 => x"832a5653",
  5039 => x"72802ebf",
  5040 => x"3876862a",
  5041 => x"b8055584",
  5042 => x"7327b438",
  5043 => x"80db1355",
  5044 => x"947327ab",
  5045 => x"38768c2a",
  5046 => x"80ee0555",
  5047 => x"80d47327",
  5048 => x"9e38768f",
  5049 => x"2a80f705",
  5050 => x"5582d473",
  5051 => x"27913876",
  5052 => x"922a80fc",
  5053 => x"05558ad4",
  5054 => x"73278438",
  5055 => x"80fe5574",
  5056 => x"10101081",
  5057 => x"d6c40588",
  5058 => x"11085556",
  5059 => x"73762e82",
  5060 => x"b3388414",
  5061 => x"08fc0653",
  5062 => x"7673278d",
  5063 => x"38881408",
  5064 => x"5473762e",
  5065 => x"098106ea",
  5066 => x"388c1408",
  5067 => x"708c1a0c",
  5068 => x"74881a0c",
  5069 => x"7888120c",
  5070 => x"56778c15",
  5071 => x"0c7a51fc",
  5072 => x"883f8c3d",
  5073 => x"0d047708",
  5074 => x"78713159",
  5075 => x"77058819",
  5076 => x"08545772",
  5077 => x"81d6cc2e",
  5078 => x"80e0388c",
  5079 => x"1808708c",
  5080 => x"150c7388",
  5081 => x"120c56fe",
  5082 => x"89398815",
  5083 => x"088c1608",
  5084 => x"708c130c",
  5085 => x"5788170c",
  5086 => x"fea33976",
  5087 => x"832a7054",
  5088 => x"55807524",
  5089 => x"81983872",
  5090 => x"822c8171",
  5091 => x"2b81d6c8",
  5092 => x"080781d6",
  5093 => x"c40b8405",
  5094 => x"0c537410",
  5095 => x"101081d6",
  5096 => x"c4058811",
  5097 => x"08555675",
  5098 => x"8c190c73",
  5099 => x"88190c77",
  5100 => x"88170c77",
  5101 => x"8c150cff",
  5102 => x"8439815a",
  5103 => x"fdb43978",
  5104 => x"17738106",
  5105 => x"54577298",
  5106 => x"38770878",
  5107 => x"71315977",
  5108 => x"058c1908",
  5109 => x"881a0871",
  5110 => x"8c120c88",
  5111 => x"120c5757",
  5112 => x"76810784",
  5113 => x"190c7781",
  5114 => x"d6c40b88",
  5115 => x"050c81d6",
  5116 => x"c0087726",
  5117 => x"fec73881",
  5118 => x"d6bc0852",
  5119 => x"7a51fafe",
  5120 => x"3f7a51fa",
  5121 => x"c43ffeba",
  5122 => x"3981788c",
  5123 => x"150c7888",
  5124 => x"150c738c",
  5125 => x"1a0c7388",
  5126 => x"1a0c5afd",
  5127 => x"80398315",
  5128 => x"70822c81",
  5129 => x"712b81d6",
  5130 => x"c8080781",
  5131 => x"d6c40b84",
  5132 => x"050c5153",
  5133 => x"74101010",
  5134 => x"81d6c405",
  5135 => x"88110855",
  5136 => x"56fee439",
  5137 => x"74538075",
  5138 => x"24a73872",
  5139 => x"822c8171",
  5140 => x"2b81d6c8",
  5141 => x"080781d6",
  5142 => x"c40b8405",
  5143 => x"0c53758c",
  5144 => x"190c7388",
  5145 => x"190c7788",
  5146 => x"170c778c",
  5147 => x"150cfdcd",
  5148 => x"39831570",
  5149 => x"822c8171",
  5150 => x"2b81d6c8",
  5151 => x"080781d6",
  5152 => x"c40b8405",
  5153 => x"0c5153d6",
  5154 => x"39810bb0",
  5155 => x"0c04803d",
  5156 => x"0d72812e",
  5157 => x"8938800b",
  5158 => x"b00c823d",
  5159 => x"0d047351",
  5160 => x"b23ffe3d",
  5161 => x"0d81f2e0",
  5162 => x"0851708a",
  5163 => x"3881f2e8",
  5164 => x"7081f2e0",
  5165 => x"0c517075",
  5166 => x"125252ff",
  5167 => x"537087fb",
  5168 => x"80802688",
  5169 => x"387081f2",
  5170 => x"e00c7153",
  5171 => x"72b00c84",
  5172 => x"3d0d0400",
  5173 => x"ff390000",
  5174 => x"00000000",
  5175 => x"00000000",
  5176 => x"00000000",
  5177 => x"00000000",
  5178 => x"00cac5ca",
  5179 => x"c5c0c0c0",
  5180 => x"c0c0c0c0",
  5181 => x"c0c0c0cf",
  5182 => x"cfcfcf00",
  5183 => x"00000f0f",
  5184 => x"0f0f8f8f",
  5185 => x"cfcfcfcf",
  5186 => x"cfcf4f0f",
  5187 => x"0f0f0000",
  5188 => x"cfcfcfcf",
  5189 => x"0f0f0f0f",
  5190 => x"0f0f0f0f",
  5191 => x"0f0ffefe",
  5192 => x"fefc0000",
  5193 => x"cfcfcfcf",
  5194 => x"cfcfcfcf",
  5195 => x"cfcfcfcf",
  5196 => x"cfffff7e",
  5197 => x"7e000000",
  5198 => x"00000000",
  5199 => x"00000000",
  5200 => x"00000000",
  5201 => x"00003f3f",
  5202 => x"3f3f0101",
  5203 => x"01010101",
  5204 => x"01010101",
  5205 => x"3f3f3f3f",
  5206 => x"0000383c",
  5207 => x"3e3e3f3f",
  5208 => x"3f3b3b39",
  5209 => x"39383838",
  5210 => x"38383800",
  5211 => x"003f3f3f",
  5212 => x"3f383838",
  5213 => x"38383838",
  5214 => x"38383c3f",
  5215 => x"3f1f0f00",
  5216 => x"003f3f3f",
  5217 => x"3f030303",
  5218 => x"03030303",
  5219 => x"03033f3f",
  5220 => x"3f3e0000",
  5221 => x"00000000",
  5222 => x"00000000",
  5223 => x"00000000",
  5224 => x"00000000",
  5225 => x"00000000",
  5226 => x"00000000",
  5227 => x"00000000",
  5228 => x"00000000",
  5229 => x"00000000",
  5230 => x"00000000",
  5231 => x"00000000",
  5232 => x"00000000",
  5233 => x"00000000",
  5234 => x"00000000",
  5235 => x"00000000",
  5236 => x"00000000",
  5237 => x"00000000",
  5238 => x"00000000",
  5239 => x"00000000",
  5240 => x"00000000",
  5241 => x"00000000",
  5242 => x"00000000",
  5243 => x"00000000",
  5244 => x"00000000",
  5245 => x"8080c0c0",
  5246 => x"e0e06000",
  5247 => x"00000000",
  5248 => x"00000000",
  5249 => x"00000000",
  5250 => x"00000000",
  5251 => x"00000000",
  5252 => x"00000000",
  5253 => x"00000000",
  5254 => x"00000000",
  5255 => x"00000000",
  5256 => x"00000000",
  5257 => x"00000000",
  5258 => x"00000000",
  5259 => x"00000000",
  5260 => x"00000000",
  5261 => x"00000000",
  5262 => x"00000000",
  5263 => x"00000000",
  5264 => x"00000000",
  5265 => x"00000000",
  5266 => x"00000000",
  5267 => x"806098ee",
  5268 => x"77bbddec",
  5269 => x"ee6e0200",
  5270 => x"00000000",
  5271 => x"00e08080",
  5272 => x"e00000e0",
  5273 => x"a0a00000",
  5274 => x"e0000000",
  5275 => x"00e0c000",
  5276 => x"c0e00000",
  5277 => x"e08080e0",
  5278 => x"0000c020",
  5279 => x"20c00000",
  5280 => x"e0000000",
  5281 => x"20e02000",
  5282 => x"0020a060",
  5283 => x"20000000",
  5284 => x"00000000",
  5285 => x"00000000",
  5286 => x"00000000",
  5287 => x"00000000",
  5288 => x"00000000",
  5289 => x"00000000",
  5290 => x"00030007",
  5291 => x"00070701",
  5292 => x"00000000",
  5293 => x"00000000",
  5294 => x"00000300",
  5295 => x"c0030000",
  5296 => x"034242c0",
  5297 => x"00c34242",
  5298 => x"0000c380",
  5299 => x"01c00340",
  5300 => x"c04300c0",
  5301 => x"43408001",
  5302 => x"c20201c0",
  5303 => x"00c38202",
  5304 => x"80c00300",
  5305 => x"00c04342",
  5306 => x"8202c040",
  5307 => x"40800000",
  5308 => x"c0404000",
  5309 => x"80404000",
  5310 => x"00c04040",
  5311 => x"8000c040",
  5312 => x"4000c080",
  5313 => x"00c00000",
  5314 => x"00000000",
  5315 => x"00000000",
  5316 => x"00000000",
  5317 => x"00000000",
  5318 => x"00ff0000",
  5319 => x"0000c645",
  5320 => x"44800785",
  5321 => x"45408007",
  5322 => x"80424700",
  5323 => x"80474000",
  5324 => x"07c14344",
  5325 => x"00c38404",
  5326 => x"c30007c1",
  5327 => x"42418700",
  5328 => x"80404784",
  5329 => x"04c34047",
  5330 => x"8101c640",
  5331 => x"40070505",
  5332 => x"00040502",
  5333 => x"00000704",
  5334 => x"04030007",
  5335 => x"05050007",
  5336 => x"00020700",
  5337 => x"00000000",
  5338 => x"00000000",
  5339 => x"00000000",
  5340 => x"00000000",
  5341 => x"0000ff00",
  5342 => x"00000007",
  5343 => x"01030500",
  5344 => x"03040403",
  5345 => x"00040502",
  5346 => x"00040502",
  5347 => x"00000705",
  5348 => x"05000700",
  5349 => x"02070000",
  5350 => x"07040403",
  5351 => x"00030404",
  5352 => x"03000701",
  5353 => x"03050007",
  5354 => x"01010000",
  5355 => x"00000000",
  5356 => x"00000000",
  5357 => x"00000000",
  5358 => x"00000000",
  5359 => x"00000000",
  5360 => x"71756974",
  5361 => x"00000000",
  5362 => x"68656c70",
  5363 => x"00000000",
  5364 => x"0a307800",
  5365 => x"69326320",
  5366 => x"464d430a",
  5367 => x"00000000",
  5368 => x"61646472",
  5369 => x"6573733a",
  5370 => x"20307800",
  5371 => x"2020202d",
  5372 => x"2d3e2020",
  5373 => x"2041434b",
  5374 => x"0a000000",
  5375 => x"72656164",
  5376 => x"20646174",
  5377 => x"61202800",
  5378 => x"20627974",
  5379 => x"65732920",
  5380 => x"66726f6d",
  5381 => x"20493243",
  5382 => x"2d616464",
  5383 => x"72657373",
  5384 => x"20307800",
  5385 => x"0a0a0000",
  5386 => x"6e6f6163",
  5387 => x"6b200000",
  5388 => x"6368726f",
  5389 => x"6e74656c",
  5390 => x"20726567",
  5391 => x"20307800",
  5392 => x"3a203078",
  5393 => x"00000000",
  5394 => x"206e6163",
  5395 => x"6b000000",
  5396 => x"6572726f",
  5397 => x"7220286e",
  5398 => x"61636b29",
  5399 => x"0a000000",
  5400 => x"0a202063",
  5401 => x"68616e6e",
  5402 => x"656c2033",
  5403 => x"20696e70",
  5404 => x"7574206f",
  5405 => x"76657266",
  5406 => x"6c6f7700",
  5407 => x"0a202063",
  5408 => x"68616e6e",
  5409 => x"656c2032",
  5410 => x"20696e70",
  5411 => x"7574206f",
  5412 => x"76657266",
  5413 => x"6c6f7700",
  5414 => x"0a202063",
  5415 => x"68616e6e",
  5416 => x"656c2031",
  5417 => x"20696e70",
  5418 => x"7574206f",
  5419 => x"76657266",
  5420 => x"6c6f7700",
  5421 => x"0a202063",
  5422 => x"68616e6e",
  5423 => x"656c2030",
  5424 => x"20696e70",
  5425 => x"7574206f",
  5426 => x"76657266",
  5427 => x"6c6f7700",
  5428 => x"0a202063",
  5429 => x"68616e6e",
  5430 => x"656c2033",
  5431 => x"20717561",
  5432 => x"6473756d",
  5433 => x"206f7665",
  5434 => x"72666c6f",
  5435 => x"77000000",
  5436 => x"0a202063",
  5437 => x"68616e6e",
  5438 => x"656c2032",
  5439 => x"20717561",
  5440 => x"6473756d",
  5441 => x"206f7665",
  5442 => x"72666c6f",
  5443 => x"77000000",
  5444 => x"0a202063",
  5445 => x"68616e6e",
  5446 => x"656c2031",
  5447 => x"20717561",
  5448 => x"6473756d",
  5449 => x"206f7665",
  5450 => x"72666c6f",
  5451 => x"77000000",
  5452 => x"0a202063",
  5453 => x"68616e6e",
  5454 => x"656c2030",
  5455 => x"20717561",
  5456 => x"6473756d",
  5457 => x"206f7665",
  5458 => x"72666c6f",
  5459 => x"77000000",
  5460 => x"0a202073",
  5461 => x"756d2076",
  5462 => x"616c7565",
  5463 => x"20637574",
  5464 => x"74656400",
  5465 => x"0a202063",
  5466 => x"68616e6e",
  5467 => x"656c2033",
  5468 => x"20646976",
  5469 => x"6964656e",
  5470 => x"64206375",
  5471 => x"74746564",
  5472 => x"00000000",
  5473 => x"0a202063",
  5474 => x"68616e6e",
  5475 => x"656c2033",
  5476 => x"206e6f69",
  5477 => x"73652063",
  5478 => x"6f6d7065",
  5479 => x"6e736174",
  5480 => x"696f6e20",
  5481 => x"746f2062",
  5482 => x"69670000",
  5483 => x"0a202063",
  5484 => x"68616e6e",
  5485 => x"656c2033",
  5486 => x"206e6f69",
  5487 => x"73652076",
  5488 => x"616c7565",
  5489 => x"20637574",
  5490 => x"74656400",
  5491 => x"0a202063",
  5492 => x"68616e6e",
  5493 => x"656c2032",
  5494 => x"20646976",
  5495 => x"6964656e",
  5496 => x"64206375",
  5497 => x"74746564",
  5498 => x"00000000",
  5499 => x"0a202063",
  5500 => x"68616e6e",
  5501 => x"656c2032",
  5502 => x"206e6f69",
  5503 => x"73652063",
  5504 => x"6f6d7065",
  5505 => x"6e736174",
  5506 => x"696f6e20",
  5507 => x"746f2062",
  5508 => x"69670000",
  5509 => x"0a202063",
  5510 => x"68616e6e",
  5511 => x"656c2032",
  5512 => x"206e6f69",
  5513 => x"73652076",
  5514 => x"616c7565",
  5515 => x"20637574",
  5516 => x"74656400",
  5517 => x"0a202063",
  5518 => x"68616e6e",
  5519 => x"656c2031",
  5520 => x"20646976",
  5521 => x"6964656e",
  5522 => x"64206375",
  5523 => x"74746564",
  5524 => x"00000000",
  5525 => x"0a202063",
  5526 => x"68616e6e",
  5527 => x"656c2031",
  5528 => x"206e6f69",
  5529 => x"73652063",
  5530 => x"6f6d7065",
  5531 => x"6e736174",
  5532 => x"696f6e20",
  5533 => x"746f2062",
  5534 => x"69670000",
  5535 => x"0a202063",
  5536 => x"68616e6e",
  5537 => x"656c2031",
  5538 => x"206e6f69",
  5539 => x"73652076",
  5540 => x"616c7565",
  5541 => x"20637574",
  5542 => x"74656400",
  5543 => x"0a202063",
  5544 => x"68616e6e",
  5545 => x"656c2030",
  5546 => x"20646976",
  5547 => x"6964656e",
  5548 => x"64206375",
  5549 => x"74746564",
  5550 => x"00000000",
  5551 => x"0a202063",
  5552 => x"68616e6e",
  5553 => x"656c2030",
  5554 => x"206e6f69",
  5555 => x"73652063",
  5556 => x"6f6d7065",
  5557 => x"6e736174",
  5558 => x"696f6e20",
  5559 => x"746f2062",
  5560 => x"69670000",
  5561 => x"0a202063",
  5562 => x"68616e6e",
  5563 => x"656c2030",
  5564 => x"206e6f69",
  5565 => x"73652076",
  5566 => x"616c7565",
  5567 => x"20637574",
  5568 => x"74656400",
  5569 => x"0a202073",
  5570 => x"6f667477",
  5571 => x"61726520",
  5572 => x"6572726f",
  5573 => x"72000000",
  5574 => x"0a657874",
  5575 => x"65726e61",
  5576 => x"6c20636c",
  5577 => x"6f636b20",
  5578 => x"20202020",
  5579 => x"2020203a",
  5580 => x"20000000",
  5581 => x"61637469",
  5582 => x"76650000",
  5583 => x"0a6d6963",
  5584 => x"726f7075",
  5585 => x"6c736520",
  5586 => x"736f7572",
  5587 => x"63652020",
  5588 => x"2020203a",
  5589 => x"20000000",
  5590 => x"65787465",
  5591 => x"726e616c",
  5592 => x"00000000",
  5593 => x"0a6d6963",
  5594 => x"726f7075",
  5595 => x"6c736520",
  5596 => x"6576656e",
  5597 => x"74206c69",
  5598 => x"6d69743a",
  5599 => x"20000000",
  5600 => x"0a6d6561",
  5601 => x"73757265",
  5602 => x"6d656e74",
  5603 => x"206c656e",
  5604 => x"67746820",
  5605 => x"2020203a",
  5606 => x"20000000",
  5607 => x"0a626561",
  5608 => x"6d20706f",
  5609 => x"73697469",
  5610 => x"6f6e206d",
  5611 => x"6f6e6974",
  5612 => x"6f722072",
  5613 => x"65676973",
  5614 => x"74657273",
  5615 => x"00000000",
  5616 => x"0a202020",
  5617 => x"20202020",
  5618 => x"20202020",
  5619 => x"20202020",
  5620 => x"20202020",
  5621 => x"20202020",
  5622 => x"20636861",
  5623 => x"6e6e656c",
  5624 => x"20302020",
  5625 => x"20636861",
  5626 => x"6e6e656c",
  5627 => x"20312020",
  5628 => x"20636861",
  5629 => x"6e6e656c",
  5630 => x"20322020",
  5631 => x"20636861",
  5632 => x"6e6e656c",
  5633 => x"20330000",
  5634 => x"0a202020",
  5635 => x"20202020",
  5636 => x"20202020",
  5637 => x"20202020",
  5638 => x"20202020",
  5639 => x"20202020",
  5640 => x"202d2d2d",
  5641 => x"2d20686f",
  5642 => x"72697a6f",
  5643 => x"6e74616c",
  5644 => x"202d2d2d",
  5645 => x"2d2d2020",
  5646 => x"202d2d2d",
  5647 => x"2d2d2d20",
  5648 => x"76657274",
  5649 => x"6963616c",
  5650 => x"202d2d2d",
  5651 => x"2d2d0000",
  5652 => x"0a736361",
  5653 => x"6c657220",
  5654 => x"76616c75",
  5655 => x"65732020",
  5656 => x"20202020",
  5657 => x"20202020",
  5658 => x"20000000",
  5659 => x"0a6e6f69",
  5660 => x"73652063",
  5661 => x"6f6d7065",
  5662 => x"6e736174",
  5663 => x"696f6e20",
  5664 => x"20202020",
  5665 => x"20000000",
  5666 => x"0a6d6561",
  5667 => x"73757265",
  5668 => x"6d656e74",
  5669 => x"20202020",
  5670 => x"20202020",
  5671 => x"20202020",
  5672 => x"20000000",
  5673 => x"0a73616d",
  5674 => x"706c6573",
  5675 => x"20286469",
  5676 => x"7629203a",
  5677 => x"20000000",
  5678 => x"0a73756d",
  5679 => x"20636861",
  5680 => x"6e6e656c",
  5681 => x"2020203a",
  5682 => x"20000000",
  5683 => x"0a0a706f",
  5684 => x"73697469",
  5685 => x"6f6e2063",
  5686 => x"6f6d7075",
  5687 => x"74617469",
  5688 => x"6f6e0000",
  5689 => x"0a202073",
  5690 => x"63616c65",
  5691 => x"72207661",
  5692 => x"6c756573",
  5693 => x"20202020",
  5694 => x"20202020",
  5695 => x"20000000",
  5696 => x"0a20206f",
  5697 => x"66667365",
  5698 => x"74202020",
  5699 => x"20202020",
  5700 => x"20202020",
  5701 => x"20202020",
  5702 => x"20000000",
  5703 => x"0a6f7574",
  5704 => x"70757420",
  5705 => x"73656c65",
  5706 => x"6374203a",
  5707 => x"20000000",
  5708 => x"74657374",
  5709 => x"67656e00",
  5710 => x"4e4f5420",
  5711 => x"00000000",
  5712 => x"6368616e",
  5713 => x"6e656c20",
  5714 => x"30000000",
  5715 => x"0a63616c",
  5716 => x"63207374",
  5717 => x"61746520",
  5718 => x"2020203a",
  5719 => x"20307800",
  5720 => x"76657274",
  5721 => x"6963616c",
  5722 => x"00000000",
  5723 => x"686f7269",
  5724 => x"7a6f6e74",
  5725 => x"616c0000",
  5726 => x"73756d00",
  5727 => x"6368616e",
  5728 => x"6e656c20",
  5729 => x"33000000",
  5730 => x"6368616e",
  5731 => x"6e656c20",
  5732 => x"32000000",
  5733 => x"6368616e",
  5734 => x"6e656c20",
  5735 => x"31000000",
  5736 => x"786d6f64",
  5737 => x"656d2074",
  5738 => x"72616e73",
  5739 => x"6d69742e",
  5740 => x"2e2e0a00",
  5741 => x"20627974",
  5742 => x"65732074",
  5743 => x"72616e73",
  5744 => x"6d697474",
  5745 => x"65640a00",
  5746 => x"63616e63",
  5747 => x"656c0a00",
  5748 => x"72657472",
  5749 => x"79206f75",
  5750 => x"740a0000",
  5751 => x"786d6f64",
  5752 => x"656d2072",
  5753 => x"65636569",
  5754 => x"76652e2e",
  5755 => x"2e0a0000",
  5756 => x"20627974",
  5757 => x"65732072",
  5758 => x"65636569",
  5759 => x"7665640a",
  5760 => x"00000000",
  5761 => x"72782062",
  5762 => x"75666665",
  5763 => x"72206675",
  5764 => x"6c6c0a00",
  5765 => x"74696d65",
  5766 => x"206f7574",
  5767 => x"0a000000",
  5768 => x"64656275",
  5769 => x"67207265",
  5770 => x"67697374",
  5771 => x"65727300",
  5772 => x"0a6d6f64",
  5773 => x"65202020",
  5774 => x"20202020",
  5775 => x"203a2000",
  5776 => x"0a616464",
  5777 => x"72657373",
  5778 => x"20302020",
  5779 => x"203a2030",
  5780 => x"78000000",
  5781 => x"0a616464",
  5782 => x"72657373",
  5783 => x"20312020",
  5784 => x"203a2030",
  5785 => x"78000000",
  5786 => x"0a627566",
  5787 => x"66657220",
  5788 => x"73697a65",
  5789 => x"203a2000",
  5790 => x"6d61783a",
  5791 => x"20000000",
  5792 => x"6d696e3a",
  5793 => x"20000000",
  5794 => x"63683a20",
  5795 => x"00000000",
  5796 => x"73706c3a",
  5797 => x"20000000",
  5798 => x"73686f77",
  5799 => x"2042504d",
  5800 => x"20726567",
  5801 => x"69737465",
  5802 => x"72730000",
  5803 => x"62706d00",
  5804 => x"73656c65",
  5805 => x"6374206f",
  5806 => x"75747075",
  5807 => x"74206368",
  5808 => x"616e6e65",
  5809 => x"6c202830",
  5810 => x"2e2e3320",
  5811 => x"73756d20",
  5812 => x"68207629",
  5813 => x"00000000",
  5814 => x"73656c65",
  5815 => x"63740000",
  5816 => x"73797374",
  5817 => x"656d2072",
  5818 => x"65736574",
  5819 => x"00000000",
  5820 => x"72657365",
  5821 => x"74000000",
  5822 => x"73686f77",
  5823 => x"20737973",
  5824 => x"74656d20",
  5825 => x"696e666f",
  5826 => x"203c7665",
  5827 => x"72626f73",
  5828 => x"653e0000",
  5829 => x"73797369",
  5830 => x"6e666f00",
  5831 => x"73686f77",
  5832 => x"2f736574",
  5833 => x"20646562",
  5834 => x"75672072",
  5835 => x"65676973",
  5836 => x"74657273",
  5837 => x"203c7365",
  5838 => x"74206d6f",
  5839 => x"64653e00",
  5840 => x"64656275",
  5841 => x"67000000",
  5842 => x"636c6b20",
  5843 => x"736f7572",
  5844 => x"63653a20",
  5845 => x"2030203d",
  5846 => x"20696e74",
  5847 => x"2c203120",
  5848 => x"3d206578",
  5849 => x"74000000",
  5850 => x"636c6b00",
  5851 => x"6d696372",
  5852 => x"6f70756c",
  5853 => x"73652073",
  5854 => x"6f757263",
  5855 => x"653a2030",
  5856 => x"203d2069",
  5857 => x"6e742c20",
  5858 => x"31203d20",
  5859 => x"65787400",
  5860 => x"6d696372",
  5861 => x"6f000000",
  5862 => x"74657374",
  5863 => x"67656e65",
  5864 => x"7261746f",
  5865 => x"72203c73",
  5866 => x"63616c65",
  5867 => x"723e203c",
  5868 => x"72657374",
  5869 => x"6172743e",
  5870 => x"00000000",
  5871 => x"3c6d7574",
  5872 => x"655f6e3e",
  5873 => x"203c7273",
  5874 => x"745f6e3e",
  5875 => x"203c6270",
  5876 => x"625f6e3e",
  5877 => x"203c6f73",
  5878 => x"72313e20",
  5879 => x"3c6f7372",
  5880 => x"323e0000",
  5881 => x"64616363",
  5882 => x"6f6e6600",
  5883 => x"3c6d756c",
  5884 => x"7469706c",
  5885 => x"6965723e",
  5886 => x"20696e69",
  5887 => x"7469616c",
  5888 => x"697a6520",
  5889 => x"62756666",
  5890 => x"65720000",
  5891 => x"64616374",
  5892 => x"65737400",
  5893 => x"72657365",
  5894 => x"74206361",
  5895 => x"6c63756c",
  5896 => x"6174696f",
  5897 => x"6e206572",
  5898 => x"726f7273",
  5899 => x"00000000",
  5900 => x"63616c63",
  5901 => x"72657300",
  5902 => x"73686f77",
  5903 => x"20646562",
  5904 => x"75672062",
  5905 => x"75666665",
  5906 => x"72203c6c",
  5907 => x"656e6774",
  5908 => x"683e0000",
  5909 => x"636c6561",
  5910 => x"72206465",
  5911 => x"62756720",
  5912 => x"62756666",
  5913 => x"65720000",
  5914 => x"62636c65",
  5915 => x"61720000",
  5916 => x"62756666",
  5917 => x"6572206f",
  5918 => x"6e204c43",
  5919 => x"44203c63",
  5920 => x"683e203c",
  5921 => x"636f6d62",
  5922 => x"3e000000",
  5923 => x"73636f70",
  5924 => x"65000000",
  5925 => x"64656275",
  5926 => x"67207472",
  5927 => x"61636520",
  5928 => x"3c636c65",
  5929 => x"61723e00",
  5930 => x"74726163",
  5931 => x"65000000",
  5932 => x"73657475",
  5933 => x"70206368",
  5934 => x"616e6e65",
  5935 => x"6c207465",
  5936 => x"7374203c",
  5937 => x"63683e20",
  5938 => x"3c76616c",
  5939 => x"302e2e37",
  5940 => x"3e000000",
  5941 => x"63687465",
  5942 => x"73740000",
  5943 => x"72756e6e",
  5944 => x"696e6720",
  5945 => x"6c696768",
  5946 => x"74000000",
  5947 => x"72756e00",
  5948 => x"72756e20",
  5949 => x"64697370",
  5950 => x"6c617920",
  5951 => x"74657374",
  5952 => x"2066756e",
  5953 => x"6374696f",
  5954 => x"6e000000",
  5955 => x"64697370",
  5956 => x"6c617900",
  5957 => x"73657420",
  5958 => x"6261636b",
  5959 => x"6c696768",
  5960 => x"74203c30",
  5961 => x"2e2e3331",
  5962 => x"3e000000",
  5963 => x"6261636b",
  5964 => x"00000000",
  5965 => x"73686f77",
  5966 => x"206c6f67",
  5967 => x"6f206f6e",
  5968 => x"20676c63",
  5969 => x"64000000",
  5970 => x"6c6f676f",
  5971 => x"00000000",
  5972 => x"63686563",
  5973 => x"6b204932",
  5974 => x"43206164",
  5975 => x"64726573",
  5976 => x"73000000",
  5977 => x"69326300",
  5978 => x"72656164",
  5979 => x"20454550",
  5980 => x"524f4d20",
  5981 => x"3c627573",
  5982 => x"3e203c69",
  5983 => x"32635f61",
  5984 => x"6464723e",
  5985 => x"203c6c65",
  5986 => x"6e677468",
  5987 => x"3e000000",
  5988 => x"65657072",
  5989 => x"6f6d0000",
  5990 => x"41444320",
  5991 => x"72656769",
  5992 => x"73746572",
  5993 => x"20747261",
  5994 => x"6e736665",
  5995 => x"72203c76",
  5996 => x"616c7565",
  5997 => x"3e000000",
  5998 => x"61747261",
  5999 => x"6e730000",
  6000 => x"696e6974",
  6001 => x"20414443",
  6002 => x"20726567",
  6003 => x"69737465",
  6004 => x"72730000",
  6005 => x"61696e69",
  6006 => x"74000000",
  6007 => x"616c6961",
  6008 => x"7320666f",
  6009 => x"72207800",
  6010 => x"6d656d00",
  6011 => x"77726974",
  6012 => x"6520776f",
  6013 => x"7264203c",
  6014 => x"61646472",
  6015 => x"3e203c6c",
  6016 => x"656e6774",
  6017 => x"683e203c",
  6018 => x"76616c75",
  6019 => x"65287329",
  6020 => x"3e000000",
  6021 => x"776d656d",
  6022 => x"00000000",
  6023 => x"6558616d",
  6024 => x"696e6520",
  6025 => x"6d656d6f",
  6026 => x"72790000",
  6027 => x"636c6561",
  6028 => x"72207363",
  6029 => x"7265656e",
  6030 => x"00000000",
  6031 => x"636c6561",
  6032 => x"72000000",
  6033 => x"0a646562",
  6034 => x"75672074",
  6035 => x"72616365",
  6036 => x"206d656d",
  6037 => x"6f727900",
  6038 => x"0a74696d",
  6039 => x"65207374",
  6040 => x"616d7020",
  6041 => x"20202073",
  6042 => x"74617465",
  6043 => x"00000000",
  6044 => x"20203078",
  6045 => x"00000000",
  6046 => x"65787465",
  6047 => x"726e616c",
  6048 => x"20636c6f",
  6049 => x"636b2000",
  6050 => x"61637469",
  6051 => x"76650a00",
  6052 => x"73656c65",
  6053 => x"63746564",
  6054 => x"0a000000",
  6055 => x"6d696372",
  6056 => x"6f70756c",
  6057 => x"73652073",
  6058 => x"6f757263",
  6059 => x"653a2000",
  6060 => x"6265616d",
  6061 => x"20706f73",
  6062 => x"6974696f",
  6063 => x"6e206d6f",
  6064 => x"6e69746f",
  6065 => x"72000000",
  6066 => x"20286f6e",
  6067 => x"2073696d",
  6068 => x"290a0000",
  6069 => x"0a485720",
  6070 => x"73796e74",
  6071 => x"68657369",
  6072 => x"7a65643a",
  6073 => x"20000000",
  6074 => x"0a535720",
  6075 => x"636f6d70",
  6076 => x"696c6564",
  6077 => x"2020203a",
  6078 => x"20417567",
  6079 => x"20313120",
  6080 => x"32303131",
  6081 => x"20203131",
  6082 => x"3a30353a",
  6083 => x"32370000",
  6084 => x"0a737973",
  6085 => x"74656d20",
  6086 => x"636c6f63",
  6087 => x"6b20203a",
  6088 => x"20000000",
  6089 => x"204d487a",
  6090 => x"0a000000",
  6091 => x"44454255",
  6092 => x"47204d4f",
  6093 => x"44450000",
  6094 => x"204f4e0a",
  6095 => x"00000000",
  6096 => x"0000117b",
  6097 => x"000011e4",
  6098 => x"000011d9",
  6099 => x"000011ce",
  6100 => x"000011c3",
  6101 => x"000011b9",
  6102 => x"000011af",
  6103 => x"000002c2",
  6104 => x"fc1902c4",
  6105 => x"fffefd3f",
  6106 => x"03e7fd3b",
  6107 => x"0000485d",
  6108 => x"999b4888",
  6109 => x"ffc4b7ce",
  6110 => x"6665b74e",
  6111 => x"3e200000",
  6112 => x"636f6d6d",
  6113 => x"616e6420",
  6114 => x"6e6f7420",
  6115 => x"666f756e",
  6116 => x"642e0a00",
  6117 => x"73757070",
  6118 => x"6f727465",
  6119 => x"6420636f",
  6120 => x"6d6d616e",
  6121 => x"64733a0a",
  6122 => x"0a000000",
  6123 => x"202d2000",
  6124 => x"76656e64",
  6125 => x"6f723f20",
  6126 => x"20000000",
  6127 => x"67616973",
  6128 => x"6c657220",
  6129 => x"20000000",
  6130 => x"756e6b6e",
  6131 => x"6f776e20",
  6132 => x"64657669",
  6133 => x"63650000",
  6134 => x"485a4452",
  6135 => x"20202020",
  6136 => x"20000000",
  6137 => x"47656e65",
  6138 => x"72616c20",
  6139 => x"50757270",
  6140 => x"6f736520",
  6141 => x"492f4f20",
  6142 => x"706f7274",
  6143 => x"00000000",
  6144 => x"56474120",
  6145 => x"636f6e74",
  6146 => x"726f6c6c",
  6147 => x"65720000",
  6148 => x"4475616c",
  6149 => x"2d706f72",
  6150 => x"74204148",
  6151 => x"42205352",
  6152 => x"414d206d",
  6153 => x"6f64756c",
  6154 => x"65000000",
  6155 => x"64656275",
  6156 => x"67206275",
  6157 => x"66666572",
  6158 => x"20636f6e",
  6159 => x"74726f6c",
  6160 => x"00000000",
  6161 => x"74726967",
  6162 => x"67657220",
  6163 => x"67656e65",
  6164 => x"7261746f",
  6165 => x"72000000",
  6166 => x"64656275",
  6167 => x"6720636f",
  6168 => x"6e736f6c",
  6169 => x"65000000",
  6170 => x"64656275",
  6171 => x"67207472",
  6172 => x"61636572",
  6173 => x"206d656d",
  6174 => x"6f727900",
  6175 => x"4541444f",
  6176 => x"47533130",
  6177 => x"32206469",
  6178 => x"73706c61",
  6179 => x"79206472",
  6180 => x"69766572",
  6181 => x"00000000",
  6182 => x"44434d20",
  6183 => x"70686173",
  6184 => x"65207368",
  6185 => x"69667420",
  6186 => x"636f6e74",
  6187 => x"726f6c00",
  6188 => x"5a505520",
  6189 => x"4d656d6f",
  6190 => x"72792077",
  6191 => x"72617070",
  6192 => x"65720000",
  6193 => x"5a505520",
  6194 => x"41484220",
  6195 => x"57726170",
  6196 => x"70657200",
  6197 => x"4148422f",
  6198 => x"41504220",
  6199 => x"42726964",
  6200 => x"67650000",
  6201 => x"4d6f6475",
  6202 => x"6c617220",
  6203 => x"54696d65",
  6204 => x"7220556e",
  6205 => x"69740000",
  6206 => x"414d4241",
  6207 => x"20577261",
  6208 => x"70706572",
  6209 => x"20666f72",
  6210 => x"204f4320",
  6211 => x"4932432d",
  6212 => x"6d617374",
  6213 => x"65720000",
  6214 => x"47656e65",
  6215 => x"72696320",
  6216 => x"55415254",
  6217 => x"00000000",
  6218 => x"20206170",
  6219 => x"62736c76",
  6220 => x"00000000",
  6221 => x"76656e64",
  6222 => x"20307800",
  6223 => x"64657620",
  6224 => x"30780000",
  6225 => x"76657220",
  6226 => x"00000000",
  6227 => x"69727120",
  6228 => x"00000000",
  6229 => x"61646472",
  6230 => x"20307800",
  6231 => x"6168626d",
  6232 => x"73740000",
  6233 => x"61686273",
  6234 => x"6c760000",
  6235 => x"00002af2",
  6236 => x"00002bb3",
  6237 => x"00002ba8",
  6238 => x"00002b9d",
  6239 => x"00002b7c",
  6240 => x"00002b71",
  6241 => x"00002b66",
  6242 => x"00002b5b",
  6243 => x"00002b92",
  6244 => x"00002b87",
  6245 => x"04580808",
  6246 => x"20ff0000",
  6247 => x"000061a4",
  6248 => x"00006284",
  6249 => x"02010305",
  6250 => x"05070501",
  6251 => x"03030505",
  6252 => x"02030104",
  6253 => x"05050505",
  6254 => x"05050505",
  6255 => x"05050101",
  6256 => x"04050404",
  6257 => x"07050505",
  6258 => x"05050505",
  6259 => x"05030405",
  6260 => x"05050505",
  6261 => x"05050505",
  6262 => x"05050505",
  6263 => x"05050503",
  6264 => x"04030505",
  6265 => x"02050504",
  6266 => x"05050405",
  6267 => x"04010204",
  6268 => x"02050404",
  6269 => x"05050404",
  6270 => x"04040507",
  6271 => x"05040404",
  6272 => x"02040500",
  6273 => x"04050200",
  6274 => x"04080303",
  6275 => x"04090003",
  6276 => x"06000000",
  6277 => x"00020204",
  6278 => x"04040400",
  6279 => x"04060003",
  6280 => x"05000000",
  6281 => x"00000404",
  6282 => x"05050204",
  6283 => x"05060305",
  6284 => x"04030705",
  6285 => x"04050303",
  6286 => x"02040502",
  6287 => x"03020405",
  6288 => x"06060604",
  6289 => x"05050505",
  6290 => x"05050504",
  6291 => x"04040404",
  6292 => x"03030303",
  6293 => x"05050505",
  6294 => x"05050505",
  6295 => x"05040404",
  6296 => x"04050404",
  6297 => x"04040404",
  6298 => x"04040503",
  6299 => x"04040404",
  6300 => x"02020303",
  6301 => x"04040404",
  6302 => x"04040405",
  6303 => x"04040404",
  6304 => x"04030303",
  6305 => x"00005f07",
  6306 => x"0007741c",
  6307 => x"771c172e",
  6308 => x"6a3e2b3a",
  6309 => x"06493608",
  6310 => x"36493036",
  6311 => x"49597648",
  6312 => x"073c4281",
  6313 => x"81423c0a",
  6314 => x"041f040a",
  6315 => x"08083e08",
  6316 => x"08806008",
  6317 => x"080840c0",
  6318 => x"300c033e",
  6319 => x"4141413e",
  6320 => x"44427f40",
  6321 => x"40466151",
  6322 => x"49462241",
  6323 => x"49493618",
  6324 => x"14127f10",
  6325 => x"27454545",
  6326 => x"393e4949",
  6327 => x"49300101",
  6328 => x"710d0336",
  6329 => x"49494936",
  6330 => x"06494929",
  6331 => x"1e36d008",
  6332 => x"14224114",
  6333 => x"14141414",
  6334 => x"41221408",
  6335 => x"02510906",
  6336 => x"3c4299a5",
  6337 => x"bd421c7c",
  6338 => x"1211127c",
  6339 => x"7f494949",
  6340 => x"363e4141",
  6341 => x"41227f41",
  6342 => x"41413e7f",
  6343 => x"49494941",
  6344 => x"7f090909",
  6345 => x"013e4149",
  6346 => x"497a7f08",
  6347 => x"08087f41",
  6348 => x"7f414041",
  6349 => x"413f7f08",
  6350 => x"1422417f",
  6351 => x"40404040",
  6352 => x"7f060c06",
  6353 => x"7f7f0608",
  6354 => x"307f3e41",
  6355 => x"41413e7f",
  6356 => x"09090906",
  6357 => x"3e4161c1",
  6358 => x"be7f0919",
  6359 => x"29462649",
  6360 => x"49493201",
  6361 => x"017f0101",
  6362 => x"3f404040",
  6363 => x"3f073840",
  6364 => x"38071f60",
  6365 => x"1f601f63",
  6366 => x"14081463",
  6367 => x"01067806",
  6368 => x"01615149",
  6369 => x"45437f41",
  6370 => x"41030c30",
  6371 => x"c041417f",
  6372 => x"04020102",
  6373 => x"04808080",
  6374 => x"80800102",
  6375 => x"20545454",
  6376 => x"787f4444",
  6377 => x"44383844",
  6378 => x"44443844",
  6379 => x"44447f38",
  6380 => x"54545458",
  6381 => x"087e0901",
  6382 => x"18a4a4a4",
  6383 => x"787f0404",
  6384 => x"787d807d",
  6385 => x"7f102844",
  6386 => x"3f407c04",
  6387 => x"7804787c",
  6388 => x"04047838",
  6389 => x"444438fc",
  6390 => x"24242418",
  6391 => x"18242424",
  6392 => x"fc7c0804",
  6393 => x"04485454",
  6394 => x"24043f44",
  6395 => x"403c4040",
  6396 => x"7c1c2040",
  6397 => x"201c1c60",
  6398 => x"601c6060",
  6399 => x"1c442810",
  6400 => x"28449ca0",
  6401 => x"601c6454",
  6402 => x"544c187e",
  6403 => x"8181ffff",
  6404 => x"81817e18",
  6405 => x"18040810",
  6406 => x"0c143e55",
  6407 => x"55ff8181",
  6408 => x"81ff8060",
  6409 => x"80608060",
  6410 => x"60600060",
  6411 => x"60006060",
  6412 => x"047f0414",
  6413 => x"7f140201",
  6414 => x"01024629",
  6415 => x"1608344a",
  6416 => x"31483000",
  6417 => x"18243e41",
  6418 => x"227f4941",
  6419 => x"03040403",
  6420 => x"03040304",
  6421 => x"04030403",
  6422 => x"183c3c18",
  6423 => x"08080808",
  6424 => x"03010203",
  6425 => x"020e020e",
  6426 => x"060e0048",
  6427 => x"30384438",
  6428 => x"54483844",
  6429 => x"fe44487e",
  6430 => x"49014438",
  6431 => x"28384403",
  6432 => x"147c1403",
  6433 => x"e7e74e55",
  6434 => x"55390101",
  6435 => x"0001011c",
  6436 => x"2a555522",
  6437 => x"1c1d151e",
  6438 => x"18240018",
  6439 => x"24080808",
  6440 => x"18080808",
  6441 => x"3c42bd95",
  6442 => x"a9423c01",
  6443 => x"01010101",
  6444 => x"06090906",
  6445 => x"44445f44",
  6446 => x"44191512",
  6447 => x"15150a02",
  6448 => x"01fc2020",
  6449 => x"1c0e7f01",
  6450 => x"7f011818",
  6451 => x"00804002",
  6452 => x"1f060909",
  6453 => x"06241800",
  6454 => x"2418824f",
  6455 => x"304c62f1",
  6456 => x"824f300c",
  6457 => x"d2b1955f",
  6458 => x"304c62f1",
  6459 => x"30484520",
  6460 => x"60392e38",
  6461 => x"6060382e",
  6462 => x"3960701d",
  6463 => x"131d7072",
  6464 => x"1d121e71",
  6465 => x"701d121d",
  6466 => x"70603b25",
  6467 => x"3b607e11",
  6468 => x"7f49411e",
  6469 => x"2161927c",
  6470 => x"5556447c",
  6471 => x"5655447c",
  6472 => x"5655467d",
  6473 => x"54544545",
  6474 => x"7e44447e",
  6475 => x"45467d46",
  6476 => x"457c4508",
  6477 => x"7f49413e",
  6478 => x"7e091222",
  6479 => x"7d384546",
  6480 => x"44383844",
  6481 => x"46453838",
  6482 => x"46454638",
  6483 => x"3a454546",
  6484 => x"39384544",
  6485 => x"45382214",
  6486 => x"081422bc",
  6487 => x"625a463d",
  6488 => x"3c41423c",
  6489 => x"3c42413c",
  6490 => x"3c42413e",
  6491 => x"3d40403d",
  6492 => x"0608f209",
  6493 => x"067f2222",
  6494 => x"1cfe0989",
  6495 => x"76205556",
  6496 => x"78205655",
  6497 => x"78225555",
  6498 => x"7a235556",
  6499 => x"7b205554",
  6500 => x"79275557",
  6501 => x"78205438",
  6502 => x"54483844",
  6503 => x"c4385556",
  6504 => x"58385655",
  6505 => x"583a5555",
  6506 => x"5a395454",
  6507 => x"59017a7a",
  6508 => x"01027902",
  6509 => x"02780260",
  6510 => x"91927c7b",
  6511 => x"090a7338",
  6512 => x"45463838",
  6513 => x"4645383a",
  6514 => x"45453a3b",
  6515 => x"45463b39",
  6516 => x"44443908",
  6517 => x"082a0808",
  6518 => x"b8644c3a",
  6519 => x"3c41427c",
  6520 => x"3c42417c",
  6521 => x"3a41417a",
  6522 => x"3d40407d",
  6523 => x"986219ff",
  6524 => x"423c9a60",
  6525 => x"1a000000",
  6526 => x"30622020",
  6527 => x"20202020",
  6528 => x"20202020",
  6529 => x"20202020",
  6530 => x"20202020",
  6531 => x"20202020",
  6532 => x"20202020",
  6533 => x"20202020",
  6534 => x"20200000",
  6535 => x"20202020",
  6536 => x"20202020",
  6537 => x"00000000",
  6538 => x"00202020",
  6539 => x"20202020",
  6540 => x"20202828",
  6541 => x"28282820",
  6542 => x"20202020",
  6543 => x"20202020",
  6544 => x"20202020",
  6545 => x"20202020",
  6546 => x"20881010",
  6547 => x"10101010",
  6548 => x"10101010",
  6549 => x"10101010",
  6550 => x"10040404",
  6551 => x"04040404",
  6552 => x"04040410",
  6553 => x"10101010",
  6554 => x"10104141",
  6555 => x"41414141",
  6556 => x"01010101",
  6557 => x"01010101",
  6558 => x"01010101",
  6559 => x"01010101",
  6560 => x"01010101",
  6561 => x"10101010",
  6562 => x"10104242",
  6563 => x"42424242",
  6564 => x"02020202",
  6565 => x"02020202",
  6566 => x"02020202",
  6567 => x"02020202",
  6568 => x"02020202",
  6569 => x"10101010",
  6570 => x"20000000",
  6571 => x"00000000",
  6572 => x"00000000",
  6573 => x"00000000",
  6574 => x"00000000",
  6575 => x"00000000",
  6576 => x"00000000",
  6577 => x"00000000",
  6578 => x"00000000",
  6579 => x"00000000",
  6580 => x"00000000",
  6581 => x"00000000",
  6582 => x"00000000",
  6583 => x"00000000",
  6584 => x"00000000",
  6585 => x"00000000",
  6586 => x"00000000",
  6587 => x"00000000",
  6588 => x"00000000",
  6589 => x"00000000",
  6590 => x"00000000",
  6591 => x"00000000",
  6592 => x"00000000",
  6593 => x"00000000",
  6594 => x"00000000",
  6595 => x"00000000",
  6596 => x"00000000",
  6597 => x"00000000",
  6598 => x"00000000",
  6599 => x"00000000",
  6600 => x"00000000",
  6601 => x"00000000",
  6602 => x"00000000",
  6603 => x"43000000",
  6604 => x"00000000",
  6605 => x"80000c00",
  6606 => x"80000b00",
  6607 => x"80000800",
  6608 => x"00000000",
  6609 => x"ff000000",
  6610 => x"00000000",
  6611 => x"00000000",
  6612 => x"00ffffff",
  6613 => x"ff00ffff",
  6614 => x"ffff00ff",
  6615 => x"ffffff00",
  6616 => x"00000000",
  6617 => x"00000000",
  6618 => x"80000a00",
  6619 => x"80000700",
  6620 => x"80000600",
  6621 => x"80000400",
  6622 => x"80000200",
  6623 => x"80000100",
  6624 => x"80000004",
  6625 => x"80000000",
  6626 => x"0000678c",
  6627 => x"00000000",
  6628 => x"000069f4",
  6629 => x"00006a50",
  6630 => x"00006aac",
  6631 => x"00000000",
  6632 => x"00000000",
  6633 => x"00000000",
  6634 => x"00000000",
  6635 => x"00000000",
  6636 => x"00000000",
  6637 => x"00000000",
  6638 => x"00000000",
  6639 => x"00000000",
  6640 => x"0000672c",
  6641 => x"00000000",
  6642 => x"00000000",
  6643 => x"00000000",
  6644 => x"00000000",
  6645 => x"00000000",
  6646 => x"00000000",
  6647 => x"00000000",
  6648 => x"00000000",
  6649 => x"00000000",
  6650 => x"00000000",
  6651 => x"00000000",
  6652 => x"00000000",
  6653 => x"00000000",
  6654 => x"00000000",
  6655 => x"00000000",
  6656 => x"00000000",
  6657 => x"00000000",
  6658 => x"00000000",
  6659 => x"00000000",
  6660 => x"00000000",
  6661 => x"00000000",
  6662 => x"00000000",
  6663 => x"00000000",
  6664 => x"00000000",
  6665 => x"00000000",
  6666 => x"00000000",
  6667 => x"00000000",
  6668 => x"00000000",
  6669 => x"00000001",
  6670 => x"330eabcd",
  6671 => x"1234e66d",
  6672 => x"deec0005",
  6673 => x"000b0000",
  6674 => x"00000000",
  6675 => x"00000000",
  6676 => x"00000000",
  6677 => x"00000000",
  6678 => x"00000000",
  6679 => x"00000000",
  6680 => x"00000000",
  6681 => x"00000000",
  6682 => x"00000000",
  6683 => x"00000000",
  6684 => x"00000000",
  6685 => x"00000000",
  6686 => x"00000000",
  6687 => x"00000000",
  6688 => x"00000000",
  6689 => x"00000000",
  6690 => x"00000000",
  6691 => x"00000000",
  6692 => x"00000000",
  6693 => x"00000000",
  6694 => x"00000000",
  6695 => x"00000000",
  6696 => x"00000000",
  6697 => x"00000000",
  6698 => x"00000000",
  6699 => x"00000000",
  6700 => x"00000000",
  6701 => x"00000000",
  6702 => x"00000000",
  6703 => x"00000000",
  6704 => x"00000000",
  6705 => x"00000000",
  6706 => x"00000000",
  6707 => x"00000000",
  6708 => x"00000000",
  6709 => x"00000000",
  6710 => x"00000000",
  6711 => x"00000000",
  6712 => x"00000000",
  6713 => x"00000000",
  6714 => x"00000000",
  6715 => x"00000000",
  6716 => x"00000000",
  6717 => x"00000000",
  6718 => x"00000000",
  6719 => x"00000000",
  6720 => x"00000000",
  6721 => x"00000000",
  6722 => x"00000000",
  6723 => x"00000000",
  6724 => x"00000000",
  6725 => x"00000000",
  6726 => x"00000000",
  6727 => x"00000000",
  6728 => x"00000000",
  6729 => x"00000000",
  6730 => x"00000000",
  6731 => x"00000000",
  6732 => x"00000000",
  6733 => x"00000000",
  6734 => x"00000000",
  6735 => x"00000000",
  6736 => x"00000000",
  6737 => x"00000000",
  6738 => x"00000000",
  6739 => x"00000000",
  6740 => x"00000000",
  6741 => x"00000000",
  6742 => x"00000000",
  6743 => x"00000000",
  6744 => x"00000000",
  6745 => x"00000000",
  6746 => x"00000000",
  6747 => x"00000000",
  6748 => x"00000000",
  6749 => x"00000000",
  6750 => x"00000000",
  6751 => x"00000000",
  6752 => x"00000000",
  6753 => x"00000000",
  6754 => x"00000000",
  6755 => x"00000000",
  6756 => x"00000000",
  6757 => x"00000000",
  6758 => x"00000000",
  6759 => x"00000000",
  6760 => x"00000000",
  6761 => x"00000000",
  6762 => x"00000000",
  6763 => x"00000000",
  6764 => x"00000000",
  6765 => x"00000000",
  6766 => x"00000000",
  6767 => x"00000000",
  6768 => x"00000000",
  6769 => x"00000000",
  6770 => x"00000000",
  6771 => x"00000000",
  6772 => x"00000000",
  6773 => x"00000000",
  6774 => x"00000000",
  6775 => x"00000000",
  6776 => x"00000000",
  6777 => x"00000000",
  6778 => x"00000000",
  6779 => x"00000000",
  6780 => x"00000000",
  6781 => x"00000000",
  6782 => x"00000000",
  6783 => x"00000000",
  6784 => x"00000000",
  6785 => x"00000000",
  6786 => x"00000000",
  6787 => x"00000000",
  6788 => x"00000000",
  6789 => x"00000000",
  6790 => x"00000000",
  6791 => x"00000000",
  6792 => x"00000000",
  6793 => x"00000000",
  6794 => x"00000000",
  6795 => x"00000000",
  6796 => x"00000000",
  6797 => x"00000000",
  6798 => x"00000000",
  6799 => x"00000000",
  6800 => x"00000000",
  6801 => x"00000000",
  6802 => x"00000000",
  6803 => x"00000000",
  6804 => x"00000000",
  6805 => x"00000000",
  6806 => x"00000000",
  6807 => x"00000000",
  6808 => x"00000000",
  6809 => x"00000000",
  6810 => x"00000000",
  6811 => x"00000000",
  6812 => x"00000000",
  6813 => x"00000000",
  6814 => x"00000000",
  6815 => x"00000000",
  6816 => x"00000000",
  6817 => x"00000000",
  6818 => x"00000000",
  6819 => x"00000000",
  6820 => x"00000000",
  6821 => x"00000000",
  6822 => x"00000000",
  6823 => x"00000000",
  6824 => x"00000000",
  6825 => x"00000000",
  6826 => x"00000000",
  6827 => x"00000000",
  6828 => x"00000000",
  6829 => x"00000000",
  6830 => x"00000000",
  6831 => x"00000000",
  6832 => x"00000000",
  6833 => x"00000000",
  6834 => x"00000000",
  6835 => x"00000000",
  6836 => x"00000000",
  6837 => x"00000000",
  6838 => x"00000000",
  6839 => x"00000000",
  6840 => x"00000000",
  6841 => x"00000000",
  6842 => x"00000000",
  6843 => x"00000000",
  6844 => x"00000000",
  6845 => x"00000000",
  6846 => x"00000000",
  6847 => x"00000000",
  6848 => x"00000000",
  6849 => x"00000000",
  6850 => x"00000000",
  6851 => x"00000000",
  6852 => x"00000000",
  6853 => x"00000000",
  6854 => x"00000000",
  6855 => x"00000000",
  6856 => x"00000000",
  6857 => x"00000000",
  6858 => x"00000000",
  6859 => x"00000000",
  6860 => x"00000000",
  6861 => x"00000000",
  6862 => x"ffffffff",
  6863 => x"00000000",
  6864 => x"00020000",
  6865 => x"00000000",
  6866 => x"00000000",
  6867 => x"00006b44",
  6868 => x"00006b44",
  6869 => x"00006b4c",
  6870 => x"00006b4c",
  6871 => x"00006b54",
  6872 => x"00006b54",
  6873 => x"00006b5c",
  6874 => x"00006b5c",
  6875 => x"00006b64",
  6876 => x"00006b64",
  6877 => x"00006b6c",
  6878 => x"00006b6c",
  6879 => x"00006b74",
  6880 => x"00006b74",
  6881 => x"00006b7c",
  6882 => x"00006b7c",
  6883 => x"00006b84",
  6884 => x"00006b84",
  6885 => x"00006b8c",
  6886 => x"00006b8c",
  6887 => x"00006b94",
  6888 => x"00006b94",
  6889 => x"00006b9c",
  6890 => x"00006b9c",
  6891 => x"00006ba4",
  6892 => x"00006ba4",
  6893 => x"00006bac",
  6894 => x"00006bac",
  6895 => x"00006bb4",
  6896 => x"00006bb4",
  6897 => x"00006bbc",
  6898 => x"00006bbc",
  6899 => x"00006bc4",
  6900 => x"00006bc4",
  6901 => x"00006bcc",
  6902 => x"00006bcc",
  6903 => x"00006bd4",
  6904 => x"00006bd4",
  6905 => x"00006bdc",
  6906 => x"00006bdc",
  6907 => x"00006be4",
  6908 => x"00006be4",
  6909 => x"00006bec",
  6910 => x"00006bec",
  6911 => x"00006bf4",
  6912 => x"00006bf4",
  6913 => x"00006bfc",
  6914 => x"00006bfc",
  6915 => x"00006c04",
  6916 => x"00006c04",
  6917 => x"00006c0c",
  6918 => x"00006c0c",
  6919 => x"00006c14",
  6920 => x"00006c14",
  6921 => x"00006c1c",
  6922 => x"00006c1c",
  6923 => x"00006c24",
  6924 => x"00006c24",
  6925 => x"00006c2c",
  6926 => x"00006c2c",
  6927 => x"00006c34",
  6928 => x"00006c34",
  6929 => x"00006c3c",
  6930 => x"00006c3c",
  6931 => x"00006c44",
  6932 => x"00006c44",
  6933 => x"00006c4c",
  6934 => x"00006c4c",
  6935 => x"00006c54",
  6936 => x"00006c54",
  6937 => x"00006c5c",
  6938 => x"00006c5c",
  6939 => x"00006c64",
  6940 => x"00006c64",
  6941 => x"00006c6c",
  6942 => x"00006c6c",
  6943 => x"00006c74",
  6944 => x"00006c74",
  6945 => x"00006c7c",
  6946 => x"00006c7c",
  6947 => x"00006c84",
  6948 => x"00006c84",
  6949 => x"00006c8c",
  6950 => x"00006c8c",
  6951 => x"00006c94",
  6952 => x"00006c94",
  6953 => x"00006c9c",
  6954 => x"00006c9c",
  6955 => x"00006ca4",
  6956 => x"00006ca4",
  6957 => x"00006cac",
  6958 => x"00006cac",
  6959 => x"00006cb4",
  6960 => x"00006cb4",
  6961 => x"00006cbc",
  6962 => x"00006cbc",
  6963 => x"00006cc4",
  6964 => x"00006cc4",
  6965 => x"00006ccc",
  6966 => x"00006ccc",
  6967 => x"00006cd4",
  6968 => x"00006cd4",
  6969 => x"00006cdc",
  6970 => x"00006cdc",
  6971 => x"00006ce4",
  6972 => x"00006ce4",
  6973 => x"00006cec",
  6974 => x"00006cec",
  6975 => x"00006cf4",
  6976 => x"00006cf4",
  6977 => x"00006cfc",
  6978 => x"00006cfc",
  6979 => x"00006d04",
  6980 => x"00006d04",
  6981 => x"00006d0c",
  6982 => x"00006d0c",
  6983 => x"00006d14",
  6984 => x"00006d14",
  6985 => x"00006d1c",
  6986 => x"00006d1c",
  6987 => x"00006d24",
  6988 => x"00006d24",
  6989 => x"00006d2c",
  6990 => x"00006d2c",
  6991 => x"00006d34",
  6992 => x"00006d34",
  6993 => x"00006d3c",
  6994 => x"00006d3c",
  6995 => x"00006d44",
  6996 => x"00006d44",
  6997 => x"00006d4c",
  6998 => x"00006d4c",
  6999 => x"00006d54",
  7000 => x"00006d54",
  7001 => x"00006d5c",
  7002 => x"00006d5c",
  7003 => x"00006d64",
  7004 => x"00006d64",
  7005 => x"00006d6c",
  7006 => x"00006d6c",
  7007 => x"00006d74",
  7008 => x"00006d74",
  7009 => x"00006d7c",
  7010 => x"00006d7c",
  7011 => x"00006d84",
  7012 => x"00006d84",
  7013 => x"00006d8c",
  7014 => x"00006d8c",
  7015 => x"00006d94",
  7016 => x"00006d94",
  7017 => x"00006d9c",
  7018 => x"00006d9c",
  7019 => x"00006da4",
  7020 => x"00006da4",
  7021 => x"00006dac",
  7022 => x"00006dac",
  7023 => x"00006db4",
  7024 => x"00006db4",
  7025 => x"00006dbc",
  7026 => x"00006dbc",
  7027 => x"00006dc4",
  7028 => x"00006dc4",
  7029 => x"00006dcc",
  7030 => x"00006dcc",
  7031 => x"00006dd4",
  7032 => x"00006dd4",
  7033 => x"00006ddc",
  7034 => x"00006ddc",
  7035 => x"00006de4",
  7036 => x"00006de4",
  7037 => x"00006dec",
  7038 => x"00006dec",
  7039 => x"00006df4",
  7040 => x"00006df4",
  7041 => x"00006dfc",
  7042 => x"00006dfc",
  7043 => x"00006e04",
  7044 => x"00006e04",
  7045 => x"00006e0c",
  7046 => x"00006e0c",
  7047 => x"00006e14",
  7048 => x"00006e14",
  7049 => x"00006e1c",
  7050 => x"00006e1c",
  7051 => x"00006e24",
  7052 => x"00006e24",
  7053 => x"00006e2c",
  7054 => x"00006e2c",
  7055 => x"00006e34",
  7056 => x"00006e34",
  7057 => x"00006e3c",
  7058 => x"00006e3c",
  7059 => x"00006e44",
  7060 => x"00006e44",
  7061 => x"00006e4c",
  7062 => x"00006e4c",
  7063 => x"00006e54",
  7064 => x"00006e54",
  7065 => x"00006e5c",
  7066 => x"00006e5c",
  7067 => x"00006e64",
  7068 => x"00006e64",
  7069 => x"00006e6c",
  7070 => x"00006e6c",
  7071 => x"00006e74",
  7072 => x"00006e74",
  7073 => x"00006e7c",
  7074 => x"00006e7c",
  7075 => x"00006e84",
  7076 => x"00006e84",
  7077 => x"00006e8c",
  7078 => x"00006e8c",
  7079 => x"00006e94",
  7080 => x"00006e94",
  7081 => x"00006e9c",
  7082 => x"00006e9c",
  7083 => x"00006ea4",
  7084 => x"00006ea4",
  7085 => x"00006eac",
  7086 => x"00006eac",
  7087 => x"00006eb4",
  7088 => x"00006eb4",
  7089 => x"00006ebc",
  7090 => x"00006ebc",
  7091 => x"00006ec4",
  7092 => x"00006ec4",
  7093 => x"00006ecc",
  7094 => x"00006ecc",
  7095 => x"00006ed4",
  7096 => x"00006ed4",
  7097 => x"00006edc",
  7098 => x"00006edc",
  7099 => x"00006ee4",
  7100 => x"00006ee4",
  7101 => x"00006eec",
  7102 => x"00006eec",
  7103 => x"00006ef4",
  7104 => x"00006ef4",
  7105 => x"00006efc",
  7106 => x"00006efc",
  7107 => x"00006f04",
  7108 => x"00006f04",
  7109 => x"00006f0c",
  7110 => x"00006f0c",
  7111 => x"00006f14",
  7112 => x"00006f14",
  7113 => x"00006f1c",
  7114 => x"00006f1c",
  7115 => x"00006f24",
  7116 => x"00006f24",
  7117 => x"00006f2c",
  7118 => x"00006f2c",
  7119 => x"00006f34",
  7120 => x"00006f34",
  7121 => x"00006f3c",
  7122 => x"00006f3c",
	--others => x"aaaaaaaa" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
