-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b80f3",
     1 => x"ea040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b80f6",
     9 => x"d1040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b80f6",
    73 => x"83040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b80f5e6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b81cc",
   162 => x"d8738306",
   163 => x"10100508",
   164 => x"060b0b80",
   165 => x"f5e90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b80f6",
   169 => x"b8040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b80f6",
   177 => x"9f040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"81cce80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053370",
   258 => x"525280f3",
   259 => x"ac3f7151",
   260 => x"80f3f63f",
   261 => x"71b00c83",
   262 => x"3d0d04ff",
   263 => x"3d0d81cc",
   264 => x"c408b811",
   265 => x"08535180",
   266 => x"0bb8120c",
   267 => x"71b00c83",
   268 => x"3d0d0480",
   269 => x"0b81eff8",
   270 => x"34800bb0",
   271 => x"0c04fb3d",
   272 => x"0d815180",
   273 => x"c7dd3fb0",
   274 => x"08538251",
   275 => x"80c7d43f",
   276 => x"b00856b0",
   277 => x"08833890",
   278 => x"5672fc06",
   279 => x"5575812e",
   280 => x"80fb3880",
   281 => x"54737627",
   282 => x"ad387383",
   283 => x"06537280",
   284 => x"2eb23881",
   285 => x"c0c85180",
   286 => x"ee983f74",
   287 => x"70840556",
   288 => x"0852a051",
   289 => x"80eeae3f",
   290 => x"a05180ed",
   291 => x"eb3f8114",
   292 => x"54757426",
   293 => x"d5388a51",
   294 => x"80eddd3f",
   295 => x"800bb00c",
   296 => x"873d0d04",
   297 => x"81a5b051",
   298 => x"80ede73f",
   299 => x"7452a051",
   300 => x"80ee823f",
   301 => x"81b29c51",
   302 => x"80edd73f",
   303 => x"81c0c851",
   304 => x"80edcf3f",
   305 => x"74708405",
   306 => x"560852a0",
   307 => x"5180ede5",
   308 => x"3fa05180",
   309 => x"eda23f81",
   310 => x"1454ffb5",
   311 => x"3981c0c8",
   312 => x"5180edae",
   313 => x"3f740852",
   314 => x"a05180ed",
   315 => x"c83f8a51",
   316 => x"80ed853f",
   317 => x"800bb00c",
   318 => x"873d0d04",
   319 => x"fc3d0d81",
   320 => x"5180c69f",
   321 => x"3fb00852",
   322 => x"825180c4",
   323 => x"e43fb008",
   324 => x"81ff0672",
   325 => x"56538354",
   326 => x"72802ea2",
   327 => x"38735180",
   328 => x"c6813f81",
   329 => x"147081ff",
   330 => x"06ff1570",
   331 => x"81ff06b0",
   332 => x"08797084",
   333 => x"055b0c56",
   334 => x"52555272",
   335 => x"e03872b0",
   336 => x"0c863d0d",
   337 => x"04803d0d",
   338 => x"8c5180ec",
   339 => x"ab3f800b",
   340 => x"b00c823d",
   341 => x"0d04fb3d",
   342 => x"0d800b81",
   343 => x"a5b45256",
   344 => x"80ecaf3f",
   345 => x"75557410",
   346 => x"81fe0653",
   347 => x"81d05281",
   348 => x"ccf00851",
   349 => x"80d2d13f",
   350 => x"b008982b",
   351 => x"54807424",
   352 => x"a23881a5",
   353 => x"c05180ec",
   354 => x"893f7452",
   355 => x"885180ec",
   356 => x"a43f81a5",
   357 => x"cc5180eb",
   358 => x"f93f8116",
   359 => x"7083ffff",
   360 => x"06575481",
   361 => x"157081ff",
   362 => x"0670982b",
   363 => x"52565473",
   364 => x"8025ffb2",
   365 => x"3875b00c",
   366 => x"873d0d04",
   367 => x"f33d0d7f",
   368 => x"02840580",
   369 => x"c3053302",
   370 => x"880580c6",
   371 => x"052281a5",
   372 => x"dc545b55",
   373 => x"5880ebba",
   374 => x"3f785180",
   375 => x"ecfe3f81",
   376 => x"a5e85180",
   377 => x"ebac3f73",
   378 => x"52885180",
   379 => x"ebc73f81",
   380 => x"a6845180",
   381 => x"eb9c3f80",
   382 => x"57767927",
   383 => x"81a13873",
   384 => x"108e3d5d",
   385 => x"5a7981ff",
   386 => x"06538190",
   387 => x"52775180",
   388 => x"d1b63f76",
   389 => x"882a5390",
   390 => x"52775180",
   391 => x"d1aa3f76",
   392 => x"81ff0653",
   393 => x"90527751",
   394 => x"80d19d3f",
   395 => x"811a7081",
   396 => x"ff065455",
   397 => x"81905277",
   398 => x"5180d18c",
   399 => x"3f805380",
   400 => x"e0527751",
   401 => x"80d1813f",
   402 => x"b008982b",
   403 => x"54807424",
   404 => x"8a388818",
   405 => x"087081ff",
   406 => x"065c567a",
   407 => x"81ff0681",
   408 => x"c0c85256",
   409 => x"80eaab3f",
   410 => x"75528851",
   411 => x"80eac63f",
   412 => x"81aff851",
   413 => x"80ea9b3f",
   414 => x"e0165480",
   415 => x"df7427b6",
   416 => x"38768706",
   417 => x"701d5755",
   418 => x"a0763474",
   419 => x"872eb938",
   420 => x"81177083",
   421 => x"ffff0658",
   422 => x"55787726",
   423 => x"fee73880",
   424 => x"e00b8c19",
   425 => x"0c8c1808",
   426 => x"70812a81",
   427 => x"06585a76",
   428 => x"f4388f3d",
   429 => x"0d047687",
   430 => x"06701d55",
   431 => x"55757434",
   432 => x"74872e09",
   433 => x"8106c938",
   434 => x"7b5180e9",
   435 => x"c53f8a51",
   436 => x"80e9a53f",
   437 => x"81177083",
   438 => x"ffff0658",
   439 => x"55787726",
   440 => x"fea338ff",
   441 => x"ba39fb3d",
   442 => x"0d815180",
   443 => x"c1833fb0",
   444 => x"0881ff06",
   445 => x"54825180",
   446 => x"c2a93fb0",
   447 => x"0881ff06",
   448 => x"56835180",
   449 => x"c0eb3fb0",
   450 => x"0883ffff",
   451 => x"0655739c",
   452 => x"3881ccf0",
   453 => x"08547484",
   454 => x"38818055",
   455 => x"74537552",
   456 => x"7351fd98",
   457 => x"3f74b00c",
   458 => x"873d0d04",
   459 => x"81ccf408",
   460 => x"54e439f8",
   461 => x"3d0d02aa",
   462 => x"052281cc",
   463 => x"cc3381f7",
   464 => x"06585876",
   465 => x"81cccc34",
   466 => x"81ccf008",
   467 => x"5580c053",
   468 => x"81905274",
   469 => x"5180cef0",
   470 => x"3f745180",
   471 => x"cf9c3fb0",
   472 => x"0881ff06",
   473 => x"5473802e",
   474 => x"84903876",
   475 => x"5380d052",
   476 => x"745180ce",
   477 => x"d33f8059",
   478 => x"8f5781cc",
   479 => x"cc3381fe",
   480 => x"06547381",
   481 => x"cccc3481",
   482 => x"ccf00874",
   483 => x"575580c0",
   484 => x"53819052",
   485 => x"745180ce",
   486 => x"af3f7451",
   487 => x"80cedb3f",
   488 => x"b00881ff",
   489 => x"06547380",
   490 => x"2e83c438",
   491 => x"755380d0",
   492 => x"52745180",
   493 => x"ce923f77",
   494 => x"772c8106",
   495 => x"5574802e",
   496 => x"83a23881",
   497 => x"cccc3382",
   498 => x"07547381",
   499 => x"cccc3481",
   500 => x"ccf00874",
   501 => x"575580c0",
   502 => x"53819052",
   503 => x"745180cd",
   504 => x"e73f7451",
   505 => x"80ce933f",
   506 => x"b00881ff",
   507 => x"06547380",
   508 => x"2e82e638",
   509 => x"755380d0",
   510 => x"52745180",
   511 => x"cdca3f81",
   512 => x"ccf00855",
   513 => x"80c15381",
   514 => x"90527451",
   515 => x"80cdb93f",
   516 => x"745180cd",
   517 => x"e53fb008",
   518 => x"81ff0656",
   519 => x"75802e82",
   520 => x"8c388053",
   521 => x"80e05274",
   522 => x"5180cd9c",
   523 => x"3f745180",
   524 => x"cdc83fb0",
   525 => x"0881ff06",
   526 => x"5473802e",
   527 => x"81ef3888",
   528 => x"15087090",
   529 => x"2b70902c",
   530 => x"56565673",
   531 => x"822a8106",
   532 => x"5473802e",
   533 => x"8d388177",
   534 => x"2b790770",
   535 => x"83ffff06",
   536 => x"5a5681cc",
   537 => x"cc338107",
   538 => x"547381cc",
   539 => x"cc3481cc",
   540 => x"f0087457",
   541 => x"5580c053",
   542 => x"81905274",
   543 => x"5180ccc8",
   544 => x"3f745180",
   545 => x"ccf43fb0",
   546 => x"0881ff06",
   547 => x"5473802e",
   548 => x"81a83875",
   549 => x"5380d052",
   550 => x"745180cc",
   551 => x"ab3f7681",
   552 => x"800a2981",
   553 => x"ff0a0570",
   554 => x"982c5856",
   555 => x"768025fd",
   556 => x"c93881cc",
   557 => x"cc338207",
   558 => x"577681cc",
   559 => x"cc3481cc",
   560 => x"f0085580",
   561 => x"c0538190",
   562 => x"52745180",
   563 => x"cbfa3f74",
   564 => x"5180cca6",
   565 => x"3fb00881",
   566 => x"ff065877",
   567 => x"802e81b8",
   568 => x"38765380",
   569 => x"d0527451",
   570 => x"80cbdd3f",
   571 => x"81cccc33",
   572 => x"88075776",
   573 => x"81cccc34",
   574 => x"81ccf008",
   575 => x"5580c053",
   576 => x"81905274",
   577 => x"5180cbc0",
   578 => x"3f745180",
   579 => x"cbec3fb0",
   580 => x"0881ff06",
   581 => x"5877802e",
   582 => x"80ef3876",
   583 => x"5380d052",
   584 => x"745180cb",
   585 => x"a33f78b0",
   586 => x"0c8a3d0d",
   587 => x"0481a688",
   588 => x"5180e4de",
   589 => x"3fff54fe",
   590 => x"923981a6",
   591 => x"885180e4",
   592 => x"d13f7681",
   593 => x"800a2981",
   594 => x"ff0a0570",
   595 => x"982c5856",
   596 => x"768025fc",
   597 => x"a538feda",
   598 => x"3981a688",
   599 => x"5180e4b2",
   600 => x"3ffd9c39",
   601 => x"81cccc33",
   602 => x"81fd0654",
   603 => x"fcdc3981",
   604 => x"a6885180",
   605 => x"e49c3ffc",
   606 => x"be3981a6",
   607 => x"885180e4",
   608 => x"913f8059",
   609 => x"8f57fbf2",
   610 => x"3981a688",
   611 => x"5180e482",
   612 => x"3f78b00c",
   613 => x"8a3d0d04",
   614 => x"81a68851",
   615 => x"80e3f33f",
   616 => x"feca39ff",
   617 => x"3d0d8151",
   618 => x"bbc73fb0",
   619 => x"0881ff06",
   620 => x"52818051",
   621 => x"fafd3f82",
   622 => x"8051faf7",
   623 => x"3f848351",
   624 => x"faf13f86",
   625 => x"f151faeb",
   626 => x"3f71832b",
   627 => x"88830751",
   628 => x"fae13f71",
   629 => x"b00c833d",
   630 => x"0d04fe3d",
   631 => x"0d029305",
   632 => x"33028405",
   633 => x"97053354",
   634 => x"52717327",
   635 => x"9438a051",
   636 => x"80e3853f",
   637 => x"81127081",
   638 => x"ff065152",
   639 => x"727226ee",
   640 => x"38843d0d",
   641 => x"04fe3d0d",
   642 => x"74708106",
   643 => x"53537185",
   644 => x"d0387281",
   645 => x"2a708106",
   646 => x"51527185",
   647 => x"ac387282",
   648 => x"2a708106",
   649 => x"51527185",
   650 => x"88387283",
   651 => x"2a708106",
   652 => x"51527184",
   653 => x"e4387284",
   654 => x"2a708106",
   655 => x"51527184",
   656 => x"c0387285",
   657 => x"2a708106",
   658 => x"51527184",
   659 => x"9c387286",
   660 => x"2a708106",
   661 => x"51527183",
   662 => x"f8387287",
   663 => x"2a708106",
   664 => x"51527183",
   665 => x"d4387288",
   666 => x"2a708106",
   667 => x"51527183",
   668 => x"b0387289",
   669 => x"2a708106",
   670 => x"51527183",
   671 => x"8c38728a",
   672 => x"2a708106",
   673 => x"51527182",
   674 => x"e838728b",
   675 => x"2a708106",
   676 => x"51527182",
   677 => x"c438728c",
   678 => x"2a708106",
   679 => x"51527182",
   680 => x"a038728d",
   681 => x"2a708106",
   682 => x"51527181",
   683 => x"fc38728e",
   684 => x"2a708106",
   685 => x"51527181",
   686 => x"d838728f",
   687 => x"2a708106",
   688 => x"51527181",
   689 => x"b4387290",
   690 => x"2a708106",
   691 => x"51527181",
   692 => x"90387291",
   693 => x"2a708106",
   694 => x"51527180",
   695 => x"ec387292",
   696 => x"2a708106",
   697 => x"51527180",
   698 => x"c8387293",
   699 => x"2a708106",
   700 => x"515271a6",
   701 => x"3872942a",
   702 => x"70810651",
   703 => x"52718b38",
   704 => x"80732483",
   705 => x"f438843d",
   706 => x"0d0481a6",
   707 => x"c05180e1",
   708 => x"813f7280",
   709 => x"25f03883",
   710 => x"e03981a6",
   711 => x"dc5180e0",
   712 => x"f13f7294",
   713 => x"2a708106",
   714 => x"51527180",
   715 => x"2ed238da",
   716 => x"3981a6f8",
   717 => x"5180e0da",
   718 => x"3f72932a",
   719 => x"70810651",
   720 => x"5271802e",
   721 => x"ffaf38d2",
   722 => x"3981a794",
   723 => x"5180e0c2",
   724 => x"3f72922a",
   725 => x"70810651",
   726 => x"5271802e",
   727 => x"ff8c38d1",
   728 => x"3981a7b0",
   729 => x"5180e0aa",
   730 => x"3f72912a",
   731 => x"70810651",
   732 => x"5271802e",
   733 => x"fee838d1",
   734 => x"3981a7d0",
   735 => x"5180e092",
   736 => x"3f72902a",
   737 => x"70810651",
   738 => x"5271802e",
   739 => x"fec438d1",
   740 => x"3981a7f0",
   741 => x"5180dffa",
   742 => x"3f728f2a",
   743 => x"70810651",
   744 => x"5271802e",
   745 => x"fea038d1",
   746 => x"3981a890",
   747 => x"5180dfe2",
   748 => x"3f728e2a",
   749 => x"70810651",
   750 => x"5271802e",
   751 => x"fdfc38d1",
   752 => x"3981a8b0",
   753 => x"5180dfca",
   754 => x"3f728d2a",
   755 => x"70810651",
   756 => x"5271802e",
   757 => x"fdd838d1",
   758 => x"3981a8c4",
   759 => x"5180dfb2",
   760 => x"3f728c2a",
   761 => x"70810651",
   762 => x"5271802e",
   763 => x"fdb438d1",
   764 => x"3981a8e4",
   765 => x"5180df9a",
   766 => x"3f728b2a",
   767 => x"70810651",
   768 => x"5271802e",
   769 => x"fd9038d1",
   770 => x"3981a98c",
   771 => x"5180df82",
   772 => x"3f728a2a",
   773 => x"70810651",
   774 => x"5271802e",
   775 => x"fcec38d1",
   776 => x"3981a9ac",
   777 => x"5180deea",
   778 => x"3f72892a",
   779 => x"70810651",
   780 => x"5271802e",
   781 => x"fcc838d1",
   782 => x"3981a9cc",
   783 => x"5180ded2",
   784 => x"3f72882a",
   785 => x"70810651",
   786 => x"5271802e",
   787 => x"fca438d1",
   788 => x"3981a9f4",
   789 => x"5180deba",
   790 => x"3f72872a",
   791 => x"70810651",
   792 => x"5271802e",
   793 => x"fc8038d1",
   794 => x"3981aa94",
   795 => x"5180dea2",
   796 => x"3f72862a",
   797 => x"70810651",
   798 => x"5271802e",
   799 => x"fbdc38d1",
   800 => x"3981aab4",
   801 => x"5180de8a",
   802 => x"3f72852a",
   803 => x"70810651",
   804 => x"5271802e",
   805 => x"fbb838d1",
   806 => x"3981aadc",
   807 => x"5180ddf2",
   808 => x"3f72842a",
   809 => x"70810651",
   810 => x"5271802e",
   811 => x"fb9438d1",
   812 => x"3981aafc",
   813 => x"5180ddda",
   814 => x"3f72832a",
   815 => x"70810651",
   816 => x"5271802e",
   817 => x"faf038d1",
   818 => x"3981ab9c",
   819 => x"5180ddc2",
   820 => x"3f72822a",
   821 => x"70810651",
   822 => x"5271802e",
   823 => x"facc38d1",
   824 => x"3981abc4",
   825 => x"5180ddaa",
   826 => x"3f72812a",
   827 => x"70810651",
   828 => x"5271802e",
   829 => x"faa838d1",
   830 => x"3981abe4",
   831 => x"5180dd92",
   832 => x"3f843d0d",
   833 => x"04fd3d0d",
   834 => x"81abf851",
   835 => x"80dd833f",
   836 => x"81ccfc08",
   837 => x"7008709e",
   838 => x"2a708106",
   839 => x"51525553",
   840 => x"81547283",
   841 => x"38725473",
   842 => x"802e88c4",
   843 => x"3881ac94",
   844 => x"5180dcde",
   845 => x"3f81ac9c",
   846 => x"5180dcd6",
   847 => x"3f81ccfc",
   848 => x"08841108",
   849 => x"709d2a81",
   850 => x"06515553",
   851 => x"73802e87",
   852 => x"b03881ac",
   853 => x"b85180dc",
   854 => x"b93f81ac",
   855 => x"c45180dc",
   856 => x"b13f81cc",
   857 => x"c40880d4",
   858 => x"11085254",
   859 => x"80dded3f",
   860 => x"81ace051",
   861 => x"80dc9b3f",
   862 => x"81ccc408",
   863 => x"80d01108",
   864 => x"525380dd",
   865 => x"d73f8a51",
   866 => x"80dbed3f",
   867 => x"81acfc51",
   868 => x"80dbff3f",
   869 => x"81ada051",
   870 => x"80dbf73f",
   871 => x"81ade851",
   872 => x"80dbef3f",
   873 => x"81aeb051",
   874 => x"80dbe73f",
   875 => x"81ccc408",
   876 => x"70085254",
   877 => x"80dda53f",
   878 => x"b00881ff",
   879 => x"0653728c",
   880 => x"279438a0",
   881 => x"5180dbb0",
   882 => x"3f811370",
   883 => x"81ff0651",
   884 => x"538c7326",
   885 => x"ee3881cc",
   886 => x"c4088411",
   887 => x"08525480",
   888 => x"dcfa3fb0",
   889 => x"0881ff06",
   890 => x"53728c27",
   891 => x"9438a051",
   892 => x"80db853f",
   893 => x"81137081",
   894 => x"ff065153",
   895 => x"8c7326ee",
   896 => x"3881ccc4",
   897 => x"08881108",
   898 => x"525480dc",
   899 => x"cf3fb008",
   900 => x"81ff0653",
   901 => x"728c2794",
   902 => x"38a05180",
   903 => x"dada3f81",
   904 => x"137081ff",
   905 => x"0651538c",
   906 => x"7326ee38",
   907 => x"81ccc408",
   908 => x"8c110852",
   909 => x"5480dca4",
   910 => x"3fb00881",
   911 => x"ff065372",
   912 => x"8c279438",
   913 => x"a05180da",
   914 => x"af3f8113",
   915 => x"7081ff06",
   916 => x"51538c73",
   917 => x"26ee3881",
   918 => x"aecc5180",
   919 => x"dab43f81",
   920 => x"ccc40890",
   921 => x"11085254",
   922 => x"80dbf13f",
   923 => x"b00881ff",
   924 => x"0653728c",
   925 => x"279438a0",
   926 => x"5180d9fc",
   927 => x"3f811370",
   928 => x"81ff0651",
   929 => x"538c7326",
   930 => x"ee3881cc",
   931 => x"c4089411",
   932 => x"08525480",
   933 => x"dbc63fb0",
   934 => x"0881ff06",
   935 => x"53728c27",
   936 => x"9438a051",
   937 => x"80d9d13f",
   938 => x"81137081",
   939 => x"ff065153",
   940 => x"8c7326ee",
   941 => x"3881ccc4",
   942 => x"08981108",
   943 => x"525480db",
   944 => x"9b3fb008",
   945 => x"81ff0653",
   946 => x"728c2794",
   947 => x"38a05180",
   948 => x"d9a63f81",
   949 => x"137081ff",
   950 => x"0651538c",
   951 => x"7326ee38",
   952 => x"81ccc408",
   953 => x"9c110852",
   954 => x"5480daf0",
   955 => x"3fb00881",
   956 => x"ff065372",
   957 => x"8c279438",
   958 => x"a05180d8",
   959 => x"fb3f8113",
   960 => x"7081ff06",
   961 => x"51538c73",
   962 => x"26ee3881",
   963 => x"aee85180",
   964 => x"d9803f81",
   965 => x"ccc40854",
   966 => x"810bb015",
   967 => x"0cb01408",
   968 => x"53728025",
   969 => x"f838a014",
   970 => x"085180da",
   971 => x"af3fb008",
   972 => x"81ff0653",
   973 => x"728c2794",
   974 => x"38a05180",
   975 => x"d8ba3f81",
   976 => x"137081ff",
   977 => x"0654548c",
   978 => x"7326ee38",
   979 => x"81ccc408",
   980 => x"a4110852",
   981 => x"5380da84",
   982 => x"3fb00881",
   983 => x"ff065372",
   984 => x"8c279438",
   985 => x"a05180d8",
   986 => x"8f3f8113",
   987 => x"7081ff06",
   988 => x"54548c73",
   989 => x"26ee3881",
   990 => x"ccc408a8",
   991 => x"11085253",
   992 => x"80d9d93f",
   993 => x"b00881ff",
   994 => x"0653728c",
   995 => x"279438a0",
   996 => x"5180d7e4",
   997 => x"3f811370",
   998 => x"81ff0654",
   999 => x"548c7326",
  1000 => x"ee3881cc",
  1001 => x"c408ac11",
  1002 => x"08525380",
  1003 => x"d9ae3fb0",
  1004 => x"0881ff06",
  1005 => x"53728c27",
  1006 => x"9438a051",
  1007 => x"80d7b93f",
  1008 => x"81137081",
  1009 => x"ff065454",
  1010 => x"8c7326ee",
  1011 => x"3881af84",
  1012 => x"5180d7be",
  1013 => x"3f81ccc4",
  1014 => x"0880e011",
  1015 => x"08525380",
  1016 => x"d8fa3f81",
  1017 => x"af985180",
  1018 => x"d7a83f81",
  1019 => x"ccc408b0",
  1020 => x"1108fe0a",
  1021 => x"06525480",
  1022 => x"d8e23f81",
  1023 => x"ccc40854",
  1024 => x"800bb015",
  1025 => x"0c81afac",
  1026 => x"5180d786",
  1027 => x"3f81afc4",
  1028 => x"5180d6fe",
  1029 => x"3f81ccc4",
  1030 => x"0880c011",
  1031 => x"08525380",
  1032 => x"d8ba3fb0",
  1033 => x"0881ff06",
  1034 => x"53729827",
  1035 => x"9438a051",
  1036 => x"80d6c53f",
  1037 => x"81137081",
  1038 => x"ff065454",
  1039 => x"987326ee",
  1040 => x"3881ccc4",
  1041 => x"0880c811",
  1042 => x"08525380",
  1043 => x"d88e3fb0",
  1044 => x"0881ff06",
  1045 => x"53729827",
  1046 => x"9438a051",
  1047 => x"80d6993f",
  1048 => x"81137081",
  1049 => x"ff065454",
  1050 => x"987326ee",
  1051 => x"3881afe0",
  1052 => x"5180d69e",
  1053 => x"3f81ccc4",
  1054 => x"0880c411",
  1055 => x"08525380",
  1056 => x"d7da3fb0",
  1057 => x"0881ff06",
  1058 => x"53729827",
  1059 => x"9438a051",
  1060 => x"80d5e53f",
  1061 => x"81137081",
  1062 => x"ff065454",
  1063 => x"987326ee",
  1064 => x"3881ccc4",
  1065 => x"0880cc11",
  1066 => x"08525380",
  1067 => x"d7ae3fb0",
  1068 => x"0881ff06",
  1069 => x"53729827",
  1070 => x"9438a051",
  1071 => x"80d5b93f",
  1072 => x"81137081",
  1073 => x"ff065454",
  1074 => x"987326ee",
  1075 => x"388a5180",
  1076 => x"d5a63f81",
  1077 => x"ccc408b4",
  1078 => x"110881af",
  1079 => x"fc535153",
  1080 => x"80d5af3f",
  1081 => x"725180d6",
  1082 => x"f33fa051",
  1083 => x"80d5893f",
  1084 => x"72862681",
  1085 => x"8e387210",
  1086 => x"1081bcb0",
  1087 => x"05547308",
  1088 => x"0481b090",
  1089 => x"5180d58a",
  1090 => x"3f81acc4",
  1091 => x"5180d582",
  1092 => x"3f81ccc4",
  1093 => x"0880d411",
  1094 => x"08525480",
  1095 => x"d6be3f81",
  1096 => x"ace05180",
  1097 => x"d4ec3f81",
  1098 => x"ccc40880",
  1099 => x"d0110852",
  1100 => x"5380d6a8",
  1101 => x"3f8a5180",
  1102 => x"d4be3f81",
  1103 => x"acfc5180",
  1104 => x"d4d03f81",
  1105 => x"ada05180",
  1106 => x"d4c83f81",
  1107 => x"ade85180",
  1108 => x"d4c03f81",
  1109 => x"aeb05180",
  1110 => x"d4b83f81",
  1111 => x"ccc40870",
  1112 => x"08525480",
  1113 => x"d5f63fb0",
  1114 => x"0881ff06",
  1115 => x"53f8cf39",
  1116 => x"81b09851",
  1117 => x"80d49b3f",
  1118 => x"f7b33981",
  1119 => x"b0a05180",
  1120 => x"d4903f81",
  1121 => x"ccc408b8",
  1122 => x"110881b0",
  1123 => x"ac535454",
  1124 => x"80d3ff3f",
  1125 => x"7252a051",
  1126 => x"80d49a3f",
  1127 => x"7251f0e5",
  1128 => x"3f8a5180",
  1129 => x"d3d23f80",
  1130 => x"0bb00c85",
  1131 => x"3d0d0481",
  1132 => x"b0c05180",
  1133 => x"d3dc3fcb",
  1134 => x"3981b0cc",
  1135 => x"5180d3d2",
  1136 => x"3fc13981",
  1137 => x"b0d85180",
  1138 => x"d3c83fff",
  1139 => x"b63981b0",
  1140 => x"dc5180d3",
  1141 => x"bd3fffab",
  1142 => x"3981b0e8",
  1143 => x"5180d3b2",
  1144 => x"3fffa039",
  1145 => x"81b0f451",
  1146 => x"80d3a73f",
  1147 => x"ff9539fe",
  1148 => x"3d0d8151",
  1149 => x"aafb3fb0",
  1150 => x"0881ff06",
  1151 => x"81ccc408",
  1152 => x"71b4120c",
  1153 => x"53b00c84",
  1154 => x"3d0d04fe",
  1155 => x"3d0d880a",
  1156 => x"53840a0b",
  1157 => x"81ccc008",
  1158 => x"8c110851",
  1159 => x"52528071",
  1160 => x"27953880",
  1161 => x"73708405",
  1162 => x"550c8072",
  1163 => x"70840554",
  1164 => x"0cff1151",
  1165 => x"70ed3880",
  1166 => x"0bb00c84",
  1167 => x"3d0d04fa",
  1168 => x"3d0d880a",
  1169 => x"57840a56",
  1170 => x"8151aaa5",
  1171 => x"3fb00883",
  1172 => x"ffff0654",
  1173 => x"73833890",
  1174 => x"54805574",
  1175 => x"742781c2",
  1176 => x"38750870",
  1177 => x"902c5253",
  1178 => x"80d3f13f",
  1179 => x"b00881ff",
  1180 => x"0652718a",
  1181 => x"279438a0",
  1182 => x"5180d1fc",
  1183 => x"3f811270",
  1184 => x"81ff0651",
  1185 => x"528a7226",
  1186 => x"ee387290",
  1187 => x"2b70902c",
  1188 => x"525280d3",
  1189 => x"c73fb008",
  1190 => x"81ff0652",
  1191 => x"718a2794",
  1192 => x"38a05180",
  1193 => x"d1d23f81",
  1194 => x"127081ff",
  1195 => x"0653538a",
  1196 => x"7226ee38",
  1197 => x"76087090",
  1198 => x"2c525380",
  1199 => x"d39e3fb0",
  1200 => x"0881ff06",
  1201 => x"52718a27",
  1202 => x"9438a051",
  1203 => x"80d1a93f",
  1204 => x"81127081",
  1205 => x"ff065152",
  1206 => x"8a7226ee",
  1207 => x"3872902b",
  1208 => x"70902c52",
  1209 => x"5280d2f4",
  1210 => x"3fb00881",
  1211 => x"ff065271",
  1212 => x"8a279438",
  1213 => x"a05180d0",
  1214 => x"ff3f8112",
  1215 => x"7081ff06",
  1216 => x"53538a72",
  1217 => x"26ee388a",
  1218 => x"5180d0ec",
  1219 => x"3f841784",
  1220 => x"17811770",
  1221 => x"83ffff06",
  1222 => x"58545757",
  1223 => x"737526fe",
  1224 => x"c03873b0",
  1225 => x"0c883d0d",
  1226 => x"04fd3d0d",
  1227 => x"8151a8c1",
  1228 => x"3fb00881",
  1229 => x"ff065473",
  1230 => x"802ea438",
  1231 => x"73842690",
  1232 => x"3881ccc0",
  1233 => x"0874710c",
  1234 => x"5373b00c",
  1235 => x"853d0d04",
  1236 => x"81ccc008",
  1237 => x"5380730c",
  1238 => x"73b00c85",
  1239 => x"3d0d0481",
  1240 => x"b2805180",
  1241 => x"d0ac3f81",
  1242 => x"b2905180",
  1243 => x"d0a43f81",
  1244 => x"ccc00870",
  1245 => x"08525380",
  1246 => x"d1e23f81",
  1247 => x"b2a05180",
  1248 => x"d0903f81",
  1249 => x"ccc00884",
  1250 => x"11085353",
  1251 => x"a05180d0",
  1252 => x"a43f81b2",
  1253 => x"b45180cf",
  1254 => x"f93f81cc",
  1255 => x"c0088811",
  1256 => x"085353a0",
  1257 => x"5180d08d",
  1258 => x"3f81b2c8",
  1259 => x"5180cfe2",
  1260 => x"3f81ccc0",
  1261 => x"088c1108",
  1262 => x"525380d1",
  1263 => x"9f3f8a51",
  1264 => x"80cfb53f",
  1265 => x"73b00c85",
  1266 => x"3d0d04bc",
  1267 => x"0802bc0c",
  1268 => x"f93d0d02",
  1269 => x"bc08fc05",
  1270 => x"0c880a0b",
  1271 => x"bc08f405",
  1272 => x"0cfc3d0d",
  1273 => x"823dbc08",
  1274 => x"f0050c81",
  1275 => x"51a7823f",
  1276 => x"b00881ff",
  1277 => x"06bc08f8",
  1278 => x"050c8251",
  1279 => x"a6f33fb0",
  1280 => x"08bc08f0",
  1281 => x"05082383",
  1282 => x"51a6e63f",
  1283 => x"b008bc08",
  1284 => x"f0050882",
  1285 => x"05238451",
  1286 => x"a6d73fb0",
  1287 => x"08bc08f0",
  1288 => x"05088405",
  1289 => x"238551a6",
  1290 => x"c83fb008",
  1291 => x"bc08f005",
  1292 => x"08860523",
  1293 => x"8651a6b9",
  1294 => x"3fb008bc",
  1295 => x"08f00508",
  1296 => x"88052387",
  1297 => x"51a6aa3f",
  1298 => x"b008bc08",
  1299 => x"f005088a",
  1300 => x"05238851",
  1301 => x"a69b3fb0",
  1302 => x"08bc08f0",
  1303 => x"05088c05",
  1304 => x"238951a6",
  1305 => x"8c3fb008",
  1306 => x"bc08f005",
  1307 => x"088e0523",
  1308 => x"800b81cc",
  1309 => x"c008708c",
  1310 => x"050851bc",
  1311 => x"08e4050c",
  1312 => x"bc08ec05",
  1313 => x"0cbc08ec",
  1314 => x"0508bc08",
  1315 => x"e4050827",
  1316 => x"818f38bc",
  1317 => x"08e40508",
  1318 => x"bc08e805",
  1319 => x"0cbc08f8",
  1320 => x"0508802e",
  1321 => x"81b638bc",
  1322 => x"08ec0508",
  1323 => x"10bc08f0",
  1324 => x"05080570",
  1325 => x"22bc08f4",
  1326 => x"05088205",
  1327 => x"2271902b",
  1328 => x"07bc08f4",
  1329 => x"05080cbc",
  1330 => x"08e4050c",
  1331 => x"bc08f805",
  1332 => x"0cbc08ec",
  1333 => x"05088105",
  1334 => x"7081ff06",
  1335 => x"bc08e405",
  1336 => x"0cbc08f8",
  1337 => x"050c860b",
  1338 => x"bc08ec05",
  1339 => x"08278838",
  1340 => x"800bbc08",
  1341 => x"e4050cbc",
  1342 => x"08e40508",
  1343 => x"bc08f405",
  1344 => x"088405bc",
  1345 => x"08e80508",
  1346 => x"ff05bc08",
  1347 => x"e8050cbc",
  1348 => x"08f4050c",
  1349 => x"bc08ec05",
  1350 => x"0cbc08e8",
  1351 => x"0508ff87",
  1352 => x"38bc08fc",
  1353 => x"05080d80",
  1354 => x"0bb00c89",
  1355 => x"3d0dbc0c",
  1356 => x"04bc08e4",
  1357 => x"0508bc08",
  1358 => x"f4050884",
  1359 => x"05bc08e8",
  1360 => x"0508ff05",
  1361 => x"bc08e805",
  1362 => x"0cbc08f4",
  1363 => x"050cbc08",
  1364 => x"ec050cbc",
  1365 => x"08e80508",
  1366 => x"802ec638",
  1367 => x"bc08ec05",
  1368 => x"0810bc08",
  1369 => x"f0050805",
  1370 => x"70227090",
  1371 => x"2bbc08f4",
  1372 => x"050808fc",
  1373 => x"80800671",
  1374 => x"902c07bc",
  1375 => x"08f40508",
  1376 => x"0c52bc08",
  1377 => x"e4050cbc",
  1378 => x"08f8050c",
  1379 => x"800bbc08",
  1380 => x"e4050cbc",
  1381 => x"08ec0508",
  1382 => x"8626ff95",
  1383 => x"38bc08ec",
  1384 => x"05088105",
  1385 => x"7081ff06",
  1386 => x"bc08f405",
  1387 => x"088405bc",
  1388 => x"08e80508",
  1389 => x"ff05bc08",
  1390 => x"e8050cbc",
  1391 => x"08f4050c",
  1392 => x"bc08ec05",
  1393 => x"0cbc08e4",
  1394 => x"050cbc08",
  1395 => x"e80508ff",
  1396 => x"8b38fecd",
  1397 => x"39fb3d0d",
  1398 => x"029f0533",
  1399 => x"79982b70",
  1400 => x"982c5154",
  1401 => x"55810a54",
  1402 => x"805672e8",
  1403 => x"25bd38e8",
  1404 => x"53751081",
  1405 => x"07738180",
  1406 => x"0a298180",
  1407 => x"0a057098",
  1408 => x"2c515456",
  1409 => x"807324e9",
  1410 => x"38807325",
  1411 => x"80c73873",
  1412 => x"812a810a",
  1413 => x"07738180",
  1414 => x"0a2981ff",
  1415 => x"0a057098",
  1416 => x"2c515454",
  1417 => x"728024e7",
  1418 => x"38ab3997",
  1419 => x"73259a38",
  1420 => x"9774812a",
  1421 => x"810a0771",
  1422 => x"81800a29",
  1423 => x"81ff0a05",
  1424 => x"70982c51",
  1425 => x"525553dc",
  1426 => x"39807324",
  1427 => x"ffa33872",
  1428 => x"8024ffbb",
  1429 => x"38745280",
  1430 => x"51b1b53f",
  1431 => x"7381ff06",
  1432 => x"51b2b33f",
  1433 => x"74528151",
  1434 => x"b1a63f73",
  1435 => x"882a7081",
  1436 => x"ff065253",
  1437 => x"b2a03f74",
  1438 => x"528251b1",
  1439 => x"933f7390",
  1440 => x"2a7081ff",
  1441 => x"065253b2",
  1442 => x"8d3f7452",
  1443 => x"8351b180",
  1444 => x"3f73982a",
  1445 => x"51b1ff3f",
  1446 => x"74528451",
  1447 => x"b0f23f75",
  1448 => x"81ff0651",
  1449 => x"b1f03f74",
  1450 => x"528551b0",
  1451 => x"e33f7588",
  1452 => x"2a7081ff",
  1453 => x"065253b1",
  1454 => x"dd3f7452",
  1455 => x"8651b0d0",
  1456 => x"3f75902a",
  1457 => x"7081ff06",
  1458 => x"5254b1ca",
  1459 => x"3f745287",
  1460 => x"51b0bd3f",
  1461 => x"75982a51",
  1462 => x"b1bc3f87",
  1463 => x"3d0d04f2",
  1464 => x"3d0d0280",
  1465 => x"c3053302",
  1466 => x"840580c7",
  1467 => x"05338180",
  1468 => x"0a712b98",
  1469 => x"2a81ccc0",
  1470 => x"088c1108",
  1471 => x"71084453",
  1472 => x"565c5557",
  1473 => x"80730c80",
  1474 => x"7071725c",
  1475 => x"5a5e5b80",
  1476 => x"56757a27",
  1477 => x"80d73881",
  1478 => x"772783ce",
  1479 => x"387783ff",
  1480 => x"ff068119",
  1481 => x"71101084",
  1482 => x"0a057930",
  1483 => x"7a823270",
  1484 => x"30728025",
  1485 => x"71802507",
  1486 => x"56585841",
  1487 => x"57595c7b",
  1488 => x"802e83d5",
  1489 => x"38821522",
  1490 => x"5372902b",
  1491 => x"70902c54",
  1492 => x"55727b25",
  1493 => x"8338725b",
  1494 => x"7c732583",
  1495 => x"38725d81",
  1496 => x"167081ff",
  1497 => x"06575e79",
  1498 => x"7626ffb1",
  1499 => x"38811970",
  1500 => x"81ff065a",
  1501 => x"5680e579",
  1502 => x"27ff9438",
  1503 => x"987d3590",
  1504 => x"2b70902c",
  1505 => x"7c309871",
  1506 => x"35902b70",
  1507 => x"902c5c5c",
  1508 => x"55565477",
  1509 => x"54777525",
  1510 => x"83387454",
  1511 => x"73902b70",
  1512 => x"902c5d55",
  1513 => x"7b54807c",
  1514 => x"2583d738",
  1515 => x"73902b70",
  1516 => x"902c5f56",
  1517 => x"80705d58",
  1518 => x"80705a56",
  1519 => x"757a2780",
  1520 => x"e4388177",
  1521 => x"27838c38",
  1522 => x"7783ffff",
  1523 => x"06811971",
  1524 => x"1010840a",
  1525 => x"0579307a",
  1526 => x"82327030",
  1527 => x"72802571",
  1528 => x"80250753",
  1529 => x"51575357",
  1530 => x"59547380",
  1531 => x"2e83a438",
  1532 => x"82152254",
  1533 => x"73902b70",
  1534 => x"902c719f",
  1535 => x"2c707232",
  1536 => x"7131799f",
  1537 => x"2c707b32",
  1538 => x"71315154",
  1539 => x"51565653",
  1540 => x"72742583",
  1541 => x"38745681",
  1542 => x"197081ff",
  1543 => x"065a5579",
  1544 => x"7926ffa4",
  1545 => x"387d7635",
  1546 => x"982b7098",
  1547 => x"2c53547b",
  1548 => x"51fba23f",
  1549 => x"811c7081",
  1550 => x"ff065d59",
  1551 => x"80e57c27",
  1552 => x"fef63881",
  1553 => x"ccc0087f",
  1554 => x"710c5880",
  1555 => x"5281c19c",
  1556 => x"51b1b33f",
  1557 => x"81f0dc08",
  1558 => x"80f3ca0b",
  1559 => x"81f0dc0c",
  1560 => x"5f805280",
  1561 => x"51ada93f",
  1562 => x"81b2d851",
  1563 => x"80c6a33f",
  1564 => x"7c5180c7",
  1565 => x"e73f8052",
  1566 => x"8751ad94",
  1567 => x"3f81b2e0",
  1568 => x"5180c68e",
  1569 => x"3f7a5180",
  1570 => x"c7d23f80",
  1571 => x"d2528051",
  1572 => x"acfe3f81",
  1573 => x"b2e85180",
  1574 => x"c5f83f76",
  1575 => x"5180c7bc",
  1576 => x"3f80c052",
  1577 => x"8751ace8",
  1578 => x"3f81b2f0",
  1579 => x"5180c5e2",
  1580 => x"3f7980e6",
  1581 => x"295180c7",
  1582 => x"a33f7e81",
  1583 => x"f0dc0c90",
  1584 => x"3d0d0474",
  1585 => x"22537290",
  1586 => x"2b70902c",
  1587 => x"545c727b",
  1588 => x"25833872",
  1589 => x"5b7c7325",
  1590 => x"8338725d",
  1591 => x"81167081",
  1592 => x"ff06575e",
  1593 => x"757a27fd",
  1594 => x"84387783",
  1595 => x"ffff0681",
  1596 => x"19711010",
  1597 => x"880a0579",
  1598 => x"307a8232",
  1599 => x"70307280",
  1600 => x"25718025",
  1601 => x"07565840",
  1602 => x"41575954",
  1603 => x"73802eff",
  1604 => x"b2388215",
  1605 => x"2253ffae",
  1606 => x"39742253",
  1607 => x"fcab3974",
  1608 => x"22547390",
  1609 => x"2b70902c",
  1610 => x"719f2c70",
  1611 => x"72327131",
  1612 => x"799f2c70",
  1613 => x"7b327131",
  1614 => x"51545156",
  1615 => x"56537274",
  1616 => x"25833874",
  1617 => x"56811970",
  1618 => x"81ff065a",
  1619 => x"55787a27",
  1620 => x"fdd33877",
  1621 => x"83ffff06",
  1622 => x"81197110",
  1623 => x"10880a05",
  1624 => x"79307a82",
  1625 => x"32703072",
  1626 => x"80257180",
  1627 => x"25075351",
  1628 => x"57535759",
  1629 => x"5473802e",
  1630 => x"ffa53882",
  1631 => x"152254ff",
  1632 => x"a1398170",
  1633 => x"902b7090",
  1634 => x"2c405754",
  1635 => x"80705d58",
  1636 => x"fca63974",
  1637 => x"2254fcdc",
  1638 => x"39fa3d0d",
  1639 => x"8a5180c3",
  1640 => x"d73f97c8",
  1641 => x"3f9a8553",
  1642 => x"81b2f852",
  1643 => x"81b38c51",
  1644 => x"97cd3fa3",
  1645 => x"ef5381b3",
  1646 => x"905281b3",
  1647 => x"b85197bf",
  1648 => x"3fbbea53",
  1649 => x"81b3c052",
  1650 => x"81b3d051",
  1651 => x"97b13fbb",
  1652 => x"d15381b3",
  1653 => x"d85281b3",
  1654 => x"f45197a3",
  1655 => x"3fa6a953",
  1656 => x"81b3fc52",
  1657 => x"81b4a051",
  1658 => x"97953fbe",
  1659 => x"ad5381b4",
  1660 => x"a85281b4",
  1661 => x"c8519787",
  1662 => x"3fbfcb53",
  1663 => x"81b4cc52",
  1664 => x"81b4f051",
  1665 => x"96f93fbc",
  1666 => x"815381b4",
  1667 => x"f85281b0",
  1668 => x"905196eb",
  1669 => x"3fbcc253",
  1670 => x"81b59c52",
  1671 => x"81b5c451",
  1672 => x"96dd3fbd",
  1673 => x"ea5381b5",
  1674 => x"cc5281b5",
  1675 => x"ec5196cf",
  1676 => x"3f889b53",
  1677 => x"81b5f452",
  1678 => x"81b69051",
  1679 => x"96c13fa4",
  1680 => x"bf5381b6",
  1681 => x"985281b5",
  1682 => x"e45196b3",
  1683 => x"3fa48b53",
  1684 => x"81b6b452",
  1685 => x"81b6c851",
  1686 => x"96a53fb9",
  1687 => x"905381b6",
  1688 => x"d05281b6",
  1689 => x"ec519697",
  1690 => x"3fb9b653",
  1691 => x"81b6f452",
  1692 => x"81b78851",
  1693 => x"96893fa7",
  1694 => x"cb5381b7",
  1695 => x"905281b7",
  1696 => x"b45195fb",
  1697 => x"3f80c0a9",
  1698 => x"5381b7bc",
  1699 => x"5281b7cc",
  1700 => x"5195ec3f",
  1701 => x"80c2f453",
  1702 => x"81b7d052",
  1703 => x"81b7ec51",
  1704 => x"95dd3fbb",
  1705 => x"975381b7",
  1706 => x"f45281b8",
  1707 => x"8c5195cf",
  1708 => x"3f80c2fc",
  1709 => x"5381b894",
  1710 => x"5281b8a8",
  1711 => x"5195c03f",
  1712 => x"8ad65381",
  1713 => x"b8b05281",
  1714 => x"b8c45195",
  1715 => x"b23f8de6",
  1716 => x"5381b8c8",
  1717 => x"5281b8f0",
  1718 => x"5195a43f",
  1719 => x"bbb35381",
  1720 => x"b8f85281",
  1721 => x"b9985195",
  1722 => x"963f93a3",
  1723 => x"5381b9a0",
  1724 => x"5281b9b4",
  1725 => x"5195883f",
  1726 => x"88be5381",
  1727 => x"b9bc5281",
  1728 => x"b9c85194",
  1729 => x"fa3f89fc",
  1730 => x"5381b9cc",
  1731 => x"5281b9f4",
  1732 => x"5194ec3f",
  1733 => x"88be5381",
  1734 => x"b9fc5281",
  1735 => x"b2b05194",
  1736 => x"de3f8ac5",
  1737 => x"5381ba9c",
  1738 => x"5281baac",
  1739 => x"5194d03f",
  1740 => x"88b35381",
  1741 => x"a5bc5281",
  1742 => x"a5a05194",
  1743 => x"c23f80d1",
  1744 => x"d55381a5",
  1745 => x"bc5281a5",
  1746 => x"a85194b3",
  1747 => x"3f9b863f",
  1748 => x"94f93f81",
  1749 => x"0b81eff8",
  1750 => x"3481dcd8",
  1751 => x"337081ff",
  1752 => x"06555573",
  1753 => x"b23880c4",
  1754 => x"9b3fb008",
  1755 => x"903894e9",
  1756 => x"3f81eff8",
  1757 => x"335675e1",
  1758 => x"38883d0d",
  1759 => x"0480c497",
  1760 => x"3fb00881",
  1761 => x"ff065195",
  1762 => x"be3f94cd",
  1763 => x"3f81eff8",
  1764 => x"335675c5",
  1765 => x"38e33980",
  1766 => x"0b81dcd8",
  1767 => x"349bd63f",
  1768 => x"81ccfc08",
  1769 => x"70087087",
  1770 => x"2a810652",
  1771 => x"57547380",
  1772 => x"2e8f3876",
  1773 => x"802e81c5",
  1774 => x"38ff1770",
  1775 => x"81ff0658",
  1776 => x"5475862a",
  1777 => x"81065574",
  1778 => x"802eaa38",
  1779 => x"7680f738",
  1780 => x"81960b81",
  1781 => x"ccfc0884",
  1782 => x"110870ef",
  1783 => x"ff0a06ae",
  1784 => x"800a0784",
  1785 => x"130c5784",
  1786 => x"110870be",
  1787 => x"800a0784",
  1788 => x"130c5755",
  1789 => x"5775852a",
  1790 => x"81065574",
  1791 => x"802e9638",
  1792 => x"76ba3881",
  1793 => x"960b81cc",
  1794 => x"c408b811",
  1795 => x"08575557",
  1796 => x"800bb815",
  1797 => x"0c75842a",
  1798 => x"81065675",
  1799 => x"802efec6",
  1800 => x"3876802e",
  1801 => x"ac38ff17",
  1802 => x"7081ff06",
  1803 => x"585580c2",
  1804 => x"d33fb008",
  1805 => x"802efeb6",
  1806 => x"38fec239",
  1807 => x"ff177081",
  1808 => x"ff065855",
  1809 => x"d039ff17",
  1810 => x"7081ff06",
  1811 => x"5854ffa5",
  1812 => x"3981960b",
  1813 => x"81ccfc08",
  1814 => x"84110884",
  1815 => x"0a078412",
  1816 => x"0c5657a6",
  1817 => x"ce3f8052",
  1818 => x"81c19c51",
  1819 => x"a9983f80",
  1820 => x"c2923fb0",
  1821 => x"08802efd",
  1822 => x"f538fe81",
  1823 => x"39819676",
  1824 => x"822a8306",
  1825 => x"53768306",
  1826 => x"5257f4d3",
  1827 => x"3ffeb239",
  1828 => x"fe3d0d81",
  1829 => x"5195da3f",
  1830 => x"b00881ff",
  1831 => x"06538251",
  1832 => x"95cf3fb0",
  1833 => x"0881ff06",
  1834 => x"527251f4",
  1835 => x"b23f800b",
  1836 => x"b00c843d",
  1837 => x"0d04f93d",
  1838 => x"0d815195",
  1839 => x"b43fb008",
  1840 => x"81ff0681",
  1841 => x"bab45257",
  1842 => x"bdc83f81",
  1843 => x"bac851bd",
  1844 => x"c13ff880",
  1845 => x"809a8054",
  1846 => x"80557370",
  1847 => x"84055508",
  1848 => x"74708405",
  1849 => x"56085456",
  1850 => x"72a03881",
  1851 => x"157081ff",
  1852 => x"06565687",
  1853 => x"7527e338",
  1854 => x"76812e80",
  1855 => x"d8388a51",
  1856 => x"bcf63f76",
  1857 => x"b00c893d",
  1858 => x"0d048a51",
  1859 => x"bcea3f72",
  1860 => x"51bec93f",
  1861 => x"b00881ff",
  1862 => x"0653728c",
  1863 => x"279338a0",
  1864 => x"51bcd53f",
  1865 => x"81137081",
  1866 => x"ff065153",
  1867 => x"8c7326ef",
  1868 => x"3881bae0",
  1869 => x"51bcdb3f",
  1870 => x"7552a051",
  1871 => x"bcf73f75",
  1872 => x"51d9c23f",
  1873 => x"81157081",
  1874 => x"ff065656",
  1875 => x"877527ff",
  1876 => x"8938ffa4",
  1877 => x"39f88080",
  1878 => x"9a805480",
  1879 => x"53807470",
  1880 => x"8405560c",
  1881 => x"80747084",
  1882 => x"05560c81",
  1883 => x"137081ff",
  1884 => x"06545572",
  1885 => x"8726ff86",
  1886 => x"38807470",
  1887 => x"8405560c",
  1888 => x"80747084",
  1889 => x"05560c81",
  1890 => x"137081ff",
  1891 => x"06545587",
  1892 => x"7327ca38",
  1893 => x"fee839fe",
  1894 => x"3d0d8151",
  1895 => x"93d33fb0",
  1896 => x"0881ff06",
  1897 => x"81ccbc08",
  1898 => x"7188120c",
  1899 => x"53b00c84",
  1900 => x"3d0d0480",
  1901 => x"3d0d8151",
  1902 => x"94e93fb0",
  1903 => x"0883ffff",
  1904 => x"0651d2ef",
  1905 => x"3fb00883",
  1906 => x"ffff06b0",
  1907 => x"0c823d0d",
  1908 => x"04803d0d",
  1909 => x"81519399",
  1910 => x"3fb00881",
  1911 => x"ff06519e",
  1912 => x"a83f800b",
  1913 => x"b00c823d",
  1914 => x"0d04803d",
  1915 => x"0d81cd88",
  1916 => x"0851f8bb",
  1917 => x"9586a171",
  1918 => x"0c810bb0",
  1919 => x"0c823d0d",
  1920 => x"04fc3d0d",
  1921 => x"815192e9",
  1922 => x"3fb00881",
  1923 => x"ff065482",
  1924 => x"5192de3f",
  1925 => x"b00881ff",
  1926 => x"0681ccfc",
  1927 => x"08841108",
  1928 => x"70fe8f0a",
  1929 => x"0677982b",
  1930 => x"07515456",
  1931 => x"5372802e",
  1932 => x"86387181",
  1933 => x"0a075271",
  1934 => x"84160c71",
  1935 => x"b00c863d",
  1936 => x"0d04fd3d",
  1937 => x"0d81ccfc",
  1938 => x"08841108",
  1939 => x"55538151",
  1940 => x"929f3fb0",
  1941 => x"0881ff06",
  1942 => x"74dfffff",
  1943 => x"06545271",
  1944 => x"802e8738",
  1945 => x"73a08080",
  1946 => x"07538251",
  1947 => x"92833fb0",
  1948 => x"0881ff06",
  1949 => x"73efff0a",
  1950 => x"06555271",
  1951 => x"802e8738",
  1952 => x"7290800a",
  1953 => x"07548351",
  1954 => x"91e73fb0",
  1955 => x"0881ff06",
  1956 => x"74f7ff0a",
  1957 => x"06545271",
  1958 => x"802e8738",
  1959 => x"7388800a",
  1960 => x"07538451",
  1961 => x"91cb3fb0",
  1962 => x"0881ff06",
  1963 => x"73fbff0a",
  1964 => x"06555271",
  1965 => x"802e8738",
  1966 => x"7284800a",
  1967 => x"07548551",
  1968 => x"91af3fb0",
  1969 => x"0881ff06",
  1970 => x"74fdff0a",
  1971 => x"06545271",
  1972 => x"802e8738",
  1973 => x"7382800a",
  1974 => x"075381cc",
  1975 => x"fc087384",
  1976 => x"120c5472",
  1977 => x"b00c853d",
  1978 => x"0d04fa3d",
  1979 => x"0d880a0b",
  1980 => x"81ccc008",
  1981 => x"8c110859",
  1982 => x"55568151",
  1983 => x"90f33fb0",
  1984 => x"08902b70",
  1985 => x"902c5653",
  1986 => x"80772799",
  1987 => x"38807754",
  1988 => x"547383ff",
  1989 => x"ff067670",
  1990 => x"8405580c",
  1991 => x"ff137515",
  1992 => x"555372ed",
  1993 => x"38800bb0",
  1994 => x"0c883d0d",
  1995 => x"04fc3d0d",
  1996 => x"81bae851",
  1997 => x"b8dc3f81",
  1998 => x"ccfc0870",
  1999 => x"08709e2a",
  2000 => x"70810651",
  2001 => x"54545481",
  2002 => x"53718338",
  2003 => x"71537280",
  2004 => x"2e80d238",
  2005 => x"81baf851",
  2006 => x"b8b83f81",
  2007 => x"5190923f",
  2008 => x"b00881ff",
  2009 => x"0681bae8",
  2010 => x"5255b8a6",
  2011 => x"3f74802e",
  2012 => x"ab3881bb",
  2013 => x"8051b89a",
  2014 => x"3f81ccfc",
  2015 => x"08841108",
  2016 => x"70fd0a06",
  2017 => x"54545474",
  2018 => x"802e8638",
  2019 => x"72820a07",
  2020 => x"52718415",
  2021 => x"0c71b00c",
  2022 => x"863d0d04",
  2023 => x"81b09851",
  2024 => x"b7f03fce",
  2025 => x"3981b098",
  2026 => x"51b7e73f",
  2027 => x"81baf851",
  2028 => x"b7e03f81",
  2029 => x"518fba3f",
  2030 => x"b00881ff",
  2031 => x"0681bae8",
  2032 => x"5255b7ce",
  2033 => x"3f74ffaa",
  2034 => x"38d239fd",
  2035 => x"3d0d8151",
  2036 => x"8f9f3fb0",
  2037 => x"0881ff06",
  2038 => x"81bb8c52",
  2039 => x"54b7b33f",
  2040 => x"73a43881",
  2041 => x"b09051b7",
  2042 => x"a93f81cc",
  2043 => x"fc088411",
  2044 => x"0870fb0a",
  2045 => x"0684130c",
  2046 => x"53538a51",
  2047 => x"b6fa3f73",
  2048 => x"b00c853d",
  2049 => x"0d0481ac",
  2050 => x"b851b786",
  2051 => x"3f81ccfc",
  2052 => x"08841108",
  2053 => x"70840a07",
  2054 => x"84130c53",
  2055 => x"538a51b6",
  2056 => x"d73f73b0",
  2057 => x"0c853d0d",
  2058 => x"04fd3d0d",
  2059 => x"81dcd408",
  2060 => x"52f881c0",
  2061 => x"8e800b81",
  2062 => x"ccfc0855",
  2063 => x"5371802e",
  2064 => x"80f73872",
  2065 => x"81ff0684",
  2066 => x"150c81cc",
  2067 => x"b8337081",
  2068 => x"ff065152",
  2069 => x"71802e80",
  2070 => x"c238729f",
  2071 => x"2a731007",
  2072 => x"5381dcd8",
  2073 => x"337081ff",
  2074 => x"06515271",
  2075 => x"802ed438",
  2076 => x"800b81dc",
  2077 => x"d83491fd",
  2078 => x"3f81ccc8",
  2079 => x"33547380",
  2080 => x"e23881cc",
  2081 => x"fc087381",
  2082 => x"ff068412",
  2083 => x"0c81ccb8",
  2084 => x"337081ff",
  2085 => x"06515354",
  2086 => x"71c03872",
  2087 => x"812a739f",
  2088 => x"2b0753ff",
  2089 => x"bc397281",
  2090 => x"2a739f2b",
  2091 => x"075380fd",
  2092 => x"51b8f23f",
  2093 => x"81ccfc08",
  2094 => x"547281ff",
  2095 => x"0684150c",
  2096 => x"81ccb833",
  2097 => x"7081ff06",
  2098 => x"53547180",
  2099 => x"2ed83872",
  2100 => x"9f2a7310",
  2101 => x"075380fd",
  2102 => x"51b8ca3f",
  2103 => x"81ccfc08",
  2104 => x"54d73980",
  2105 => x"0bb00c85",
  2106 => x"3d0d04f7",
  2107 => x"3d0d853d",
  2108 => x"54965381",
  2109 => x"bba05273",
  2110 => x"51bbe83f",
  2111 => x"9ea63f81",
  2112 => x"518cee3f",
  2113 => x"80528051",
  2114 => x"9c863f73",
  2115 => x"53805281",
  2116 => x"c19c51b0",
  2117 => x"c53f8052",
  2118 => x"81519bf4",
  2119 => x"3f735382",
  2120 => x"5281c19c",
  2121 => x"51b0b33f",
  2122 => x"80528251",
  2123 => x"9be23f73",
  2124 => x"53815281",
  2125 => x"c19c51b0",
  2126 => x"a13f8052",
  2127 => x"84519bd0",
  2128 => x"3f735384",
  2129 => x"5281c19c",
  2130 => x"51b08f3f",
  2131 => x"80528551",
  2132 => x"9bbe3f73",
  2133 => x"53905281",
  2134 => x"c19c51af",
  2135 => x"fd3f8052",
  2136 => x"86519bac",
  2137 => x"3f735383",
  2138 => x"5281c19c",
  2139 => x"51afeb3f",
  2140 => x"8b3d0d04",
  2141 => x"fef53f80",
  2142 => x"0bb00c04",
  2143 => x"fc3d0d81",
  2144 => x"9fb85480",
  2145 => x"55845274",
  2146 => x"519b853f",
  2147 => x"80537370",
  2148 => x"81055533",
  2149 => x"519bff3f",
  2150 => x"81137081",
  2151 => x"ff065153",
  2152 => x"80dc7327",
  2153 => x"e9388115",
  2154 => x"7081ff06",
  2155 => x"56538775",
  2156 => x"27d33880",
  2157 => x"0bb00c86",
  2158 => x"3d0d04fd",
  2159 => x"3d0d81cc",
  2160 => x"b8337081",
  2161 => x"ff065454",
  2162 => x"72bf26ac",
  2163 => x"3881ccb8",
  2164 => x"337081ff",
  2165 => x"0681ccbc",
  2166 => x"08528812",
  2167 => x"0c5480e4",
  2168 => x"5280c3bb",
  2169 => x"518fee3f",
  2170 => x"81ccb833",
  2171 => x"81055372",
  2172 => x"81ccb834",
  2173 => x"853d0d04",
  2174 => x"80e45280",
  2175 => x"c492518f",
  2176 => x"d43f81cc",
  2177 => x"b8338105",
  2178 => x"537281cc",
  2179 => x"b834853d",
  2180 => x"0d04fd3d",
  2181 => x"0d81ccb8",
  2182 => x"337081ff",
  2183 => x"06545472",
  2184 => x"bf2680c9",
  2185 => x"3881ccb8",
  2186 => x"337081ff",
  2187 => x"0681ccbc",
  2188 => x"08568816",
  2189 => x"0c5381cc",
  2190 => x"b8337081",
  2191 => x"ff065553",
  2192 => x"73bf2e80",
  2193 => x"d13880e4",
  2194 => x"5280c492",
  2195 => x"518f863f",
  2196 => x"81ccb833",
  2197 => x"81055372",
  2198 => x"81ccb834",
  2199 => x"81ccb833",
  2200 => x"80ff0653",
  2201 => x"7281ccb8",
  2202 => x"34853d0d",
  2203 => x"0481ccb8",
  2204 => x"337081ff",
  2205 => x"0680ff71",
  2206 => x"3181ccbc",
  2207 => x"08528812",
  2208 => x"0c555381",
  2209 => x"ccb83370",
  2210 => x"81ff0655",
  2211 => x"5373bf2e",
  2212 => x"098106ff",
  2213 => x"b13880ce",
  2214 => x"905280c4",
  2215 => x"92518eb5",
  2216 => x"3f81ccb8",
  2217 => x"33810553",
  2218 => x"7281ccb8",
  2219 => x"3481ccb8",
  2220 => x"3380ff06",
  2221 => x"537281cc",
  2222 => x"b834853d",
  2223 => x"0d04810b",
  2224 => x"81ccc834",
  2225 => x"04fe3d0d",
  2226 => x"81cd8008",
  2227 => x"98110870",
  2228 => x"842a7081",
  2229 => x"06515353",
  2230 => x"5370802e",
  2231 => x"8d3871ef",
  2232 => x"0698140c",
  2233 => x"810b81dc",
  2234 => x"d834843d",
  2235 => x"0d04fb3d",
  2236 => x"0d81ccfc",
  2237 => x"08700881",
  2238 => x"0a0681dc",
  2239 => x"d40c54b4",
  2240 => x"c73fb4ea",
  2241 => x"3f8f8b3f",
  2242 => x"81cd8008",
  2243 => x"98110888",
  2244 => x"0798120c",
  2245 => x"5481dcd4",
  2246 => x"0880f6e2",
  2247 => x"55537284",
  2248 => x"38888054",
  2249 => x"7381f0dc",
  2250 => x"0c72802e",
  2251 => x"84b03881",
  2252 => x"a68451b0",
  2253 => x"dd3f8c51",
  2254 => x"b0be3f81",
  2255 => x"bba051b0",
  2256 => x"d13f81dc",
  2257 => x"d408802e",
  2258 => x"81e83881",
  2259 => x"bbb851b0",
  2260 => x"c13f81dc",
  2261 => x"d4085473",
  2262 => x"802e82d3",
  2263 => x"3881ccc0",
  2264 => x"08548174",
  2265 => x"0c81ccfc",
  2266 => x"08841108",
  2267 => x"70565755",
  2268 => x"805373fe",
  2269 => x"8f0a0673",
  2270 => x"982b0770",
  2271 => x"84170c81",
  2272 => x"147081ff",
  2273 => x"06515454",
  2274 => x"8f7327e6",
  2275 => x"38758416",
  2276 => x"0c81ccc4",
  2277 => x"0854800b",
  2278 => x"b8150c80",
  2279 => x"0bf88080",
  2280 => x"9e800ca0",
  2281 => x"808d0a08",
  2282 => x"51b1b13f",
  2283 => x"8a51afc8",
  2284 => x"3f825280",
  2285 => x"c5be518c",
  2286 => x"9c3ff881",
  2287 => x"c08e800b",
  2288 => x"81ccfc08",
  2289 => x"565481dc",
  2290 => x"d408802e",
  2291 => x"81b73873",
  2292 => x"81ff0684",
  2293 => x"160c81cc",
  2294 => x"b8337081",
  2295 => x"ff065456",
  2296 => x"72802e80",
  2297 => x"c238739f",
  2298 => x"2a741007",
  2299 => x"5481dcd8",
  2300 => x"337081ff",
  2301 => x"06575375",
  2302 => x"802ed438",
  2303 => x"800b81dc",
  2304 => x"d8348af1",
  2305 => x"3f81ccc8",
  2306 => x"33557482",
  2307 => x"dc3881cc",
  2308 => x"fc087481",
  2309 => x"ff068412",
  2310 => x"0c81ccb8",
  2311 => x"337081ff",
  2312 => x"06555755",
  2313 => x"72c03873",
  2314 => x"812a749f",
  2315 => x"2b0754ff",
  2316 => x"bc3981bb",
  2317 => x"c451aeda",
  2318 => x"3f810a51",
  2319 => x"aed43f81",
  2320 => x"bbd851ae",
  2321 => x"cd3f81bc",
  2322 => x"8051aec6",
  2323 => x"3fb451b0",
  2324 => x"8b3f81bc",
  2325 => x"9451aeba",
  2326 => x"3f81bc9c",
  2327 => x"51aeb33f",
  2328 => x"81bca851",
  2329 => x"aeac3f81",
  2330 => x"dcd40854",
  2331 => x"73fdee38",
  2332 => x"be397381",
  2333 => x"2a749f2b",
  2334 => x"075480fd",
  2335 => x"51b1a63f",
  2336 => x"81ccfc08",
  2337 => x"557381ff",
  2338 => x"0684160c",
  2339 => x"81ccb833",
  2340 => x"7081ff06",
  2341 => x"56567480",
  2342 => x"2ed83873",
  2343 => x"9f2a7410",
  2344 => x"075480fd",
  2345 => x"51b0fe3f",
  2346 => x"81ccfc08",
  2347 => x"55d73981",
  2348 => x"ccc40874",
  2349 => x"b4120c56",
  2350 => x"818051c4",
  2351 => x"f63f8280",
  2352 => x"51c4f03f",
  2353 => x"848351c4",
  2354 => x"ea3f86f1",
  2355 => x"51c4e43f",
  2356 => x"888351c4",
  2357 => x"de3f81cc",
  2358 => x"fc087008",
  2359 => x"709e2a70",
  2360 => x"81065155",
  2361 => x"56548155",
  2362 => x"72802e80",
  2363 => x"f7387481",
  2364 => x"ff068415",
  2365 => x"0870fd0a",
  2366 => x"06585653",
  2367 => x"72802e86",
  2368 => x"3874820a",
  2369 => x"07567584",
  2370 => x"150c8414",
  2371 => x"08be800a",
  2372 => x"0784150c",
  2373 => x"84140884",
  2374 => x"0a078415",
  2375 => x"0c81ccc4",
  2376 => x"0855800b",
  2377 => x"b8160c81",
  2378 => x"ccc00854",
  2379 => x"81740c93",
  2380 => x"c45280c2",
  2381 => x"fc51899d",
  2382 => x"3f87e852",
  2383 => x"80c3bb51",
  2384 => x"89933fe8",
  2385 => x"d43f81cc",
  2386 => x"c0085481",
  2387 => x"740c81cc",
  2388 => x"fc088411",
  2389 => x"08705657",
  2390 => x"558053fc",
  2391 => x"953995c4",
  2392 => x"3ffbcc39",
  2393 => x"7255ff86",
  2394 => x"39b2eb3f",
  2395 => x"800b81ef",
  2396 => x"f034800b",
  2397 => x"81efec34",
  2398 => x"800b81ef",
  2399 => x"f40c04fc",
  2400 => x"3d0d7652",
  2401 => x"81efec33",
  2402 => x"70101010",
  2403 => x"71100581",
  2404 => x"dcdc0552",
  2405 => x"54b7da3f",
  2406 => x"775281ef",
  2407 => x"ec337090",
  2408 => x"29713170",
  2409 => x"101081df",
  2410 => x"9c055355",
  2411 => x"55b7c23f",
  2412 => x"81efec33",
  2413 => x"70101081",
  2414 => x"ee9c057a",
  2415 => x"710c5481",
  2416 => x"05537281",
  2417 => x"efec3486",
  2418 => x"3d0d0480",
  2419 => x"3d0d81bc",
  2420 => x"ec51abbe",
  2421 => x"3f823d0d",
  2422 => x"04fe3d0d",
  2423 => x"81eff408",
  2424 => x"53728538",
  2425 => x"843d0d04",
  2426 => x"722db008",
  2427 => x"53800b81",
  2428 => x"eff40cb0",
  2429 => x"088c3881",
  2430 => x"bcec51ab",
  2431 => x"953f843d",
  2432 => x"0d0481c0",
  2433 => x"c851ab8a",
  2434 => x"3f7283ff",
  2435 => x"ff26aa38",
  2436 => x"81ff7327",
  2437 => x"96387252",
  2438 => x"9051ab99",
  2439 => x"3f8a51aa",
  2440 => x"d73f81bc",
  2441 => x"ec51aaea",
  2442 => x"3fd43972",
  2443 => x"528851ab",
  2444 => x"843f8a51",
  2445 => x"aac23fea",
  2446 => x"397252a0",
  2447 => x"51aaf63f",
  2448 => x"8a51aab4",
  2449 => x"3fdc39fa",
  2450 => x"3d0d02a3",
  2451 => x"05335675",
  2452 => x"8d2e80f4",
  2453 => x"38758832",
  2454 => x"70307780",
  2455 => x"ff327030",
  2456 => x"72802571",
  2457 => x"80250754",
  2458 => x"51565855",
  2459 => x"7495389f",
  2460 => x"76278c38",
  2461 => x"81eff033",
  2462 => x"5580ce75",
  2463 => x"27ae3888",
  2464 => x"3d0d0481",
  2465 => x"eff03356",
  2466 => x"75802ef3",
  2467 => x"388851a9",
  2468 => x"e73fa051",
  2469 => x"a9e23f88",
  2470 => x"51a9dd3f",
  2471 => x"81eff033",
  2472 => x"ff055776",
  2473 => x"81eff034",
  2474 => x"883d0d04",
  2475 => x"7551a9c8",
  2476 => x"3f81eff0",
  2477 => x"33811155",
  2478 => x"577381ef",
  2479 => x"f0347581",
  2480 => x"ef9c1834",
  2481 => x"883d0d04",
  2482 => x"8a51a9ac",
  2483 => x"3f81eff0",
  2484 => x"33811156",
  2485 => x"547481ef",
  2486 => x"f034800b",
  2487 => x"81ef9c15",
  2488 => x"34805680",
  2489 => x"0b81ef9c",
  2490 => x"17335654",
  2491 => x"74a02e83",
  2492 => x"38815474",
  2493 => x"802e9038",
  2494 => x"73802e8b",
  2495 => x"38811670",
  2496 => x"81ff0657",
  2497 => x"57dd3975",
  2498 => x"802ebf38",
  2499 => x"800b81ef",
  2500 => x"ec335555",
  2501 => x"747427ab",
  2502 => x"38735774",
  2503 => x"10101075",
  2504 => x"10057654",
  2505 => x"81ef9c53",
  2506 => x"81dcdc05",
  2507 => x"51b68e3f",
  2508 => x"b008802e",
  2509 => x"a6388115",
  2510 => x"7081ff06",
  2511 => x"56547675",
  2512 => x"26d93881",
  2513 => x"bcf051a8",
  2514 => x"c93f81bc",
  2515 => x"ec51a8c2",
  2516 => x"3f800b81",
  2517 => x"eff03488",
  2518 => x"3d0d0474",
  2519 => x"101081ee",
  2520 => x"9c057008",
  2521 => x"81eff40c",
  2522 => x"56800b81",
  2523 => x"eff034e7",
  2524 => x"39f73d0d",
  2525 => x"02af0533",
  2526 => x"59800b81",
  2527 => x"ef9c3381",
  2528 => x"ef9c5955",
  2529 => x"5673a02e",
  2530 => x"09810696",
  2531 => x"38811670",
  2532 => x"81ff0681",
  2533 => x"ef9c1170",
  2534 => x"33535957",
  2535 => x"5473a02e",
  2536 => x"ec388058",
  2537 => x"77792780",
  2538 => x"ea388077",
  2539 => x"33565474",
  2540 => x"742e8338",
  2541 => x"815474a0",
  2542 => x"2e9a3873",
  2543 => x"80c53874",
  2544 => x"a02e9138",
  2545 => x"81187081",
  2546 => x"ff065955",
  2547 => x"787826da",
  2548 => x"3880c039",
  2549 => x"81167081",
  2550 => x"ff0681ef",
  2551 => x"9c117033",
  2552 => x"57525757",
  2553 => x"73a02e09",
  2554 => x"8106d938",
  2555 => x"81167081",
  2556 => x"ff0681ef",
  2557 => x"9c117033",
  2558 => x"57525757",
  2559 => x"73a02ed4",
  2560 => x"38c23981",
  2561 => x"167081ff",
  2562 => x"0681ef9c",
  2563 => x"11595755",
  2564 => x"ff98398a",
  2565 => x"538b3dfc",
  2566 => x"05527651",
  2567 => x"b8e43f8b",
  2568 => x"3d0d04f7",
  2569 => x"3d0d02af",
  2570 => x"05335980",
  2571 => x"0b81ef9c",
  2572 => x"3381ef9c",
  2573 => x"59555673",
  2574 => x"a02e0981",
  2575 => x"06963881",
  2576 => x"167081ff",
  2577 => x"0681ef9c",
  2578 => x"11703353",
  2579 => x"59575473",
  2580 => x"a02eec38",
  2581 => x"80587779",
  2582 => x"2780ea38",
  2583 => x"80773356",
  2584 => x"5474742e",
  2585 => x"83388154",
  2586 => x"74a02e9a",
  2587 => x"387380c5",
  2588 => x"3874a02e",
  2589 => x"91388118",
  2590 => x"7081ff06",
  2591 => x"59557878",
  2592 => x"26da3880",
  2593 => x"c0398116",
  2594 => x"7081ff06",
  2595 => x"81ef9c11",
  2596 => x"70335752",
  2597 => x"575773a0",
  2598 => x"2e098106",
  2599 => x"d9388116",
  2600 => x"7081ff06",
  2601 => x"81ef9c11",
  2602 => x"70335752",
  2603 => x"575773a0",
  2604 => x"2ed438c2",
  2605 => x"39811670",
  2606 => x"81ff0681",
  2607 => x"ef9c1159",
  2608 => x"5755ff98",
  2609 => x"3990538b",
  2610 => x"3dfc0552",
  2611 => x"7651bacf",
  2612 => x"3f8b3d0d",
  2613 => x"04fc3d0d",
  2614 => x"8a51a59c",
  2615 => x"3f81bd84",
  2616 => x"51a5af3f",
  2617 => x"800b81ef",
  2618 => x"ec335353",
  2619 => x"72722780",
  2620 => x"f5387210",
  2621 => x"10107310",
  2622 => x"0581dcdc",
  2623 => x"05705254",
  2624 => x"a5903f72",
  2625 => x"842b7074",
  2626 => x"31822b81",
  2627 => x"df9c1133",
  2628 => x"51535571",
  2629 => x"802eb738",
  2630 => x"7351b1c2",
  2631 => x"3fb00881",
  2632 => x"ff065271",
  2633 => x"89269338",
  2634 => x"a051a4cc",
  2635 => x"3f811270",
  2636 => x"81ff0653",
  2637 => x"54897227",
  2638 => x"ef3881bd",
  2639 => x"9c51a4d2",
  2640 => x"3f747331",
  2641 => x"822b81df",
  2642 => x"9c0551a4",
  2643 => x"c53f8a51",
  2644 => x"a4a63f81",
  2645 => x"137081ff",
  2646 => x"0681efec",
  2647 => x"33545455",
  2648 => x"717326ff",
  2649 => x"8d388a51",
  2650 => x"a48e3f81",
  2651 => x"efec33b0",
  2652 => x"0c863d0d",
  2653 => x"04fe3d0d",
  2654 => x"81f0cc22",
  2655 => x"ff055170",
  2656 => x"81f0cc23",
  2657 => x"7083ffff",
  2658 => x"06517080",
  2659 => x"c43881f0",
  2660 => x"d0335170",
  2661 => x"81ff2eb9",
  2662 => x"38701010",
  2663 => x"1081effc",
  2664 => x"05527133",
  2665 => x"81f0d034",
  2666 => x"fe723481",
  2667 => x"f0d03370",
  2668 => x"10101081",
  2669 => x"effc0552",
  2670 => x"53821122",
  2671 => x"81f0cc23",
  2672 => x"84120853",
  2673 => x"722d81f0",
  2674 => x"cc225170",
  2675 => x"802effbe",
  2676 => x"38843d0d",
  2677 => x"04f93d0d",
  2678 => x"02aa0522",
  2679 => x"56805574",
  2680 => x"10101081",
  2681 => x"effc0570",
  2682 => x"33525270",
  2683 => x"81fe2e99",
  2684 => x"38811570",
  2685 => x"81ff0656",
  2686 => x"52748a2e",
  2687 => x"098106df",
  2688 => x"38810bb0",
  2689 => x"0c893d0d",
  2690 => x"0481f0d0",
  2691 => x"337081ff",
  2692 => x"0681f0cc",
  2693 => x"22535458",
  2694 => x"7281ff2e",
  2695 => x"b0387283",
  2696 => x"2b547076",
  2697 => x"2780de38",
  2698 => x"75713170",
  2699 => x"83ffff06",
  2700 => x"7481effc",
  2701 => x"17337083",
  2702 => x"2b81effe",
  2703 => x"11225658",
  2704 => x"56525757",
  2705 => x"7281ff2e",
  2706 => x"098106d6",
  2707 => x"38727234",
  2708 => x"75821323",
  2709 => x"7984130c",
  2710 => x"7781ff06",
  2711 => x"5473732e",
  2712 => x"96387610",
  2713 => x"101081ef",
  2714 => x"fc055374",
  2715 => x"73348051",
  2716 => x"70b00c89",
  2717 => x"3d0d0474",
  2718 => x"81f0d034",
  2719 => x"7581f0cc",
  2720 => x"238051ec",
  2721 => x"39707631",
  2722 => x"517081ef",
  2723 => x"fe1523ff",
  2724 => x"bc39ff3d",
  2725 => x"0d8a5271",
  2726 => x"10101081",
  2727 => x"eff40551",
  2728 => x"fe7134ff",
  2729 => x"127081ff",
  2730 => x"06535171",
  2731 => x"ea38ff0b",
  2732 => x"81f0d034",
  2733 => x"833d0d04",
  2734 => x"fe3d0d02",
  2735 => x"93053302",
  2736 => x"84059705",
  2737 => x"33545271",
  2738 => x"812e9238",
  2739 => x"7180d52e",
  2740 => x"bb3881bd",
  2741 => x"a051a1ba",
  2742 => x"3f843d0d",
  2743 => x"0481bdac",
  2744 => x"51a1af3f",
  2745 => x"72912e81",
  2746 => x"f6387291",
  2747 => x"24b53872",
  2748 => x"8c2e81f6",
  2749 => x"38728c24",
  2750 => x"80e33872",
  2751 => x"862e81d4",
  2752 => x"3881bdb8",
  2753 => x"51a18b3f",
  2754 => x"843d0d04",
  2755 => x"81bdc851",
  2756 => x"a1803f72",
  2757 => x"8926ea38",
  2758 => x"72101081",
  2759 => x"c0f40552",
  2760 => x"71080472",
  2761 => x"a82e81cd",
  2762 => x"38a87325",
  2763 => x"9c387280",
  2764 => x"c52e81cc",
  2765 => x"387280e1",
  2766 => x"2e098106",
  2767 => x"c43881bd",
  2768 => x"d451a0ce",
  2769 => x"3f843d0d",
  2770 => x"04729a2e",
  2771 => x"098106ff",
  2772 => x"b03881bd",
  2773 => x"e451a0ba",
  2774 => x"3f843d0d",
  2775 => x"04728f2e",
  2776 => x"098106ff",
  2777 => x"9c3881be",
  2778 => x"8051a0a6",
  2779 => x"3f843d0d",
  2780 => x"0481be9c",
  2781 => x"51a09b3f",
  2782 => x"843d0d04",
  2783 => x"81bba051",
  2784 => x"a0903f84",
  2785 => x"3d0d0481",
  2786 => x"beb451a0",
  2787 => x"853f843d",
  2788 => x"0d0481be",
  2789 => x"c8519ffa",
  2790 => x"3f843d0d",
  2791 => x"0481bed8",
  2792 => x"519fef3f",
  2793 => x"843d0d04",
  2794 => x"81beec51",
  2795 => x"9fe43f84",
  2796 => x"3d0d0481",
  2797 => x"bf88519f",
  2798 => x"d93f843d",
  2799 => x"0d0481bf",
  2800 => x"a0519fce",
  2801 => x"3f843d0d",
  2802 => x"0481bfb4",
  2803 => x"519fc33f",
  2804 => x"843d0d04",
  2805 => x"81bfc451",
  2806 => x"9fb83f84",
  2807 => x"3d0d0481",
  2808 => x"bfd4519f",
  2809 => x"ad3f843d",
  2810 => x"0d0481bf",
  2811 => x"e8519fa2",
  2812 => x"3f843d0d",
  2813 => x"0481bff8",
  2814 => x"519f973f",
  2815 => x"843d0d04",
  2816 => x"81c09851",
  2817 => x"9f8c3f84",
  2818 => x"3d0d04f7",
  2819 => x"3d0d02b3",
  2820 => x"05337c70",
  2821 => x"08c08080",
  2822 => x"0659545a",
  2823 => x"80567583",
  2824 => x"2b7707bf",
  2825 => x"e0800770",
  2826 => x"70840552",
  2827 => x"0871088c",
  2828 => x"2abffe80",
  2829 => x"06790771",
  2830 => x"982a728c",
  2831 => x"2a9fff06",
  2832 => x"73852a70",
  2833 => x"8f06759f",
  2834 => x"06565158",
  2835 => x"5d585255",
  2836 => x"58748d38",
  2837 => x"8116568f",
  2838 => x"7627c338",
  2839 => x"8b3d0d04",
  2840 => x"81c0b051",
  2841 => x"9eac3f75",
  2842 => x"519ff13f",
  2843 => x"8452b008",
  2844 => x"51ffbae6",
  2845 => x"3f81c0bc",
  2846 => x"519e973f",
  2847 => x"74528851",
  2848 => x"9eb33f84",
  2849 => x"52b00851",
  2850 => x"ffbacf3f",
  2851 => x"81c0c451",
  2852 => x"9e803f78",
  2853 => x"5290519e",
  2854 => x"9c3f8652",
  2855 => x"b00851ff",
  2856 => x"bab83f81",
  2857 => x"c0cc519d",
  2858 => x"e93f7251",
  2859 => x"9fae3f84",
  2860 => x"52b00851",
  2861 => x"ffbaa33f",
  2862 => x"81c0d451",
  2863 => x"9dd43f73",
  2864 => x"519f993f",
  2865 => x"8452b008",
  2866 => x"51ffba8e",
  2867 => x"3f81c0dc",
  2868 => x"519dbf3f",
  2869 => x"7752a051",
  2870 => x"9ddb3f8a",
  2871 => x"52b00851",
  2872 => x"ffb9f73f",
  2873 => x"7992388a",
  2874 => x"519d8d3f",
  2875 => x"8116568f",
  2876 => x"7627feaa",
  2877 => x"38fee539",
  2878 => x"7881ff06",
  2879 => x"527451fb",
  2880 => x"b73f8a51",
  2881 => x"9cf23fe4",
  2882 => x"39f83d0d",
  2883 => x"02ab0533",
  2884 => x"59805675",
  2885 => x"852be090",
  2886 => x"11e08012",
  2887 => x"0870982a",
  2888 => x"718c2a9f",
  2889 => x"ff067285",
  2890 => x"2a708f06",
  2891 => x"749f0655",
  2892 => x"51585b53",
  2893 => x"56595574",
  2894 => x"802e81a7",
  2895 => x"3875bf26",
  2896 => x"81af3881",
  2897 => x"c0e4519c",
  2898 => x"c93f7551",
  2899 => x"9e8e3f86",
  2900 => x"52b00851",
  2901 => x"ffb9833f",
  2902 => x"81c0bc51",
  2903 => x"9cb43f74",
  2904 => x"5288519c",
  2905 => x"d03f8452",
  2906 => x"b00851ff",
  2907 => x"b8ec3f81",
  2908 => x"c0c4519c",
  2909 => x"9d3f7652",
  2910 => x"90519cb9",
  2911 => x"3f8652b0",
  2912 => x"0851ffb8",
  2913 => x"d53f81c0",
  2914 => x"cc519c86",
  2915 => x"3f72519d",
  2916 => x"cb3f8452",
  2917 => x"b00851ff",
  2918 => x"b8c03f81",
  2919 => x"c0d4519b",
  2920 => x"f13f7351",
  2921 => x"9db63f84",
  2922 => x"52b00851",
  2923 => x"ffb8ab3f",
  2924 => x"81c0dc51",
  2925 => x"9bdc3f77",
  2926 => x"08c08080",
  2927 => x"0652a051",
  2928 => x"9bf33f8a",
  2929 => x"52b00851",
  2930 => x"ffb88f3f",
  2931 => x"7881b238",
  2932 => x"8a519ba4",
  2933 => x"3f805374",
  2934 => x"812e81df",
  2935 => x"3876862e",
  2936 => x"81bb3881",
  2937 => x"165680ff",
  2938 => x"7627fea7",
  2939 => x"388a3d0d",
  2940 => x"0481c0ec",
  2941 => x"519b9b3f",
  2942 => x"c016519c",
  2943 => x"df3f8652",
  2944 => x"b00851ff",
  2945 => x"b7d43f81",
  2946 => x"c0bc519b",
  2947 => x"853f7452",
  2948 => x"88519ba1",
  2949 => x"3f8452b0",
  2950 => x"0851ffb7",
  2951 => x"bd3f81c0",
  2952 => x"c4519aee",
  2953 => x"3f765290",
  2954 => x"519b8a3f",
  2955 => x"8652b008",
  2956 => x"51ffb7a6",
  2957 => x"3f81c0cc",
  2958 => x"519ad73f",
  2959 => x"72519c9c",
  2960 => x"3f8452b0",
  2961 => x"0851ffb7",
  2962 => x"913f81c0",
  2963 => x"d4519ac2",
  2964 => x"3f73519c",
  2965 => x"873f8452",
  2966 => x"b00851ff",
  2967 => x"b6fc3f81",
  2968 => x"c0dc519a",
  2969 => x"ad3f7708",
  2970 => x"c0808006",
  2971 => x"52a0519a",
  2972 => x"c43f8a52",
  2973 => x"b00851ff",
  2974 => x"b6e03f78",
  2975 => x"802efed0",
  2976 => x"387681ff",
  2977 => x"06527451",
  2978 => x"f8ae3f8a",
  2979 => x"5199e93f",
  2980 => x"80537481",
  2981 => x"2e098106",
  2982 => x"fec3389f",
  2983 => x"39728106",
  2984 => x"5776802e",
  2985 => x"febd3878",
  2986 => x"527751fa",
  2987 => x"de3f8116",
  2988 => x"5680ff76",
  2989 => x"27fcdc38",
  2990 => x"feb33974",
  2991 => x"5376862e",
  2992 => x"098106fe",
  2993 => x"9e38d639",
  2994 => x"fe3d0d74",
  2995 => x"02840597",
  2996 => x"05330288",
  2997 => x"059b0533",
  2998 => x"88130c8c",
  2999 => x"120c538c",
  3000 => x"13087081",
  3001 => x"2a810651",
  3002 => x"5271f438",
  3003 => x"8c130870",
  3004 => x"81ff06b0",
  3005 => x"0c51843d",
  3006 => x"0d04803d",
  3007 => x"0d728c11",
  3008 => x"0870872a",
  3009 => x"81328106",
  3010 => x"b00c5151",
  3011 => x"823d0d04",
  3012 => x"fd3d0d02",
  3013 => x"97053302",
  3014 => x"84059b05",
  3015 => x"337181b0",
  3016 => x"0781bf06",
  3017 => x"535454f8",
  3018 => x"80809880",
  3019 => x"71710c73",
  3020 => x"842a9007",
  3021 => x"710c738f",
  3022 => x"06710c52",
  3023 => x"7281ccd0",
  3024 => x"347381cc",
  3025 => x"d434853d",
  3026 => x"0d04fd3d",
  3027 => x"0d029705",
  3028 => x"3381ccd4",
  3029 => x"33547305",
  3030 => x"87060284",
  3031 => x"059a0522",
  3032 => x"81ccd033",
  3033 => x"54730570",
  3034 => x"81ff0672",
  3035 => x"81b00754",
  3036 => x"515454f8",
  3037 => x"80809880",
  3038 => x"71710c73",
  3039 => x"842a9007",
  3040 => x"710c738f",
  3041 => x"06710c52",
  3042 => x"7281ccd0",
  3043 => x"347381cc",
  3044 => x"d434853d",
  3045 => x"0d04ff3d",
  3046 => x"0d028f05",
  3047 => x"33f88080",
  3048 => x"98840c81",
  3049 => x"ccd03381",
  3050 => x"05517081",
  3051 => x"ccd03483",
  3052 => x"3d0d04ff",
  3053 => x"3d0d8052",
  3054 => x"7181b007",
  3055 => x"81bf06f8",
  3056 => x"80809880",
  3057 => x"0c900bf8",
  3058 => x"80809880",
  3059 => x"0c800bf8",
  3060 => x"80809880",
  3061 => x"0c805180",
  3062 => x"0bf88080",
  3063 => x"98840c81",
  3064 => x"117081ff",
  3065 => x"06515180",
  3066 => x"e57127eb",
  3067 => x"38811270",
  3068 => x"81ff0653",
  3069 => x"51877227",
  3070 => x"ffbe3881",
  3071 => x"b00bf880",
  3072 => x"8098800c",
  3073 => x"900bf880",
  3074 => x"8098800c",
  3075 => x"800bf880",
  3076 => x"8098800c",
  3077 => x"800b81cc",
  3078 => x"d034800b",
  3079 => x"81ccd434",
  3080 => x"833d0d04",
  3081 => x"ff3d0d80",
  3082 => x"c00bf880",
  3083 => x"8098800c",
  3084 => x"81a10bf8",
  3085 => x"80809880",
  3086 => x"0c81c00b",
  3087 => x"f8808098",
  3088 => x"800c81a4",
  3089 => x"0bf88080",
  3090 => x"98800c81",
  3091 => x"a60bf880",
  3092 => x"8098800c",
  3093 => x"81a20bf8",
  3094 => x"80809880",
  3095 => x"0caf0bf8",
  3096 => x"80809880",
  3097 => x"0ca50bf8",
  3098 => x"80809880",
  3099 => x"0c81810b",
  3100 => x"f8808098",
  3101 => x"800c9d0b",
  3102 => x"f8808098",
  3103 => x"800c81fa",
  3104 => x"0bf88080",
  3105 => x"98800c80",
  3106 => x"0bf88080",
  3107 => x"98800c80",
  3108 => x"527181b0",
  3109 => x"0781bf06",
  3110 => x"f8808098",
  3111 => x"800c900b",
  3112 => x"f8808098",
  3113 => x"800c800b",
  3114 => x"f8808098",
  3115 => x"800c8051",
  3116 => x"800bf880",
  3117 => x"8098840c",
  3118 => x"81117081",
  3119 => x"ff065151",
  3120 => x"80e57127",
  3121 => x"eb388112",
  3122 => x"7081ff06",
  3123 => x"53518772",
  3124 => x"27ffbe38",
  3125 => x"81b00bf8",
  3126 => x"80809880",
  3127 => x"0c900bf8",
  3128 => x"80809880",
  3129 => x"0c800bf8",
  3130 => x"80809880",
  3131 => x"0c800b81",
  3132 => x"ccd03480",
  3133 => x"0b81ccd4",
  3134 => x"3481af0b",
  3135 => x"f8808098",
  3136 => x"800c833d",
  3137 => x"0d04803d",
  3138 => x"0d028f05",
  3139 => x"337381f0",
  3140 => x"d40c5170",
  3141 => x"81f0d834",
  3142 => x"823d0d04",
  3143 => x"ee3d0d64",
  3144 => x"02840580",
  3145 => x"d7053302",
  3146 => x"880580db",
  3147 => x"05335957",
  3148 => x"59807681",
  3149 => x"0677812a",
  3150 => x"81067883",
  3151 => x"2b818006",
  3152 => x"79822a81",
  3153 => x"06575e41",
  3154 => x"5f5d81ff",
  3155 => x"42727d2e",
  3156 => x"09810683",
  3157 => x"387c4276",
  3158 => x"8a2e83b9",
  3159 => x"38881908",
  3160 => x"5574802e",
  3161 => x"83a43885",
  3162 => x"19335aff",
  3163 => x"53767a26",
  3164 => x"8e388419",
  3165 => x"33547377",
  3166 => x"26853876",
  3167 => x"74315374",
  3168 => x"13703354",
  3169 => x"587281ff",
  3170 => x"06831a33",
  3171 => x"70982b81",
  3172 => x"ff0a119b",
  3173 => x"2a81055b",
  3174 => x"45424081",
  3175 => x"53748338",
  3176 => x"74537281",
  3177 => x"ff064380",
  3178 => x"7a81ff06",
  3179 => x"545cff54",
  3180 => x"7673268b",
  3181 => x"38841933",
  3182 => x"53767327",
  3183 => x"83f43873",
  3184 => x"7481ff06",
  3185 => x"5553805a",
  3186 => x"797324ab",
  3187 => x"38747a2e",
  3188 => x"09810682",
  3189 => x"e1386098",
  3190 => x"2b81ff0a",
  3191 => x"119b2a82",
  3192 => x"1b337171",
  3193 => x"29117081",
  3194 => x"ff067871",
  3195 => x"298c1f08",
  3196 => x"0552455d",
  3197 => x"575d537f",
  3198 => x"63057081",
  3199 => x"ff067061",
  3200 => x"2b7081ff",
  3201 => x"067b622b",
  3202 => x"7081ff06",
  3203 => x"7b832a81",
  3204 => x"065f5358",
  3205 => x"525e4255",
  3206 => x"78802e8f",
  3207 => x"3881ccd0",
  3208 => x"33610556",
  3209 => x"7580e624",
  3210 => x"83c5387f",
  3211 => x"78296130",
  3212 => x"41577c7e",
  3213 => x"2c982b70",
  3214 => x"982c5555",
  3215 => x"73772581",
  3216 => x"8238ff1c",
  3217 => x"7d81065a",
  3218 => x"537c732e",
  3219 => x"83c4387e",
  3220 => x"86a63861",
  3221 => x"84eb387d",
  3222 => x"802e82a4",
  3223 => x"38791470",
  3224 => x"33705854",
  3225 => x"55805578",
  3226 => x"752e8538",
  3227 => x"72842a56",
  3228 => x"75832a70",
  3229 => x"81065153",
  3230 => x"72802e84",
  3231 => x"3881c055",
  3232 => x"75822a70",
  3233 => x"81065153",
  3234 => x"72802e85",
  3235 => x"3874b007",
  3236 => x"5575812a",
  3237 => x"70810651",
  3238 => x"5372802e",
  3239 => x"8538748c",
  3240 => x"07557581",
  3241 => x"06537280",
  3242 => x"2e853874",
  3243 => x"83075574",
  3244 => x"51f9e33f",
  3245 => x"7714982b",
  3246 => x"70982c55",
  3247 => x"56767424",
  3248 => x"ff9b3862",
  3249 => x"802e9538",
  3250 => x"61ff1d54",
  3251 => x"547c732e",
  3252 => x"81fb3873",
  3253 => x"51f9bf3f",
  3254 => x"7e81ea38",
  3255 => x"7f528151",
  3256 => x"f8e83f81",
  3257 => x"1d7081ff",
  3258 => x"065e547b",
  3259 => x"7d26fec2",
  3260 => x"3860527b",
  3261 => x"3070982b",
  3262 => x"70982c53",
  3263 => x"585bf8ca",
  3264 => x"3f605372",
  3265 => x"b00c943d",
  3266 => x"0d048219",
  3267 => x"33851a33",
  3268 => x"5b53fcf1",
  3269 => x"3981ccd4",
  3270 => x"33537287",
  3271 => x"26819a38",
  3272 => x"81135680",
  3273 => x"527581ff",
  3274 => x"0651f7e4",
  3275 => x"3f805372",
  3276 => x"b00c943d",
  3277 => x"0d047380",
  3278 => x"2eaf38ff",
  3279 => x"147081ff",
  3280 => x"06555a73",
  3281 => x"81ff2ea1",
  3282 => x"38747081",
  3283 => x"0556337c",
  3284 => x"057083ff",
  3285 => x"ff06ff16",
  3286 => x"7081ff06",
  3287 => x"575c5d53",
  3288 => x"7381ff2e",
  3289 => x"098106e1",
  3290 => x"3860982b",
  3291 => x"81ff0a11",
  3292 => x"9b2a707e",
  3293 => x"291e8c1c",
  3294 => x"08055c42",
  3295 => x"55fcf839",
  3296 => x"79147033",
  3297 => x"5259f88e",
  3298 => x"3f771498",
  3299 => x"2b70982c",
  3300 => x"55567377",
  3301 => x"25feac38",
  3302 => x"79147033",
  3303 => x"5259f7f6",
  3304 => x"3f771498",
  3305 => x"2b70982c",
  3306 => x"55567674",
  3307 => x"24d238fe",
  3308 => x"92397673",
  3309 => x"3154fc87",
  3310 => x"39805280",
  3311 => x"51f6d13f",
  3312 => x"8053feeb",
  3313 => x"397351f7",
  3314 => x"cd3ffe90",
  3315 => x"39617b32",
  3316 => x"7081ff06",
  3317 => x"55557d80",
  3318 => x"2efdf838",
  3319 => x"7a812a74",
  3320 => x"32705254",
  3321 => x"f7b03f7e",
  3322 => x"802efdf0",
  3323 => x"38d73981",
  3324 => x"ccd4337c",
  3325 => x"05538052",
  3326 => x"7281ff06",
  3327 => x"51f6913f",
  3328 => x"805376a0",
  3329 => x"2efdfc38",
  3330 => x"7f782961",
  3331 => x"304157fc",
  3332 => x"a1397e87",
  3333 => x"ad386185",
  3334 => x"eb387d80",
  3335 => x"2e80ec38",
  3336 => x"79147033",
  3337 => x"7c077052",
  3338 => x"54568055",
  3339 => x"78752e85",
  3340 => x"3872842a",
  3341 => x"5675832a",
  3342 => x"70810651",
  3343 => x"5372802e",
  3344 => x"843881c0",
  3345 => x"5575822a",
  3346 => x"70810651",
  3347 => x"5372802e",
  3348 => x"853874b0",
  3349 => x"07557581",
  3350 => x"2a708106",
  3351 => x"51537280",
  3352 => x"2e853874",
  3353 => x"8c075575",
  3354 => x"81065372",
  3355 => x"802e8538",
  3356 => x"74830755",
  3357 => x"7451f69e",
  3358 => x"3f771498",
  3359 => x"2b70982c",
  3360 => x"55537674",
  3361 => x"24ff9938",
  3362 => x"fcb93979",
  3363 => x"1470337c",
  3364 => x"075256f6",
  3365 => x"813f7714",
  3366 => x"982b7098",
  3367 => x"2c555973",
  3368 => x"7725fc9f",
  3369 => x"38791470",
  3370 => x"337c0752",
  3371 => x"56f5e73f",
  3372 => x"7714982b",
  3373 => x"70982c55",
  3374 => x"59767424",
  3375 => x"ce38fc83",
  3376 => x"397d802e",
  3377 => x"80f03879",
  3378 => x"14703370",
  3379 => x"58545580",
  3380 => x"5578752e",
  3381 => x"85387284",
  3382 => x"2a567583",
  3383 => x"2a708106",
  3384 => x"51537280",
  3385 => x"2e843881",
  3386 => x"c0557582",
  3387 => x"2a708106",
  3388 => x"51537280",
  3389 => x"2e853874",
  3390 => x"b0075575",
  3391 => x"812a7081",
  3392 => x"06515372",
  3393 => x"802e8538",
  3394 => x"748c0755",
  3395 => x"75810653",
  3396 => x"72802e85",
  3397 => x"38748307",
  3398 => x"55740970",
  3399 => x"81ff0652",
  3400 => x"53f4f33f",
  3401 => x"7714982b",
  3402 => x"70982c55",
  3403 => x"56767424",
  3404 => x"ff9538fb",
  3405 => x"8e397914",
  3406 => x"70337009",
  3407 => x"7081ff06",
  3408 => x"54585455",
  3409 => x"f4d03f77",
  3410 => x"14982b70",
  3411 => x"982c5559",
  3412 => x"737725fa",
  3413 => x"ee387914",
  3414 => x"70337009",
  3415 => x"7081ff06",
  3416 => x"54585455",
  3417 => x"f4b03f77",
  3418 => x"14982b70",
  3419 => x"982c5559",
  3420 => x"767424c2",
  3421 => x"38facc39",
  3422 => x"61802e81",
  3423 => x"ce387d80",
  3424 => x"2e80f738",
  3425 => x"79147033",
  3426 => x"70585455",
  3427 => x"80557875",
  3428 => x"2e853872",
  3429 => x"842a5675",
  3430 => x"832a7081",
  3431 => x"06515372",
  3432 => x"802e8438",
  3433 => x"81c05575",
  3434 => x"822a7081",
  3435 => x"06515372",
  3436 => x"802e8538",
  3437 => x"74b00755",
  3438 => x"75812a70",
  3439 => x"81065153",
  3440 => x"72802e85",
  3441 => x"38748c07",
  3442 => x"55758106",
  3443 => x"5372802e",
  3444 => x"85387483",
  3445 => x"07557409",
  3446 => x"7081ff06",
  3447 => x"70535753",
  3448 => x"f3b43f75",
  3449 => x"51f3af3f",
  3450 => x"7714982b",
  3451 => x"70982c55",
  3452 => x"55767424",
  3453 => x"ff8e38f9",
  3454 => x"ca397914",
  3455 => x"70337009",
  3456 => x"7081ff06",
  3457 => x"70555955",
  3458 => x"5659f38a",
  3459 => x"3f7551f3",
  3460 => x"853f7714",
  3461 => x"982b7098",
  3462 => x"2c555973",
  3463 => x"7725f9a3",
  3464 => x"38791470",
  3465 => x"33700970",
  3466 => x"81ff0670",
  3467 => x"55595556",
  3468 => x"59f2e33f",
  3469 => x"7551f2de",
  3470 => x"3f771498",
  3471 => x"2b70982c",
  3472 => x"55597674",
  3473 => x"24ffb338",
  3474 => x"f8f9397d",
  3475 => x"802e80f4",
  3476 => x"38791470",
  3477 => x"33705854",
  3478 => x"55805578",
  3479 => x"752e8538",
  3480 => x"72842a56",
  3481 => x"75832a70",
  3482 => x"81065153",
  3483 => x"72802e84",
  3484 => x"3881c055",
  3485 => x"75822a70",
  3486 => x"81065153",
  3487 => x"72802e85",
  3488 => x"3874b007",
  3489 => x"5575812a",
  3490 => x"70810651",
  3491 => x"5372802e",
  3492 => x"8538748c",
  3493 => x"07557581",
  3494 => x"06537280",
  3495 => x"2e853874",
  3496 => x"83075574",
  3497 => x"81ff0670",
  3498 => x"5256f1ea",
  3499 => x"3f7551f1",
  3500 => x"e53f7714",
  3501 => x"982b7098",
  3502 => x"2c555576",
  3503 => x"7424ff91",
  3504 => x"38f88039",
  3505 => x"79147033",
  3506 => x"70535753",
  3507 => x"f1c83f75",
  3508 => x"51f1c33f",
  3509 => x"7714982b",
  3510 => x"70982c55",
  3511 => x"59737725",
  3512 => x"f7e13879",
  3513 => x"14703370",
  3514 => x"535753f1",
  3515 => x"a93f7551",
  3516 => x"f1a43f77",
  3517 => x"14982b70",
  3518 => x"982c5559",
  3519 => x"767424c4",
  3520 => x"38f7c039",
  3521 => x"7d802e80",
  3522 => x"f2387914",
  3523 => x"70337c07",
  3524 => x"70525456",
  3525 => x"80557875",
  3526 => x"2e853872",
  3527 => x"842a5675",
  3528 => x"832a7081",
  3529 => x"06515372",
  3530 => x"802e8438",
  3531 => x"81c05575",
  3532 => x"822a7081",
  3533 => x"06515372",
  3534 => x"802e8538",
  3535 => x"74b00755",
  3536 => x"75812a70",
  3537 => x"81065153",
  3538 => x"72802e85",
  3539 => x"38748c07",
  3540 => x"55758106",
  3541 => x"5372802e",
  3542 => x"85387483",
  3543 => x"07557409",
  3544 => x"7081ff06",
  3545 => x"5256f0ae",
  3546 => x"3f771498",
  3547 => x"2b70982c",
  3548 => x"55537674",
  3549 => x"24ff9338",
  3550 => x"f6c93979",
  3551 => x"1470337c",
  3552 => x"07700970",
  3553 => x"81ff0654",
  3554 => x"555659f0",
  3555 => x"893f7714",
  3556 => x"982b7098",
  3557 => x"2c555973",
  3558 => x"7725f6a7",
  3559 => x"38791470",
  3560 => x"337c0770",
  3561 => x"097081ff",
  3562 => x"06545556",
  3563 => x"59efe73f",
  3564 => x"7714982b",
  3565 => x"70982c55",
  3566 => x"59767424",
  3567 => x"ffbd38f6",
  3568 => x"82396180",
  3569 => x"2e81d438",
  3570 => x"7d802e80",
  3571 => x"f9387914",
  3572 => x"70337c07",
  3573 => x"70525456",
  3574 => x"80557875",
  3575 => x"2e853872",
  3576 => x"842a5675",
  3577 => x"832a7081",
  3578 => x"06515372",
  3579 => x"802e8438",
  3580 => x"81c05575",
  3581 => x"822a7081",
  3582 => x"06515372",
  3583 => x"802e8538",
  3584 => x"74b00755",
  3585 => x"75812a70",
  3586 => x"81065153",
  3587 => x"72802e85",
  3588 => x"38748c07",
  3589 => x"55758106",
  3590 => x"5372802e",
  3591 => x"85387483",
  3592 => x"07557409",
  3593 => x"7081ff06",
  3594 => x"70535456",
  3595 => x"eee83f72",
  3596 => x"51eee33f",
  3597 => x"7714982b",
  3598 => x"70982c55",
  3599 => x"56767424",
  3600 => x"ff8c38f4",
  3601 => x"fe397914",
  3602 => x"70337c07",
  3603 => x"70097081",
  3604 => x"ff067055",
  3605 => x"53575753",
  3606 => x"eebc3f72",
  3607 => x"51eeb73f",
  3608 => x"7714982b",
  3609 => x"70982c55",
  3610 => x"59737725",
  3611 => x"f4d53879",
  3612 => x"1470337c",
  3613 => x"07700970",
  3614 => x"81ff0670",
  3615 => x"55535757",
  3616 => x"53ee933f",
  3617 => x"7251ee8e",
  3618 => x"3f771498",
  3619 => x"2b70982c",
  3620 => x"55597674",
  3621 => x"24ffaf38",
  3622 => x"f4a9397d",
  3623 => x"802e80f6",
  3624 => x"38791470",
  3625 => x"337c0770",
  3626 => x"52545680",
  3627 => x"5578752e",
  3628 => x"85387284",
  3629 => x"2a567583",
  3630 => x"2a708106",
  3631 => x"51537280",
  3632 => x"2e843881",
  3633 => x"c0557582",
  3634 => x"2a708106",
  3635 => x"51537280",
  3636 => x"2e853874",
  3637 => x"b0075575",
  3638 => x"812a7081",
  3639 => x"06515372",
  3640 => x"802e8538",
  3641 => x"748c0755",
  3642 => x"75810653",
  3643 => x"72802e85",
  3644 => x"38748307",
  3645 => x"557481ff",
  3646 => x"06705256",
  3647 => x"ed983f75",
  3648 => x"51ed933f",
  3649 => x"7714982b",
  3650 => x"70982c55",
  3651 => x"53767424",
  3652 => x"ff8f38f3",
  3653 => x"ae397914",
  3654 => x"70337c07",
  3655 => x"70535456",
  3656 => x"ecf43f72",
  3657 => x"51ecef3f",
  3658 => x"7714982b",
  3659 => x"70982c55",
  3660 => x"59737725",
  3661 => x"f38d3879",
  3662 => x"1470337c",
  3663 => x"07705354",
  3664 => x"56ecd33f",
  3665 => x"7251ecce",
  3666 => x"3f771498",
  3667 => x"2b70982c",
  3668 => x"55597674",
  3669 => x"24c038f2",
  3670 => x"ea39f83d",
  3671 => x"0d7a7d02",
  3672 => x"8805af05",
  3673 => x"335a5559",
  3674 => x"80747081",
  3675 => x"05563375",
  3676 => x"58565774",
  3677 => x"772e0981",
  3678 => x"06883876",
  3679 => x"b00c8a3d",
  3680 => x"0d047453",
  3681 => x"77527851",
  3682 => x"ef923fb0",
  3683 => x"0881ff06",
  3684 => x"77057083",
  3685 => x"ffff0677",
  3686 => x"70810559",
  3687 => x"33525855",
  3688 => x"74802ed7",
  3689 => x"38745377",
  3690 => x"527851ee",
  3691 => x"ef3fb008",
  3692 => x"81ff0677",
  3693 => x"057083ff",
  3694 => x"ff067770",
  3695 => x"81055933",
  3696 => x"52585574",
  3697 => x"ffbc38ff",
  3698 => x"b239fe3d",
  3699 => x"0d029305",
  3700 => x"335381f0",
  3701 => x"d8335281",
  3702 => x"f0d40851",
  3703 => x"eebe3fb0",
  3704 => x"0881ff06",
  3705 => x"b00c843d",
  3706 => x"0d04d282",
  3707 => x"3f04fb3d",
  3708 => x"0d777955",
  3709 => x"55805675",
  3710 => x"7524ab38",
  3711 => x"8074249d",
  3712 => x"38805373",
  3713 => x"52745180",
  3714 => x"e13fb008",
  3715 => x"5475802e",
  3716 => x"8538b008",
  3717 => x"305473b0",
  3718 => x"0c873d0d",
  3719 => x"04733076",
  3720 => x"81325754",
  3721 => x"dc397430",
  3722 => x"55815673",
  3723 => x"8025d238",
  3724 => x"ec39fa3d",
  3725 => x"0d787a57",
  3726 => x"55805776",
  3727 => x"7524a438",
  3728 => x"759f2c54",
  3729 => x"81537574",
  3730 => x"32743152",
  3731 => x"74519b3f",
  3732 => x"b0085476",
  3733 => x"802e8538",
  3734 => x"b0083054",
  3735 => x"73b00c88",
  3736 => x"3d0d0474",
  3737 => x"30558157",
  3738 => x"d739fc3d",
  3739 => x"0d767853",
  3740 => x"54815380",
  3741 => x"74732652",
  3742 => x"5572802e",
  3743 => x"98387080",
  3744 => x"2ea93880",
  3745 => x"7224a438",
  3746 => x"71107310",
  3747 => x"75722653",
  3748 => x"545272ea",
  3749 => x"38735178",
  3750 => x"83387451",
  3751 => x"70b00c86",
  3752 => x"3d0d0472",
  3753 => x"812a7281",
  3754 => x"2a535372",
  3755 => x"802ee638",
  3756 => x"717426ef",
  3757 => x"38737231",
  3758 => x"75740774",
  3759 => x"812a7481",
  3760 => x"2a555556",
  3761 => x"54e53910",
  3762 => x"10101010",
  3763 => x"10101010",
  3764 => x"10101010",
  3765 => x"10101010",
  3766 => x"10101010",
  3767 => x"10101010",
  3768 => x"10101010",
  3769 => x"10105351",
  3770 => x"047381ff",
  3771 => x"06738306",
  3772 => x"09810583",
  3773 => x"05101010",
  3774 => x"2b0772fc",
  3775 => x"060c5151",
  3776 => x"043c0472",
  3777 => x"72807281",
  3778 => x"06ff0509",
  3779 => x"72060571",
  3780 => x"1052720a",
  3781 => x"100a5372",
  3782 => x"ed385151",
  3783 => x"535104b0",
  3784 => x"08b408b8",
  3785 => x"08757580",
  3786 => x"f4b22d50",
  3787 => x"50b00856",
  3788 => x"b80cb40c",
  3789 => x"b00c5104",
  3790 => x"b008b408",
  3791 => x"b8087575",
  3792 => x"80f3ee2d",
  3793 => x"5050b008",
  3794 => x"56b80cb4",
  3795 => x"0cb00c51",
  3796 => x"04b008b4",
  3797 => x"08b80880",
  3798 => x"c5c52db8",
  3799 => x"0cb40cb0",
  3800 => x"0c04ff3d",
  3801 => x"0d028f05",
  3802 => x"3381cd8c",
  3803 => x"0852710c",
  3804 => x"800bb00c",
  3805 => x"833d0d04",
  3806 => x"ff3d0d02",
  3807 => x"8f053351",
  3808 => x"81f0dc08",
  3809 => x"52712db0",
  3810 => x"0881ff06",
  3811 => x"b00c833d",
  3812 => x"0d04fe3d",
  3813 => x"0d747033",
  3814 => x"53537180",
  3815 => x"2e933881",
  3816 => x"13725281",
  3817 => x"f0dc0853",
  3818 => x"53712d72",
  3819 => x"335271ef",
  3820 => x"38843d0d",
  3821 => x"04f43d0d",
  3822 => x"7f028405",
  3823 => x"bb053355",
  3824 => x"57880b8c",
  3825 => x"3d5b5989",
  3826 => x"5381caa4",
  3827 => x"52795186",
  3828 => x"923f7379",
  3829 => x"2e80ff38",
  3830 => x"78567390",
  3831 => x"2e80ec38",
  3832 => x"02a70558",
  3833 => x"768f0654",
  3834 => x"73892680",
  3835 => x"c2387518",
  3836 => x"b0155555",
  3837 => x"73753476",
  3838 => x"842aff17",
  3839 => x"7081ff06",
  3840 => x"58555775",
  3841 => x"df38781a",
  3842 => x"55757534",
  3843 => x"79703355",
  3844 => x"5573802e",
  3845 => x"93388115",
  3846 => x"745281f0",
  3847 => x"dc085755",
  3848 => x"752d7433",
  3849 => x"5473ef38",
  3850 => x"78b00c8e",
  3851 => x"3d0d0475",
  3852 => x"18b71555",
  3853 => x"55737534",
  3854 => x"76842aff",
  3855 => x"177081ff",
  3856 => x"06585557",
  3857 => x"75ff9d38",
  3858 => x"ffbc3984",
  3859 => x"70575902",
  3860 => x"a70558ff",
  3861 => x"8f398270",
  3862 => x"5759f439",
  3863 => x"f13d0d61",
  3864 => x"8d3d705b",
  3865 => x"5c5a807a",
  3866 => x"5657767a",
  3867 => x"24818538",
  3868 => x"7817548a",
  3869 => x"52745184",
  3870 => x"b83fb008",
  3871 => x"b0055372",
  3872 => x"74348117",
  3873 => x"578a5274",
  3874 => x"5184813f",
  3875 => x"b00855b0",
  3876 => x"08de38b0",
  3877 => x"08779f2a",
  3878 => x"1870812c",
  3879 => x"5a565680",
  3880 => x"78259e38",
  3881 => x"7817ff05",
  3882 => x"55751970",
  3883 => x"33555374",
  3884 => x"33733473",
  3885 => x"75348116",
  3886 => x"ff165656",
  3887 => x"777624e9",
  3888 => x"38761958",
  3889 => x"80783480",
  3890 => x"7a241770",
  3891 => x"81ff067c",
  3892 => x"70335657",
  3893 => x"55567280",
  3894 => x"2e933881",
  3895 => x"15735281",
  3896 => x"f0dc0858",
  3897 => x"55762d74",
  3898 => x"335372ef",
  3899 => x"3873b00c",
  3900 => x"913d0d04",
  3901 => x"ad7b3402",
  3902 => x"ad057a30",
  3903 => x"71195656",
  3904 => x"598a5274",
  3905 => x"5183aa3f",
  3906 => x"b008b005",
  3907 => x"53727434",
  3908 => x"8117578a",
  3909 => x"52745182",
  3910 => x"f33fb008",
  3911 => x"55b008fe",
  3912 => x"cf38feef",
  3913 => x"39fd3d0d",
  3914 => x"81cd8008",
  3915 => x"76b2e429",
  3916 => x"94120c54",
  3917 => x"850b9815",
  3918 => x"0c981408",
  3919 => x"70810651",
  3920 => x"5372f638",
  3921 => x"853d0d04",
  3922 => x"803d0d81",
  3923 => x"cd800851",
  3924 => x"870b8412",
  3925 => x"0cff0ba4",
  3926 => x"120ca70b",
  3927 => x"a8120cb2",
  3928 => x"e40b9412",
  3929 => x"0c870b98",
  3930 => x"120c823d",
  3931 => x"0d04803d",
  3932 => x"0d81cd84",
  3933 => x"0851b80b",
  3934 => x"8c120c83",
  3935 => x"0b88120c",
  3936 => x"823d0d04",
  3937 => x"803d0d81",
  3938 => x"cd840884",
  3939 => x"11088106",
  3940 => x"b00c5182",
  3941 => x"3d0d04ff",
  3942 => x"3d0d81cd",
  3943 => x"84085284",
  3944 => x"12087081",
  3945 => x"06515170",
  3946 => x"802ef438",
  3947 => x"71087081",
  3948 => x"ff06b00c",
  3949 => x"51833d0d",
  3950 => x"04fe3d0d",
  3951 => x"02930533",
  3952 => x"53728a2e",
  3953 => x"9c3881cd",
  3954 => x"84085284",
  3955 => x"12087089",
  3956 => x"2a708106",
  3957 => x"51515170",
  3958 => x"f2387272",
  3959 => x"0c843d0d",
  3960 => x"0481cd84",
  3961 => x"08528412",
  3962 => x"0870892a",
  3963 => x"70810651",
  3964 => x"515170f2",
  3965 => x"388d720c",
  3966 => x"84120870",
  3967 => x"892a7081",
  3968 => x"06515151",
  3969 => x"70c538d2",
  3970 => x"39fa3d0d",
  3971 => x"02a30533",
  3972 => x"81ccf808",
  3973 => x"81f0e033",
  3974 => x"7081ff06",
  3975 => x"70101011",
  3976 => x"81f0e433",
  3977 => x"7081ff06",
  3978 => x"72902911",
  3979 => x"70882b78",
  3980 => x"07770c53",
  3981 => x"5b5b5555",
  3982 => x"59545473",
  3983 => x"8a2e9838",
  3984 => x"7480cf2e",
  3985 => x"9238738c",
  3986 => x"2ea43881",
  3987 => x"16537281",
  3988 => x"f0e43488",
  3989 => x"3d0d0471",
  3990 => x"a326a338",
  3991 => x"81175271",
  3992 => x"81f0e034",
  3993 => x"800b81f0",
  3994 => x"e434883d",
  3995 => x"0d048052",
  3996 => x"71882b73",
  3997 => x"0c811252",
  3998 => x"97907226",
  3999 => x"f338800b",
  4000 => x"81f0e034",
  4001 => x"800b81f0",
  4002 => x"e434df39",
  4003 => x"bc0802bc",
  4004 => x"0cfd3d0d",
  4005 => x"8053bc08",
  4006 => x"8c050852",
  4007 => x"bc088805",
  4008 => x"0851f7c6",
  4009 => x"3fb00870",
  4010 => x"b00c5485",
  4011 => x"3d0dbc0c",
  4012 => x"04bc0802",
  4013 => x"bc0cfd3d",
  4014 => x"0d8153bc",
  4015 => x"088c0508",
  4016 => x"52bc0888",
  4017 => x"050851f7",
  4018 => x"a13fb008",
  4019 => x"70b00c54",
  4020 => x"853d0dbc",
  4021 => x"0c04803d",
  4022 => x"0d865184",
  4023 => x"963f8151",
  4024 => x"a1d33ffc",
  4025 => x"3d0d7670",
  4026 => x"797b5555",
  4027 => x"55558f72",
  4028 => x"278c3872",
  4029 => x"75078306",
  4030 => x"5170802e",
  4031 => x"a738ff12",
  4032 => x"5271ff2e",
  4033 => x"98387270",
  4034 => x"81055433",
  4035 => x"74708105",
  4036 => x"5634ff12",
  4037 => x"5271ff2e",
  4038 => x"098106ea",
  4039 => x"3874b00c",
  4040 => x"863d0d04",
  4041 => x"74517270",
  4042 => x"84055408",
  4043 => x"71708405",
  4044 => x"530c7270",
  4045 => x"84055408",
  4046 => x"71708405",
  4047 => x"530c7270",
  4048 => x"84055408",
  4049 => x"71708405",
  4050 => x"530c7270",
  4051 => x"84055408",
  4052 => x"71708405",
  4053 => x"530cf012",
  4054 => x"52718f26",
  4055 => x"c9388372",
  4056 => x"27953872",
  4057 => x"70840554",
  4058 => x"08717084",
  4059 => x"05530cfc",
  4060 => x"12527183",
  4061 => x"26ed3870",
  4062 => x"54ff8339",
  4063 => x"fd3d0d75",
  4064 => x"5384d813",
  4065 => x"08802e8a",
  4066 => x"38805372",
  4067 => x"b00c853d",
  4068 => x"0d048180",
  4069 => x"5272518d",
  4070 => x"9b3fb008",
  4071 => x"84d8140c",
  4072 => x"ff53b008",
  4073 => x"802ee438",
  4074 => x"b008549f",
  4075 => x"53807470",
  4076 => x"8405560c",
  4077 => x"ff135380",
  4078 => x"7324ce38",
  4079 => x"80747084",
  4080 => x"05560cff",
  4081 => x"13537280",
  4082 => x"25e338ff",
  4083 => x"bc39fd3d",
  4084 => x"0d757755",
  4085 => x"539f7427",
  4086 => x"8d389673",
  4087 => x"0cff5271",
  4088 => x"b00c853d",
  4089 => x"0d0484d8",
  4090 => x"13085271",
  4091 => x"802e9338",
  4092 => x"73101012",
  4093 => x"70087972",
  4094 => x"0c515271",
  4095 => x"b00c853d",
  4096 => x"0d047251",
  4097 => x"fef63fff",
  4098 => x"52b008d3",
  4099 => x"3884d813",
  4100 => x"08741010",
  4101 => x"1170087a",
  4102 => x"720c5151",
  4103 => x"52dd39f9",
  4104 => x"3d0d797b",
  4105 => x"5856769f",
  4106 => x"2680e838",
  4107 => x"84d81608",
  4108 => x"5473802e",
  4109 => x"aa387610",
  4110 => x"10147008",
  4111 => x"55557380",
  4112 => x"2eba3880",
  4113 => x"5873812e",
  4114 => x"8f3873ff",
  4115 => x"2ea33880",
  4116 => x"750c7651",
  4117 => x"732d8058",
  4118 => x"77b00c89",
  4119 => x"3d0d0475",
  4120 => x"51fe993f",
  4121 => x"ff58b008",
  4122 => x"ef3884d8",
  4123 => x"160854c6",
  4124 => x"3996760c",
  4125 => x"810bb00c",
  4126 => x"893d0d04",
  4127 => x"755181ed",
  4128 => x"3f7653b0",
  4129 => x"08527551",
  4130 => x"81ad3fb0",
  4131 => x"08b00c89",
  4132 => x"3d0d0496",
  4133 => x"760cff0b",
  4134 => x"b00c893d",
  4135 => x"0d04fc3d",
  4136 => x"0d767856",
  4137 => x"53ff5474",
  4138 => x"9f26b138",
  4139 => x"84d81308",
  4140 => x"5271802e",
  4141 => x"ae387410",
  4142 => x"10127008",
  4143 => x"53538154",
  4144 => x"71802e98",
  4145 => x"38825471",
  4146 => x"ff2e9138",
  4147 => x"83547181",
  4148 => x"2e8a3880",
  4149 => x"730c7451",
  4150 => x"712d8054",
  4151 => x"73b00c86",
  4152 => x"3d0d0472",
  4153 => x"51fd953f",
  4154 => x"b008f138",
  4155 => x"84d81308",
  4156 => x"52c439ff",
  4157 => x"3d0d7352",
  4158 => x"81cd9008",
  4159 => x"51fea03f",
  4160 => x"833d0d04",
  4161 => x"fe3d0d75",
  4162 => x"53745281",
  4163 => x"cd900851",
  4164 => x"fdbc3f84",
  4165 => x"3d0d0480",
  4166 => x"3d0d81cd",
  4167 => x"900851fc",
  4168 => x"db3f823d",
  4169 => x"0d04ff3d",
  4170 => x"0d735281",
  4171 => x"cd900851",
  4172 => x"feec3f83",
  4173 => x"3d0d04fc",
  4174 => x"3d0d800b",
  4175 => x"81f0ec0c",
  4176 => x"78527751",
  4177 => x"9caa3fb0",
  4178 => x"0854b008",
  4179 => x"ff2e8838",
  4180 => x"73b00c86",
  4181 => x"3d0d0481",
  4182 => x"f0ec0855",
  4183 => x"74802ef0",
  4184 => x"38767571",
  4185 => x"0c5373b0",
  4186 => x"0c863d0d",
  4187 => x"049bfc3f",
  4188 => x"04fc3d0d",
  4189 => x"76707970",
  4190 => x"73078306",
  4191 => x"54545455",
  4192 => x"7080c338",
  4193 => x"71700870",
  4194 => x"0970f7fb",
  4195 => x"fdff1306",
  4196 => x"70f88482",
  4197 => x"81800651",
  4198 => x"51535354",
  4199 => x"70a63884",
  4200 => x"14727470",
  4201 => x"8405560c",
  4202 => x"70087009",
  4203 => x"70f7fbfd",
  4204 => x"ff130670",
  4205 => x"f8848281",
  4206 => x"80065151",
  4207 => x"53535470",
  4208 => x"802edc38",
  4209 => x"73527170",
  4210 => x"81055333",
  4211 => x"51707370",
  4212 => x"81055534",
  4213 => x"70f03874",
  4214 => x"b00c863d",
  4215 => x"0d04fd3d",
  4216 => x"0d757071",
  4217 => x"83065355",
  4218 => x"5270b838",
  4219 => x"71700870",
  4220 => x"09f7fbfd",
  4221 => x"ff120670",
  4222 => x"f8848281",
  4223 => x"80065151",
  4224 => x"5253709d",
  4225 => x"38841370",
  4226 => x"087009f7",
  4227 => x"fbfdff12",
  4228 => x"0670f884",
  4229 => x"82818006",
  4230 => x"51515253",
  4231 => x"70802ee5",
  4232 => x"38725271",
  4233 => x"33517080",
  4234 => x"2e8a3881",
  4235 => x"12703352",
  4236 => x"5270f838",
  4237 => x"717431b0",
  4238 => x"0c853d0d",
  4239 => x"04fa3d0d",
  4240 => x"787a7c70",
  4241 => x"54555552",
  4242 => x"72802e80",
  4243 => x"d9387174",
  4244 => x"07830651",
  4245 => x"70802e80",
  4246 => x"d438ff13",
  4247 => x"5372ff2e",
  4248 => x"b1387133",
  4249 => x"74335651",
  4250 => x"74712e09",
  4251 => x"8106a938",
  4252 => x"72802e81",
  4253 => x"87387081",
  4254 => x"ff065170",
  4255 => x"802e80fc",
  4256 => x"38811281",
  4257 => x"15ff1555",
  4258 => x"555272ff",
  4259 => x"2e098106",
  4260 => x"d1387133",
  4261 => x"74335651",
  4262 => x"7081ff06",
  4263 => x"7581ff06",
  4264 => x"71713151",
  4265 => x"525270b0",
  4266 => x"0c883d0d",
  4267 => x"04717457",
  4268 => x"55837327",
  4269 => x"88387108",
  4270 => x"74082e88",
  4271 => x"38747655",
  4272 => x"52ff9739",
  4273 => x"fc135372",
  4274 => x"802eb138",
  4275 => x"74087009",
  4276 => x"f7fbfdff",
  4277 => x"120670f8",
  4278 => x"84828180",
  4279 => x"06515151",
  4280 => x"709a3884",
  4281 => x"15841757",
  4282 => x"55837327",
  4283 => x"d0387408",
  4284 => x"76082ed0",
  4285 => x"38747655",
  4286 => x"52fedf39",
  4287 => x"800bb00c",
  4288 => x"883d0d04",
  4289 => x"f33d0d60",
  4290 => x"6264725a",
  4291 => x"5a5e5e80",
  4292 => x"5c767081",
  4293 => x"05583381",
  4294 => x"cab11133",
  4295 => x"70832a70",
  4296 => x"81065155",
  4297 => x"555672e9",
  4298 => x"3875ad2e",
  4299 => x"82883875",
  4300 => x"ab2e8284",
  4301 => x"38773070",
  4302 => x"79078025",
  4303 => x"79903270",
  4304 => x"30707207",
  4305 => x"80257307",
  4306 => x"53575751",
  4307 => x"5372802e",
  4308 => x"873875b0",
  4309 => x"2e81eb38",
  4310 => x"778a3888",
  4311 => x"5875b02e",
  4312 => x"83388a58",
  4313 => x"810a5a7b",
  4314 => x"8438fe0a",
  4315 => x"5a775279",
  4316 => x"51f6be3f",
  4317 => x"b0087853",
  4318 => x"7a525bf6",
  4319 => x"8f3fb008",
  4320 => x"5a807081",
  4321 => x"cab11833",
  4322 => x"70822a70",
  4323 => x"81065156",
  4324 => x"565a5572",
  4325 => x"802e80c1",
  4326 => x"38d01656",
  4327 => x"75782580",
  4328 => x"d7388079",
  4329 => x"24757b26",
  4330 => x"07537293",
  4331 => x"38747a2e",
  4332 => x"80eb387a",
  4333 => x"762580ed",
  4334 => x"3872802e",
  4335 => x"80e738ff",
  4336 => x"77708105",
  4337 => x"59335759",
  4338 => x"81cab116",
  4339 => x"3370822a",
  4340 => x"70810651",
  4341 => x"545472c1",
  4342 => x"38738306",
  4343 => x"5372802e",
  4344 => x"97387381",
  4345 => x"06c91755",
  4346 => x"53728538",
  4347 => x"ffa91654",
  4348 => x"73567776",
  4349 => x"24ffab38",
  4350 => x"80792480",
  4351 => x"f0387b80",
  4352 => x"2e843874",
  4353 => x"30557c80",
  4354 => x"2e8c38ff",
  4355 => x"17537883",
  4356 => x"387d5372",
  4357 => x"7d0c74b0",
  4358 => x"0c8f3d0d",
  4359 => x"04815375",
  4360 => x"7b24ff95",
  4361 => x"38817579",
  4362 => x"29177870",
  4363 => x"81055a33",
  4364 => x"585659ff",
  4365 => x"9339815c",
  4366 => x"76708105",
  4367 => x"583356fd",
  4368 => x"f4398077",
  4369 => x"33545472",
  4370 => x"80f82eb2",
  4371 => x"387280d8",
  4372 => x"32703070",
  4373 => x"80257607",
  4374 => x"51515372",
  4375 => x"802efdf8",
  4376 => x"38811733",
  4377 => x"82185856",
  4378 => x"9058fdf8",
  4379 => x"39810a55",
  4380 => x"7b8438fe",
  4381 => x"0a557f53",
  4382 => x"a2730cff",
  4383 => x"89398154",
  4384 => x"cc39fd3d",
  4385 => x"0d775476",
  4386 => x"53755281",
  4387 => x"cd900851",
  4388 => x"fcf23f85",
  4389 => x"3d0d04f3",
  4390 => x"3d0d6062",
  4391 => x"64725a5a",
  4392 => x"5d5d805e",
  4393 => x"76708105",
  4394 => x"583381ca",
  4395 => x"b1113370",
  4396 => x"832a7081",
  4397 => x"06515555",
  4398 => x"5672e938",
  4399 => x"75ad2e81",
  4400 => x"ff3875ab",
  4401 => x"2e81fb38",
  4402 => x"77307079",
  4403 => x"07802579",
  4404 => x"90327030",
  4405 => x"70720780",
  4406 => x"25730753",
  4407 => x"57575153",
  4408 => x"72802e87",
  4409 => x"3875b02e",
  4410 => x"81e23877",
  4411 => x"8a388858",
  4412 => x"75b02e83",
  4413 => x"388a5877",
  4414 => x"52ff51f3",
  4415 => x"8f3fb008",
  4416 => x"78535aff",
  4417 => x"51f3aa3f",
  4418 => x"b0085b80",
  4419 => x"705a5581",
  4420 => x"cab11633",
  4421 => x"70822a70",
  4422 => x"81065154",
  4423 => x"5472802e",
  4424 => x"80c138d0",
  4425 => x"16567578",
  4426 => x"2580d738",
  4427 => x"80792475",
  4428 => x"7b260753",
  4429 => x"72933874",
  4430 => x"7a2e80eb",
  4431 => x"387a7625",
  4432 => x"80ed3872",
  4433 => x"802e80e7",
  4434 => x"38ff7770",
  4435 => x"81055933",
  4436 => x"575981ca",
  4437 => x"b1163370",
  4438 => x"822a7081",
  4439 => x"06515454",
  4440 => x"72c13873",
  4441 => x"83065372",
  4442 => x"802e9738",
  4443 => x"738106c9",
  4444 => x"17555372",
  4445 => x"8538ffa9",
  4446 => x"16547356",
  4447 => x"777624ff",
  4448 => x"ab388079",
  4449 => x"24818938",
  4450 => x"7d802e84",
  4451 => x"38743055",
  4452 => x"7b802e8c",
  4453 => x"38ff1753",
  4454 => x"7883387c",
  4455 => x"53727c0c",
  4456 => x"74b00c8f",
  4457 => x"3d0d0481",
  4458 => x"53757b24",
  4459 => x"ff953881",
  4460 => x"75792917",
  4461 => x"78708105",
  4462 => x"5a335856",
  4463 => x"59ff9339",
  4464 => x"815e7670",
  4465 => x"81055833",
  4466 => x"56fdfd39",
  4467 => x"80773354",
  4468 => x"547280f8",
  4469 => x"2e80c338",
  4470 => x"7280d832",
  4471 => x"70307080",
  4472 => x"25760751",
  4473 => x"51537280",
  4474 => x"2efe8038",
  4475 => x"81173382",
  4476 => x"18585690",
  4477 => x"705358ff",
  4478 => x"51f1913f",
  4479 => x"b0087853",
  4480 => x"5aff51f1",
  4481 => x"ac3fb008",
  4482 => x"5b80705a",
  4483 => x"55fe8039",
  4484 => x"ff605455",
  4485 => x"a2730cfe",
  4486 => x"f7398154",
  4487 => x"ffba39fd",
  4488 => x"3d0d7754",
  4489 => x"76537552",
  4490 => x"81cd9008",
  4491 => x"51fce83f",
  4492 => x"853d0d04",
  4493 => x"f33d0d7f",
  4494 => x"618b1170",
  4495 => x"f8065c55",
  4496 => x"555e7296",
  4497 => x"26833890",
  4498 => x"59807924",
  4499 => x"747a2607",
  4500 => x"53805472",
  4501 => x"742e0981",
  4502 => x"0680cb38",
  4503 => x"7d518bca",
  4504 => x"3f7883f7",
  4505 => x"2680c638",
  4506 => x"78832a70",
  4507 => x"10101081",
  4508 => x"d4cc058c",
  4509 => x"11085959",
  4510 => x"5a76782e",
  4511 => x"83b03884",
  4512 => x"1708fc06",
  4513 => x"568c1708",
  4514 => x"88180871",
  4515 => x"8c120c88",
  4516 => x"120c5875",
  4517 => x"17841108",
  4518 => x"81078412",
  4519 => x"0c537d51",
  4520 => x"8b893f88",
  4521 => x"175473b0",
  4522 => x"0c8f3d0d",
  4523 => x"0478892a",
  4524 => x"79832a5b",
  4525 => x"5372802e",
  4526 => x"bf387886",
  4527 => x"2ab8055a",
  4528 => x"847327b4",
  4529 => x"3880db13",
  4530 => x"5a947327",
  4531 => x"ab38788c",
  4532 => x"2a80ee05",
  4533 => x"5a80d473",
  4534 => x"279e3878",
  4535 => x"8f2a80f7",
  4536 => x"055a82d4",
  4537 => x"73279138",
  4538 => x"78922a80",
  4539 => x"fc055a8a",
  4540 => x"d4732784",
  4541 => x"3880fe5a",
  4542 => x"79101010",
  4543 => x"81d4cc05",
  4544 => x"8c110858",
  4545 => x"5576752e",
  4546 => x"a3388417",
  4547 => x"08fc0670",
  4548 => x"7a315556",
  4549 => x"738f2488",
  4550 => x"d5387380",
  4551 => x"25fee638",
  4552 => x"8c170857",
  4553 => x"76752e09",
  4554 => x"8106df38",
  4555 => x"811a5a81",
  4556 => x"d4dc0857",
  4557 => x"7681d4d4",
  4558 => x"2e82c038",
  4559 => x"841708fc",
  4560 => x"06707a31",
  4561 => x"5556738f",
  4562 => x"2481f938",
  4563 => x"81d4d40b",
  4564 => x"81d4e00c",
  4565 => x"81d4d40b",
  4566 => x"81d4dc0c",
  4567 => x"738025fe",
  4568 => x"b23883ff",
  4569 => x"762783df",
  4570 => x"3875892a",
  4571 => x"76832a55",
  4572 => x"5372802e",
  4573 => x"bf387586",
  4574 => x"2ab80554",
  4575 => x"847327b4",
  4576 => x"3880db13",
  4577 => x"54947327",
  4578 => x"ab38758c",
  4579 => x"2a80ee05",
  4580 => x"5480d473",
  4581 => x"279e3875",
  4582 => x"8f2a80f7",
  4583 => x"055482d4",
  4584 => x"73279138",
  4585 => x"75922a80",
  4586 => x"fc05548a",
  4587 => x"d4732784",
  4588 => x"3880fe54",
  4589 => x"73101010",
  4590 => x"81d4cc05",
  4591 => x"88110856",
  4592 => x"5874782e",
  4593 => x"86cf3884",
  4594 => x"1508fc06",
  4595 => x"53757327",
  4596 => x"8d388815",
  4597 => x"08557478",
  4598 => x"2e098106",
  4599 => x"ea388c15",
  4600 => x"0881d4cc",
  4601 => x"0b840508",
  4602 => x"718c1a0c",
  4603 => x"76881a0c",
  4604 => x"7888130c",
  4605 => x"788c180c",
  4606 => x"5d587953",
  4607 => x"807a2483",
  4608 => x"e6387282",
  4609 => x"2c81712b",
  4610 => x"5c537a7c",
  4611 => x"26819838",
  4612 => x"7b7b0653",
  4613 => x"7282f138",
  4614 => x"79fc0684",
  4615 => x"055a7a10",
  4616 => x"707d0654",
  4617 => x"5b7282e0",
  4618 => x"38841a5a",
  4619 => x"f1398817",
  4620 => x"8c110858",
  4621 => x"5876782e",
  4622 => x"098106fc",
  4623 => x"c238821a",
  4624 => x"5afdec39",
  4625 => x"78177981",
  4626 => x"0784190c",
  4627 => x"7081d4e0",
  4628 => x"0c7081d4",
  4629 => x"dc0c81d4",
  4630 => x"d40b8c12",
  4631 => x"0c8c1108",
  4632 => x"88120c74",
  4633 => x"81078412",
  4634 => x"0c741175",
  4635 => x"710c5153",
  4636 => x"7d5187b7",
  4637 => x"3f881754",
  4638 => x"fcac3981",
  4639 => x"d4cc0b84",
  4640 => x"05087a54",
  4641 => x"5c798025",
  4642 => x"fef83882",
  4643 => x"da397a09",
  4644 => x"7c067081",
  4645 => x"d4cc0b84",
  4646 => x"050c5c7a",
  4647 => x"105b7a7c",
  4648 => x"2685387a",
  4649 => x"85b83881",
  4650 => x"d4cc0b88",
  4651 => x"05087084",
  4652 => x"1208fc06",
  4653 => x"707c317c",
  4654 => x"72268f72",
  4655 => x"25075757",
  4656 => x"5c5d5572",
  4657 => x"802e80db",
  4658 => x"38797a16",
  4659 => x"81d4c408",
  4660 => x"1b90115a",
  4661 => x"55575b81",
  4662 => x"d4c008ff",
  4663 => x"2e8838a0",
  4664 => x"8f13e080",
  4665 => x"06577652",
  4666 => x"7d5186c0",
  4667 => x"3fb00854",
  4668 => x"b008ff2e",
  4669 => x"9038b008",
  4670 => x"76278299",
  4671 => x"387481d4",
  4672 => x"cc2e8291",
  4673 => x"3881d4cc",
  4674 => x"0b880508",
  4675 => x"55841508",
  4676 => x"fc06707a",
  4677 => x"317a7226",
  4678 => x"8f722507",
  4679 => x"52555372",
  4680 => x"83e63874",
  4681 => x"79810784",
  4682 => x"170c7916",
  4683 => x"7081d4cc",
  4684 => x"0b88050c",
  4685 => x"75810784",
  4686 => x"120c547e",
  4687 => x"525785eb",
  4688 => x"3f881754",
  4689 => x"fae03975",
  4690 => x"832a7054",
  4691 => x"54807424",
  4692 => x"819b3872",
  4693 => x"822c8171",
  4694 => x"2b81d4d0",
  4695 => x"08077081",
  4696 => x"d4cc0b84",
  4697 => x"050c7510",
  4698 => x"101081d4",
  4699 => x"cc058811",
  4700 => x"08585a5d",
  4701 => x"53778c18",
  4702 => x"0c748818",
  4703 => x"0c768819",
  4704 => x"0c768c16",
  4705 => x"0cfcf339",
  4706 => x"797a1010",
  4707 => x"1081d4cc",
  4708 => x"05705759",
  4709 => x"5d8c1508",
  4710 => x"5776752e",
  4711 => x"a3388417",
  4712 => x"08fc0670",
  4713 => x"7a315556",
  4714 => x"738f2483",
  4715 => x"ca387380",
  4716 => x"25848138",
  4717 => x"8c170857",
  4718 => x"76752e09",
  4719 => x"8106df38",
  4720 => x"8815811b",
  4721 => x"70830655",
  4722 => x"5b5572c9",
  4723 => x"387c8306",
  4724 => x"5372802e",
  4725 => x"fdb838ff",
  4726 => x"1df81959",
  4727 => x"5d881808",
  4728 => x"782eea38",
  4729 => x"fdb53983",
  4730 => x"1a53fc96",
  4731 => x"39831470",
  4732 => x"822c8171",
  4733 => x"2b81d4d0",
  4734 => x"08077081",
  4735 => x"d4cc0b84",
  4736 => x"050c7610",
  4737 => x"101081d4",
  4738 => x"cc058811",
  4739 => x"08595b5e",
  4740 => x"5153fee1",
  4741 => x"3981d490",
  4742 => x"081758b0",
  4743 => x"08762e81",
  4744 => x"8d3881d4",
  4745 => x"c008ff2e",
  4746 => x"83ec3873",
  4747 => x"76311881",
  4748 => x"d4900c73",
  4749 => x"87067057",
  4750 => x"5372802e",
  4751 => x"88388873",
  4752 => x"31701555",
  4753 => x"5676149f",
  4754 => x"ff06a080",
  4755 => x"71311770",
  4756 => x"547f5357",
  4757 => x"5383d53f",
  4758 => x"b00853b0",
  4759 => x"08ff2e81",
  4760 => x"a03881d4",
  4761 => x"90081670",
  4762 => x"81d4900c",
  4763 => x"747581d4",
  4764 => x"cc0b8805",
  4765 => x"0c747631",
  4766 => x"18708107",
  4767 => x"51555658",
  4768 => x"7b81d4cc",
  4769 => x"2e839c38",
  4770 => x"798f2682",
  4771 => x"cb38810b",
  4772 => x"84150c84",
  4773 => x"1508fc06",
  4774 => x"707a317a",
  4775 => x"72268f72",
  4776 => x"25075255",
  4777 => x"5372802e",
  4778 => x"fcf93880",
  4779 => x"db39b008",
  4780 => x"9fff0653",
  4781 => x"72feeb38",
  4782 => x"7781d490",
  4783 => x"0c81d4cc",
  4784 => x"0b880508",
  4785 => x"7b188107",
  4786 => x"84120c55",
  4787 => x"81d4bc08",
  4788 => x"78278638",
  4789 => x"7781d4bc",
  4790 => x"0c81d4b8",
  4791 => x"087827fc",
  4792 => x"ac387781",
  4793 => x"d4b80c84",
  4794 => x"1508fc06",
  4795 => x"707a317a",
  4796 => x"72268f72",
  4797 => x"25075255",
  4798 => x"5372802e",
  4799 => x"fca53888",
  4800 => x"39807454",
  4801 => x"56fedb39",
  4802 => x"7d51829f",
  4803 => x"3f800bb0",
  4804 => x"0c8f3d0d",
  4805 => x"04735380",
  4806 => x"7424a938",
  4807 => x"72822c81",
  4808 => x"712b81d4",
  4809 => x"d0080770",
  4810 => x"81d4cc0b",
  4811 => x"84050c5d",
  4812 => x"53778c18",
  4813 => x"0c748818",
  4814 => x"0c768819",
  4815 => x"0c768c16",
  4816 => x"0cf9b739",
  4817 => x"83147082",
  4818 => x"2c81712b",
  4819 => x"81d4d008",
  4820 => x"077081d4",
  4821 => x"cc0b8405",
  4822 => x"0c5e5153",
  4823 => x"d4397b7b",
  4824 => x"065372fc",
  4825 => x"a338841a",
  4826 => x"7b105c5a",
  4827 => x"f139ff1a",
  4828 => x"8111515a",
  4829 => x"f7b93978",
  4830 => x"17798107",
  4831 => x"84190c8c",
  4832 => x"18088819",
  4833 => x"08718c12",
  4834 => x"0c88120c",
  4835 => x"597081d4",
  4836 => x"e00c7081",
  4837 => x"d4dc0c81",
  4838 => x"d4d40b8c",
  4839 => x"120c8c11",
  4840 => x"0888120c",
  4841 => x"74810784",
  4842 => x"120c7411",
  4843 => x"75710c51",
  4844 => x"53f9bd39",
  4845 => x"75178411",
  4846 => x"08810784",
  4847 => x"120c538c",
  4848 => x"17088818",
  4849 => x"08718c12",
  4850 => x"0c88120c",
  4851 => x"587d5180",
  4852 => x"da3f8817",
  4853 => x"54f5cf39",
  4854 => x"7284150c",
  4855 => x"f41af806",
  4856 => x"70841e08",
  4857 => x"81060784",
  4858 => x"1e0c701d",
  4859 => x"545b850b",
  4860 => x"84140c85",
  4861 => x"0b88140c",
  4862 => x"8f7b27fd",
  4863 => x"cf38881c",
  4864 => x"527d5182",
  4865 => x"903f81d4",
  4866 => x"cc0b8805",
  4867 => x"0881d490",
  4868 => x"085955fd",
  4869 => x"b7397781",
  4870 => x"d4900c73",
  4871 => x"81d4c00c",
  4872 => x"fc913972",
  4873 => x"84150cfd",
  4874 => x"a3390404",
  4875 => x"fd3d0d80",
  4876 => x"0b81f0ec",
  4877 => x"0c765186",
  4878 => x"cb3fb008",
  4879 => x"53b008ff",
  4880 => x"2e883872",
  4881 => x"b00c853d",
  4882 => x"0d0481f0",
  4883 => x"ec085473",
  4884 => x"802ef038",
  4885 => x"7574710c",
  4886 => x"5272b00c",
  4887 => x"853d0d04",
  4888 => x"fb3d0d77",
  4889 => x"705256c2",
  4890 => x"3f81d4cc",
  4891 => x"0b880508",
  4892 => x"841108fc",
  4893 => x"06707b31",
  4894 => x"9fef05e0",
  4895 => x"8006e080",
  4896 => x"05565653",
  4897 => x"a0807424",
  4898 => x"94388052",
  4899 => x"7551ff9c",
  4900 => x"3f81d4d4",
  4901 => x"08155372",
  4902 => x"b0082e8f",
  4903 => x"387551ff",
  4904 => x"8a3f8053",
  4905 => x"72b00c87",
  4906 => x"3d0d0473",
  4907 => x"30527551",
  4908 => x"fefa3fb0",
  4909 => x"08ff2ea8",
  4910 => x"3881d4cc",
  4911 => x"0b880508",
  4912 => x"75753181",
  4913 => x"0784120c",
  4914 => x"5381d490",
  4915 => x"08743181",
  4916 => x"d4900c75",
  4917 => x"51fed43f",
  4918 => x"810bb00c",
  4919 => x"873d0d04",
  4920 => x"80527551",
  4921 => x"fec63f81",
  4922 => x"d4cc0b88",
  4923 => x"0508b008",
  4924 => x"71315653",
  4925 => x"8f7525ff",
  4926 => x"a438b008",
  4927 => x"81d4c008",
  4928 => x"3181d490",
  4929 => x"0c748107",
  4930 => x"84140c75",
  4931 => x"51fe9c3f",
  4932 => x"8053ff90",
  4933 => x"39f63d0d",
  4934 => x"7c7e545b",
  4935 => x"72802e82",
  4936 => x"83387a51",
  4937 => x"fe843ff8",
  4938 => x"13841108",
  4939 => x"70fe0670",
  4940 => x"13841108",
  4941 => x"fc065d58",
  4942 => x"59545881",
  4943 => x"d4d40875",
  4944 => x"2e82de38",
  4945 => x"7884160c",
  4946 => x"80738106",
  4947 => x"545a727a",
  4948 => x"2e81d538",
  4949 => x"78158411",
  4950 => x"08810651",
  4951 => x"5372a038",
  4952 => x"78175779",
  4953 => x"81e63888",
  4954 => x"15085372",
  4955 => x"81d4d42e",
  4956 => x"82f9388c",
  4957 => x"1508708c",
  4958 => x"150c7388",
  4959 => x"120c5676",
  4960 => x"81078419",
  4961 => x"0c761877",
  4962 => x"710c5379",
  4963 => x"81913883",
  4964 => x"ff772781",
  4965 => x"c8387689",
  4966 => x"2a77832a",
  4967 => x"56537280",
  4968 => x"2ebf3876",
  4969 => x"862ab805",
  4970 => x"55847327",
  4971 => x"b43880db",
  4972 => x"13559473",
  4973 => x"27ab3876",
  4974 => x"8c2a80ee",
  4975 => x"055580d4",
  4976 => x"73279e38",
  4977 => x"768f2a80",
  4978 => x"f7055582",
  4979 => x"d4732791",
  4980 => x"3876922a",
  4981 => x"80fc0555",
  4982 => x"8ad47327",
  4983 => x"843880fe",
  4984 => x"55741010",
  4985 => x"1081d4cc",
  4986 => x"05881108",
  4987 => x"55567376",
  4988 => x"2e82b338",
  4989 => x"841408fc",
  4990 => x"06537673",
  4991 => x"278d3888",
  4992 => x"14085473",
  4993 => x"762e0981",
  4994 => x"06ea388c",
  4995 => x"1408708c",
  4996 => x"1a0c7488",
  4997 => x"1a0c7888",
  4998 => x"120c5677",
  4999 => x"8c150c7a",
  5000 => x"51fc883f",
  5001 => x"8c3d0d04",
  5002 => x"77087871",
  5003 => x"31597705",
  5004 => x"88190854",
  5005 => x"577281d4",
  5006 => x"d42e80e0",
  5007 => x"388c1808",
  5008 => x"708c150c",
  5009 => x"7388120c",
  5010 => x"56fe8939",
  5011 => x"8815088c",
  5012 => x"1608708c",
  5013 => x"130c5788",
  5014 => x"170cfea3",
  5015 => x"3976832a",
  5016 => x"70545580",
  5017 => x"75248198",
  5018 => x"3872822c",
  5019 => x"81712b81",
  5020 => x"d4d00807",
  5021 => x"81d4cc0b",
  5022 => x"84050c53",
  5023 => x"74101010",
  5024 => x"81d4cc05",
  5025 => x"88110855",
  5026 => x"56758c19",
  5027 => x"0c738819",
  5028 => x"0c778817",
  5029 => x"0c778c15",
  5030 => x"0cff8439",
  5031 => x"815afdb4",
  5032 => x"39781773",
  5033 => x"81065457",
  5034 => x"72983877",
  5035 => x"08787131",
  5036 => x"5977058c",
  5037 => x"1908881a",
  5038 => x"08718c12",
  5039 => x"0c88120c",
  5040 => x"57577681",
  5041 => x"0784190c",
  5042 => x"7781d4cc",
  5043 => x"0b88050c",
  5044 => x"81d4c808",
  5045 => x"7726fec7",
  5046 => x"3881d4c4",
  5047 => x"08527a51",
  5048 => x"fafe3f7a",
  5049 => x"51fac43f",
  5050 => x"feba3981",
  5051 => x"788c150c",
  5052 => x"7888150c",
  5053 => x"738c1a0c",
  5054 => x"73881a0c",
  5055 => x"5afd8039",
  5056 => x"83157082",
  5057 => x"2c81712b",
  5058 => x"81d4d008",
  5059 => x"0781d4cc",
  5060 => x"0b84050c",
  5061 => x"51537410",
  5062 => x"101081d4",
  5063 => x"cc058811",
  5064 => x"085556fe",
  5065 => x"e4397453",
  5066 => x"807524a7",
  5067 => x"3872822c",
  5068 => x"81712b81",
  5069 => x"d4d00807",
  5070 => x"81d4cc0b",
  5071 => x"84050c53",
  5072 => x"758c190c",
  5073 => x"7388190c",
  5074 => x"7788170c",
  5075 => x"778c150c",
  5076 => x"fdcd3983",
  5077 => x"1570822c",
  5078 => x"81712b81",
  5079 => x"d4d00807",
  5080 => x"81d4cc0b",
  5081 => x"84050c51",
  5082 => x"53d63981",
  5083 => x"0bb00c04",
  5084 => x"803d0d72",
  5085 => x"812e8938",
  5086 => x"800bb00c",
  5087 => x"823d0d04",
  5088 => x"7351b23f",
  5089 => x"fe3d0d81",
  5090 => x"f0e80851",
  5091 => x"708a3881",
  5092 => x"f0f07081",
  5093 => x"f0e80c51",
  5094 => x"70751252",
  5095 => x"52ff5370",
  5096 => x"87fb8080",
  5097 => x"26883870",
  5098 => x"81f0e80c",
  5099 => x"715372b0",
  5100 => x"0c843d0d",
  5101 => x"0400ff39",
  5102 => x"00000000",
  5103 => x"00000000",
  5104 => x"00000000",
  5105 => x"00000000",
  5106 => x"00cac5ca",
  5107 => x"c5c0c0c0",
  5108 => x"c0c0c0c0",
  5109 => x"c0c0c0cf",
  5110 => x"cfcfcf00",
  5111 => x"00000f0f",
  5112 => x"0f0f8f8f",
  5113 => x"cfcfcfcf",
  5114 => x"cfcf4f0f",
  5115 => x"0f0f0000",
  5116 => x"cfcfcfcf",
  5117 => x"0f0f0f0f",
  5118 => x"0f0f0f0f",
  5119 => x"0f0ffefe",
  5120 => x"fefc0000",
  5121 => x"cfcfcfcf",
  5122 => x"cfcfcfcf",
  5123 => x"cfcfcfcf",
  5124 => x"cfffff7e",
  5125 => x"7e000000",
  5126 => x"00000000",
  5127 => x"00000000",
  5128 => x"00000000",
  5129 => x"00003f3f",
  5130 => x"3f3f0101",
  5131 => x"01010101",
  5132 => x"01010101",
  5133 => x"3f3f3f3f",
  5134 => x"0000383c",
  5135 => x"3e3e3f3f",
  5136 => x"3f3b3b39",
  5137 => x"39383838",
  5138 => x"38383800",
  5139 => x"003f3f3f",
  5140 => x"3f383838",
  5141 => x"38383838",
  5142 => x"38383c3f",
  5143 => x"3f1f0f00",
  5144 => x"003f3f3f",
  5145 => x"3f030303",
  5146 => x"03030303",
  5147 => x"03033f3f",
  5148 => x"3f3e0000",
  5149 => x"00000000",
  5150 => x"00000000",
  5151 => x"00000000",
  5152 => x"00000000",
  5153 => x"00000000",
  5154 => x"00000000",
  5155 => x"00000000",
  5156 => x"00000000",
  5157 => x"00000000",
  5158 => x"00000000",
  5159 => x"00000000",
  5160 => x"00000000",
  5161 => x"00000000",
  5162 => x"00000000",
  5163 => x"00000000",
  5164 => x"00000000",
  5165 => x"00000000",
  5166 => x"00000000",
  5167 => x"00000000",
  5168 => x"00000000",
  5169 => x"00000000",
  5170 => x"00000000",
  5171 => x"00000000",
  5172 => x"00000000",
  5173 => x"8080c0c0",
  5174 => x"e0e06000",
  5175 => x"00000000",
  5176 => x"00000000",
  5177 => x"00000000",
  5178 => x"00000000",
  5179 => x"00000000",
  5180 => x"00000000",
  5181 => x"00000000",
  5182 => x"00000000",
  5183 => x"00000000",
  5184 => x"00000000",
  5185 => x"00000000",
  5186 => x"00000000",
  5187 => x"00000000",
  5188 => x"00000000",
  5189 => x"00000000",
  5190 => x"00000000",
  5191 => x"00000000",
  5192 => x"00000000",
  5193 => x"00000000",
  5194 => x"00000000",
  5195 => x"806098ee",
  5196 => x"77bbddec",
  5197 => x"ee6e0200",
  5198 => x"00000000",
  5199 => x"00e08080",
  5200 => x"e00000e0",
  5201 => x"a0a00000",
  5202 => x"e0000000",
  5203 => x"00e0c000",
  5204 => x"c0e00000",
  5205 => x"e08080e0",
  5206 => x"0000c020",
  5207 => x"20c00000",
  5208 => x"e0000000",
  5209 => x"20e02000",
  5210 => x"0020a060",
  5211 => x"20000000",
  5212 => x"00000000",
  5213 => x"00000000",
  5214 => x"00000000",
  5215 => x"00000000",
  5216 => x"00000000",
  5217 => x"00000000",
  5218 => x"00030007",
  5219 => x"00070701",
  5220 => x"00000000",
  5221 => x"00000000",
  5222 => x"00000300",
  5223 => x"c0030000",
  5224 => x"034242c0",
  5225 => x"00c34242",
  5226 => x"0000c380",
  5227 => x"01c00340",
  5228 => x"c04300c0",
  5229 => x"43408001",
  5230 => x"c20201c0",
  5231 => x"00c38202",
  5232 => x"80c00300",
  5233 => x"00c04342",
  5234 => x"8202c040",
  5235 => x"40800000",
  5236 => x"c0404000",
  5237 => x"80404000",
  5238 => x"00c04040",
  5239 => x"8000c040",
  5240 => x"4000c080",
  5241 => x"00c00000",
  5242 => x"00000000",
  5243 => x"00000000",
  5244 => x"00000000",
  5245 => x"00000000",
  5246 => x"00ff0000",
  5247 => x"0000c645",
  5248 => x"44800785",
  5249 => x"45408007",
  5250 => x"80424700",
  5251 => x"80474000",
  5252 => x"07c14344",
  5253 => x"00c38404",
  5254 => x"c30007c1",
  5255 => x"42418700",
  5256 => x"80404784",
  5257 => x"04c34047",
  5258 => x"8101c640",
  5259 => x"40070505",
  5260 => x"00040502",
  5261 => x"00000704",
  5262 => x"04030007",
  5263 => x"05050007",
  5264 => x"00020700",
  5265 => x"00000000",
  5266 => x"00000000",
  5267 => x"00000000",
  5268 => x"00000000",
  5269 => x"0000ff00",
  5270 => x"00000007",
  5271 => x"01030500",
  5272 => x"03040403",
  5273 => x"00040502",
  5274 => x"00040502",
  5275 => x"00000705",
  5276 => x"05000700",
  5277 => x"02070000",
  5278 => x"07040403",
  5279 => x"00030404",
  5280 => x"03000701",
  5281 => x"03050007",
  5282 => x"01010000",
  5283 => x"00000000",
  5284 => x"00000000",
  5285 => x"00000000",
  5286 => x"00000000",
  5287 => x"00000000",
  5288 => x"71756974",
  5289 => x"00000000",
  5290 => x"68656c70",
  5291 => x"00000000",
  5292 => x"0a307800",
  5293 => x"69326320",
  5294 => x"464d430a",
  5295 => x"00000000",
  5296 => x"61646472",
  5297 => x"6573733a",
  5298 => x"20307800",
  5299 => x"2020202d",
  5300 => x"2d3e2020",
  5301 => x"2041434b",
  5302 => x"0a000000",
  5303 => x"72656164",
  5304 => x"20646174",
  5305 => x"61202800",
  5306 => x"20627974",
  5307 => x"65732920",
  5308 => x"66726f6d",
  5309 => x"20493243",
  5310 => x"2d616464",
  5311 => x"72657373",
  5312 => x"20307800",
  5313 => x"0a0a0000",
  5314 => x"6e6f6163",
  5315 => x"6b200000",
  5316 => x"6368726f",
  5317 => x"6e74656c",
  5318 => x"20726567",
  5319 => x"20307800",
  5320 => x"3a203078",
  5321 => x"00000000",
  5322 => x"206e6163",
  5323 => x"6b000000",
  5324 => x"6572726f",
  5325 => x"7220286e",
  5326 => x"61636b29",
  5327 => x"0a000000",
  5328 => x"0a202063",
  5329 => x"68616e6e",
  5330 => x"656c2033",
  5331 => x"20696e70",
  5332 => x"7574206f",
  5333 => x"76657266",
  5334 => x"6c6f7700",
  5335 => x"0a202063",
  5336 => x"68616e6e",
  5337 => x"656c2032",
  5338 => x"20696e70",
  5339 => x"7574206f",
  5340 => x"76657266",
  5341 => x"6c6f7700",
  5342 => x"0a202063",
  5343 => x"68616e6e",
  5344 => x"656c2031",
  5345 => x"20696e70",
  5346 => x"7574206f",
  5347 => x"76657266",
  5348 => x"6c6f7700",
  5349 => x"0a202063",
  5350 => x"68616e6e",
  5351 => x"656c2030",
  5352 => x"20696e70",
  5353 => x"7574206f",
  5354 => x"76657266",
  5355 => x"6c6f7700",
  5356 => x"0a202063",
  5357 => x"68616e6e",
  5358 => x"656c2033",
  5359 => x"20717561",
  5360 => x"6473756d",
  5361 => x"206f7665",
  5362 => x"72666c6f",
  5363 => x"77000000",
  5364 => x"0a202063",
  5365 => x"68616e6e",
  5366 => x"656c2032",
  5367 => x"20717561",
  5368 => x"6473756d",
  5369 => x"206f7665",
  5370 => x"72666c6f",
  5371 => x"77000000",
  5372 => x"0a202063",
  5373 => x"68616e6e",
  5374 => x"656c2031",
  5375 => x"20717561",
  5376 => x"6473756d",
  5377 => x"206f7665",
  5378 => x"72666c6f",
  5379 => x"77000000",
  5380 => x"0a202063",
  5381 => x"68616e6e",
  5382 => x"656c2030",
  5383 => x"20717561",
  5384 => x"6473756d",
  5385 => x"206f7665",
  5386 => x"72666c6f",
  5387 => x"77000000",
  5388 => x"0a202073",
  5389 => x"756d2076",
  5390 => x"616c7565",
  5391 => x"20637574",
  5392 => x"74656400",
  5393 => x"0a202063",
  5394 => x"68616e6e",
  5395 => x"656c2033",
  5396 => x"20646976",
  5397 => x"6964656e",
  5398 => x"64206375",
  5399 => x"74746564",
  5400 => x"00000000",
  5401 => x"0a202063",
  5402 => x"68616e6e",
  5403 => x"656c2033",
  5404 => x"206e6f69",
  5405 => x"73652063",
  5406 => x"6f6d7065",
  5407 => x"6e736174",
  5408 => x"696f6e20",
  5409 => x"746f2062",
  5410 => x"69670000",
  5411 => x"0a202063",
  5412 => x"68616e6e",
  5413 => x"656c2033",
  5414 => x"206e6f69",
  5415 => x"73652076",
  5416 => x"616c7565",
  5417 => x"20637574",
  5418 => x"74656400",
  5419 => x"0a202063",
  5420 => x"68616e6e",
  5421 => x"656c2032",
  5422 => x"20646976",
  5423 => x"6964656e",
  5424 => x"64206375",
  5425 => x"74746564",
  5426 => x"00000000",
  5427 => x"0a202063",
  5428 => x"68616e6e",
  5429 => x"656c2032",
  5430 => x"206e6f69",
  5431 => x"73652063",
  5432 => x"6f6d7065",
  5433 => x"6e736174",
  5434 => x"696f6e20",
  5435 => x"746f2062",
  5436 => x"69670000",
  5437 => x"0a202063",
  5438 => x"68616e6e",
  5439 => x"656c2032",
  5440 => x"206e6f69",
  5441 => x"73652076",
  5442 => x"616c7565",
  5443 => x"20637574",
  5444 => x"74656400",
  5445 => x"0a202063",
  5446 => x"68616e6e",
  5447 => x"656c2031",
  5448 => x"20646976",
  5449 => x"6964656e",
  5450 => x"64206375",
  5451 => x"74746564",
  5452 => x"00000000",
  5453 => x"0a202063",
  5454 => x"68616e6e",
  5455 => x"656c2031",
  5456 => x"206e6f69",
  5457 => x"73652063",
  5458 => x"6f6d7065",
  5459 => x"6e736174",
  5460 => x"696f6e20",
  5461 => x"746f2062",
  5462 => x"69670000",
  5463 => x"0a202063",
  5464 => x"68616e6e",
  5465 => x"656c2031",
  5466 => x"206e6f69",
  5467 => x"73652076",
  5468 => x"616c7565",
  5469 => x"20637574",
  5470 => x"74656400",
  5471 => x"0a202063",
  5472 => x"68616e6e",
  5473 => x"656c2030",
  5474 => x"20646976",
  5475 => x"6964656e",
  5476 => x"64206375",
  5477 => x"74746564",
  5478 => x"00000000",
  5479 => x"0a202063",
  5480 => x"68616e6e",
  5481 => x"656c2030",
  5482 => x"206e6f69",
  5483 => x"73652063",
  5484 => x"6f6d7065",
  5485 => x"6e736174",
  5486 => x"696f6e20",
  5487 => x"746f2062",
  5488 => x"69670000",
  5489 => x"0a202063",
  5490 => x"68616e6e",
  5491 => x"656c2030",
  5492 => x"206e6f69",
  5493 => x"73652076",
  5494 => x"616c7565",
  5495 => x"20637574",
  5496 => x"74656400",
  5497 => x"0a202073",
  5498 => x"6f667477",
  5499 => x"61726520",
  5500 => x"6572726f",
  5501 => x"72000000",
  5502 => x"0a657874",
  5503 => x"65726e61",
  5504 => x"6c20636c",
  5505 => x"6f636b20",
  5506 => x"20202020",
  5507 => x"2020203a",
  5508 => x"20000000",
  5509 => x"61637469",
  5510 => x"76650000",
  5511 => x"0a6d6963",
  5512 => x"726f7075",
  5513 => x"6c736520",
  5514 => x"736f7572",
  5515 => x"63652020",
  5516 => x"2020203a",
  5517 => x"20000000",
  5518 => x"65787465",
  5519 => x"726e616c",
  5520 => x"00000000",
  5521 => x"0a6d6963",
  5522 => x"726f7075",
  5523 => x"6c736520",
  5524 => x"6576656e",
  5525 => x"74206c69",
  5526 => x"6d69743a",
  5527 => x"20000000",
  5528 => x"0a6d6561",
  5529 => x"73757265",
  5530 => x"6d656e74",
  5531 => x"206c656e",
  5532 => x"67746820",
  5533 => x"2020203a",
  5534 => x"20000000",
  5535 => x"0a626561",
  5536 => x"6d20706f",
  5537 => x"73697469",
  5538 => x"6f6e206d",
  5539 => x"6f6e6974",
  5540 => x"6f722072",
  5541 => x"65676973",
  5542 => x"74657273",
  5543 => x"00000000",
  5544 => x"0a202020",
  5545 => x"20202020",
  5546 => x"20202020",
  5547 => x"20202020",
  5548 => x"20202020",
  5549 => x"20202020",
  5550 => x"20636861",
  5551 => x"6e6e656c",
  5552 => x"20302020",
  5553 => x"20636861",
  5554 => x"6e6e656c",
  5555 => x"20312020",
  5556 => x"20636861",
  5557 => x"6e6e656c",
  5558 => x"20322020",
  5559 => x"20636861",
  5560 => x"6e6e656c",
  5561 => x"20330000",
  5562 => x"0a202020",
  5563 => x"20202020",
  5564 => x"20202020",
  5565 => x"20202020",
  5566 => x"20202020",
  5567 => x"20202020",
  5568 => x"202d2d2d",
  5569 => x"2d20686f",
  5570 => x"72697a6f",
  5571 => x"6e74616c",
  5572 => x"202d2d2d",
  5573 => x"2d2d2020",
  5574 => x"202d2d2d",
  5575 => x"2d2d2d20",
  5576 => x"76657274",
  5577 => x"6963616c",
  5578 => x"202d2d2d",
  5579 => x"2d2d0000",
  5580 => x"0a736361",
  5581 => x"6c657220",
  5582 => x"76616c75",
  5583 => x"65732020",
  5584 => x"20202020",
  5585 => x"20202020",
  5586 => x"20000000",
  5587 => x"0a6e6f69",
  5588 => x"73652063",
  5589 => x"6f6d7065",
  5590 => x"6e736174",
  5591 => x"696f6e20",
  5592 => x"20202020",
  5593 => x"20000000",
  5594 => x"0a6d6561",
  5595 => x"73757265",
  5596 => x"6d656e74",
  5597 => x"20202020",
  5598 => x"20202020",
  5599 => x"20202020",
  5600 => x"20000000",
  5601 => x"0a73616d",
  5602 => x"706c6573",
  5603 => x"20286469",
  5604 => x"7629203a",
  5605 => x"20000000",
  5606 => x"0a73756d",
  5607 => x"20636861",
  5608 => x"6e6e656c",
  5609 => x"2020203a",
  5610 => x"20000000",
  5611 => x"0a0a706f",
  5612 => x"73697469",
  5613 => x"6f6e2063",
  5614 => x"6f6d7075",
  5615 => x"74617469",
  5616 => x"6f6e0000",
  5617 => x"0a202073",
  5618 => x"63616c65",
  5619 => x"72207661",
  5620 => x"6c756573",
  5621 => x"20202020",
  5622 => x"20202020",
  5623 => x"20000000",
  5624 => x"0a20206f",
  5625 => x"66667365",
  5626 => x"74202020",
  5627 => x"20202020",
  5628 => x"20202020",
  5629 => x"20202020",
  5630 => x"20000000",
  5631 => x"0a6f7574",
  5632 => x"70757420",
  5633 => x"73656c65",
  5634 => x"6374203a",
  5635 => x"20000000",
  5636 => x"74657374",
  5637 => x"67656e00",
  5638 => x"4e4f5420",
  5639 => x"00000000",
  5640 => x"6368616e",
  5641 => x"6e656c20",
  5642 => x"30000000",
  5643 => x"0a63616c",
  5644 => x"63207374",
  5645 => x"61746520",
  5646 => x"2020203a",
  5647 => x"20307800",
  5648 => x"76657274",
  5649 => x"6963616c",
  5650 => x"00000000",
  5651 => x"686f7269",
  5652 => x"7a6f6e74",
  5653 => x"616c0000",
  5654 => x"73756d00",
  5655 => x"6368616e",
  5656 => x"6e656c20",
  5657 => x"33000000",
  5658 => x"6368616e",
  5659 => x"6e656c20",
  5660 => x"32000000",
  5661 => x"6368616e",
  5662 => x"6e656c20",
  5663 => x"31000000",
  5664 => x"786d6f64",
  5665 => x"656d2074",
  5666 => x"72616e73",
  5667 => x"6d69742e",
  5668 => x"2e2e0a00",
  5669 => x"20627974",
  5670 => x"65732074",
  5671 => x"72616e73",
  5672 => x"6d697474",
  5673 => x"65640a00",
  5674 => x"63616e63",
  5675 => x"656c0a00",
  5676 => x"72657472",
  5677 => x"79206f75",
  5678 => x"740a0000",
  5679 => x"786d6f64",
  5680 => x"656d2072",
  5681 => x"65636569",
  5682 => x"76652e2e",
  5683 => x"2e0a0000",
  5684 => x"20627974",
  5685 => x"65732072",
  5686 => x"65636569",
  5687 => x"7665640a",
  5688 => x"00000000",
  5689 => x"72782062",
  5690 => x"75666665",
  5691 => x"72206675",
  5692 => x"6c6c0a00",
  5693 => x"74696d65",
  5694 => x"206f7574",
  5695 => x"0a000000",
  5696 => x"64656275",
  5697 => x"67207265",
  5698 => x"67697374",
  5699 => x"65727300",
  5700 => x"0a6d6f64",
  5701 => x"65202020",
  5702 => x"20202020",
  5703 => x"203a2000",
  5704 => x"0a616464",
  5705 => x"72657373",
  5706 => x"20302020",
  5707 => x"203a2030",
  5708 => x"78000000",
  5709 => x"0a616464",
  5710 => x"72657373",
  5711 => x"20312020",
  5712 => x"203a2030",
  5713 => x"78000000",
  5714 => x"0a627566",
  5715 => x"66657220",
  5716 => x"73697a65",
  5717 => x"203a2000",
  5718 => x"6d61783a",
  5719 => x"20000000",
  5720 => x"6d696e3a",
  5721 => x"20000000",
  5722 => x"63683a20",
  5723 => x"00000000",
  5724 => x"73706c3a",
  5725 => x"20000000",
  5726 => x"73686f77",
  5727 => x"2042504d",
  5728 => x"20726567",
  5729 => x"69737465",
  5730 => x"72730000",
  5731 => x"62706d00",
  5732 => x"73656c65",
  5733 => x"6374206f",
  5734 => x"75747075",
  5735 => x"74206368",
  5736 => x"616e6e65",
  5737 => x"6c202830",
  5738 => x"2e2e3320",
  5739 => x"73756d20",
  5740 => x"68207629",
  5741 => x"00000000",
  5742 => x"73656c65",
  5743 => x"63740000",
  5744 => x"73797374",
  5745 => x"656d2072",
  5746 => x"65736574",
  5747 => x"00000000",
  5748 => x"72657365",
  5749 => x"74000000",
  5750 => x"73686f77",
  5751 => x"20737973",
  5752 => x"74656d20",
  5753 => x"696e666f",
  5754 => x"203c7665",
  5755 => x"72626f73",
  5756 => x"653e0000",
  5757 => x"73797369",
  5758 => x"6e666f00",
  5759 => x"73686f77",
  5760 => x"2f736574",
  5761 => x"20646562",
  5762 => x"75672072",
  5763 => x"65676973",
  5764 => x"74657273",
  5765 => x"203c7365",
  5766 => x"74206d6f",
  5767 => x"64653e00",
  5768 => x"64656275",
  5769 => x"67000000",
  5770 => x"636c6b20",
  5771 => x"736f7572",
  5772 => x"63653a20",
  5773 => x"2030203d",
  5774 => x"20696e74",
  5775 => x"2c203120",
  5776 => x"3d206578",
  5777 => x"74000000",
  5778 => x"636c6b00",
  5779 => x"6d696372",
  5780 => x"6f70756c",
  5781 => x"73652073",
  5782 => x"6f757263",
  5783 => x"653a2030",
  5784 => x"203d2069",
  5785 => x"6e742c20",
  5786 => x"31203d20",
  5787 => x"65787400",
  5788 => x"6d696372",
  5789 => x"6f000000",
  5790 => x"74657374",
  5791 => x"67656e65",
  5792 => x"7261746f",
  5793 => x"72203c73",
  5794 => x"63616c65",
  5795 => x"723e203c",
  5796 => x"72657374",
  5797 => x"6172743e",
  5798 => x"00000000",
  5799 => x"3c6d7574",
  5800 => x"655f6e3e",
  5801 => x"203c7273",
  5802 => x"745f6e3e",
  5803 => x"203c6270",
  5804 => x"625f6e3e",
  5805 => x"203c6f73",
  5806 => x"72313e20",
  5807 => x"3c6f7372",
  5808 => x"323e0000",
  5809 => x"64616363",
  5810 => x"6f6e6600",
  5811 => x"3c6d756c",
  5812 => x"7469706c",
  5813 => x"6965723e",
  5814 => x"20696e69",
  5815 => x"7469616c",
  5816 => x"697a6520",
  5817 => x"62756666",
  5818 => x"65720000",
  5819 => x"64616374",
  5820 => x"65737400",
  5821 => x"72657365",
  5822 => x"74206361",
  5823 => x"6c63756c",
  5824 => x"6174696f",
  5825 => x"6e206572",
  5826 => x"726f7273",
  5827 => x"00000000",
  5828 => x"63616c63",
  5829 => x"72657300",
  5830 => x"73686f77",
  5831 => x"20646562",
  5832 => x"75672062",
  5833 => x"75666665",
  5834 => x"72203c6c",
  5835 => x"656e6774",
  5836 => x"683e0000",
  5837 => x"636c6561",
  5838 => x"72206465",
  5839 => x"62756720",
  5840 => x"62756666",
  5841 => x"65720000",
  5842 => x"62636c65",
  5843 => x"61720000",
  5844 => x"62756666",
  5845 => x"6572206f",
  5846 => x"6e204c43",
  5847 => x"44203c63",
  5848 => x"683e203c",
  5849 => x"636f6d62",
  5850 => x"3e000000",
  5851 => x"73636f70",
  5852 => x"65000000",
  5853 => x"64656275",
  5854 => x"67207472",
  5855 => x"61636520",
  5856 => x"3c636c65",
  5857 => x"61723e00",
  5858 => x"74726163",
  5859 => x"65000000",
  5860 => x"73657475",
  5861 => x"70206368",
  5862 => x"616e6e65",
  5863 => x"6c207465",
  5864 => x"7374203c",
  5865 => x"63683e20",
  5866 => x"3c76616c",
  5867 => x"302e2e37",
  5868 => x"3e000000",
  5869 => x"63687465",
  5870 => x"73740000",
  5871 => x"72756e6e",
  5872 => x"696e6720",
  5873 => x"6c696768",
  5874 => x"74000000",
  5875 => x"72756e00",
  5876 => x"72756e20",
  5877 => x"64697370",
  5878 => x"6c617920",
  5879 => x"74657374",
  5880 => x"2066756e",
  5881 => x"6374696f",
  5882 => x"6e000000",
  5883 => x"64697370",
  5884 => x"6c617900",
  5885 => x"73657420",
  5886 => x"6261636b",
  5887 => x"6c696768",
  5888 => x"74203c30",
  5889 => x"2e2e3331",
  5890 => x"3e000000",
  5891 => x"6261636b",
  5892 => x"00000000",
  5893 => x"73686f77",
  5894 => x"206c6f67",
  5895 => x"6f206f6e",
  5896 => x"20676c63",
  5897 => x"64000000",
  5898 => x"6c6f676f",
  5899 => x"00000000",
  5900 => x"63686563",
  5901 => x"6b204932",
  5902 => x"43206164",
  5903 => x"64726573",
  5904 => x"73000000",
  5905 => x"69326300",
  5906 => x"72656164",
  5907 => x"20454550",
  5908 => x"524f4d20",
  5909 => x"3c627573",
  5910 => x"3e203c69",
  5911 => x"32635f61",
  5912 => x"6464723e",
  5913 => x"203c6c65",
  5914 => x"6e677468",
  5915 => x"3e000000",
  5916 => x"65657072",
  5917 => x"6f6d0000",
  5918 => x"41444320",
  5919 => x"72656769",
  5920 => x"73746572",
  5921 => x"20747261",
  5922 => x"6e736665",
  5923 => x"72203c76",
  5924 => x"616c7565",
  5925 => x"3e000000",
  5926 => x"61747261",
  5927 => x"6e730000",
  5928 => x"696e6974",
  5929 => x"20414443",
  5930 => x"20726567",
  5931 => x"69737465",
  5932 => x"72730000",
  5933 => x"61696e69",
  5934 => x"74000000",
  5935 => x"616c6961",
  5936 => x"7320666f",
  5937 => x"72207800",
  5938 => x"6d656d00",
  5939 => x"77726974",
  5940 => x"6520776f",
  5941 => x"7264203c",
  5942 => x"61646472",
  5943 => x"3e203c6c",
  5944 => x"656e6774",
  5945 => x"683e203c",
  5946 => x"76616c75",
  5947 => x"65287329",
  5948 => x"3e000000",
  5949 => x"776d656d",
  5950 => x"00000000",
  5951 => x"6558616d",
  5952 => x"696e6520",
  5953 => x"6d656d6f",
  5954 => x"7279203c",
  5955 => x"61646472",
  5956 => x"3e203c6c",
  5957 => x"656e6774",
  5958 => x"683e0000",
  5959 => x"636c6561",
  5960 => x"72207363",
  5961 => x"7265656e",
  5962 => x"00000000",
  5963 => x"636c6561",
  5964 => x"72000000",
  5965 => x"0a646562",
  5966 => x"75672074",
  5967 => x"72616365",
  5968 => x"206d656d",
  5969 => x"6f727900",
  5970 => x"0a74696d",
  5971 => x"65207374",
  5972 => x"616d7020",
  5973 => x"20202073",
  5974 => x"74617465",
  5975 => x"00000000",
  5976 => x"20203078",
  5977 => x"00000000",
  5978 => x"65787465",
  5979 => x"726e616c",
  5980 => x"20636c6f",
  5981 => x"636b2000",
  5982 => x"61637469",
  5983 => x"76650a00",
  5984 => x"73656c65",
  5985 => x"63746564",
  5986 => x"0a000000",
  5987 => x"6d696372",
  5988 => x"6f70756c",
  5989 => x"73652073",
  5990 => x"6f757263",
  5991 => x"653a2000",
  5992 => x"6265616d",
  5993 => x"20706f73",
  5994 => x"6974696f",
  5995 => x"6e206d6f",
  5996 => x"6e69746f",
  5997 => x"72000000",
  5998 => x"20286f6e",
  5999 => x"2073696d",
  6000 => x"290a0000",
  6001 => x"0a485720",
  6002 => x"73796e74",
  6003 => x"68657369",
  6004 => x"7a65643a",
  6005 => x"20000000",
  6006 => x"0a535720",
  6007 => x"636f6d70",
  6008 => x"696c6564",
  6009 => x"2020203a",
  6010 => x"20417567",
  6011 => x"20313820",
  6012 => x"32303131",
  6013 => x"20203131",
  6014 => x"3a32323a",
  6015 => x"35300000",
  6016 => x"0a737973",
  6017 => x"74656d20",
  6018 => x"636c6f63",
  6019 => x"6b20203a",
  6020 => x"20000000",
  6021 => x"204d487a",
  6022 => x"0a000000",
  6023 => x"44454255",
  6024 => x"47204d4f",
  6025 => x"44450000",
  6026 => x"204f4e0a",
  6027 => x"00000000",
  6028 => x"0000117b",
  6029 => x"000011e4",
  6030 => x"000011d9",
  6031 => x"000011ce",
  6032 => x"000011c3",
  6033 => x"000011b9",
  6034 => x"000011af",
  6035 => x"000002c2",
  6036 => x"fc1902c4",
  6037 => x"fffefd3f",
  6038 => x"03e7fd3b",
  6039 => x"0000485d",
  6040 => x"999b4888",
  6041 => x"ffc4b7ce",
  6042 => x"6665b74e",
  6043 => x"3e200000",
  6044 => x"636f6d6d",
  6045 => x"616e6420",
  6046 => x"6e6f7420",
  6047 => x"666f756e",
  6048 => x"642e0a00",
  6049 => x"73757070",
  6050 => x"6f727465",
  6051 => x"6420636f",
  6052 => x"6d6d616e",
  6053 => x"64733a0a",
  6054 => x"0a000000",
  6055 => x"202d2000",
  6056 => x"76656e64",
  6057 => x"6f723f20",
  6058 => x"20000000",
  6059 => x"67616973",
  6060 => x"6c657220",
  6061 => x"20000000",
  6062 => x"756e6b6e",
  6063 => x"6f776e20",
  6064 => x"64657669",
  6065 => x"63650000",
  6066 => x"485a4452",
  6067 => x"20202020",
  6068 => x"20000000",
  6069 => x"56474120",
  6070 => x"636f6e74",
  6071 => x"726f6c6c",
  6072 => x"65720000",
  6073 => x"47656e65",
  6074 => x"72616c20",
  6075 => x"50757270",
  6076 => x"6f736520",
  6077 => x"492f4f20",
  6078 => x"706f7274",
  6079 => x"00000000",
  6080 => x"4475616c",
  6081 => x"2d706f72",
  6082 => x"74204148",
  6083 => x"42205352",
  6084 => x"414d206d",
  6085 => x"6f64756c",
  6086 => x"65000000",
  6087 => x"64656275",
  6088 => x"67206275",
  6089 => x"66666572",
  6090 => x"20636f6e",
  6091 => x"74726f6c",
  6092 => x"00000000",
  6093 => x"74726967",
  6094 => x"67657220",
  6095 => x"67656e65",
  6096 => x"7261746f",
  6097 => x"72000000",
  6098 => x"64656275",
  6099 => x"6720636f",
  6100 => x"6e736f6c",
  6101 => x"65000000",
  6102 => x"64656275",
  6103 => x"67207472",
  6104 => x"61636572",
  6105 => x"206d656d",
  6106 => x"6f727900",
  6107 => x"4541444f",
  6108 => x"47533130",
  6109 => x"32206469",
  6110 => x"73706c61",
  6111 => x"79206472",
  6112 => x"69766572",
  6113 => x"00000000",
  6114 => x"44434d20",
  6115 => x"70686173",
  6116 => x"65207368",
  6117 => x"69667420",
  6118 => x"636f6e74",
  6119 => x"726f6c00",
  6120 => x"5a505520",
  6121 => x"4d656d6f",
  6122 => x"72792077",
  6123 => x"72617070",
  6124 => x"65720000",
  6125 => x"5a505520",
  6126 => x"41484220",
  6127 => x"57726170",
  6128 => x"70657200",
  6129 => x"4148422f",
  6130 => x"41504220",
  6131 => x"42726964",
  6132 => x"67650000",
  6133 => x"4d6f6475",
  6134 => x"6c617220",
  6135 => x"54696d65",
  6136 => x"7220556e",
  6137 => x"69740000",
  6138 => x"47656e65",
  6139 => x"72696320",
  6140 => x"55415254",
  6141 => x"00000000",
  6142 => x"414d4241",
  6143 => x"20577261",
  6144 => x"70706572",
  6145 => x"20666f72",
  6146 => x"204f4320",
  6147 => x"4932432d",
  6148 => x"6d617374",
  6149 => x"65720000",
  6150 => x"53504920",
  6151 => x"4d656d6f",
  6152 => x"72792043",
  6153 => x"6f6e7472",
  6154 => x"6f6c6c65",
  6155 => x"72000000",
  6156 => x"20206170",
  6157 => x"62736c76",
  6158 => x"00000000",
  6159 => x"76656e64",
  6160 => x"20307800",
  6161 => x"64657620",
  6162 => x"30780000",
  6163 => x"76657220",
  6164 => x"00000000",
  6165 => x"69727120",
  6166 => x"00000000",
  6167 => x"61646472",
  6168 => x"20307800",
  6169 => x"6168626d",
  6170 => x"73740000",
  6171 => x"61686273",
  6172 => x"6c760000",
  6173 => x"00002b01",
  6174 => x"00002bc9",
  6175 => x"00002bbe",
  6176 => x"00002bb3",
  6177 => x"00002b92",
  6178 => x"00002b87",
  6179 => x"00002b7c",
  6180 => x"00002b71",
  6181 => x"00002ba8",
  6182 => x"00002b9d",
  6183 => x"04580808",
  6184 => x"20ff0000",
  6185 => x"000060ac",
  6186 => x"0000618c",
  6187 => x"02010305",
  6188 => x"05070501",
  6189 => x"03030505",
  6190 => x"02030104",
  6191 => x"05050505",
  6192 => x"05050505",
  6193 => x"05050101",
  6194 => x"04050404",
  6195 => x"07050505",
  6196 => x"05050505",
  6197 => x"05030405",
  6198 => x"05050505",
  6199 => x"05050505",
  6200 => x"05050505",
  6201 => x"05050503",
  6202 => x"04030505",
  6203 => x"02050504",
  6204 => x"05050405",
  6205 => x"04010204",
  6206 => x"02050404",
  6207 => x"05050404",
  6208 => x"04040507",
  6209 => x"05040404",
  6210 => x"02040500",
  6211 => x"04050200",
  6212 => x"04080303",
  6213 => x"04090003",
  6214 => x"06000000",
  6215 => x"00020204",
  6216 => x"04040400",
  6217 => x"04060003",
  6218 => x"05000000",
  6219 => x"00000404",
  6220 => x"05050204",
  6221 => x"05060305",
  6222 => x"04030705",
  6223 => x"04050303",
  6224 => x"02040502",
  6225 => x"03020405",
  6226 => x"06060604",
  6227 => x"05050505",
  6228 => x"05050504",
  6229 => x"04040404",
  6230 => x"03030303",
  6231 => x"05050505",
  6232 => x"05050505",
  6233 => x"05040404",
  6234 => x"04050404",
  6235 => x"04040404",
  6236 => x"04040503",
  6237 => x"04040404",
  6238 => x"02020303",
  6239 => x"04040404",
  6240 => x"04040405",
  6241 => x"04040404",
  6242 => x"04030303",
  6243 => x"00005f07",
  6244 => x"0007741c",
  6245 => x"771c172e",
  6246 => x"6a3e2b3a",
  6247 => x"06493608",
  6248 => x"36493036",
  6249 => x"49597648",
  6250 => x"073c4281",
  6251 => x"81423c0a",
  6252 => x"041f040a",
  6253 => x"08083e08",
  6254 => x"08806008",
  6255 => x"080840c0",
  6256 => x"300c033e",
  6257 => x"4141413e",
  6258 => x"44427f40",
  6259 => x"40466151",
  6260 => x"49462241",
  6261 => x"49493618",
  6262 => x"14127f10",
  6263 => x"27454545",
  6264 => x"393e4949",
  6265 => x"49300101",
  6266 => x"710d0336",
  6267 => x"49494936",
  6268 => x"06494929",
  6269 => x"1e36d008",
  6270 => x"14224114",
  6271 => x"14141414",
  6272 => x"41221408",
  6273 => x"02510906",
  6274 => x"3c4299a5",
  6275 => x"bd421c7c",
  6276 => x"1211127c",
  6277 => x"7f494949",
  6278 => x"363e4141",
  6279 => x"41227f41",
  6280 => x"41413e7f",
  6281 => x"49494941",
  6282 => x"7f090909",
  6283 => x"013e4149",
  6284 => x"497a7f08",
  6285 => x"08087f41",
  6286 => x"7f414041",
  6287 => x"413f7f08",
  6288 => x"1422417f",
  6289 => x"40404040",
  6290 => x"7f060c06",
  6291 => x"7f7f0608",
  6292 => x"307f3e41",
  6293 => x"41413e7f",
  6294 => x"09090906",
  6295 => x"3e4161c1",
  6296 => x"be7f0919",
  6297 => x"29462649",
  6298 => x"49493201",
  6299 => x"017f0101",
  6300 => x"3f404040",
  6301 => x"3f073840",
  6302 => x"38071f60",
  6303 => x"1f601f63",
  6304 => x"14081463",
  6305 => x"01067806",
  6306 => x"01615149",
  6307 => x"45437f41",
  6308 => x"41030c30",
  6309 => x"c041417f",
  6310 => x"04020102",
  6311 => x"04808080",
  6312 => x"80800102",
  6313 => x"20545454",
  6314 => x"787f4444",
  6315 => x"44383844",
  6316 => x"44443844",
  6317 => x"44447f38",
  6318 => x"54545458",
  6319 => x"087e0901",
  6320 => x"18a4a4a4",
  6321 => x"787f0404",
  6322 => x"787d807d",
  6323 => x"7f102844",
  6324 => x"3f407c04",
  6325 => x"7804787c",
  6326 => x"04047838",
  6327 => x"444438fc",
  6328 => x"24242418",
  6329 => x"18242424",
  6330 => x"fc7c0804",
  6331 => x"04485454",
  6332 => x"24043f44",
  6333 => x"403c4040",
  6334 => x"7c1c2040",
  6335 => x"201c1c60",
  6336 => x"601c6060",
  6337 => x"1c442810",
  6338 => x"28449ca0",
  6339 => x"601c6454",
  6340 => x"544c187e",
  6341 => x"8181ffff",
  6342 => x"81817e18",
  6343 => x"18040810",
  6344 => x"0c143e55",
  6345 => x"55ff8181",
  6346 => x"81ff8060",
  6347 => x"80608060",
  6348 => x"60600060",
  6349 => x"60006060",
  6350 => x"047f0414",
  6351 => x"7f140201",
  6352 => x"01024629",
  6353 => x"1608344a",
  6354 => x"31483000",
  6355 => x"18243e41",
  6356 => x"227f4941",
  6357 => x"03040403",
  6358 => x"03040304",
  6359 => x"04030403",
  6360 => x"183c3c18",
  6361 => x"08080808",
  6362 => x"03010203",
  6363 => x"020e020e",
  6364 => x"060e0048",
  6365 => x"30384438",
  6366 => x"54483844",
  6367 => x"fe44487e",
  6368 => x"49014438",
  6369 => x"28384403",
  6370 => x"147c1403",
  6371 => x"e7e74e55",
  6372 => x"55390101",
  6373 => x"0001011c",
  6374 => x"2a555522",
  6375 => x"1c1d151e",
  6376 => x"18240018",
  6377 => x"24080808",
  6378 => x"18080808",
  6379 => x"3c42bd95",
  6380 => x"a9423c01",
  6381 => x"01010101",
  6382 => x"06090906",
  6383 => x"44445f44",
  6384 => x"44191512",
  6385 => x"15150a02",
  6386 => x"01fc2020",
  6387 => x"1c0e7f01",
  6388 => x"7f011818",
  6389 => x"00804002",
  6390 => x"1f060909",
  6391 => x"06241800",
  6392 => x"2418824f",
  6393 => x"304c62f1",
  6394 => x"824f300c",
  6395 => x"d2b1955f",
  6396 => x"304c62f1",
  6397 => x"30484520",
  6398 => x"60392e38",
  6399 => x"6060382e",
  6400 => x"3960701d",
  6401 => x"131d7072",
  6402 => x"1d121e71",
  6403 => x"701d121d",
  6404 => x"70603b25",
  6405 => x"3b607e11",
  6406 => x"7f49411e",
  6407 => x"2161927c",
  6408 => x"5556447c",
  6409 => x"5655447c",
  6410 => x"5655467d",
  6411 => x"54544545",
  6412 => x"7e44447e",
  6413 => x"45467d46",
  6414 => x"457c4508",
  6415 => x"7f49413e",
  6416 => x"7e091222",
  6417 => x"7d384546",
  6418 => x"44383844",
  6419 => x"46453838",
  6420 => x"46454638",
  6421 => x"3a454546",
  6422 => x"39384544",
  6423 => x"45382214",
  6424 => x"081422bc",
  6425 => x"625a463d",
  6426 => x"3c41423c",
  6427 => x"3c42413c",
  6428 => x"3c42413e",
  6429 => x"3d40403d",
  6430 => x"0608f209",
  6431 => x"067f2222",
  6432 => x"1cfe0989",
  6433 => x"76205556",
  6434 => x"78205655",
  6435 => x"78225555",
  6436 => x"7a235556",
  6437 => x"7b205554",
  6438 => x"79275557",
  6439 => x"78205438",
  6440 => x"54483844",
  6441 => x"c4385556",
  6442 => x"58385655",
  6443 => x"583a5555",
  6444 => x"5a395454",
  6445 => x"59017a7a",
  6446 => x"01027902",
  6447 => x"02780260",
  6448 => x"91927c7b",
  6449 => x"090a7338",
  6450 => x"45463838",
  6451 => x"4645383a",
  6452 => x"45453a3b",
  6453 => x"45463b39",
  6454 => x"44443908",
  6455 => x"082a0808",
  6456 => x"b8644c3a",
  6457 => x"3c41427c",
  6458 => x"3c42417c",
  6459 => x"3a41417a",
  6460 => x"3d40407d",
  6461 => x"986219ff",
  6462 => x"423c9a60",
  6463 => x"1a000000",
  6464 => x"30622020",
  6465 => x"20202020",
  6466 => x"20202020",
  6467 => x"20202020",
  6468 => x"20202020",
  6469 => x"20202020",
  6470 => x"20202020",
  6471 => x"20202020",
  6472 => x"20200000",
  6473 => x"20202020",
  6474 => x"20202020",
  6475 => x"00000000",
  6476 => x"00202020",
  6477 => x"20202020",
  6478 => x"20202828",
  6479 => x"28282820",
  6480 => x"20202020",
  6481 => x"20202020",
  6482 => x"20202020",
  6483 => x"20202020",
  6484 => x"20881010",
  6485 => x"10101010",
  6486 => x"10101010",
  6487 => x"10101010",
  6488 => x"10040404",
  6489 => x"04040404",
  6490 => x"04040410",
  6491 => x"10101010",
  6492 => x"10104141",
  6493 => x"41414141",
  6494 => x"01010101",
  6495 => x"01010101",
  6496 => x"01010101",
  6497 => x"01010101",
  6498 => x"01010101",
  6499 => x"10101010",
  6500 => x"10104242",
  6501 => x"42424242",
  6502 => x"02020202",
  6503 => x"02020202",
  6504 => x"02020202",
  6505 => x"02020202",
  6506 => x"02020202",
  6507 => x"10101010",
  6508 => x"20000000",
  6509 => x"00000000",
  6510 => x"00000000",
  6511 => x"00000000",
  6512 => x"00000000",
  6513 => x"00000000",
  6514 => x"00000000",
  6515 => x"00000000",
  6516 => x"00000000",
  6517 => x"00000000",
  6518 => x"00000000",
  6519 => x"00000000",
  6520 => x"00000000",
  6521 => x"00000000",
  6522 => x"00000000",
  6523 => x"00000000",
  6524 => x"00000000",
  6525 => x"00000000",
  6526 => x"00000000",
  6527 => x"00000000",
  6528 => x"00000000",
  6529 => x"00000000",
  6530 => x"00000000",
  6531 => x"00000000",
  6532 => x"00000000",
  6533 => x"00000000",
  6534 => x"00000000",
  6535 => x"00000000",
  6536 => x"00000000",
  6537 => x"00000000",
  6538 => x"00000000",
  6539 => x"00000000",
  6540 => x"00000000",
  6541 => x"43000000",
  6542 => x"00000000",
  6543 => x"80000c00",
  6544 => x"80000b00",
  6545 => x"80000800",
  6546 => x"00000000",
  6547 => x"ff000000",
  6548 => x"00000000",
  6549 => x"00000000",
  6550 => x"00ffffff",
  6551 => x"ff00ffff",
  6552 => x"ffff00ff",
  6553 => x"ffffff00",
  6554 => x"00000000",
  6555 => x"00000000",
  6556 => x"80000a00",
  6557 => x"80000700",
  6558 => x"80000600",
  6559 => x"80000400",
  6560 => x"80000200",
  6561 => x"80000100",
  6562 => x"80000004",
  6563 => x"80000000",
  6564 => x"00006694",
  6565 => x"00000000",
  6566 => x"000068fc",
  6567 => x"00006958",
  6568 => x"000069b4",
  6569 => x"00000000",
  6570 => x"00000000",
  6571 => x"00000000",
  6572 => x"00000000",
  6573 => x"00000000",
  6574 => x"00000000",
  6575 => x"00000000",
  6576 => x"00000000",
  6577 => x"00000000",
  6578 => x"00006634",
  6579 => x"00000000",
  6580 => x"00000000",
  6581 => x"00000000",
  6582 => x"00000000",
  6583 => x"00000000",
  6584 => x"00000000",
  6585 => x"00000000",
  6586 => x"00000000",
  6587 => x"00000000",
  6588 => x"00000000",
  6589 => x"00000000",
  6590 => x"00000000",
  6591 => x"00000000",
  6592 => x"00000000",
  6593 => x"00000000",
  6594 => x"00000000",
  6595 => x"00000000",
  6596 => x"00000000",
  6597 => x"00000000",
  6598 => x"00000000",
  6599 => x"00000000",
  6600 => x"00000000",
  6601 => x"00000000",
  6602 => x"00000000",
  6603 => x"00000000",
  6604 => x"00000000",
  6605 => x"00000000",
  6606 => x"00000000",
  6607 => x"00000001",
  6608 => x"330eabcd",
  6609 => x"1234e66d",
  6610 => x"deec0005",
  6611 => x"000b0000",
  6612 => x"00000000",
  6613 => x"00000000",
  6614 => x"00000000",
  6615 => x"00000000",
  6616 => x"00000000",
  6617 => x"00000000",
  6618 => x"00000000",
  6619 => x"00000000",
  6620 => x"00000000",
  6621 => x"00000000",
  6622 => x"00000000",
  6623 => x"00000000",
  6624 => x"00000000",
  6625 => x"00000000",
  6626 => x"00000000",
  6627 => x"00000000",
  6628 => x"00000000",
  6629 => x"00000000",
  6630 => x"00000000",
  6631 => x"00000000",
  6632 => x"00000000",
  6633 => x"00000000",
  6634 => x"00000000",
  6635 => x"00000000",
  6636 => x"00000000",
  6637 => x"00000000",
  6638 => x"00000000",
  6639 => x"00000000",
  6640 => x"00000000",
  6641 => x"00000000",
  6642 => x"00000000",
  6643 => x"00000000",
  6644 => x"00000000",
  6645 => x"00000000",
  6646 => x"00000000",
  6647 => x"00000000",
  6648 => x"00000000",
  6649 => x"00000000",
  6650 => x"00000000",
  6651 => x"00000000",
  6652 => x"00000000",
  6653 => x"00000000",
  6654 => x"00000000",
  6655 => x"00000000",
  6656 => x"00000000",
  6657 => x"00000000",
  6658 => x"00000000",
  6659 => x"00000000",
  6660 => x"00000000",
  6661 => x"00000000",
  6662 => x"00000000",
  6663 => x"00000000",
  6664 => x"00000000",
  6665 => x"00000000",
  6666 => x"00000000",
  6667 => x"00000000",
  6668 => x"00000000",
  6669 => x"00000000",
  6670 => x"00000000",
  6671 => x"00000000",
  6672 => x"00000000",
  6673 => x"00000000",
  6674 => x"00000000",
  6675 => x"00000000",
  6676 => x"00000000",
  6677 => x"00000000",
  6678 => x"00000000",
  6679 => x"00000000",
  6680 => x"00000000",
  6681 => x"00000000",
  6682 => x"00000000",
  6683 => x"00000000",
  6684 => x"00000000",
  6685 => x"00000000",
  6686 => x"00000000",
  6687 => x"00000000",
  6688 => x"00000000",
  6689 => x"00000000",
  6690 => x"00000000",
  6691 => x"00000000",
  6692 => x"00000000",
  6693 => x"00000000",
  6694 => x"00000000",
  6695 => x"00000000",
  6696 => x"00000000",
  6697 => x"00000000",
  6698 => x"00000000",
  6699 => x"00000000",
  6700 => x"00000000",
  6701 => x"00000000",
  6702 => x"00000000",
  6703 => x"00000000",
  6704 => x"00000000",
  6705 => x"00000000",
  6706 => x"00000000",
  6707 => x"00000000",
  6708 => x"00000000",
  6709 => x"00000000",
  6710 => x"00000000",
  6711 => x"00000000",
  6712 => x"00000000",
  6713 => x"00000000",
  6714 => x"00000000",
  6715 => x"00000000",
  6716 => x"00000000",
  6717 => x"00000000",
  6718 => x"00000000",
  6719 => x"00000000",
  6720 => x"00000000",
  6721 => x"00000000",
  6722 => x"00000000",
  6723 => x"00000000",
  6724 => x"00000000",
  6725 => x"00000000",
  6726 => x"00000000",
  6727 => x"00000000",
  6728 => x"00000000",
  6729 => x"00000000",
  6730 => x"00000000",
  6731 => x"00000000",
  6732 => x"00000000",
  6733 => x"00000000",
  6734 => x"00000000",
  6735 => x"00000000",
  6736 => x"00000000",
  6737 => x"00000000",
  6738 => x"00000000",
  6739 => x"00000000",
  6740 => x"00000000",
  6741 => x"00000000",
  6742 => x"00000000",
  6743 => x"00000000",
  6744 => x"00000000",
  6745 => x"00000000",
  6746 => x"00000000",
  6747 => x"00000000",
  6748 => x"00000000",
  6749 => x"00000000",
  6750 => x"00000000",
  6751 => x"00000000",
  6752 => x"00000000",
  6753 => x"00000000",
  6754 => x"00000000",
  6755 => x"00000000",
  6756 => x"00000000",
  6757 => x"00000000",
  6758 => x"00000000",
  6759 => x"00000000",
  6760 => x"00000000",
  6761 => x"00000000",
  6762 => x"00000000",
  6763 => x"00000000",
  6764 => x"00000000",
  6765 => x"00000000",
  6766 => x"00000000",
  6767 => x"00000000",
  6768 => x"00000000",
  6769 => x"00000000",
  6770 => x"00000000",
  6771 => x"00000000",
  6772 => x"00000000",
  6773 => x"00000000",
  6774 => x"00000000",
  6775 => x"00000000",
  6776 => x"00000000",
  6777 => x"00000000",
  6778 => x"00000000",
  6779 => x"00000000",
  6780 => x"00000000",
  6781 => x"00000000",
  6782 => x"00000000",
  6783 => x"00000000",
  6784 => x"00000000",
  6785 => x"00000000",
  6786 => x"00000000",
  6787 => x"00000000",
  6788 => x"00000000",
  6789 => x"00000000",
  6790 => x"00000000",
  6791 => x"00000000",
  6792 => x"00000000",
  6793 => x"00000000",
  6794 => x"00000000",
  6795 => x"00000000",
  6796 => x"00000000",
  6797 => x"00000000",
  6798 => x"00000000",
  6799 => x"00000000",
  6800 => x"ffffffff",
  6801 => x"00000000",
  6802 => x"00020000",
  6803 => x"00000000",
  6804 => x"00000000",
  6805 => x"00006a4c",
  6806 => x"00006a4c",
  6807 => x"00006a54",
  6808 => x"00006a54",
  6809 => x"00006a5c",
  6810 => x"00006a5c",
  6811 => x"00006a64",
  6812 => x"00006a64",
  6813 => x"00006a6c",
  6814 => x"00006a6c",
  6815 => x"00006a74",
  6816 => x"00006a74",
  6817 => x"00006a7c",
  6818 => x"00006a7c",
  6819 => x"00006a84",
  6820 => x"00006a84",
  6821 => x"00006a8c",
  6822 => x"00006a8c",
  6823 => x"00006a94",
  6824 => x"00006a94",
  6825 => x"00006a9c",
  6826 => x"00006a9c",
  6827 => x"00006aa4",
  6828 => x"00006aa4",
  6829 => x"00006aac",
  6830 => x"00006aac",
  6831 => x"00006ab4",
  6832 => x"00006ab4",
  6833 => x"00006abc",
  6834 => x"00006abc",
  6835 => x"00006ac4",
  6836 => x"00006ac4",
  6837 => x"00006acc",
  6838 => x"00006acc",
  6839 => x"00006ad4",
  6840 => x"00006ad4",
  6841 => x"00006adc",
  6842 => x"00006adc",
  6843 => x"00006ae4",
  6844 => x"00006ae4",
  6845 => x"00006aec",
  6846 => x"00006aec",
  6847 => x"00006af4",
  6848 => x"00006af4",
  6849 => x"00006afc",
  6850 => x"00006afc",
  6851 => x"00006b04",
  6852 => x"00006b04",
  6853 => x"00006b0c",
  6854 => x"00006b0c",
  6855 => x"00006b14",
  6856 => x"00006b14",
  6857 => x"00006b1c",
  6858 => x"00006b1c",
  6859 => x"00006b24",
  6860 => x"00006b24",
  6861 => x"00006b2c",
  6862 => x"00006b2c",
  6863 => x"00006b34",
  6864 => x"00006b34",
  6865 => x"00006b3c",
  6866 => x"00006b3c",
  6867 => x"00006b44",
  6868 => x"00006b44",
  6869 => x"00006b4c",
  6870 => x"00006b4c",
  6871 => x"00006b54",
  6872 => x"00006b54",
  6873 => x"00006b5c",
  6874 => x"00006b5c",
  6875 => x"00006b64",
  6876 => x"00006b64",
  6877 => x"00006b6c",
  6878 => x"00006b6c",
  6879 => x"00006b74",
  6880 => x"00006b74",
  6881 => x"00006b7c",
  6882 => x"00006b7c",
  6883 => x"00006b84",
  6884 => x"00006b84",
  6885 => x"00006b8c",
  6886 => x"00006b8c",
  6887 => x"00006b94",
  6888 => x"00006b94",
  6889 => x"00006b9c",
  6890 => x"00006b9c",
  6891 => x"00006ba4",
  6892 => x"00006ba4",
  6893 => x"00006bac",
  6894 => x"00006bac",
  6895 => x"00006bb4",
  6896 => x"00006bb4",
  6897 => x"00006bbc",
  6898 => x"00006bbc",
  6899 => x"00006bc4",
  6900 => x"00006bc4",
  6901 => x"00006bcc",
  6902 => x"00006bcc",
  6903 => x"00006bd4",
  6904 => x"00006bd4",
  6905 => x"00006bdc",
  6906 => x"00006bdc",
  6907 => x"00006be4",
  6908 => x"00006be4",
  6909 => x"00006bec",
  6910 => x"00006bec",
  6911 => x"00006bf4",
  6912 => x"00006bf4",
  6913 => x"00006bfc",
  6914 => x"00006bfc",
  6915 => x"00006c04",
  6916 => x"00006c04",
  6917 => x"00006c0c",
  6918 => x"00006c0c",
  6919 => x"00006c14",
  6920 => x"00006c14",
  6921 => x"00006c1c",
  6922 => x"00006c1c",
  6923 => x"00006c24",
  6924 => x"00006c24",
  6925 => x"00006c2c",
  6926 => x"00006c2c",
  6927 => x"00006c34",
  6928 => x"00006c34",
  6929 => x"00006c3c",
  6930 => x"00006c3c",
  6931 => x"00006c44",
  6932 => x"00006c44",
  6933 => x"00006c4c",
  6934 => x"00006c4c",
  6935 => x"00006c54",
  6936 => x"00006c54",
  6937 => x"00006c5c",
  6938 => x"00006c5c",
  6939 => x"00006c64",
  6940 => x"00006c64",
  6941 => x"00006c6c",
  6942 => x"00006c6c",
  6943 => x"00006c74",
  6944 => x"00006c74",
  6945 => x"00006c7c",
  6946 => x"00006c7c",
  6947 => x"00006c84",
  6948 => x"00006c84",
  6949 => x"00006c8c",
  6950 => x"00006c8c",
  6951 => x"00006c94",
  6952 => x"00006c94",
  6953 => x"00006c9c",
  6954 => x"00006c9c",
  6955 => x"00006ca4",
  6956 => x"00006ca4",
  6957 => x"00006cac",
  6958 => x"00006cac",
  6959 => x"00006cb4",
  6960 => x"00006cb4",
  6961 => x"00006cbc",
  6962 => x"00006cbc",
  6963 => x"00006cc4",
  6964 => x"00006cc4",
  6965 => x"00006ccc",
  6966 => x"00006ccc",
  6967 => x"00006cd4",
  6968 => x"00006cd4",
  6969 => x"00006cdc",
  6970 => x"00006cdc",
  6971 => x"00006ce4",
  6972 => x"00006ce4",
  6973 => x"00006cec",
  6974 => x"00006cec",
  6975 => x"00006cf4",
  6976 => x"00006cf4",
  6977 => x"00006cfc",
  6978 => x"00006cfc",
  6979 => x"00006d04",
  6980 => x"00006d04",
  6981 => x"00006d0c",
  6982 => x"00006d0c",
  6983 => x"00006d14",
  6984 => x"00006d14",
  6985 => x"00006d1c",
  6986 => x"00006d1c",
  6987 => x"00006d24",
  6988 => x"00006d24",
  6989 => x"00006d2c",
  6990 => x"00006d2c",
  6991 => x"00006d34",
  6992 => x"00006d34",
  6993 => x"00006d3c",
  6994 => x"00006d3c",
  6995 => x"00006d44",
  6996 => x"00006d44",
  6997 => x"00006d4c",
  6998 => x"00006d4c",
  6999 => x"00006d54",
  7000 => x"00006d54",
  7001 => x"00006d5c",
  7002 => x"00006d5c",
  7003 => x"00006d64",
  7004 => x"00006d64",
  7005 => x"00006d6c",
  7006 => x"00006d6c",
  7007 => x"00006d74",
  7008 => x"00006d74",
  7009 => x"00006d7c",
  7010 => x"00006d7c",
  7011 => x"00006d84",
  7012 => x"00006d84",
  7013 => x"00006d8c",
  7014 => x"00006d8c",
  7015 => x"00006d94",
  7016 => x"00006d94",
  7017 => x"00006d9c",
  7018 => x"00006d9c",
  7019 => x"00006da4",
  7020 => x"00006da4",
  7021 => x"00006dac",
  7022 => x"00006dac",
  7023 => x"00006db4",
  7024 => x"00006db4",
  7025 => x"00006dbc",
  7026 => x"00006dbc",
  7027 => x"00006dc4",
  7028 => x"00006dc4",
  7029 => x"00006dcc",
  7030 => x"00006dcc",
  7031 => x"00006dd4",
  7032 => x"00006dd4",
  7033 => x"00006ddc",
  7034 => x"00006ddc",
  7035 => x"00006de4",
  7036 => x"00006de4",
  7037 => x"00006dec",
  7038 => x"00006dec",
  7039 => x"00006df4",
  7040 => x"00006df4",
  7041 => x"00006dfc",
  7042 => x"00006dfc",
  7043 => x"00006e04",
  7044 => x"00006e04",
  7045 => x"00006e0c",
  7046 => x"00006e0c",
  7047 => x"00006e14",
  7048 => x"00006e14",
  7049 => x"00006e1c",
  7050 => x"00006e1c",
  7051 => x"00006e24",
  7052 => x"00006e24",
  7053 => x"00006e2c",
  7054 => x"00006e2c",
  7055 => x"00006e34",
  7056 => x"00006e34",
  7057 => x"00006e3c",
  7058 => x"00006e3c",
  7059 => x"00006e44",
  7060 => x"00006e44",
	others => x"00dead00" -- mask for mem check
	--others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
