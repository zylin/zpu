-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"0b0b0b0b",
1 => x"82700b0b",
2 => x"80cfe00c",
3 => x"3a0b0b80",
4 => x"c6e00400",
5 => x"00000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"0b8af02d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"04000000",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"53510400",
38 => x"00000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"51040000",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"53510400",
55 => x"00000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"51040000",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c4040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a535104",
82 => x"00000000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"06075351",
101 => x"04000000",
102 => x"00000000",
103 => x"00000000",
104 => x"71715351",
105 => x"020d0406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"51040000",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"53510400",
125 => x"00000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"52040000",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"05055351",
138 => x"04000000",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07535104",
147 => x"00000000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"04000000",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80cf",
162 => x"cc738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88aa0400",
166 => x"00000000",
167 => x"00000000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0b8b",
171 => x"ab2d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0b8b",
179 => x"ef2d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70547106",
188 => x"73097274",
189 => x"05ff0506",
190 => x"07515151",
191 => x"04000000",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"05705471",
196 => x"06730972",
197 => x"7405ff05",
198 => x"06075151",
199 => x"51040000",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80cfdc0c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"04000000",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"04000000",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"05715351",
250 => x"020d0400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"82c53f80",
257 => x"c6e63f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"51047381",
267 => x"ff067383",
268 => x"06098105",
269 => x"83051010",
270 => x"102b0772",
271 => x"fc060c51",
272 => x"51043c04",
273 => x"72728072",
274 => x"8106ff05",
275 => x"09720605",
276 => x"71105272",
277 => x"0a100a53",
278 => x"72ed3851",
279 => x"51535104",
280 => x"fe3d0d0b",
281 => x"0b80dfc8",
282 => x"08538413",
283 => x"0870882a",
284 => x"70810651",
285 => x"52527080",
286 => x"2ef03871",
287 => x"81ff0680",
288 => x"0c843d0d",
289 => x"04ff3d0d",
290 => x"0b0b80df",
291 => x"c8085271",
292 => x"0870882a",
293 => x"81327081",
294 => x"06515151",
295 => x"70f13873",
296 => x"720c833d",
297 => x"0d0480cf",
298 => x"dc08802e",
299 => x"a43880cf",
300 => x"e008822e",
301 => x"bd388380",
302 => x"800b0b0b",
303 => x"80dfc80c",
304 => x"82a0800b",
305 => x"80dfcc0c",
306 => x"8290800b",
307 => x"80dfd00c",
308 => x"04f88080",
309 => x"80a40b0b",
310 => x"0b80dfc8",
311 => x"0cf88080",
312 => x"82800b80",
313 => x"dfcc0cf8",
314 => x"80808480",
315 => x"0b80dfd0",
316 => x"0c0480c0",
317 => x"a8808c0b",
318 => x"0b0b80df",
319 => x"c80c80c0",
320 => x"a880940b",
321 => x"80dfcc0c",
322 => x"0b0b80cf",
323 => x"980b80df",
324 => x"d00c0470",
325 => x"7080dfd4",
326 => x"335170a7",
327 => x"3880cfe8",
328 => x"08700852",
329 => x"5270802e",
330 => x"94388412",
331 => x"80cfe80c",
332 => x"702d80cf",
333 => x"e8087008",
334 => x"525270ee",
335 => x"38810b80",
336 => x"dfd43450",
337 => x"50040470",
338 => x"0b0b80df",
339 => x"c408802e",
340 => x"8e380b0b",
341 => x"0b0b800b",
342 => x"802e0981",
343 => x"06833850",
344 => x"040b0b80",
345 => x"dfc4510b",
346 => x"0b0bf594",
347 => x"3f500404",
348 => x"803d0d80",
349 => x"dfe00881",
350 => x"1180dfe0",
351 => x"0c51823d",
352 => x"0d04fe3d",
353 => x"0d80dfe0",
354 => x"085380df",
355 => x"e0085272",
356 => x"722e8f38",
357 => x"80cf9c51",
358 => x"82b03f80",
359 => x"dfe00853",
360 => x"e93980cf",
361 => x"ac5182a2",
362 => x"3fe039fb",
363 => x"3d0d7779",
364 => x"55558056",
365 => x"757524ab",
366 => x"38807424",
367 => x"9d388053",
368 => x"73527451",
369 => x"80e13f80",
370 => x"08547580",
371 => x"2e853880",
372 => x"08305473",
373 => x"800c873d",
374 => x"0d047330",
375 => x"76813257",
376 => x"54dc3974",
377 => x"30558156",
378 => x"738025d2",
379 => x"38ec39fa",
380 => x"3d0d787a",
381 => x"57558057",
382 => x"767524a4",
383 => x"38759f2c",
384 => x"54815375",
385 => x"74327431",
386 => x"5274519b",
387 => x"3f800854",
388 => x"76802e85",
389 => x"38800830",
390 => x"5473800c",
391 => x"883d0d04",
392 => x"74305581",
393 => x"57d739fc",
394 => x"3d0d7678",
395 => x"53548153",
396 => x"80747326",
397 => x"52557280",
398 => x"2e983870",
399 => x"802eab38",
400 => x"807224a6",
401 => x"38711073",
402 => x"10757226",
403 => x"53545272",
404 => x"ea387351",
405 => x"78833874",
406 => x"5170800c",
407 => x"863d0d04",
408 => x"720a100a",
409 => x"720a100a",
410 => x"53537280",
411 => x"2ee43871",
412 => x"7426ed38",
413 => x"73723175",
414 => x"7407740a",
415 => x"100a740a",
416 => x"100a5555",
417 => x"5654e339",
418 => x"f73d0d7c",
419 => x"70525380",
420 => x"fd3f7254",
421 => x"8008550b",
422 => x"0b80cfb8",
423 => x"56815780",
424 => x"0881055a",
425 => x"8b3de411",
426 => x"59538259",
427 => x"f413527b",
428 => x"88110852",
429 => x"5381b43f",
430 => x"80083070",
431 => x"8008079f",
432 => x"2c8a0780",
433 => x"0c538b3d",
434 => x"0d04f63d",
435 => x"0d7c80cf",
436 => x"ec087153",
437 => x"5553b73f",
438 => x"72558008",
439 => x"560b0b80",
440 => x"cfb85781",
441 => x"58800881",
442 => x"055b8c3d",
443 => x"e4115a53",
444 => x"825af413",
445 => x"52881408",
446 => x"5180f03f",
447 => x"80083070",
448 => x"8008079f",
449 => x"2c8a0780",
450 => x"0c548c3d",
451 => x"0d047070",
452 => x"70707570",
453 => x"71830653",
454 => x"555270b4",
455 => x"38717008",
456 => x"7009f7fb",
457 => x"fdff1206",
458 => x"f8848281",
459 => x"80065452",
460 => x"53719b38",
461 => x"84137008",
462 => x"7009f7fb",
463 => x"fdff1206",
464 => x"f8848281",
465 => x"80065452",
466 => x"5371802e",
467 => x"e7387252",
468 => x"71335372",
469 => x"802e8a38",
470 => x"81127033",
471 => x"545272f8",
472 => x"38717431",
473 => x"800c5050",
474 => x"505004f2",
475 => x"3d0d6062",
476 => x"88110870",
477 => x"58565f5a",
478 => x"73802e81",
479 => x"8c388c1a",
480 => x"2270832a",
481 => x"81328106",
482 => x"56587486",
483 => x"38901a08",
484 => x"91387951",
485 => x"90b73fff",
486 => x"55800880",
487 => x"ec388c1a",
488 => x"22587d08",
489 => x"55807883",
490 => x"ffff0670",
491 => x"0a100a81",
492 => x"06415c57",
493 => x"7e772e80",
494 => x"d7387690",
495 => x"38740884",
496 => x"16088817",
497 => x"57585676",
498 => x"802ef238",
499 => x"76548880",
500 => x"77278438",
501 => x"88805473",
502 => x"5375529c",
503 => x"1a0851a4",
504 => x"1a085877",
505 => x"2d800b80",
506 => x"082582e0",
507 => x"38800816",
508 => x"77800831",
509 => x"7f880508",
510 => x"80083170",
511 => x"6188050c",
512 => x"5b585678",
513 => x"ffb43880",
514 => x"5574800c",
515 => x"903d0d04",
516 => x"7a813281",
517 => x"06774056",
518 => x"75802e81",
519 => x"bd387690",
520 => x"38740884",
521 => x"16088817",
522 => x"57585976",
523 => x"802ef238",
524 => x"881a0878",
525 => x"83ffff06",
526 => x"70892a81",
527 => x"06565956",
528 => x"73802e82",
529 => x"f8387577",
530 => x"278b3877",
531 => x"872a8106",
532 => x"5c7b82b5",
533 => x"38767627",
534 => x"83387656",
535 => x"75537852",
536 => x"79085185",
537 => x"833f881a",
538 => x"08763188",
539 => x"1b0c7908",
540 => x"167a0c76",
541 => x"56751977",
542 => x"77317f88",
543 => x"05087831",
544 => x"70618805",
545 => x"0c415859",
546 => x"7e802efe",
547 => x"fa388c1a",
548 => x"2258ff8a",
549 => x"39787954",
550 => x"7c537b52",
551 => x"5684c93f",
552 => x"881a0879",
553 => x"31881b0c",
554 => x"7908197a",
555 => x"0c7c7631",
556 => x"5d7c8e38",
557 => x"79518ff2",
558 => x"3f800881",
559 => x"8f388008",
560 => x"5f751c77",
561 => x"77317f88",
562 => x"05087831",
563 => x"70618805",
564 => x"0c5d585c",
565 => x"7a802efe",
566 => x"ae387681",
567 => x"83387408",
568 => x"84160888",
569 => x"1757585c",
570 => x"76802ef2",
571 => x"3876538a",
572 => x"527b5182",
573 => x"d33f8008",
574 => x"7c318105",
575 => x"5d800884",
576 => x"3881175d",
577 => x"815f7c59",
578 => x"767d2783",
579 => x"38765994",
580 => x"1a08881b",
581 => x"08115758",
582 => x"807a085c",
583 => x"54901a08",
584 => x"7b278338",
585 => x"81547579",
586 => x"25843873",
587 => x"ba387779",
588 => x"24fee238",
589 => x"77537b52",
590 => x"9c1a0851",
591 => x"a41a0859",
592 => x"782d8008",
593 => x"56800880",
594 => x"24fee238",
595 => x"8c1a2280",
596 => x"c0075e7d",
597 => x"8c1b23ff",
598 => x"5574800c",
599 => x"903d0d04",
600 => x"7effa338",
601 => x"ff873975",
602 => x"537b527a",
603 => x"5182f93f",
604 => x"7908167a",
605 => x"0c79518e",
606 => x"b13f8008",
607 => x"cf387c76",
608 => x"315d7cfe",
609 => x"bc38feac",
610 => x"39901a08",
611 => x"7a087131",
612 => x"78117056",
613 => x"5a575280",
614 => x"cfec0851",
615 => x"84943f80",
616 => x"08802eff",
617 => x"a7388008",
618 => x"901b0c80",
619 => x"08167a0c",
620 => x"77941b0c",
621 => x"76881b0c",
622 => x"7656fd99",
623 => x"39790858",
624 => x"901a0878",
625 => x"27833881",
626 => x"54757727",
627 => x"843873b3",
628 => x"38941a08",
629 => x"54737726",
630 => x"80d33873",
631 => x"5378529c",
632 => x"1a0851a4",
633 => x"1a085877",
634 => x"2d800856",
635 => x"80088024",
636 => x"fd83388c",
637 => x"1a2280c0",
638 => x"075e7d8c",
639 => x"1b23ff55",
640 => x"fed73975",
641 => x"53785277",
642 => x"5181dd3f",
643 => x"7908167a",
644 => x"0c79518d",
645 => x"953f8008",
646 => x"802efcd9",
647 => x"388c1a22",
648 => x"80c0075e",
649 => x"7d8c1b23",
650 => x"ff55fead",
651 => x"39767754",
652 => x"79537852",
653 => x"5681b13f",
654 => x"881a0877",
655 => x"31881b0c",
656 => x"7908177a",
657 => x"0cfcae39",
658 => x"fa3d0d7a",
659 => x"79028805",
660 => x"a7053355",
661 => x"53548374",
662 => x"2780df38",
663 => x"71830651",
664 => x"7080d738",
665 => x"71715755",
666 => x"83517582",
667 => x"802913ff",
668 => x"12525670",
669 => x"8025f338",
670 => x"837427bc",
671 => x"38740876",
672 => x"327009f7",
673 => x"fbfdff12",
674 => x"06f88482",
675 => x"81800651",
676 => x"5170802e",
677 => x"98387451",
678 => x"80527033",
679 => x"5772772e",
680 => x"b9388111",
681 => x"81135351",
682 => x"837227ee",
683 => x"38fc1484",
684 => x"16565473",
685 => x"8326c638",
686 => x"7452ff14",
687 => x"5170ff2e",
688 => x"97387133",
689 => x"5472742e",
690 => x"98388112",
691 => x"ff125252",
692 => x"70ff2e09",
693 => x"8106eb38",
694 => x"80517080",
695 => x"0c883d0d",
696 => x"0471800c",
697 => x"883d0d04",
698 => x"fa3d0d78",
699 => x"7a7c7272",
700 => x"72595755",
701 => x"58565774",
702 => x"7727b238",
703 => x"75155176",
704 => x"7127aa38",
705 => x"707618ff",
706 => x"18535353",
707 => x"70ff2e96",
708 => x"38ff12ff",
709 => x"14545272",
710 => x"337234ff",
711 => x"115170ff",
712 => x"2e098106",
713 => x"ec387680",
714 => x"0c883d0d",
715 => x"048f7627",
716 => x"80e63874",
717 => x"77078306",
718 => x"517080dc",
719 => x"38767552",
720 => x"53707084",
721 => x"05520873",
722 => x"70840555",
723 => x"0c727170",
724 => x"84055308",
725 => x"71708405",
726 => x"530c7170",
727 => x"84055308",
728 => x"71708405",
729 => x"530c7170",
730 => x"84055308",
731 => x"71708405",
732 => x"530cf015",
733 => x"5553738f",
734 => x"26c73883",
735 => x"74279538",
736 => x"70708405",
737 => x"52087370",
738 => x"8405550c",
739 => x"fc145473",
740 => x"8326ed38",
741 => x"72715452",
742 => x"ff145170",
743 => x"ff2eff86",
744 => x"38727081",
745 => x"05543372",
746 => x"70810554",
747 => x"34ff1151",
748 => x"ea39ef3d",
749 => x"0d636567",
750 => x"405d427b",
751 => x"802e8582",
752 => x"386151a9",
753 => x"e73ff81c",
754 => x"70841208",
755 => x"70fc0670",
756 => x"628b0570",
757 => x"f8064159",
758 => x"455c5f41",
759 => x"57967427",
760 => x"82c53880",
761 => x"7b247e7c",
762 => x"26075880",
763 => x"5477742e",
764 => x"09810682",
765 => x"ab38787b",
766 => x"2581fe38",
767 => x"781780d7",
768 => x"a80b8805",
769 => x"085b5679",
770 => x"762e84c5",
771 => x"38841608",
772 => x"70fe0617",
773 => x"84110881",
774 => x"06415555",
775 => x"7e828d38",
776 => x"74fc0658",
777 => x"79762e84",
778 => x"e3387818",
779 => x"5f7e7b25",
780 => x"81ff387c",
781 => x"81065473",
782 => x"82c13876",
783 => x"77083184",
784 => x"1108fc06",
785 => x"56577580",
786 => x"2e913879",
787 => x"762e84f0",
788 => x"38741819",
789 => x"58777b25",
790 => x"84913876",
791 => x"802e829b",
792 => x"38781556",
793 => x"7a762482",
794 => x"92388c17",
795 => x"08881808",
796 => x"718c120c",
797 => x"88120c5e",
798 => x"75598817",
799 => x"61fc055b",
800 => x"5679a426",
801 => x"85ff387b",
802 => x"76595593",
803 => x"7a2780c9",
804 => x"387b7084",
805 => x"055d087c",
806 => x"56760c74",
807 => x"70840556",
808 => x"088c180c",
809 => x"9017589b",
810 => x"7a27ae38",
811 => x"74708405",
812 => x"5608780c",
813 => x"74708405",
814 => x"56089418",
815 => x"0c981758",
816 => x"a37a2795",
817 => x"38747084",
818 => x"05560878",
819 => x"0c747084",
820 => x"0556089c",
821 => x"180ca017",
822 => x"58747084",
823 => x"05560875",
824 => x"5f787084",
825 => x"055a0c77",
826 => x"7e708405",
827 => x"40087170",
828 => x"8405530c",
829 => x"7e08710c",
830 => x"5d787b31",
831 => x"56758f26",
832 => x"80c93884",
833 => x"17088106",
834 => x"79078418",
835 => x"0c781784",
836 => x"11088107",
837 => x"84120c5b",
838 => x"6151a791",
839 => x"3f881754",
840 => x"73800c93",
841 => x"3d0d0490",
842 => x"5bfdb839",
843 => x"7756fe83",
844 => x"398c1608",
845 => x"88170871",
846 => x"8c120c88",
847 => x"120c587e",
848 => x"707c3157",
849 => x"598f7627",
850 => x"ffb9387a",
851 => x"17841808",
852 => x"81067c07",
853 => x"84190c76",
854 => x"81078412",
855 => x"0c761184",
856 => x"11088107",
857 => x"84120c5b",
858 => x"88055261",
859 => x"518fda3f",
860 => x"6151a6b9",
861 => x"3f881754",
862 => x"ffa6397d",
863 => x"52615197",
864 => x"d73f8008",
865 => x"5a800880",
866 => x"2e81ab38",
867 => x"8008f805",
868 => x"60840508",
869 => x"fe066105",
870 => x"58557477",
871 => x"2e83f238",
872 => x"fc195877",
873 => x"a42681b0",
874 => x"387b8008",
875 => x"56579378",
876 => x"2780dc38",
877 => x"7b707084",
878 => x"05520880",
879 => x"08708405",
880 => x"800c0c80",
881 => x"08717084",
882 => x"0553085d",
883 => x"567b7670",
884 => x"8405580c",
885 => x"579b7827",
886 => x"b6387670",
887 => x"84055808",
888 => x"75708405",
889 => x"570c7670",
890 => x"84055808",
891 => x"75708405",
892 => x"570ca378",
893 => x"27993876",
894 => x"70840558",
895 => x"08757084",
896 => x"05570c76",
897 => x"70840558",
898 => x"08757084",
899 => x"05570c76",
900 => x"70840558",
901 => x"08775e75",
902 => x"70840557",
903 => x"0c747d70",
904 => x"84055f08",
905 => x"71708405",
906 => x"530c7d08",
907 => x"710c5f7b",
908 => x"5261518e",
909 => x"943f6151",
910 => x"a4f33f79",
911 => x"800c933d",
912 => x"0d047d52",
913 => x"61519690",
914 => x"3f800880",
915 => x"0c933d0d",
916 => x"04841608",
917 => x"55fbc939",
918 => x"77537b52",
919 => x"800851a2",
920 => x"a53f7b52",
921 => x"61518de1",
922 => x"3fcc398c",
923 => x"16088817",
924 => x"08718c12",
925 => x"0c88120c",
926 => x"5d8c1708",
927 => x"88180871",
928 => x"8c120c88",
929 => x"120c5977",
930 => x"59fbef39",
931 => x"7818901c",
932 => x"40557e75",
933 => x"24fb9c38",
934 => x"7a177080",
935 => x"d7a80b88",
936 => x"050c757c",
937 => x"31810784",
938 => x"120c5684",
939 => x"17088106",
940 => x"7b078418",
941 => x"0c6151a3",
942 => x"f43f8817",
943 => x"54fce139",
944 => x"74181990",
945 => x"1c5e5a7c",
946 => x"7a24fb8f",
947 => x"388c1708",
948 => x"88180871",
949 => x"8c120c88",
950 => x"120c5e88",
951 => x"1761fc05",
952 => x"575975a4",
953 => x"2681b638",
954 => x"7b795955",
955 => x"93762780",
956 => x"c9387b70",
957 => x"84055d08",
958 => x"7c56790c",
959 => x"74708405",
960 => x"56088c18",
961 => x"0c901758",
962 => x"9b7627ae",
963 => x"38747084",
964 => x"05560878",
965 => x"0c747084",
966 => x"05560894",
967 => x"180c9817",
968 => x"58a37627",
969 => x"95387470",
970 => x"84055608",
971 => x"780c7470",
972 => x"84055608",
973 => x"9c180ca0",
974 => x"17587470",
975 => x"84055608",
976 => x"75417870",
977 => x"84055a0c",
978 => x"77607084",
979 => x"05420871",
980 => x"70840553",
981 => x"0c600871",
982 => x"0c5e7a17",
983 => x"7080d7a8",
984 => x"0b88050c",
985 => x"7a7c3181",
986 => x"0784120c",
987 => x"58841708",
988 => x"81067b07",
989 => x"84180c61",
990 => x"51a2b23f",
991 => x"78547380",
992 => x"0c933d0d",
993 => x"0479537b",
994 => x"5275519f",
995 => x"f93ffae9",
996 => x"39841508",
997 => x"fc061960",
998 => x"5859fadd",
999 => x"3975537b",
1000 => x"5278519f",
1001 => x"e13f7a17",
1002 => x"7080d7a8",
1003 => x"0b88050c",
1004 => x"7a7c3181",
1005 => x"0784120c",
1006 => x"58841708",
1007 => x"81067b07",
1008 => x"84180c61",
1009 => x"51a1e63f",
1010 => x"7854ffb2",
1011 => x"39fa3d0d",
1012 => x"7880cfec",
1013 => x"085455b8",
1014 => x"1308802e",
1015 => x"81af388c",
1016 => x"15227083",
1017 => x"ffff0670",
1018 => x"832a8132",
1019 => x"81065555",
1020 => x"5672802e",
1021 => x"80da3873",
1022 => x"842a8132",
1023 => x"810657ff",
1024 => x"537680f2",
1025 => x"3873822a",
1026 => x"81065473",
1027 => x"802eb938",
1028 => x"b0150854",
1029 => x"73802e9c",
1030 => x"3880c015",
1031 => x"5373732e",
1032 => x"8f387352",
1033 => x"80cfec08",
1034 => x"518a9e3f",
1035 => x"8c152256",
1036 => x"76b0160c",
1037 => x"75db0657",
1038 => x"768c1623",
1039 => x"800b8416",
1040 => x"0c901508",
1041 => x"750c7656",
1042 => x"75880754",
1043 => x"738c1623",
1044 => x"90150880",
1045 => x"2ebf388c",
1046 => x"15227081",
1047 => x"06555373",
1048 => x"9c38720a",
1049 => x"100a8106",
1050 => x"56758538",
1051 => x"94150854",
1052 => x"7388160c",
1053 => x"80537280",
1054 => x"0c883d0d",
1055 => x"04800b88",
1056 => x"160c9415",
1057 => x"08309816",
1058 => x"0c8053ea",
1059 => x"39725182",
1060 => x"a63ffecb",
1061 => x"3974518f",
1062 => x"bc3f8c15",
1063 => x"22708106",
1064 => x"55537380",
1065 => x"2effbb38",
1066 => x"d439f83d",
1067 => x"0d7a5776",
1068 => x"802e8197",
1069 => x"3880cfec",
1070 => x"0854b814",
1071 => x"08802e80",
1072 => x"eb388c17",
1073 => x"2270902b",
1074 => x"70902c70",
1075 => x"832a8132",
1076 => x"81065b5b",
1077 => x"57557780",
1078 => x"cb389017",
1079 => x"08567580",
1080 => x"2e80c138",
1081 => x"76087631",
1082 => x"76780c79",
1083 => x"83065555",
1084 => x"73853894",
1085 => x"17085877",
1086 => x"88180c80",
1087 => x"7525a538",
1088 => x"74537552",
1089 => x"9c170851",
1090 => x"a4170854",
1091 => x"732d800b",
1092 => x"80082580",
1093 => x"c9388008",
1094 => x"16758008",
1095 => x"31565674",
1096 => x"8024dd38",
1097 => x"800b800c",
1098 => x"8a3d0d04",
1099 => x"73518187",
1100 => x"3f8c1722",
1101 => x"70902b70",
1102 => x"902c7083",
1103 => x"2a813281",
1104 => x"065b5b57",
1105 => x"5577dd38",
1106 => x"ff9039a1",
1107 => x"aa5280cf",
1108 => x"ec08518c",
1109 => x"d03f8008",
1110 => x"800c8a3d",
1111 => x"0d048c17",
1112 => x"2280c007",
1113 => x"58778c18",
1114 => x"23ff0b80",
1115 => x"0c8a3d0d",
1116 => x"04fa3d0d",
1117 => x"797080dc",
1118 => x"298c1154",
1119 => x"7a535657",
1120 => x"8fd63f80",
1121 => x"08800855",
1122 => x"56800880",
1123 => x"2ea23880",
1124 => x"088c0554",
1125 => x"800b8008",
1126 => x"0c768008",
1127 => x"84050c73",
1128 => x"80088805",
1129 => x"0c745380",
1130 => x"5273519c",
1131 => x"f53f7554",
1132 => x"73800c88",
1133 => x"3d0d0470",
1134 => x"707074a8",
1135 => x"f60bbc12",
1136 => x"0c53810b",
1137 => x"b8140c80",
1138 => x"0b84dc14",
1139 => x"0c830b84",
1140 => x"e0140c84",
1141 => x"e81384e4",
1142 => x"140c8413",
1143 => x"08518070",
1144 => x"720c7084",
1145 => x"130c7088",
1146 => x"130c5284",
1147 => x"0b8c1223",
1148 => x"718e1223",
1149 => x"7190120c",
1150 => x"7194120c",
1151 => x"7198120c",
1152 => x"709c120c",
1153 => x"80c1e50b",
1154 => x"a0120c80",
1155 => x"c2b10ba4",
1156 => x"120c80c3",
1157 => x"ad0ba812",
1158 => x"0c80c3fe",
1159 => x"0bac120c",
1160 => x"88130872",
1161 => x"710c7284",
1162 => x"120c7288",
1163 => x"120c5189",
1164 => x"0b8c1223",
1165 => x"810b8e12",
1166 => x"23719012",
1167 => x"0c719412",
1168 => x"0c719812",
1169 => x"0c709c12",
1170 => x"0c80c1e5",
1171 => x"0ba0120c",
1172 => x"80c2b10b",
1173 => x"a4120c80",
1174 => x"c3ad0ba8",
1175 => x"120c80c3",
1176 => x"fe0bac12",
1177 => x"0c8c1308",
1178 => x"72710c72",
1179 => x"84120c72",
1180 => x"88120c51",
1181 => x"8a0b8c12",
1182 => x"23820b8e",
1183 => x"12237190",
1184 => x"120c7194",
1185 => x"120c7198",
1186 => x"120c709c",
1187 => x"120c80c1",
1188 => x"e50ba012",
1189 => x"0c80c2b1",
1190 => x"0ba4120c",
1191 => x"80c3ad0b",
1192 => x"a8120c80",
1193 => x"c3fe0bac",
1194 => x"120c5050",
1195 => x"5004f83d",
1196 => x"0d7a80cf",
1197 => x"ec08b811",
1198 => x"08575758",
1199 => x"7481ec38",
1200 => x"a8f60bbc",
1201 => x"170c810b",
1202 => x"b8170c74",
1203 => x"84dc170c",
1204 => x"830b84e0",
1205 => x"170c84e8",
1206 => x"1684e417",
1207 => x"0c841608",
1208 => x"75710c75",
1209 => x"84120c75",
1210 => x"88120c59",
1211 => x"840b8c1a",
1212 => x"23748e1a",
1213 => x"2374901a",
1214 => x"0c74941a",
1215 => x"0c74981a",
1216 => x"0c789c1a",
1217 => x"0c80c1e5",
1218 => x"0ba01a0c",
1219 => x"80c2b10b",
1220 => x"a41a0c80",
1221 => x"c3ad0ba8",
1222 => x"1a0c80c3",
1223 => x"fe0bac1a",
1224 => x"0c881608",
1225 => x"75710c75",
1226 => x"84120c75",
1227 => x"88120c57",
1228 => x"890b8c18",
1229 => x"23810b8e",
1230 => x"18237490",
1231 => x"180c7494",
1232 => x"180c7498",
1233 => x"180c769c",
1234 => x"180c80c1",
1235 => x"e50ba018",
1236 => x"0c80c2b1",
1237 => x"0ba4180c",
1238 => x"80c3ad0b",
1239 => x"a8180c80",
1240 => x"c3fe0bac",
1241 => x"180c8c16",
1242 => x"0875710c",
1243 => x"7584120c",
1244 => x"7588120c",
1245 => x"548a0b8c",
1246 => x"1523820b",
1247 => x"8e152374",
1248 => x"90150c74",
1249 => x"94150c74",
1250 => x"98150c73",
1251 => x"9c150c80",
1252 => x"c1e50ba0",
1253 => x"150c80c2",
1254 => x"b10ba415",
1255 => x"0c80c3ad",
1256 => x"0ba8150c",
1257 => x"80c3fe0b",
1258 => x"ac150c84",
1259 => x"dc168811",
1260 => x"08841208",
1261 => x"ff055757",
1262 => x"57807524",
1263 => x"9f388c16",
1264 => x"2270902b",
1265 => x"70902c51",
1266 => x"55597380",
1267 => x"2e80ed38",
1268 => x"80dc16ff",
1269 => x"16565674",
1270 => x"8025e338",
1271 => x"76085574",
1272 => x"802e8f38",
1273 => x"74881108",
1274 => x"841208ff",
1275 => x"05575757",
1276 => x"c83982fc",
1277 => x"5277518a",
1278 => x"df3f8008",
1279 => x"80085556",
1280 => x"8008802e",
1281 => x"a3388008",
1282 => x"8c057580",
1283 => x"080c5484",
1284 => x"0b800884",
1285 => x"050c7380",
1286 => x"0888050c",
1287 => x"82f05374",
1288 => x"52735197",
1289 => x"fd3f7554",
1290 => x"7374780c",
1291 => x"5573ffb4",
1292 => x"388c780c",
1293 => x"800b800c",
1294 => x"8a3d0d04",
1295 => x"810b8c17",
1296 => x"2373760c",
1297 => x"7388170c",
1298 => x"7384170c",
1299 => x"7390170c",
1300 => x"7394170c",
1301 => x"7398170c",
1302 => x"ff0b8e17",
1303 => x"2373b017",
1304 => x"0c73b417",
1305 => x"0c7380c4",
1306 => x"170c7380",
1307 => x"c8170c75",
1308 => x"800c8a3d",
1309 => x"0d047070",
1310 => x"a1aa5273",
1311 => x"5186a63f",
1312 => x"50500470",
1313 => x"70a1aa52",
1314 => x"80cfec08",
1315 => x"5186963f",
1316 => x"505004fb",
1317 => x"3d0d7770",
1318 => x"52569890",
1319 => x"3f80d7a8",
1320 => x"0b880508",
1321 => x"841108fc",
1322 => x"06707b31",
1323 => x"9fef05e0",
1324 => x"8006e080",
1325 => x"05525555",
1326 => x"a0807524",
1327 => x"94388052",
1328 => x"755197ea",
1329 => x"3f80d7b0",
1330 => x"08145372",
1331 => x"80082e8f",
1332 => x"38755197",
1333 => x"d83f8053",
1334 => x"72800c87",
1335 => x"3d0d0474",
1336 => x"30527551",
1337 => x"97c83f80",
1338 => x"08ff2ea8",
1339 => x"3880d7a8",
1340 => x"0b880508",
1341 => x"74763181",
1342 => x"0784120c",
1343 => x"5380d6ec",
1344 => x"08753180",
1345 => x"d6ec0c75",
1346 => x"5197a23f",
1347 => x"810b800c",
1348 => x"873d0d04",
1349 => x"80527551",
1350 => x"97943f80",
1351 => x"d7a80b88",
1352 => x"05088008",
1353 => x"71315454",
1354 => x"8f7325ff",
1355 => x"a4388008",
1356 => x"80d79c08",
1357 => x"3180d6ec",
1358 => x"0c728107",
1359 => x"84150c75",
1360 => x"5196ea3f",
1361 => x"8053ff90",
1362 => x"39f73d0d",
1363 => x"7b7d545a",
1364 => x"72802e82",
1365 => x"83387951",
1366 => x"96d23ff8",
1367 => x"13841108",
1368 => x"70fe0670",
1369 => x"13841108",
1370 => x"fc065c57",
1371 => x"58545780",
1372 => x"d7b00874",
1373 => x"2e82de38",
1374 => x"7784150c",
1375 => x"80738106",
1376 => x"56597479",
1377 => x"2e81d538",
1378 => x"77148411",
1379 => x"08810656",
1380 => x"5374a038",
1381 => x"77165678",
1382 => x"81e63888",
1383 => x"14085574",
1384 => x"80d7b02e",
1385 => x"82f9388c",
1386 => x"1408708c",
1387 => x"170c7588",
1388 => x"120c5875",
1389 => x"81078418",
1390 => x"0c751776",
1391 => x"710c5478",
1392 => x"81913883",
1393 => x"ff762781",
1394 => x"c8387589",
1395 => x"2a76832a",
1396 => x"54547380",
1397 => x"2ebf3875",
1398 => x"862ab805",
1399 => x"53847427",
1400 => x"b43880db",
1401 => x"14539474",
1402 => x"27ab3875",
1403 => x"8c2a80ee",
1404 => x"055380d4",
1405 => x"74279e38",
1406 => x"758f2a80",
1407 => x"f7055382",
1408 => x"d4742791",
1409 => x"3875922a",
1410 => x"80fc0553",
1411 => x"8ad47427",
1412 => x"843880fe",
1413 => x"53721010",
1414 => x"1080d7a8",
1415 => x"05881108",
1416 => x"55557375",
1417 => x"2e82bf38",
1418 => x"841408fc",
1419 => x"06597579",
1420 => x"278d3888",
1421 => x"14085473",
1422 => x"752e0981",
1423 => x"06ea388c",
1424 => x"1408708c",
1425 => x"190c7488",
1426 => x"190c7788",
1427 => x"120c5576",
1428 => x"8c150c79",
1429 => x"5194d63f",
1430 => x"8b3d0d04",
1431 => x"76087771",
1432 => x"31587605",
1433 => x"88180856",
1434 => x"567480d7",
1435 => x"b02e80e0",
1436 => x"388c1708",
1437 => x"708c170c",
1438 => x"7588120c",
1439 => x"53fe8939",
1440 => x"8814088c",
1441 => x"1508708c",
1442 => x"130c5988",
1443 => x"190cfea3",
1444 => x"3975832a",
1445 => x"70545480",
1446 => x"74248198",
1447 => x"3872822c",
1448 => x"81712b80",
1449 => x"d7ac0807",
1450 => x"80d7a80b",
1451 => x"84050c74",
1452 => x"10101080",
1453 => x"d7a80588",
1454 => x"1108718c",
1455 => x"1b0c7088",
1456 => x"1b0c7988",
1457 => x"130c565a",
1458 => x"55768c15",
1459 => x"0cff8439",
1460 => x"8159fdb4",
1461 => x"39771673",
1462 => x"81065455",
1463 => x"72983876",
1464 => x"08777131",
1465 => x"5875058c",
1466 => x"18088819",
1467 => x"08718c12",
1468 => x"0c88120c",
1469 => x"55557481",
1470 => x"0784180c",
1471 => x"7680d7a8",
1472 => x"0b88050c",
1473 => x"80d7a408",
1474 => x"7526fec7",
1475 => x"3880d7a0",
1476 => x"08527951",
1477 => x"fafd3f79",
1478 => x"5193923f",
1479 => x"feba3981",
1480 => x"778c170c",
1481 => x"7788170c",
1482 => x"758c190c",
1483 => x"7588190c",
1484 => x"59fd8039",
1485 => x"83147082",
1486 => x"2c81712b",
1487 => x"80d7ac08",
1488 => x"0780d7a8",
1489 => x"0b84050c",
1490 => x"75101010",
1491 => x"80d7a805",
1492 => x"88110871",
1493 => x"8c1c0c70",
1494 => x"881c0c7a",
1495 => x"88130c57",
1496 => x"5b5653fe",
1497 => x"e4398073",
1498 => x"24a33872",
1499 => x"822c8171",
1500 => x"2b80d7ac",
1501 => x"080780d7",
1502 => x"a80b8405",
1503 => x"0c58748c",
1504 => x"180c7388",
1505 => x"180c7688",
1506 => x"160cfdc3",
1507 => x"39831370",
1508 => x"822c8171",
1509 => x"2b80d7ac",
1510 => x"080780d7",
1511 => x"a80b8405",
1512 => x"0c5953da",
1513 => x"39f93d0d",
1514 => x"797b5853",
1515 => x"800b80cf",
1516 => x"ec085356",
1517 => x"72722ebc",
1518 => x"3884dc13",
1519 => x"5574762e",
1520 => x"b3388815",
1521 => x"08841608",
1522 => x"ff055454",
1523 => x"80732499",
1524 => x"388c1422",
1525 => x"70902b53",
1526 => x"587180d4",
1527 => x"3880dc14",
1528 => x"ff145454",
1529 => x"728025e9",
1530 => x"38740855",
1531 => x"74d43880",
1532 => x"cfec0852",
1533 => x"84dc1255",
1534 => x"74802ead",
1535 => x"38881508",
1536 => x"841608ff",
1537 => x"05545480",
1538 => x"73249838",
1539 => x"8c142270",
1540 => x"902b5358",
1541 => x"71ad3880",
1542 => x"dc14ff14",
1543 => x"54547280",
1544 => x"25ea3874",
1545 => x"085574d5",
1546 => x"3875800c",
1547 => x"893d0d04",
1548 => x"7351762d",
1549 => x"75800807",
1550 => x"80dc15ff",
1551 => x"15555556",
1552 => x"ffa23973",
1553 => x"51762d75",
1554 => x"80080780",
1555 => x"dc15ff15",
1556 => x"555556ca",
1557 => x"39ea3d0d",
1558 => x"688c1122",
1559 => x"700a100a",
1560 => x"81065758",
1561 => x"567480e4",
1562 => x"388e1622",
1563 => x"70902b70",
1564 => x"902c5155",
1565 => x"58807424",
1566 => x"b138983d",
1567 => x"c4055373",
1568 => x"5280cfec",
1569 => x"08519481",
1570 => x"3f800b80",
1571 => x"08249738",
1572 => x"7983e080",
1573 => x"06547380",
1574 => x"c0802e81",
1575 => x"8f387382",
1576 => x"80802e81",
1577 => x"91388c16",
1578 => x"22577690",
1579 => x"80075473",
1580 => x"8c172388",
1581 => x"805280cf",
1582 => x"ec085181",
1583 => x"9b3f8008",
1584 => x"9d388c16",
1585 => x"22820755",
1586 => x"748c1723",
1587 => x"80c31670",
1588 => x"770c9017",
1589 => x"0c810b94",
1590 => x"170c983d",
1591 => x"0d0480cf",
1592 => x"ec08a8f6",
1593 => x"0bbc120c",
1594 => x"588c1622",
1595 => x"81800754",
1596 => x"738c1723",
1597 => x"8008760c",
1598 => x"80089017",
1599 => x"0c88800b",
1600 => x"94170c74",
1601 => x"802ed338",
1602 => x"8e162270",
1603 => x"902b7090",
1604 => x"2c535654",
1605 => x"9afb3f80",
1606 => x"08802eff",
1607 => x"bd388c16",
1608 => x"22810757",
1609 => x"768c1723",
1610 => x"983d0d04",
1611 => x"810b8c17",
1612 => x"225855fe",
1613 => x"f539a816",
1614 => x"0880c3ad",
1615 => x"2e098106",
1616 => x"fee4388c",
1617 => x"16228880",
1618 => x"0754738c",
1619 => x"17238880",
1620 => x"0b80cc17",
1621 => x"0cfedc39",
1622 => x"f43d0d7e",
1623 => x"608b1170",
1624 => x"f8065b55",
1625 => x"555d7296",
1626 => x"26833890",
1627 => x"58807824",
1628 => x"74792607",
1629 => x"55805474",
1630 => x"742e0981",
1631 => x"0680ca38",
1632 => x"7c518ea8",
1633 => x"3f7783f7",
1634 => x"2680c538",
1635 => x"77832a70",
1636 => x"10101080",
1637 => x"d7a8058c",
1638 => x"11085858",
1639 => x"5475772e",
1640 => x"81f03884",
1641 => x"1608fc06",
1642 => x"8c170888",
1643 => x"1808718c",
1644 => x"120c8812",
1645 => x"0c5b7605",
1646 => x"84110881",
1647 => x"0784120c",
1648 => x"537c518d",
1649 => x"e83f8816",
1650 => x"5473800c",
1651 => x"8e3d0d04",
1652 => x"77892a78",
1653 => x"832a5854",
1654 => x"73802ebf",
1655 => x"3877862a",
1656 => x"b8055784",
1657 => x"7427b438",
1658 => x"80db1457",
1659 => x"947427ab",
1660 => x"38778c2a",
1661 => x"80ee0557",
1662 => x"80d47427",
1663 => x"9e38778f",
1664 => x"2a80f705",
1665 => x"5782d474",
1666 => x"27913877",
1667 => x"922a80fc",
1668 => x"05578ad4",
1669 => x"74278438",
1670 => x"80fe5776",
1671 => x"10101080",
1672 => x"d7a8058c",
1673 => x"11085653",
1674 => x"74732ea3",
1675 => x"38841508",
1676 => x"fc067079",
1677 => x"31555673",
1678 => x"8f2488e4",
1679 => x"38738025",
1680 => x"88e6388c",
1681 => x"15085574",
1682 => x"732e0981",
1683 => x"06df3881",
1684 => x"175980d7",
1685 => x"b8085675",
1686 => x"80d7b02e",
1687 => x"82cc3884",
1688 => x"1608fc06",
1689 => x"70793155",
1690 => x"55738f24",
1691 => x"bb3880d7",
1692 => x"b00b80d7",
1693 => x"bc0c80d7",
1694 => x"b00b80d7",
1695 => x"b80c8074",
1696 => x"2480db38",
1697 => x"74168411",
1698 => x"08810784",
1699 => x"120c53fe",
1700 => x"b0398816",
1701 => x"8c110857",
1702 => x"5975792e",
1703 => x"098106fe",
1704 => x"82388214",
1705 => x"59ffab39",
1706 => x"77167881",
1707 => x"0784180c",
1708 => x"7080d7bc",
1709 => x"0c7080d7",
1710 => x"b80c80d7",
1711 => x"b00b8c12",
1712 => x"0c8c1108",
1713 => x"88120c74",
1714 => x"81078412",
1715 => x"0c740574",
1716 => x"710c5b7c",
1717 => x"518bd63f",
1718 => x"881654fd",
1719 => x"ec3983ff",
1720 => x"75278391",
1721 => x"3874892a",
1722 => x"75832a54",
1723 => x"5473802e",
1724 => x"bf387486",
1725 => x"2ab80553",
1726 => x"847427b4",
1727 => x"3880db14",
1728 => x"53947427",
1729 => x"ab38748c",
1730 => x"2a80ee05",
1731 => x"5380d474",
1732 => x"279e3874",
1733 => x"8f2a80f7",
1734 => x"055382d4",
1735 => x"74279138",
1736 => x"74922a80",
1737 => x"fc05538a",
1738 => x"d4742784",
1739 => x"3880fe53",
1740 => x"72101010",
1741 => x"80d7a805",
1742 => x"88110855",
1743 => x"5773772e",
1744 => x"868b3884",
1745 => x"1408fc06",
1746 => x"5b747b27",
1747 => x"8d388814",
1748 => x"08547377",
1749 => x"2e098106",
1750 => x"ea388c14",
1751 => x"0880d7a8",
1752 => x"0b840508",
1753 => x"718c190c",
1754 => x"7588190c",
1755 => x"7788130c",
1756 => x"5c57758c",
1757 => x"150c7853",
1758 => x"80792483",
1759 => x"98387282",
1760 => x"2c81712b",
1761 => x"5656747b",
1762 => x"2680ca38",
1763 => x"7a750657",
1764 => x"7682a338",
1765 => x"78fc0684",
1766 => x"05597410",
1767 => x"707c0655",
1768 => x"55738292",
1769 => x"38841959",
1770 => x"f13980d7",
1771 => x"a80b8405",
1772 => x"0879545b",
1773 => x"788025c6",
1774 => x"3882da39",
1775 => x"74097b06",
1776 => x"7080d7a8",
1777 => x"0b84050c",
1778 => x"5b741055",
1779 => x"747b2685",
1780 => x"387485bc",
1781 => x"3880d7a8",
1782 => x"0b880508",
1783 => x"70841208",
1784 => x"fc06707b",
1785 => x"317b7226",
1786 => x"8f722507",
1787 => x"5d575c5c",
1788 => x"5578802e",
1789 => x"80d93879",
1790 => x"1580d7a0",
1791 => x"08199011",
1792 => x"59545680",
1793 => x"d79c08ff",
1794 => x"2e8838a0",
1795 => x"8f13e080",
1796 => x"06577652",
1797 => x"7c518996",
1798 => x"3f800854",
1799 => x"8008ff2e",
1800 => x"90388008",
1801 => x"762782a7",
1802 => x"387480d7",
1803 => x"a82e829f",
1804 => x"3880d7a8",
1805 => x"0b880508",
1806 => x"55841508",
1807 => x"fc067079",
1808 => x"31797226",
1809 => x"8f722507",
1810 => x"5d555a7a",
1811 => x"83f23877",
1812 => x"81078416",
1813 => x"0c771570",
1814 => x"80d7a80b",
1815 => x"88050c74",
1816 => x"81078412",
1817 => x"0c567c51",
1818 => x"88c33f88",
1819 => x"15547380",
1820 => x"0c8e3d0d",
1821 => x"0474832a",
1822 => x"70545480",
1823 => x"7424819b",
1824 => x"3872822c",
1825 => x"81712b80",
1826 => x"d7ac0807",
1827 => x"7080d7a8",
1828 => x"0b84050c",
1829 => x"75101010",
1830 => x"80d7a805",
1831 => x"88110871",
1832 => x"8c1b0c70",
1833 => x"881b0c79",
1834 => x"88130c57",
1835 => x"555c5575",
1836 => x"8c150cfd",
1837 => x"c1397879",
1838 => x"10101080",
1839 => x"d7a80570",
1840 => x"565b5c8c",
1841 => x"14085675",
1842 => x"742ea338",
1843 => x"841608fc",
1844 => x"06707931",
1845 => x"5853768f",
1846 => x"2483f138",
1847 => x"76802584",
1848 => x"af388c16",
1849 => x"08567574",
1850 => x"2e098106",
1851 => x"df388814",
1852 => x"811a7083",
1853 => x"06555a54",
1854 => x"72c9387b",
1855 => x"83065675",
1856 => x"802efdb8",
1857 => x"38ff1cf8",
1858 => x"1b5b5c88",
1859 => x"1a087a2e",
1860 => x"ea38fdb5",
1861 => x"39831953",
1862 => x"fce43983",
1863 => x"1470822c",
1864 => x"81712b80",
1865 => x"d7ac0807",
1866 => x"7080d7a8",
1867 => x"0b84050c",
1868 => x"76101010",
1869 => x"80d7a805",
1870 => x"88110871",
1871 => x"8c1c0c70",
1872 => x"881c0c7a",
1873 => x"88130c58",
1874 => x"535d5653",
1875 => x"fee13980",
1876 => x"d6ec0817",
1877 => x"59800876",
1878 => x"2e818b38",
1879 => x"80d79c08",
1880 => x"ff2e848e",
1881 => x"38737631",
1882 => x"1980d6ec",
1883 => x"0c738706",
1884 => x"70565372",
1885 => x"802e8838",
1886 => x"88733170",
1887 => x"15555576",
1888 => x"149fff06",
1889 => x"a0807131",
1890 => x"1670547e",
1891 => x"53515386",
1892 => x"9d3f8008",
1893 => x"568008ff",
1894 => x"2e819e38",
1895 => x"80d6ec08",
1896 => x"137080d6",
1897 => x"ec0c7475",
1898 => x"80d7a80b",
1899 => x"88050c77",
1900 => x"76311581",
1901 => x"07555659",
1902 => x"7a80d7a8",
1903 => x"2e83c038",
1904 => x"798f2682",
1905 => x"ef38810b",
1906 => x"84150c84",
1907 => x"1508fc06",
1908 => x"70793179",
1909 => x"72268f72",
1910 => x"25075d55",
1911 => x"5a7a802e",
1912 => x"fced3880",
1913 => x"db398008",
1914 => x"9fff0655",
1915 => x"74feed38",
1916 => x"7880d6ec",
1917 => x"0c80d7a8",
1918 => x"0b880508",
1919 => x"7a188107",
1920 => x"84120c55",
1921 => x"80d79808",
1922 => x"79278638",
1923 => x"7880d798",
1924 => x"0c80d794",
1925 => x"087927fc",
1926 => x"a0387880",
1927 => x"d7940c84",
1928 => x"1508fc06",
1929 => x"70793179",
1930 => x"72268f72",
1931 => x"25075d55",
1932 => x"5a7a802e",
1933 => x"fc993888",
1934 => x"39807457",
1935 => x"53fedd39",
1936 => x"7c5184e9",
1937 => x"3f800b80",
1938 => x"0c8e3d0d",
1939 => x"04807324",
1940 => x"a5387282",
1941 => x"2c81712b",
1942 => x"80d7ac08",
1943 => x"077080d7",
1944 => x"a80b8405",
1945 => x"0c5c5a76",
1946 => x"8c170c73",
1947 => x"88170c75",
1948 => x"88180cf9",
1949 => x"fd398313",
1950 => x"70822c81",
1951 => x"712b80d7",
1952 => x"ac080770",
1953 => x"80d7a80b",
1954 => x"84050c5d",
1955 => x"5b53d839",
1956 => x"7a75065c",
1957 => x"7bfc9f38",
1958 => x"84197510",
1959 => x"5659f139",
1960 => x"ff178105",
1961 => x"59f7ab39",
1962 => x"8c150888",
1963 => x"1608718c",
1964 => x"120c8812",
1965 => x"0c597515",
1966 => x"84110881",
1967 => x"0784120c",
1968 => x"587c5183",
1969 => x"e83f8815",
1970 => x"54fba339",
1971 => x"77167881",
1972 => x"0784180c",
1973 => x"8c170888",
1974 => x"1808718c",
1975 => x"120c8812",
1976 => x"0c5c7080",
1977 => x"d7bc0c70",
1978 => x"80d7b80c",
1979 => x"80d7b00b",
1980 => x"8c120c8c",
1981 => x"11088812",
1982 => x"0c778107",
1983 => x"84120c77",
1984 => x"0577710c",
1985 => x"557c5183",
1986 => x"a43f8816",
1987 => x"54f5ba39",
1988 => x"72168411",
1989 => x"08810784",
1990 => x"120c588c",
1991 => x"16088817",
1992 => x"08718c12",
1993 => x"0c88120c",
1994 => x"577c5183",
1995 => x"803f8816",
1996 => x"54f59639",
1997 => x"7284150c",
1998 => x"f41af806",
1999 => x"70841d08",
2000 => x"81060784",
2001 => x"1d0c701c",
2002 => x"5556850b",
2003 => x"84150c85",
2004 => x"0b88150c",
2005 => x"8f7627fd",
2006 => x"ab38881b",
2007 => x"527c51eb",
2008 => x"e83f80d7",
2009 => x"a80b8805",
2010 => x"0880d6ec",
2011 => x"085a55fd",
2012 => x"93397880",
2013 => x"d6ec0c73",
2014 => x"80d79c0c",
2015 => x"fbef3972",
2016 => x"84150cfc",
2017 => x"ff39fb3d",
2018 => x"0d77707a",
2019 => x"7c585553",
2020 => x"568f7527",
2021 => x"80e63872",
2022 => x"76078306",
2023 => x"517080dc",
2024 => x"38757352",
2025 => x"54707084",
2026 => x"05520874",
2027 => x"70840556",
2028 => x"0c737170",
2029 => x"84055308",
2030 => x"71708405",
2031 => x"530c7170",
2032 => x"84055308",
2033 => x"71708405",
2034 => x"530c7170",
2035 => x"84055308",
2036 => x"71708405",
2037 => x"530cf016",
2038 => x"5654748f",
2039 => x"26c73883",
2040 => x"75279538",
2041 => x"70708405",
2042 => x"52087470",
2043 => x"8405560c",
2044 => x"fc155574",
2045 => x"8326ed38",
2046 => x"73715452",
2047 => x"ff155170",
2048 => x"ff2e9838",
2049 => x"72708105",
2050 => x"54337270",
2051 => x"81055434",
2052 => x"ff115170",
2053 => x"ff2e0981",
2054 => x"06ea3875",
2055 => x"800c873d",
2056 => x"0d04fb3d",
2057 => x"0d777a71",
2058 => x"028c05a3",
2059 => x"05335854",
2060 => x"54568373",
2061 => x"2780d438",
2062 => x"75830651",
2063 => x"7080cc38",
2064 => x"74882b75",
2065 => x"07707190",
2066 => x"2b075551",
2067 => x"8f7327a7",
2068 => x"38737270",
2069 => x"8405540c",
2070 => x"71747170",
2071 => x"8405530c",
2072 => x"74717084",
2073 => x"05530c74",
2074 => x"71708405",
2075 => x"530cf014",
2076 => x"5452728f",
2077 => x"26db3883",
2078 => x"73279038",
2079 => x"73727084",
2080 => x"05540cfc",
2081 => x"13537283",
2082 => x"26f238ff",
2083 => x"135170ff",
2084 => x"2e933874",
2085 => x"72708105",
2086 => x"5434ff11",
2087 => x"5170ff2e",
2088 => x"098106ef",
2089 => x"3875800c",
2090 => x"873d0d04",
2091 => x"04047070",
2092 => x"7070800b",
2093 => x"80dfe40c",
2094 => x"765184f3",
2095 => x"3f800853",
2096 => x"8008ff2e",
2097 => x"89387280",
2098 => x"0c505050",
2099 => x"500480df",
2100 => x"e4085473",
2101 => x"802eef38",
2102 => x"7574710c",
2103 => x"5272800c",
2104 => x"50505050",
2105 => x"04f93d0d",
2106 => x"797c557b",
2107 => x"548e1122",
2108 => x"70902b70",
2109 => x"902c5557",
2110 => x"80cfec08",
2111 => x"53585683",
2112 => x"f63f8008",
2113 => x"57800b80",
2114 => x"08249338",
2115 => x"80d01608",
2116 => x"80080580",
2117 => x"d0170c76",
2118 => x"800c893d",
2119 => x"0d048c16",
2120 => x"2283dfff",
2121 => x"0655748c",
2122 => x"17237680",
2123 => x"0c893d0d",
2124 => x"04fa3d0d",
2125 => x"788c1122",
2126 => x"70882a70",
2127 => x"81065157",
2128 => x"585674a9",
2129 => x"388c1622",
2130 => x"83dfff06",
2131 => x"55748c17",
2132 => x"237a5479",
2133 => x"538e1622",
2134 => x"70902b70",
2135 => x"902c5456",
2136 => x"80cfec08",
2137 => x"525681b2",
2138 => x"3f883d0d",
2139 => x"04825480",
2140 => x"538e1622",
2141 => x"70902b70",
2142 => x"902c5456",
2143 => x"80cfec08",
2144 => x"525782bb",
2145 => x"3f8c1622",
2146 => x"83dfff06",
2147 => x"55748c17",
2148 => x"237a5479",
2149 => x"538e1622",
2150 => x"70902b70",
2151 => x"902c5456",
2152 => x"80cfec08",
2153 => x"525680f2",
2154 => x"3f883d0d",
2155 => x"04f93d0d",
2156 => x"797c557b",
2157 => x"548e1122",
2158 => x"70902b70",
2159 => x"902c5557",
2160 => x"80cfec08",
2161 => x"53585681",
2162 => x"f63f8008",
2163 => x"578008ff",
2164 => x"2e99388c",
2165 => x"1622a080",
2166 => x"0755748c",
2167 => x"17238008",
2168 => x"80d0170c",
2169 => x"76800c89",
2170 => x"3d0d048c",
2171 => x"162283df",
2172 => x"ff065574",
2173 => x"8c172376",
2174 => x"800c893d",
2175 => x"0d047070",
2176 => x"70748e11",
2177 => x"2270902b",
2178 => x"70902c55",
2179 => x"51515380",
2180 => x"cfec0851",
2181 => x"bd3f5050",
2182 => x"5004fb3d",
2183 => x"0d800b80",
2184 => x"dfe40c7a",
2185 => x"53795278",
2186 => x"5182fc3f",
2187 => x"80085580",
2188 => x"08ff2e88",
2189 => x"3874800c",
2190 => x"873d0d04",
2191 => x"80dfe408",
2192 => x"5675802e",
2193 => x"f0387776",
2194 => x"710c5474",
2195 => x"800c873d",
2196 => x"0d047070",
2197 => x"7070800b",
2198 => x"80dfe40c",
2199 => x"765184c9",
2200 => x"3f800853",
2201 => x"8008ff2e",
2202 => x"89387280",
2203 => x"0c505050",
2204 => x"500480df",
2205 => x"e4085473",
2206 => x"802eef38",
2207 => x"7574710c",
2208 => x"5272800c",
2209 => x"50505050",
2210 => x"04fc3d0d",
2211 => x"800b80df",
2212 => x"e40c7852",
2213 => x"775187b0",
2214 => x"3f800854",
2215 => x"8008ff2e",
2216 => x"88387380",
2217 => x"0c863d0d",
2218 => x"0480dfe4",
2219 => x"08557480",
2220 => x"2ef03876",
2221 => x"75710c53",
2222 => x"73800c86",
2223 => x"3d0d04fb",
2224 => x"3d0d800b",
2225 => x"80dfe40c",
2226 => x"7a537952",
2227 => x"7851848b",
2228 => x"3f800855",
2229 => x"8008ff2e",
2230 => x"88387480",
2231 => x"0c873d0d",
2232 => x"0480dfe4",
2233 => x"08567580",
2234 => x"2ef03877",
2235 => x"76710c54",
2236 => x"74800c87",
2237 => x"3d0d04fb",
2238 => x"3d0d800b",
2239 => x"80dfe40c",
2240 => x"7a537952",
2241 => x"78518293",
2242 => x"3f800855",
2243 => x"8008ff2e",
2244 => x"88387480",
2245 => x"0c873d0d",
2246 => x"0480dfe4",
2247 => x"08567580",
2248 => x"2ef03877",
2249 => x"76710c54",
2250 => x"74800c87",
2251 => x"3d0d0470",
2252 => x"707080df",
2253 => x"d8088938",
2254 => x"80dfe80b",
2255 => x"80dfd80c",
2256 => x"80dfd808",
2257 => x"75115252",
2258 => x"ff537087",
2259 => x"fb808026",
2260 => x"88387080",
2261 => x"dfd80c71",
2262 => x"5372800c",
2263 => x"50505004",
2264 => x"fd3d0d80",
2265 => x"0b80cfe0",
2266 => x"08545472",
2267 => x"812e9b38",
2268 => x"7380dfdc",
2269 => x"0cc2af3f",
2270 => x"c1863f80",
2271 => x"dfb05281",
2272 => x"51c3ff3f",
2273 => x"80085186",
2274 => x"bf3f7280",
2275 => x"dfdc0cc2",
2276 => x"953fc0ec",
2277 => x"3f80dfb0",
2278 => x"528151c3",
2279 => x"e53f8008",
2280 => x"5186a53f",
2281 => x"00ff39f5",
2282 => x"3d0d7e60",
2283 => x"80dfdc08",
2284 => x"705b585b",
2285 => x"5b7580c2",
2286 => x"38777a25",
2287 => x"a138771b",
2288 => x"70337081",
2289 => x"ff065858",
2290 => x"59758a2e",
2291 => x"98387681",
2292 => x"ff0651c1",
2293 => x"b03f8118",
2294 => x"58797824",
2295 => x"e1387980",
2296 => x"0c8d3d0d",
2297 => x"048d51c1",
2298 => x"9c3f7833",
2299 => x"7081ff06",
2300 => x"5257c191",
2301 => x"3f811858",
2302 => x"e0397955",
2303 => x"7a547d53",
2304 => x"85528d3d",
2305 => x"fc0551c0",
2306 => x"b93f8008",
2307 => x"5685b23f",
2308 => x"7b80080c",
2309 => x"75800c8d",
2310 => x"3d0d04f6",
2311 => x"3d0d7d7f",
2312 => x"80dfdc08",
2313 => x"705b585a",
2314 => x"5a7580c1",
2315 => x"38777925",
2316 => x"b338c0ac",
2317 => x"3f800881",
2318 => x"ff06708d",
2319 => x"32703070",
2320 => x"9f2a5151",
2321 => x"5757768a",
2322 => x"2e80c438",
2323 => x"75802ebf",
2324 => x"38771a56",
2325 => x"76763476",
2326 => x"51c0aa3f",
2327 => x"81185878",
2328 => x"7824cf38",
2329 => x"77567580",
2330 => x"0c8c3d0d",
2331 => x"04785579",
2332 => x"547c5384",
2333 => x"528c3dfc",
2334 => x"0551ffbf",
2335 => x"c53f8008",
2336 => x"5684be3f",
2337 => x"7a80080c",
2338 => x"75800c8c",
2339 => x"3d0d0477",
2340 => x"1a598a79",
2341 => x"34811858",
2342 => x"8d51ffbf",
2343 => x"e83f8a51",
2344 => x"ffbfe23f",
2345 => x"7756ffbe",
2346 => x"39fb3d0d",
2347 => x"80dfdc08",
2348 => x"70565473",
2349 => x"88387480",
2350 => x"0c873d0d",
2351 => x"04775383",
2352 => x"52873dfc",
2353 => x"0551ffbe",
2354 => x"f93f8008",
2355 => x"5483f23f",
2356 => x"7580080c",
2357 => x"73800c87",
2358 => x"3d0d04fa",
2359 => x"3d0d80df",
2360 => x"dc08802e",
2361 => x"a3387a55",
2362 => x"79547853",
2363 => x"8652883d",
2364 => x"fc0551ff",
2365 => x"becc3f80",
2366 => x"085683c5",
2367 => x"3f768008",
2368 => x"0c75800c",
2369 => x"883d0d04",
2370 => x"83b73f9d",
2371 => x"0b80080c",
2372 => x"ff0b800c",
2373 => x"883d0d04",
2374 => x"f73d0d7b",
2375 => x"7d5b59bc",
2376 => x"53805279",
2377 => x"51f5fb3f",
2378 => x"80705657",
2379 => x"98567419",
2380 => x"70337078",
2381 => x"2b790781",
2382 => x"18f81a5a",
2383 => x"58595558",
2384 => x"847524ea",
2385 => x"38767a23",
2386 => x"84195880",
2387 => x"70565798",
2388 => x"56741870",
2389 => x"3370782b",
2390 => x"79078118",
2391 => x"f81a5a58",
2392 => x"59515484",
2393 => x"7524ea38",
2394 => x"76821b23",
2395 => x"88195880",
2396 => x"70565798",
2397 => x"56741870",
2398 => x"3370782b",
2399 => x"79078118",
2400 => x"f81a5a58",
2401 => x"59515484",
2402 => x"7524ea38",
2403 => x"76841b0c",
2404 => x"8c195880",
2405 => x"70565798",
2406 => x"56741870",
2407 => x"3370782b",
2408 => x"79078118",
2409 => x"f81a5a58",
2410 => x"59515484",
2411 => x"7524ea38",
2412 => x"76881b23",
2413 => x"90195880",
2414 => x"70565798",
2415 => x"56741870",
2416 => x"3370782b",
2417 => x"79078118",
2418 => x"f81a5a58",
2419 => x"59515484",
2420 => x"7524ea38",
2421 => x"768a1b23",
2422 => x"94195880",
2423 => x"70565798",
2424 => x"56741870",
2425 => x"3370782b",
2426 => x"79078118",
2427 => x"f81a5a58",
2428 => x"59515484",
2429 => x"7524ea38",
2430 => x"768c1b23",
2431 => x"98195880",
2432 => x"70565798",
2433 => x"56741870",
2434 => x"3370782b",
2435 => x"79078118",
2436 => x"f81a5a58",
2437 => x"59515484",
2438 => x"7524ea38",
2439 => x"768e1b23",
2440 => x"9c195880",
2441 => x"705657b8",
2442 => x"56741870",
2443 => x"3370782b",
2444 => x"79078118",
2445 => x"f81a5a58",
2446 => x"595a5488",
2447 => x"7524ea38",
2448 => x"76901b0c",
2449 => x"8b3d0d04",
2450 => x"e93d0d6a",
2451 => x"80dfdc08",
2452 => x"57577593",
2453 => x"3880c080",
2454 => x"0b84180c",
2455 => x"75ac180c",
2456 => x"75800c99",
2457 => x"3d0d0489",
2458 => x"3d70556a",
2459 => x"54558a52",
2460 => x"993dffbc",
2461 => x"0551ffbb",
2462 => x"c93f8008",
2463 => x"77537552",
2464 => x"56fd953f",
2465 => x"bc3f7780",
2466 => x"080c7580",
2467 => x"0c993d0d",
2468 => x"04fc3d0d",
2469 => x"815480df",
2470 => x"dc088838",
2471 => x"73800c86",
2472 => x"3d0d0476",
2473 => x"5397b952",
2474 => x"863dfc05",
2475 => x"51ffbb92",
2476 => x"3f800854",
2477 => x"8c3f7480",
2478 => x"080c7380",
2479 => x"0c863d0d",
2480 => x"0480cfec",
2481 => x"08800c04",
2482 => x"f73d0d7b",
2483 => x"80cfec08",
2484 => x"82c81108",
2485 => x"5a545a77",
2486 => x"802e80da",
2487 => x"38818818",
2488 => x"841908ff",
2489 => x"0581712b",
2490 => x"59555980",
2491 => x"742480ea",
2492 => x"38807424",
2493 => x"b5387382",
2494 => x"2b781188",
2495 => x"05565681",
2496 => x"80190877",
2497 => x"06537280",
2498 => x"2eb63878",
2499 => x"16700853",
2500 => x"53795174",
2501 => x"0853722d",
2502 => x"ff14fc17",
2503 => x"fc177981",
2504 => x"2c5a5757",
2505 => x"54738025",
2506 => x"d6387708",
2507 => x"5877ffad",
2508 => x"3880cfec",
2509 => x"0853bc13",
2510 => x"08a53879",
2511 => x"51f8e53f",
2512 => x"74085372",
2513 => x"2dff14fc",
2514 => x"17fc1779",
2515 => x"812c5a57",
2516 => x"57547380",
2517 => x"25ffa838",
2518 => x"d1398057",
2519 => x"ff933972",
2520 => x"51bc1308",
2521 => x"54732d79",
2522 => x"51f8b93f",
2523 => x"707080df",
2524 => x"b80bfc05",
2525 => x"70085252",
2526 => x"70ff2e91",
2527 => x"38702dfc",
2528 => x"12700852",
2529 => x"5270ff2e",
2530 => x"098106f1",
2531 => x"38505004",
2532 => x"04ffbaff",
2533 => x"3f040000",
2534 => x"00000040",
2535 => x"476f7420",
2536 => x"696e7465",
2537 => x"72727570",
2538 => x"740a0000",
2539 => x"4e6f2069",
2540 => x"6e746572",
2541 => x"72757074",
2542 => x"0a000000",
2543 => x"43000000",
2544 => x"64756d6d",
2545 => x"792e6578",
2546 => x"65000000",
2547 => x"00ffffff",
2548 => x"ff00ffff",
2549 => x"ffff00ff",
2550 => x"ffffff00",
2551 => x"00000000",
2552 => x"00000000",
2553 => x"00000000",
2554 => x"00002fc0",
2555 => x"000027f0",
2556 => x"00000000",
2557 => x"00002a58",
2558 => x"00002ab4",
2559 => x"00002b10",
2560 => x"00000000",
2561 => x"00000000",
2562 => x"00000000",
2563 => x"00000000",
2564 => x"00000000",
2565 => x"00000000",
2566 => x"00000000",
2567 => x"00000000",
2568 => x"00000000",
2569 => x"000027bc",
2570 => x"00000000",
2571 => x"00000000",
2572 => x"00000000",
2573 => x"00000000",
2574 => x"00000000",
2575 => x"00000000",
2576 => x"00000000",
2577 => x"00000000",
2578 => x"00000000",
2579 => x"00000000",
2580 => x"00000000",
2581 => x"00000000",
2582 => x"00000000",
2583 => x"00000000",
2584 => x"00000000",
2585 => x"00000000",
2586 => x"00000000",
2587 => x"00000000",
2588 => x"00000000",
2589 => x"00000000",
2590 => x"00000000",
2591 => x"00000000",
2592 => x"00000000",
2593 => x"00000000",
2594 => x"00000000",
2595 => x"00000000",
2596 => x"00000000",
2597 => x"00000000",
2598 => x"00000001",
2599 => x"330eabcd",
2600 => x"1234e66d",
2601 => x"deec0005",
2602 => x"000b0000",
2603 => x"00000000",
2604 => x"00000000",
2605 => x"00000000",
2606 => x"00000000",
2607 => x"00000000",
2608 => x"00000000",
2609 => x"00000000",
2610 => x"00000000",
2611 => x"00000000",
2612 => x"00000000",
2613 => x"00000000",
2614 => x"00000000",
2615 => x"00000000",
2616 => x"00000000",
2617 => x"00000000",
2618 => x"00000000",
2619 => x"00000000",
2620 => x"00000000",
2621 => x"00000000",
2622 => x"00000000",
2623 => x"00000000",
2624 => x"00000000",
2625 => x"00000000",
2626 => x"00000000",
2627 => x"00000000",
2628 => x"00000000",
2629 => x"00000000",
2630 => x"00000000",
2631 => x"00000000",
2632 => x"00000000",
2633 => x"00000000",
2634 => x"00000000",
2635 => x"00000000",
2636 => x"00000000",
2637 => x"00000000",
2638 => x"00000000",
2639 => x"00000000",
2640 => x"00000000",
2641 => x"00000000",
2642 => x"00000000",
2643 => x"00000000",
2644 => x"00000000",
2645 => x"00000000",
2646 => x"00000000",
2647 => x"00000000",
2648 => x"00000000",
2649 => x"00000000",
2650 => x"00000000",
2651 => x"00000000",
2652 => x"00000000",
2653 => x"00000000",
2654 => x"00000000",
2655 => x"00000000",
2656 => x"00000000",
2657 => x"00000000",
2658 => x"00000000",
2659 => x"00000000",
2660 => x"00000000",
2661 => x"00000000",
2662 => x"00000000",
2663 => x"00000000",
2664 => x"00000000",
2665 => x"00000000",
2666 => x"00000000",
2667 => x"00000000",
2668 => x"00000000",
2669 => x"00000000",
2670 => x"00000000",
2671 => x"00000000",
2672 => x"00000000",
2673 => x"00000000",
2674 => x"00000000",
2675 => x"00000000",
2676 => x"00000000",
2677 => x"00000000",
2678 => x"00000000",
2679 => x"00000000",
2680 => x"00000000",
2681 => x"00000000",
2682 => x"00000000",
2683 => x"00000000",
2684 => x"00000000",
2685 => x"00000000",
2686 => x"00000000",
2687 => x"00000000",
2688 => x"00000000",
2689 => x"00000000",
2690 => x"00000000",
2691 => x"00000000",
2692 => x"00000000",
2693 => x"00000000",
2694 => x"00000000",
2695 => x"00000000",
2696 => x"00000000",
2697 => x"00000000",
2698 => x"00000000",
2699 => x"00000000",
2700 => x"00000000",
2701 => x"00000000",
2702 => x"00000000",
2703 => x"00000000",
2704 => x"00000000",
2705 => x"00000000",
2706 => x"00000000",
2707 => x"00000000",
2708 => x"00000000",
2709 => x"00000000",
2710 => x"00000000",
2711 => x"00000000",
2712 => x"00000000",
2713 => x"00000000",
2714 => x"00000000",
2715 => x"00000000",
2716 => x"00000000",
2717 => x"00000000",
2718 => x"00000000",
2719 => x"00000000",
2720 => x"00000000",
2721 => x"00000000",
2722 => x"00000000",
2723 => x"00000000",
2724 => x"00000000",
2725 => x"00000000",
2726 => x"00000000",
2727 => x"00000000",
2728 => x"00000000",
2729 => x"00000000",
2730 => x"00000000",
2731 => x"00000000",
2732 => x"00000000",
2733 => x"00000000",
2734 => x"00000000",
2735 => x"00000000",
2736 => x"00000000",
2737 => x"00000000",
2738 => x"00000000",
2739 => x"00000000",
2740 => x"00000000",
2741 => x"00000000",
2742 => x"00000000",
2743 => x"00000000",
2744 => x"00000000",
2745 => x"00000000",
2746 => x"00000000",
2747 => x"00000000",
2748 => x"00000000",
2749 => x"00000000",
2750 => x"00000000",
2751 => x"00000000",
2752 => x"00000000",
2753 => x"00000000",
2754 => x"00000000",
2755 => x"00000000",
2756 => x"00000000",
2757 => x"00000000",
2758 => x"00000000",
2759 => x"00000000",
2760 => x"00000000",
2761 => x"00000000",
2762 => x"00000000",
2763 => x"00000000",
2764 => x"00000000",
2765 => x"00000000",
2766 => x"00000000",
2767 => x"00000000",
2768 => x"00000000",
2769 => x"00000000",
2770 => x"00000000",
2771 => x"00000000",
2772 => x"00000000",
2773 => x"00000000",
2774 => x"00000000",
2775 => x"00000000",
2776 => x"00000000",
2777 => x"00000000",
2778 => x"00000000",
2779 => x"00000000",
2780 => x"00000000",
2781 => x"00000000",
2782 => x"00000000",
2783 => x"00000000",
2784 => x"00000000",
2785 => x"00000000",
2786 => x"00000000",
2787 => x"00000000",
2788 => x"00000000",
2789 => x"00000000",
2790 => x"00000000",
2791 => x"ffffffff",
2792 => x"00000000",
2793 => x"00020000",
2794 => x"00000000",
2795 => x"00000000",
2796 => x"00002ba8",
2797 => x"00002ba8",
2798 => x"00002bb0",
2799 => x"00002bb0",
2800 => x"00002bb8",
2801 => x"00002bb8",
2802 => x"00002bc0",
2803 => x"00002bc0",
2804 => x"00002bc8",
2805 => x"00002bc8",
2806 => x"00002bd0",
2807 => x"00002bd0",
2808 => x"00002bd8",
2809 => x"00002bd8",
2810 => x"00002be0",
2811 => x"00002be0",
2812 => x"00002be8",
2813 => x"00002be8",
2814 => x"00002bf0",
2815 => x"00002bf0",
2816 => x"00002bf8",
2817 => x"00002bf8",
2818 => x"00002c00",
2819 => x"00002c00",
2820 => x"00002c08",
2821 => x"00002c08",
2822 => x"00002c10",
2823 => x"00002c10",
2824 => x"00002c18",
2825 => x"00002c18",
2826 => x"00002c20",
2827 => x"00002c20",
2828 => x"00002c28",
2829 => x"00002c28",
2830 => x"00002c30",
2831 => x"00002c30",
2832 => x"00002c38",
2833 => x"00002c38",
2834 => x"00002c40",
2835 => x"00002c40",
2836 => x"00002c48",
2837 => x"00002c48",
2838 => x"00002c50",
2839 => x"00002c50",
2840 => x"00002c58",
2841 => x"00002c58",
2842 => x"00002c60",
2843 => x"00002c60",
2844 => x"00002c68",
2845 => x"00002c68",
2846 => x"00002c70",
2847 => x"00002c70",
2848 => x"00002c78",
2849 => x"00002c78",
2850 => x"00002c80",
2851 => x"00002c80",
2852 => x"00002c88",
2853 => x"00002c88",
2854 => x"00002c90",
2855 => x"00002c90",
2856 => x"00002c98",
2857 => x"00002c98",
2858 => x"00002ca0",
2859 => x"00002ca0",
2860 => x"00002ca8",
2861 => x"00002ca8",
2862 => x"00002cb0",
2863 => x"00002cb0",
2864 => x"00002cb8",
2865 => x"00002cb8",
2866 => x"00002cc0",
2867 => x"00002cc0",
2868 => x"00002cc8",
2869 => x"00002cc8",
2870 => x"00002cd0",
2871 => x"00002cd0",
2872 => x"00002cd8",
2873 => x"00002cd8",
2874 => x"00002ce0",
2875 => x"00002ce0",
2876 => x"00002ce8",
2877 => x"00002ce8",
2878 => x"00002cf0",
2879 => x"00002cf0",
2880 => x"00002cf8",
2881 => x"00002cf8",
2882 => x"00002d00",
2883 => x"00002d00",
2884 => x"00002d08",
2885 => x"00002d08",
2886 => x"00002d10",
2887 => x"00002d10",
2888 => x"00002d18",
2889 => x"00002d18",
2890 => x"00002d20",
2891 => x"00002d20",
2892 => x"00002d28",
2893 => x"00002d28",
2894 => x"00002d30",
2895 => x"00002d30",
2896 => x"00002d38",
2897 => x"00002d38",
2898 => x"00002d40",
2899 => x"00002d40",
2900 => x"00002d48",
2901 => x"00002d48",
2902 => x"00002d50",
2903 => x"00002d50",
2904 => x"00002d58",
2905 => x"00002d58",
2906 => x"00002d60",
2907 => x"00002d60",
2908 => x"00002d68",
2909 => x"00002d68",
2910 => x"00002d70",
2911 => x"00002d70",
2912 => x"00002d78",
2913 => x"00002d78",
2914 => x"00002d80",
2915 => x"00002d80",
2916 => x"00002d88",
2917 => x"00002d88",
2918 => x"00002d90",
2919 => x"00002d90",
2920 => x"00002d98",
2921 => x"00002d98",
2922 => x"00002da0",
2923 => x"00002da0",
2924 => x"00002da8",
2925 => x"00002da8",
2926 => x"00002db0",
2927 => x"00002db0",
2928 => x"00002db8",
2929 => x"00002db8",
2930 => x"00002dc0",
2931 => x"00002dc0",
2932 => x"00002dc8",
2933 => x"00002dc8",
2934 => x"00002dd0",
2935 => x"00002dd0",
2936 => x"00002dd8",
2937 => x"00002dd8",
2938 => x"00002de0",
2939 => x"00002de0",
2940 => x"00002de8",
2941 => x"00002de8",
2942 => x"00002df0",
2943 => x"00002df0",
2944 => x"00002df8",
2945 => x"00002df8",
2946 => x"00002e00",
2947 => x"00002e00",
2948 => x"00002e08",
2949 => x"00002e08",
2950 => x"00002e10",
2951 => x"00002e10",
2952 => x"00002e18",
2953 => x"00002e18",
2954 => x"00002e20",
2955 => x"00002e20",
2956 => x"00002e28",
2957 => x"00002e28",
2958 => x"00002e30",
2959 => x"00002e30",
2960 => x"00002e38",
2961 => x"00002e38",
2962 => x"00002e40",
2963 => x"00002e40",
2964 => x"00002e48",
2965 => x"00002e48",
2966 => x"00002e50",
2967 => x"00002e50",
2968 => x"00002e58",
2969 => x"00002e58",
2970 => x"00002e60",
2971 => x"00002e60",
2972 => x"00002e68",
2973 => x"00002e68",
2974 => x"00002e70",
2975 => x"00002e70",
2976 => x"00002e78",
2977 => x"00002e78",
2978 => x"00002e80",
2979 => x"00002e80",
2980 => x"00002e88",
2981 => x"00002e88",
2982 => x"00002e90",
2983 => x"00002e90",
2984 => x"00002e98",
2985 => x"00002e98",
2986 => x"00002ea0",
2987 => x"00002ea0",
2988 => x"00002ea8",
2989 => x"00002ea8",
2990 => x"00002eb0",
2991 => x"00002eb0",
2992 => x"00002eb8",
2993 => x"00002eb8",
2994 => x"00002ec0",
2995 => x"00002ec0",
2996 => x"00002ec8",
2997 => x"00002ec8",
2998 => x"00002ed0",
2999 => x"00002ed0",
3000 => x"00002ed8",
3001 => x"00002ed8",
3002 => x"00002ee0",
3003 => x"00002ee0",
3004 => x"00002ee8",
3005 => x"00002ee8",
3006 => x"00002ef0",
3007 => x"00002ef0",
3008 => x"00002ef8",
3009 => x"00002ef8",
3010 => x"00002f00",
3011 => x"00002f00",
3012 => x"00002f08",
3013 => x"00002f08",
3014 => x"00002f10",
3015 => x"00002f10",
3016 => x"00002f18",
3017 => x"00002f18",
3018 => x"00002f20",
3019 => x"00002f20",
3020 => x"00002f28",
3021 => x"00002f28",
3022 => x"00002f30",
3023 => x"00002f30",
3024 => x"00002f38",
3025 => x"00002f38",
3026 => x"00002f40",
3027 => x"00002f40",
3028 => x"00002f48",
3029 => x"00002f48",
3030 => x"00002f50",
3031 => x"00002f50",
3032 => x"00002f58",
3033 => x"00002f58",
3034 => x"00002f60",
3035 => x"00002f60",
3036 => x"00002f68",
3037 => x"00002f68",
3038 => x"00002f70",
3039 => x"00002f70",
3040 => x"00002f78",
3041 => x"00002f78",
3042 => x"00002f80",
3043 => x"00002f80",
3044 => x"00002f88",
3045 => x"00002f88",
3046 => x"00002f90",
3047 => x"00002f90",
3048 => x"00002f98",
3049 => x"00002f98",
3050 => x"00002fa0",
3051 => x"00002fa0",
3052 => x"000027c0",
3053 => x"ffffffff",
3054 => x"00000000",
3055 => x"ffffffff",
3056 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
