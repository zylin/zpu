-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80f0ac0c",
     3 => x"3a0b0b80",
     4 => x"e2d80400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"92040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80f0",
   162 => x"98738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f9040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"e0040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80f0a80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82c43f80",
   257 => x"dcc23f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80088408",
   281 => x"88087575",
   282 => x"80c1c12d",
   283 => x"50508008",
   284 => x"56880c84",
   285 => x"0c800c51",
   286 => x"04800884",
   287 => x"08880875",
   288 => x"7580c08f",
   289 => x"2d505080",
   290 => x"0856880c",
   291 => x"840c800c",
   292 => x"51048008",
   293 => x"84088808",
   294 => x"80e3a12d",
   295 => x"880c840c",
   296 => x"800c0480",
   297 => x"f0a80880",
   298 => x"2ea43880",
   299 => x"f0ac0882",
   300 => x"2ebd3883",
   301 => x"80800b0b",
   302 => x"0b8180b4",
   303 => x"0c82a080",
   304 => x"0b8180b8",
   305 => x"0c829080",
   306 => x"0b8180bc",
   307 => x"0c04f880",
   308 => x"8080a40b",
   309 => x"0b0b8180",
   310 => x"b40cf880",
   311 => x"8082800b",
   312 => x"8180b80c",
   313 => x"f8808084",
   314 => x"800b8180",
   315 => x"bc0c0480",
   316 => x"c0a8808c",
   317 => x"0b0b0b81",
   318 => x"80b40c80",
   319 => x"c0a88094",
   320 => x"0b8180b8",
   321 => x"0c0b0b80",
   322 => x"e4f40b81",
   323 => x"80bc0c04",
   324 => x"ff3d0d81",
   325 => x"80c03351",
   326 => x"70a73880",
   327 => x"f0b40870",
   328 => x"08525270",
   329 => x"802e9438",
   330 => x"841280f0",
   331 => x"b40c702d",
   332 => x"80f0b408",
   333 => x"70085252",
   334 => x"70ee3881",
   335 => x"0b8180c0",
   336 => x"34833d0d",
   337 => x"0404803d",
   338 => x"0d0b0b81",
   339 => x"80b00880",
   340 => x"2e8e380b",
   341 => x"0b0b0b80",
   342 => x"0b802e09",
   343 => x"81068538",
   344 => x"823d0d04",
   345 => x"0b0b8180",
   346 => x"b0510b0b",
   347 => x"0bf5913f",
   348 => x"823d0d04",
   349 => x"04ff3d0d",
   350 => x"028f0533",
   351 => x"705252b2",
   352 => x"cd3f7151",
   353 => x"b3bc3f71",
   354 => x"800c833d",
   355 => x"0d04fa3d",
   356 => x"0d02a305",
   357 => x"3356758d",
   358 => x"2e80f438",
   359 => x"75883270",
   360 => x"307780ff",
   361 => x"32703072",
   362 => x"80257180",
   363 => x"25075451",
   364 => x"56585574",
   365 => x"95389f76",
   366 => x"278c3881",
   367 => x"8abc3355",
   368 => x"80ce7527",
   369 => x"ae38883d",
   370 => x"0d04818a",
   371 => x"bc335675",
   372 => x"802ef338",
   373 => x"8851adb4",
   374 => x"3fa051ad",
   375 => x"af3f8851",
   376 => x"adaa3f81",
   377 => x"8abc33ff",
   378 => x"05577681",
   379 => x"8abc3488",
   380 => x"3d0d0475",
   381 => x"51ad953f",
   382 => x"818abc33",
   383 => x"81115557",
   384 => x"73818abc",
   385 => x"34758189",
   386 => x"e8183488",
   387 => x"3d0d048a",
   388 => x"51acf93f",
   389 => x"818abc33",
   390 => x"81115654",
   391 => x"74818abc",
   392 => x"34800b81",
   393 => x"89e81534",
   394 => x"8056800b",
   395 => x"8189e817",
   396 => x"33565474",
   397 => x"a02e8338",
   398 => x"81547480",
   399 => x"2e903873",
   400 => x"802e8b38",
   401 => x"81167081",
   402 => x"ff065757",
   403 => x"dd397580",
   404 => x"2ebf3880",
   405 => x"0b818ab8",
   406 => x"33555574",
   407 => x"7427ab38",
   408 => x"73577410",
   409 => x"10107510",
   410 => x"05765481",
   411 => x"89e85381",
   412 => x"80c80551",
   413 => x"bdfc3f80",
   414 => x"08802ea6",
   415 => x"38811570",
   416 => x"81ff0656",
   417 => x"54767526",
   418 => x"d93880e5",
   419 => x"8451ac96",
   420 => x"3f80e580",
   421 => x"51ac8f3f",
   422 => x"800b818a",
   423 => x"bc34883d",
   424 => x"0d047410",
   425 => x"108189a8",
   426 => x"05700881",
   427 => x"8ac00c56",
   428 => x"800b818a",
   429 => x"bc34e739",
   430 => x"800b818a",
   431 => x"c43404fc",
   432 => x"3d0d8a51",
   433 => x"abc63f80",
   434 => x"e59851ab",
   435 => x"d93f800b",
   436 => x"818ab833",
   437 => x"53537272",
   438 => x"2780f538",
   439 => x"72101010",
   440 => x"73100581",
   441 => x"80c80570",
   442 => x"5254abba",
   443 => x"3f72842b",
   444 => x"70743182",
   445 => x"2b8181e8",
   446 => x"11335153",
   447 => x"5571802e",
   448 => x"b7387351",
   449 => x"bc8d3f80",
   450 => x"0881ff06",
   451 => x"52718926",
   452 => x"9338a051",
   453 => x"aaf63f81",
   454 => x"127081ff",
   455 => x"06535489",
   456 => x"7227ef38",
   457 => x"80e5b051",
   458 => x"aafc3f74",
   459 => x"7331822b",
   460 => x"8181e805",
   461 => x"51aaef3f",
   462 => x"8a51aad0",
   463 => x"3f811370",
   464 => x"81ff0681",
   465 => x"8ab83354",
   466 => x"54557173",
   467 => x"26ff8d38",
   468 => x"8a51aab8",
   469 => x"3f863d0d",
   470 => x"04fc3d0d",
   471 => x"8a51aaac",
   472 => x"3f800b81",
   473 => x"8abc3480",
   474 => x"0b818ab8",
   475 => x"34800b81",
   476 => x"8ac00c80",
   477 => x"e5b45281",
   478 => x"80c851ba",
   479 => x"a93f80e5",
   480 => x"b852818a",
   481 => x"b8337090",
   482 => x"29713170",
   483 => x"10108181",
   484 => x"e8055356",
   485 => x"54ba8f3f",
   486 => x"818ab833",
   487 => x"70101081",
   488 => x"89a805ab",
   489 => x"94710c54",
   490 => x"81115155",
   491 => x"74818ab8",
   492 => x"3480e5cc",
   493 => x"527481ff",
   494 => x"06708a29",
   495 => x"8180c805",
   496 => x"5253b9e2",
   497 => x"3f80e5d4",
   498 => x"52818ab8",
   499 => x"33709029",
   500 => x"71317010",
   501 => x"108181e8",
   502 => x"05535555",
   503 => x"b9c83f81",
   504 => x"8ab83370",
   505 => x"10108189",
   506 => x"a8059cae",
   507 => x"710c5481",
   508 => x"11515473",
   509 => x"818ab834",
   510 => x"80e5e852",
   511 => x"7381ff06",
   512 => x"708a2981",
   513 => x"80c80552",
   514 => x"53b99b3f",
   515 => x"80e5f052",
   516 => x"818ab833",
   517 => x"70902971",
   518 => x"31701010",
   519 => x"8181e805",
   520 => x"535654b9",
   521 => x"813f818a",
   522 => x"b8337010",
   523 => x"108189a8",
   524 => x"059e8971",
   525 => x"0c548111",
   526 => x"51557481",
   527 => x"8ab83480",
   528 => x"e6885274",
   529 => x"81ff0670",
   530 => x"8a298180",
   531 => x"c8055253",
   532 => x"b8d43f80",
   533 => x"e6905281",
   534 => x"8ab83370",
   535 => x"90297131",
   536 => x"70101081",
   537 => x"81e80553",
   538 => x"5555b8ba",
   539 => x"3f818ab8",
   540 => x"33701010",
   541 => x"8189a805",
   542 => x"a0bf710c",
   543 => x"54811151",
   544 => x"5473818a",
   545 => x"b83480e6",
   546 => x"a8527381",
   547 => x"ff06708a",
   548 => x"298180c8",
   549 => x"055253b8",
   550 => x"8d3f80e6",
   551 => x"b052818a",
   552 => x"b8337090",
   553 => x"29713170",
   554 => x"10108181",
   555 => x"e8055356",
   556 => x"54b7f33f",
   557 => x"818ab833",
   558 => x"70101081",
   559 => x"89a805a6",
   560 => x"e8710c54",
   561 => x"81115155",
   562 => x"74818ab8",
   563 => x"3480e6c8",
   564 => x"527481ff",
   565 => x"06708a29",
   566 => x"8180c805",
   567 => x"5253b7c6",
   568 => x"3f80e6d0",
   569 => x"52818ab8",
   570 => x"33709029",
   571 => x"71317010",
   572 => x"108181e8",
   573 => x"05535555",
   574 => x"b7ac3f81",
   575 => x"8ab83370",
   576 => x"10108189",
   577 => x"a805a28f",
   578 => x"710c5481",
   579 => x"11515473",
   580 => x"818ab834",
   581 => x"80e6f852",
   582 => x"7381ff06",
   583 => x"708a2981",
   584 => x"80c80552",
   585 => x"53b6ff3f",
   586 => x"80e6fc52",
   587 => x"818ab833",
   588 => x"70902971",
   589 => x"31701010",
   590 => x"8181e805",
   591 => x"535654b6",
   592 => x"e53f818a",
   593 => x"b8337010",
   594 => x"108189a8",
   595 => x"05969071",
   596 => x"0c548111",
   597 => x"51557481",
   598 => x"8ab83480",
   599 => x"e7885274",
   600 => x"81ff0670",
   601 => x"8a298180",
   602 => x"c8055253",
   603 => x"b6b83f80",
   604 => x"e7905281",
   605 => x"8ab83370",
   606 => x"90297131",
   607 => x"70101081",
   608 => x"81e80553",
   609 => x"5555b69e",
   610 => x"3f818ab8",
   611 => x"33701010",
   612 => x"8189a805",
   613 => x"99d2710c",
   614 => x"54811151",
   615 => x"5473818a",
   616 => x"b83480e8",
   617 => x"ec527381",
   618 => x"ff06708a",
   619 => x"298180c8",
   620 => x"055253b5",
   621 => x"f13f80e7",
   622 => x"9c52818a",
   623 => x"b8337090",
   624 => x"29713170",
   625 => x"10108181",
   626 => x"e8055356",
   627 => x"54b5d73f",
   628 => x"818ab833",
   629 => x"70101081",
   630 => x"89a80596",
   631 => x"90710c54",
   632 => x"81115155",
   633 => x"74818ab8",
   634 => x"3480e7ac",
   635 => x"527481ff",
   636 => x"06708a29",
   637 => x"8180c805",
   638 => x"5253b5aa",
   639 => x"3f80e7b4",
   640 => x"52818ab8",
   641 => x"33709029",
   642 => x"71317010",
   643 => x"108181e8",
   644 => x"05535555",
   645 => x"b5903f81",
   646 => x"8ab83370",
   647 => x"10108189",
   648 => x"a8059ca2",
   649 => x"710c5481",
   650 => x"11515473",
   651 => x"818ab834",
   652 => x"80e7c452",
   653 => x"7381ff06",
   654 => x"708a2981",
   655 => x"80c80552",
   656 => x"53b4e33f",
   657 => x"80e7ec52",
   658 => x"818ab833",
   659 => x"70902971",
   660 => x"31701010",
   661 => x"8181e805",
   662 => x"535654b4",
   663 => x"c93f818a",
   664 => x"b8337010",
   665 => x"108189a8",
   666 => x"058db871",
   667 => x"0c548111",
   668 => x"51557481",
   669 => x"8ab83480",
   670 => x"e4f85274",
   671 => x"81ff0670",
   672 => x"8a298180",
   673 => x"c8055253",
   674 => x"b49c3f80",
   675 => x"e7ec5281",
   676 => x"8ab83370",
   677 => x"90297131",
   678 => x"70101081",
   679 => x"81e80553",
   680 => x"5555b482",
   681 => x"3f818ab8",
   682 => x"33701010",
   683 => x"8189a805",
   684 => x"8dbf710c",
   685 => x"54810553",
   686 => x"72818ab8",
   687 => x"34f8803f",
   688 => x"80e58051",
   689 => x"a3e03f81",
   690 => x"0b818ac4",
   691 => x"34a7ca3f",
   692 => x"8008ae38",
   693 => x"818ac008",
   694 => x"53728d38",
   695 => x"818ac433",
   696 => x"5372ea38",
   697 => x"863d0d04",
   698 => x"722d800b",
   699 => x"818ac00c",
   700 => x"80e58051",
   701 => x"a3b03f81",
   702 => x"8ac43353",
   703 => x"72cf38e4",
   704 => x"39a7a93f",
   705 => x"800881ff",
   706 => x"0651f582",
   707 => x"3fffbe39",
   708 => x"f63d0d80",
   709 => x"0b8189e8",
   710 => x"338189e8",
   711 => x"59555673",
   712 => x"a02e0981",
   713 => x"06963881",
   714 => x"167081ff",
   715 => x"068189e8",
   716 => x"11703353",
   717 => x"59575473",
   718 => x"a02eec38",
   719 => x"80588077",
   720 => x"33565474",
   721 => x"742e8338",
   722 => x"815474a0",
   723 => x"2e81ce38",
   724 => x"7381fb38",
   725 => x"74a02e81",
   726 => x"c4388118",
   727 => x"7081ff06",
   728 => x"59548178",
   729 => x"26d83890",
   730 => x"538c3dfc",
   731 => x"05527651",
   732 => x"b8cf3f80",
   733 => x"0859800b",
   734 => x"8189e833",
   735 => x"8189e859",
   736 => x"555673a0",
   737 => x"2e098106",
   738 => x"96388116",
   739 => x"7081ff06",
   740 => x"8189e811",
   741 => x"70335759",
   742 => x"575873a0",
   743 => x"2eec3880",
   744 => x"58807733",
   745 => x"56547474",
   746 => x"2e833881",
   747 => x"5474a02e",
   748 => x"81ac3873",
   749 => x"828c3874",
   750 => x"a02e81a2",
   751 => x"38811870",
   752 => x"81ff0659",
   753 => x"55827826",
   754 => x"d8389053",
   755 => x"8c3df805",
   756 => x"527651b7",
   757 => x"ec3f8008",
   758 => x"57800883",
   759 => x"38905778",
   760 => x"fc065580",
   761 => x"56757727",
   762 => x"ab387583",
   763 => x"06597880",
   764 => x"2e819c38",
   765 => x"80e7cc51",
   766 => x"a1ac3f74",
   767 => x"70840556",
   768 => x"0852a051",
   769 => x"a1c33fa0",
   770 => x"51a1813f",
   771 => x"81165676",
   772 => x"7626d738",
   773 => x"8a51a0f4",
   774 => x"3f8c3d0d",
   775 => x"04811670",
   776 => x"81ff0681",
   777 => x"89e81170",
   778 => x"335c5257",
   779 => x"5778a02e",
   780 => x"098106fe",
   781 => x"a5388116",
   782 => x"7081ff06",
   783 => x"8189e811",
   784 => x"70335c52",
   785 => x"575778a0",
   786 => x"2ed338fe",
   787 => x"8d398116",
   788 => x"7081ff06",
   789 => x"8189e811",
   790 => x"595755fd",
   791 => x"e1398116",
   792 => x"7081ff06",
   793 => x"8189e811",
   794 => x"70335752",
   795 => x"575773a0",
   796 => x"2e098106",
   797 => x"fec73881",
   798 => x"167081ff",
   799 => x"068189e8",
   800 => x"11703357",
   801 => x"52575773",
   802 => x"a02ed338",
   803 => x"feaf3980",
   804 => x"e7d051a0",
   805 => x"913f7452",
   806 => x"a051a0ad",
   807 => x"3f80e7d4",
   808 => x"51a0833f",
   809 => x"80e7cc51",
   810 => x"9ffc3f74",
   811 => x"70840556",
   812 => x"0852a051",
   813 => x"a0933fa0",
   814 => x"519fd13f",
   815 => x"811656fe",
   816 => x"ce398116",
   817 => x"7081ff06",
   818 => x"8189e811",
   819 => x"595755fd",
   820 => x"d039f63d",
   821 => x"0d800b81",
   822 => x"89e83381",
   823 => x"89e85955",
   824 => x"5673a02e",
   825 => x"09810696",
   826 => x"38811670",
   827 => x"81ff0681",
   828 => x"89e81170",
   829 => x"33535957",
   830 => x"5473a02e",
   831 => x"ec388058",
   832 => x"80773356",
   833 => x"5474742e",
   834 => x"83388154",
   835 => x"74a02e81",
   836 => x"8f387381",
   837 => x"bc3874a0",
   838 => x"2e818538",
   839 => x"81187081",
   840 => x"ff065954",
   841 => x"817826d8",
   842 => x"3890538c",
   843 => x"3dfc0552",
   844 => x"7651b58d",
   845 => x"3f800859",
   846 => x"800b8189",
   847 => x"e8338189",
   848 => x"e8595556",
   849 => x"73a02e09",
   850 => x"81069638",
   851 => x"81167081",
   852 => x"ff068189",
   853 => x"e8117033",
   854 => x"57595758",
   855 => x"73a02eec",
   856 => x"38805880",
   857 => x"77335654",
   858 => x"74742e83",
   859 => x"38815474",
   860 => x"a02e80ed",
   861 => x"3873819a",
   862 => x"3874a02e",
   863 => x"80e33881",
   864 => x"187081ff",
   865 => x"06595582",
   866 => x"7826d838",
   867 => x"90538c3d",
   868 => x"f8055276",
   869 => x"51b4aa3f",
   870 => x"8008790c",
   871 => x"8c3d0d04",
   872 => x"81167081",
   873 => x"ff068189",
   874 => x"e8117033",
   875 => x"5c525757",
   876 => x"78a02e09",
   877 => x"8106fee4",
   878 => x"38811670",
   879 => x"81ff0681",
   880 => x"89e81170",
   881 => x"335c5257",
   882 => x"5778a02e",
   883 => x"d338fecc",
   884 => x"39811670",
   885 => x"81ff0681",
   886 => x"89e81159",
   887 => x"5755fea0",
   888 => x"39811670",
   889 => x"81ff0681",
   890 => x"89e81170",
   891 => x"33575257",
   892 => x"5773a02e",
   893 => x"098106ff",
   894 => x"86388116",
   895 => x"7081ff06",
   896 => x"8189e811",
   897 => x"70335752",
   898 => x"575773a0",
   899 => x"2ed338fe",
   900 => x"ee398116",
   901 => x"7081ff06",
   902 => x"8189e811",
   903 => x"595755fe",
   904 => x"c239803d",
   905 => x"0d8c519c",
   906 => x"e33f823d",
   907 => x"0d04fb3d",
   908 => x"0d80e7d8",
   909 => x"519cef3f",
   910 => x"805680f0",
   911 => x"bc087610",
   912 => x"81fe0688",
   913 => x"120c5481",
   914 => x"d00b8c15",
   915 => x"0c8c1408",
   916 => x"70812a81",
   917 => x"06515574",
   918 => x"f4388c14",
   919 => x"0870872a",
   920 => x"81065553",
   921 => x"73802e80",
   922 => x"de388116",
   923 => x"7081ff06",
   924 => x"70982b56",
   925 => x"57537380",
   926 => x"25c03880",
   927 => x"e7e4519c",
   928 => x"a53f80f0",
   929 => x"b8087510",
   930 => x"81fe0688",
   931 => x"120c5481",
   932 => x"d00b8c15",
   933 => x"0c8c1408",
   934 => x"70812a81",
   935 => x"06515372",
   936 => x"f4388c14",
   937 => x"0870872a",
   938 => x"81065553",
   939 => x"73802e80",
   940 => x"c0388115",
   941 => x"7081ff06",
   942 => x"70982b56",
   943 => x"56567380",
   944 => x"25c03887",
   945 => x"3d0d0480",
   946 => x"e7f0519b",
   947 => x"d93f7552",
   948 => x"88519bf5",
   949 => x"3f80e880",
   950 => x"519bcb3f",
   951 => x"81167081",
   952 => x"ff067098",
   953 => x"2b565753",
   954 => x"738025fe",
   955 => x"cd38ff8b",
   956 => x"3980e7f0",
   957 => x"519baf3f",
   958 => x"74528851",
   959 => x"9bcb3f80",
   960 => x"e880519b",
   961 => x"a13fffaa",
   962 => x"39f83d0d",
   963 => x"80e89051",
   964 => x"9b943f82",
   965 => x"80519cd3",
   966 => x"3f80e8a4",
   967 => x"519b873f",
   968 => x"80d05288",
   969 => x"519ba23f",
   970 => x"80e8c051",
   971 => x"9af83f80",
   972 => x"5780f0bc",
   973 => x"085581a1",
   974 => x"0b88160c",
   975 => x"81900b8c",
   976 => x"160c8c15",
   977 => x"0870812a",
   978 => x"81065154",
   979 => x"73f4388c",
   980 => x"15087488",
   981 => x"170c5380",
   982 => x"e00b8c16",
   983 => x"0c8c1508",
   984 => x"70812a81",
   985 => x"06575475",
   986 => x"f4388c15",
   987 => x"0870872a",
   988 => x"81067887",
   989 => x"06565156",
   990 => x"75802eb3",
   991 => x"3873872e",
   992 => x"81803881",
   993 => x"177083ff",
   994 => x"ff065855",
   995 => x"82807726",
   996 => x"ff9f3880",
   997 => x"f0bc0854",
   998 => x"80e00b8c",
   999 => x"150c8c14",
  1000 => x"0870812a",
  1001 => x"81065856",
  1002 => x"76f4388a",
  1003 => x"3d0d0488",
  1004 => x"15087081",
  1005 => x"ff0680e7",
  1006 => x"cc535654",
  1007 => x"99e83f74",
  1008 => x"5288519a",
  1009 => x"843f80eb",
  1010 => x"e45199da",
  1011 => x"3f755474",
  1012 => x"80e62ebe",
  1013 => x"38748d32",
  1014 => x"70307080",
  1015 => x"25760752",
  1016 => x"57537280",
  1017 => x"c138748a",
  1018 => x"2ebc3876",
  1019 => x"87068b3d",
  1020 => x"7105f805",
  1021 => x"54547473",
  1022 => x"3473872e",
  1023 => x"098106ff",
  1024 => x"82388a3d",
  1025 => x"f8055199",
  1026 => x"9d3f8a51",
  1027 => x"98fe3ffe",
  1028 => x"f2398175",
  1029 => x"8d327030",
  1030 => x"70802573",
  1031 => x"07525854",
  1032 => x"5472802e",
  1033 => x"c1387687",
  1034 => x"068b3d71",
  1035 => x"05f80557",
  1036 => x"54a07634",
  1037 => x"73872e09",
  1038 => x"8106fec7",
  1039 => x"38c439fb",
  1040 => x"3d0d9c56",
  1041 => x"80e8c451",
  1042 => x"98dc3f75",
  1043 => x"52885198",
  1044 => x"f83f80f0",
  1045 => x"bc085481",
  1046 => x"ec0b8815",
  1047 => x"0c81900b",
  1048 => x"8c150c8c",
  1049 => x"14087081",
  1050 => x"2a810651",
  1051 => x"5372f438",
  1052 => x"8c140876",
  1053 => x"88160c53",
  1054 => x"900b8c15",
  1055 => x"0c8c1408",
  1056 => x"70812a81",
  1057 => x"06515574",
  1058 => x"f4388c14",
  1059 => x"085381ed",
  1060 => x"0b88150c",
  1061 => x"81900b8c",
  1062 => x"150c8c14",
  1063 => x"0870812a",
  1064 => x"81065155",
  1065 => x"74f4388c",
  1066 => x"14087588",
  1067 => x"160c5380",
  1068 => x"e00b8c15",
  1069 => x"0c8c1408",
  1070 => x"70812a81",
  1071 => x"06515372",
  1072 => x"f4388c14",
  1073 => x"08881508",
  1074 => x"7081ff06",
  1075 => x"8c170870",
  1076 => x"872a8132",
  1077 => x"81065852",
  1078 => x"57515373",
  1079 => x"802ea738",
  1080 => x"80e8d451",
  1081 => x"97c03f74",
  1082 => x"52885197",
  1083 => x"dc3f8a51",
  1084 => x"979a3f81",
  1085 => x"167081ff",
  1086 => x"06575580",
  1087 => x"d57627fe",
  1088 => x"c338873d",
  1089 => x"0d0480e8",
  1090 => x"dc51979a",
  1091 => x"3fe039f6",
  1092 => x"3d0d800b",
  1093 => x"8189e833",
  1094 => x"8189e859",
  1095 => x"555673a0",
  1096 => x"2e098106",
  1097 => x"96388116",
  1098 => x"7081ff06",
  1099 => x"8189e811",
  1100 => x"70335359",
  1101 => x"575473a0",
  1102 => x"2eec3880",
  1103 => x"58807733",
  1104 => x"56547474",
  1105 => x"2e833881",
  1106 => x"5474a02e",
  1107 => x"83883873",
  1108 => x"83b53874",
  1109 => x"a02e82fe",
  1110 => x"38811870",
  1111 => x"81ff0659",
  1112 => x"54817826",
  1113 => x"d8389053",
  1114 => x"8c3dfc05",
  1115 => x"527651ac",
  1116 => x"d03f8008",
  1117 => x"81ff0659",
  1118 => x"800b8189",
  1119 => x"e8338189",
  1120 => x"e8595556",
  1121 => x"73a02e09",
  1122 => x"81069638",
  1123 => x"81167081",
  1124 => x"ff068189",
  1125 => x"e8117033",
  1126 => x"57595758",
  1127 => x"73a02eec",
  1128 => x"38805880",
  1129 => x"77335654",
  1130 => x"74742e83",
  1131 => x"38815474",
  1132 => x"a02e82e3",
  1133 => x"38738390",
  1134 => x"3874a02e",
  1135 => x"82d93881",
  1136 => x"187081ff",
  1137 => x"06595582",
  1138 => x"7826d838",
  1139 => x"90538c3d",
  1140 => x"f8055276",
  1141 => x"51abea3f",
  1142 => x"800881ff",
  1143 => x"0680f0bc",
  1144 => x"08565681",
  1145 => x"ec0b8816",
  1146 => x"0c81900b",
  1147 => x"8c160c8c",
  1148 => x"15087081",
  1149 => x"2a810659",
  1150 => x"5777f438",
  1151 => x"8c150879",
  1152 => x"88170c54",
  1153 => x"900b8c16",
  1154 => x"0c8c1508",
  1155 => x"70812a81",
  1156 => x"06595777",
  1157 => x"f4388c15",
  1158 => x"08768817",
  1159 => x"0c5480d0",
  1160 => x"0b8c160c",
  1161 => x"8c150870",
  1162 => x"812a8106",
  1163 => x"575475f4",
  1164 => x"388c1508",
  1165 => x"5481ec0b",
  1166 => x"88160c81",
  1167 => x"900b8c16",
  1168 => x"0c8c1508",
  1169 => x"70812a81",
  1170 => x"06585876",
  1171 => x"f4388c15",
  1172 => x"08798817",
  1173 => x"0c54900b",
  1174 => x"8c160c8c",
  1175 => x"15087081",
  1176 => x"2a81065a",
  1177 => x"5778f438",
  1178 => x"8c150854",
  1179 => x"81ed0b88",
  1180 => x"160c8190",
  1181 => x"0b8c160c",
  1182 => x"8c150870",
  1183 => x"812a8106",
  1184 => x"515675f4",
  1185 => x"388c1508",
  1186 => x"7688170c",
  1187 => x"5480e00b",
  1188 => x"8c160c8c",
  1189 => x"15087081",
  1190 => x"2a81065a",
  1191 => x"5778f438",
  1192 => x"8c150888",
  1193 => x"16087081",
  1194 => x"ff068c18",
  1195 => x"0870872a",
  1196 => x"81328106",
  1197 => x"595c5851",
  1198 => x"5474802e",
  1199 => x"819a3880",
  1200 => x"e8e45193",
  1201 => x"e13f7552",
  1202 => x"885193fd",
  1203 => x"3f8a5193",
  1204 => x"bb3f8c3d",
  1205 => x"0d048116",
  1206 => x"7081ff06",
  1207 => x"8189e811",
  1208 => x"70335c52",
  1209 => x"575778a0",
  1210 => x"2e098106",
  1211 => x"fceb3881",
  1212 => x"167081ff",
  1213 => x"068189e8",
  1214 => x"1170335c",
  1215 => x"52575778",
  1216 => x"a02ed338",
  1217 => x"fcd33981",
  1218 => x"167081ff",
  1219 => x"068189e8",
  1220 => x"11595755",
  1221 => x"fca73981",
  1222 => x"167081ff",
  1223 => x"068189e8",
  1224 => x"11703357",
  1225 => x"52575773",
  1226 => x"a02e0981",
  1227 => x"06fd9038",
  1228 => x"81167081",
  1229 => x"ff068189",
  1230 => x"e8117033",
  1231 => x"57525757",
  1232 => x"73a02ed3",
  1233 => x"38fcf839",
  1234 => x"81167081",
  1235 => x"ff068189",
  1236 => x"e8115957",
  1237 => x"55fccc39",
  1238 => x"80e8f051",
  1239 => x"92c83f8a",
  1240 => x"5192a93f",
  1241 => x"8c3d0d04",
  1242 => x"ff3d0d80",
  1243 => x"f0bc0852",
  1244 => x"81ec0b88",
  1245 => x"130c8190",
  1246 => x"0b8c130c",
  1247 => x"8c120870",
  1248 => x"812a7081",
  1249 => x"06515151",
  1250 => x"70f2388c",
  1251 => x"1208519d",
  1252 => x"0b88130c",
  1253 => x"900b8c13",
  1254 => x"0c8c1208",
  1255 => x"70812a70",
  1256 => x"81065151",
  1257 => x"5170f238",
  1258 => x"8c120851",
  1259 => x"80c50b88",
  1260 => x"130c80d0",
  1261 => x"0b8c130c",
  1262 => x"8c120870",
  1263 => x"812a7081",
  1264 => x"06515151",
  1265 => x"70f2388c",
  1266 => x"12085181",
  1267 => x"ec0b8813",
  1268 => x"0c81900b",
  1269 => x"8c130c8c",
  1270 => x"12087081",
  1271 => x"2a708106",
  1272 => x"51515170",
  1273 => x"f2388c12",
  1274 => x"0851a10b",
  1275 => x"88130c90",
  1276 => x"0b8c130c",
  1277 => x"8c120870",
  1278 => x"812a7081",
  1279 => x"06515151",
  1280 => x"70f2388c",
  1281 => x"12085189",
  1282 => x"0b88130c",
  1283 => x"80d00b8c",
  1284 => x"130c8c12",
  1285 => x"0870812a",
  1286 => x"70810651",
  1287 => x"515170f2",
  1288 => x"388c1208",
  1289 => x"5181ec0b",
  1290 => x"88130c81",
  1291 => x"900b8c13",
  1292 => x"0c8c1208",
  1293 => x"70812a70",
  1294 => x"81065151",
  1295 => x"5170f238",
  1296 => x"8c120851",
  1297 => x"b30b8813",
  1298 => x"0c900b8c",
  1299 => x"130c8c12",
  1300 => x"0870812a",
  1301 => x"70810651",
  1302 => x"515170f2",
  1303 => x"388c1208",
  1304 => x"51880b88",
  1305 => x"130c80d0",
  1306 => x"0b8c130c",
  1307 => x"8c120870",
  1308 => x"812a7081",
  1309 => x"06515151",
  1310 => x"70f2388c",
  1311 => x"12085181",
  1312 => x"ec0b8813",
  1313 => x"0c81900b",
  1314 => x"8c130c8c",
  1315 => x"12087081",
  1316 => x"2a708106",
  1317 => x"51515170",
  1318 => x"f2388c12",
  1319 => x"0851b40b",
  1320 => x"88130c90",
  1321 => x"0b8c130c",
  1322 => x"8c120870",
  1323 => x"812a7081",
  1324 => x"06515151",
  1325 => x"70f2388c",
  1326 => x"12085196",
  1327 => x"0b88130c",
  1328 => x"80d00b8c",
  1329 => x"130c8c12",
  1330 => x"0870812a",
  1331 => x"70810651",
  1332 => x"515170f2",
  1333 => x"388c1208",
  1334 => x"5181ec0b",
  1335 => x"88130c81",
  1336 => x"900b8c13",
  1337 => x"0c8c1208",
  1338 => x"70812a70",
  1339 => x"81065151",
  1340 => x"5170f238",
  1341 => x"8c120851",
  1342 => x"b60b8813",
  1343 => x"0c900b8c",
  1344 => x"130c8c12",
  1345 => x"0870812a",
  1346 => x"70810651",
  1347 => x"515170f2",
  1348 => x"388c1208",
  1349 => x"5180e00b",
  1350 => x"88130c80",
  1351 => x"d00b8c13",
  1352 => x"0c8c1208",
  1353 => x"70812a70",
  1354 => x"81065151",
  1355 => x"5170f238",
  1356 => x"8c120851",
  1357 => x"81ec0b88",
  1358 => x"130c8190",
  1359 => x"0b8c130c",
  1360 => x"8c120870",
  1361 => x"812a7081",
  1362 => x"06515151",
  1363 => x"70f2388c",
  1364 => x"12085180",
  1365 => x"c90b8813",
  1366 => x"0c900b8c",
  1367 => x"130c8c12",
  1368 => x"0870812a",
  1369 => x"70810651",
  1370 => x"515170f2",
  1371 => x"388c1208",
  1372 => x"5181c00b",
  1373 => x"88130c80",
  1374 => x"d00b8c13",
  1375 => x"0c8c1208",
  1376 => x"70812a70",
  1377 => x"81065151",
  1378 => x"5170f238",
  1379 => x"8c120851",
  1380 => x"833d0d04",
  1381 => x"fe3d0d80",
  1382 => x"e980518e",
  1383 => x"893f80e9",
  1384 => x"a0518e82",
  1385 => x"3f80e9e8",
  1386 => x"518dfb3f",
  1387 => x"80eab051",
  1388 => x"8df43f80",
  1389 => x"f0c00870",
  1390 => x"0852528f",
  1391 => x"ae3f8008",
  1392 => x"81ff0652",
  1393 => x"718c2793",
  1394 => x"38a0518d",
  1395 => x"bf3f8112",
  1396 => x"7081ff06",
  1397 => x"53538c72",
  1398 => x"26ef3880",
  1399 => x"f0c00884",
  1400 => x"11085252",
  1401 => x"8f853f80",
  1402 => x"0881ff06",
  1403 => x"52718c27",
  1404 => x"9338a051",
  1405 => x"8d963f81",
  1406 => x"127081ff",
  1407 => x"0653538c",
  1408 => x"7226ef38",
  1409 => x"80f0c008",
  1410 => x"88110852",
  1411 => x"528edc3f",
  1412 => x"800881ff",
  1413 => x"0652718c",
  1414 => x"279338a0",
  1415 => x"518ced3f",
  1416 => x"81127081",
  1417 => x"ff065353",
  1418 => x"8c7226ef",
  1419 => x"3880f0c0",
  1420 => x"088c1108",
  1421 => x"52528eb3",
  1422 => x"3f800881",
  1423 => x"ff065271",
  1424 => x"8c279338",
  1425 => x"a0518cc4",
  1426 => x"3f811270",
  1427 => x"81ff0653",
  1428 => x"538c7226",
  1429 => x"ef3880ea",
  1430 => x"cc518cca",
  1431 => x"3f80f0c0",
  1432 => x"08901108",
  1433 => x"52528e83",
  1434 => x"3f800881",
  1435 => x"ff065271",
  1436 => x"8c279338",
  1437 => x"a0518c94",
  1438 => x"3f811270",
  1439 => x"81ff0653",
  1440 => x"538c7226",
  1441 => x"ef3880f0",
  1442 => x"c0089411",
  1443 => x"0852528d",
  1444 => x"da3f8008",
  1445 => x"81ff0652",
  1446 => x"718c2793",
  1447 => x"38a0518b",
  1448 => x"eb3f8112",
  1449 => x"7081ff06",
  1450 => x"53538c72",
  1451 => x"26ef3880",
  1452 => x"f0c00898",
  1453 => x"11085252",
  1454 => x"8db13f80",
  1455 => x"0881ff06",
  1456 => x"52718c27",
  1457 => x"9338a051",
  1458 => x"8bc23f81",
  1459 => x"127081ff",
  1460 => x"0653538c",
  1461 => x"7226ef38",
  1462 => x"80f0c008",
  1463 => x"9c110852",
  1464 => x"528d883f",
  1465 => x"800881ff",
  1466 => x"0652718c",
  1467 => x"279338a0",
  1468 => x"518b993f",
  1469 => x"81127081",
  1470 => x"ff065353",
  1471 => x"8c7226ef",
  1472 => x"3880eae8",
  1473 => x"518b9f3f",
  1474 => x"80f0c008",
  1475 => x"53810bb0",
  1476 => x"140cb013",
  1477 => x"08527180",
  1478 => x"25f838a0",
  1479 => x"1308518c",
  1480 => x"ca3f8008",
  1481 => x"81ff0652",
  1482 => x"718c2793",
  1483 => x"38a0518a",
  1484 => x"db3f8112",
  1485 => x"7081ff06",
  1486 => x"53538c72",
  1487 => x"26ef3880",
  1488 => x"f0c008a4",
  1489 => x"11085252",
  1490 => x"8ca13f80",
  1491 => x"0881ff06",
  1492 => x"52718c27",
  1493 => x"9338a051",
  1494 => x"8ab23f81",
  1495 => x"127081ff",
  1496 => x"0653538c",
  1497 => x"7226ef38",
  1498 => x"80f0c008",
  1499 => x"a8110852",
  1500 => x"528bf83f",
  1501 => x"800881ff",
  1502 => x"0652718c",
  1503 => x"279338a0",
  1504 => x"518a893f",
  1505 => x"81127081",
  1506 => x"ff065353",
  1507 => x"8c7226ef",
  1508 => x"3880f0c0",
  1509 => x"08ac1108",
  1510 => x"52528bcf",
  1511 => x"3f800881",
  1512 => x"ff065271",
  1513 => x"8c279338",
  1514 => x"a05189e0",
  1515 => x"3f811270",
  1516 => x"81ff0653",
  1517 => x"538c7226",
  1518 => x"ef3880eb",
  1519 => x"845189e6",
  1520 => x"3f80f0c0",
  1521 => x"08b01108",
  1522 => x"fe0a0652",
  1523 => x"538b9c3f",
  1524 => x"80f0c008",
  1525 => x"53800bb0",
  1526 => x"140c80eb",
  1527 => x"985189c6",
  1528 => x"3f80ebb0",
  1529 => x"5189bf3f",
  1530 => x"80f0c008",
  1531 => x"80c01108",
  1532 => x"52528af7",
  1533 => x"3f800881",
  1534 => x"ff065271",
  1535 => x"98279338",
  1536 => x"a0518988",
  1537 => x"3f811270",
  1538 => x"81ff0651",
  1539 => x"52987226",
  1540 => x"ef3880f0",
  1541 => x"c00880c8",
  1542 => x"11085253",
  1543 => x"8acd3f80",
  1544 => x"0881ff06",
  1545 => x"52719827",
  1546 => x"9338a051",
  1547 => x"88de3f81",
  1548 => x"127081ff",
  1549 => x"06515298",
  1550 => x"7226ef38",
  1551 => x"80ebcc51",
  1552 => x"88e43f80",
  1553 => x"f0c00880",
  1554 => x"c4110852",
  1555 => x"538a9c3f",
  1556 => x"800881ff",
  1557 => x"06527198",
  1558 => x"279338a0",
  1559 => x"5188ad3f",
  1560 => x"81127081",
  1561 => x"ff065152",
  1562 => x"987226ef",
  1563 => x"3880f0c0",
  1564 => x"0880cc11",
  1565 => x"08525389",
  1566 => x"f23f8008",
  1567 => x"81ff0652",
  1568 => x"71982793",
  1569 => x"38a05188",
  1570 => x"833f8112",
  1571 => x"7081ff06",
  1572 => x"51529872",
  1573 => x"26ef388a",
  1574 => x"5187f13f",
  1575 => x"80f0c008",
  1576 => x"b4110870",
  1577 => x"81ff0680",
  1578 => x"ebe85452",
  1579 => x"545287f6",
  1580 => x"3f715189",
  1581 => x"b63fa051",
  1582 => x"87d23f71",
  1583 => x"86269338",
  1584 => x"71101080",
  1585 => x"edb80553",
  1586 => x"72080480",
  1587 => x"ebfc5187",
  1588 => x"d53f8a51",
  1589 => x"87b63f84",
  1590 => x"3d0d0480",
  1591 => x"ec885187",
  1592 => x"c53fef39",
  1593 => x"80ec9451",
  1594 => x"87bc3fe6",
  1595 => x"3980eca0",
  1596 => x"5187b33f",
  1597 => x"dd3980ec",
  1598 => x"a45187aa",
  1599 => x"3fd43980",
  1600 => x"ecb05187",
  1601 => x"a13fcb39",
  1602 => x"80ecbc51",
  1603 => x"87983fc2",
  1604 => x"39fc3d0d",
  1605 => x"80f0c808",
  1606 => x"7008810a",
  1607 => x"068180c4",
  1608 => x"0c538aae",
  1609 => x"3f8adc3f",
  1610 => x"8180c408",
  1611 => x"b8f65452",
  1612 => x"7184388a",
  1613 => x"f5537281",
  1614 => x"8acc0c71",
  1615 => x"802e8298",
  1616 => x"3880e8c0",
  1617 => x"5186df3f",
  1618 => x"8c5186c0",
  1619 => x"3f80ecc8",
  1620 => x"5186d33f",
  1621 => x"8180c408",
  1622 => x"802e80f2",
  1623 => x"3880ece0",
  1624 => x"5186c33f",
  1625 => x"8180c408",
  1626 => x"802e81c4",
  1627 => x"3880f0c0",
  1628 => x"0853800b",
  1629 => x"b4140cf8",
  1630 => x"9b3ff881",
  1631 => x"c08e8053",
  1632 => x"9f0b80f0",
  1633 => x"c8085555",
  1634 => x"8180c408",
  1635 => x"802e80fb",
  1636 => x"387281ff",
  1637 => x"0684150c",
  1638 => x"818ac808",
  1639 => x"5271802e",
  1640 => x"9f38729f",
  1641 => x"2a731007",
  1642 => x"5374802e",
  1643 => x"9e38ff15",
  1644 => x"7381ff06",
  1645 => x"84160c81",
  1646 => x"8ac80853",
  1647 => x"5571e338",
  1648 => x"72812a73",
  1649 => x"9f2b0753",
  1650 => x"74e43890",
  1651 => x"be3f80ec",
  1652 => x"ec5185d2",
  1653 => x"3f80ed90",
  1654 => x"5185cb3f",
  1655 => x"b451878b",
  1656 => x"3f80eda0",
  1657 => x"5185bf3f",
  1658 => x"80eda851",
  1659 => x"85b83f81",
  1660 => x"80c408fe",
  1661 => x"f838b939",
  1662 => x"72812a73",
  1663 => x"9f2b0753",
  1664 => x"80fd5188",
  1665 => x"aa3f80f0",
  1666 => x"c8085472",
  1667 => x"81ff0684",
  1668 => x"150c818a",
  1669 => x"c8085574",
  1670 => x"802edd38",
  1671 => x"729f2a73",
  1672 => x"10075380",
  1673 => x"fd518887",
  1674 => x"3f80f0c8",
  1675 => x"0854dc39",
  1676 => x"daa73f80",
  1677 => x"f0c00853",
  1678 => x"800bb414",
  1679 => x"0cf6d53f",
  1680 => x"f881c08e",
  1681 => x"80539f0b",
  1682 => x"80f0c808",
  1683 => x"55558180",
  1684 => x"c408febd",
  1685 => x"38ffb439",
  1686 => x"89c43f80",
  1687 => x"f0bc0853",
  1688 => x"99730c81",
  1689 => x"800b8414",
  1690 => x"0c80f0b8",
  1691 => x"08549974",
  1692 => x"0c81800b",
  1693 => x"84150c81",
  1694 => x"ec0b8814",
  1695 => x"0c81900b",
  1696 => x"8c140c8c",
  1697 => x"13087081",
  1698 => x"2a810656",
  1699 => x"5474f438",
  1700 => x"8c130852",
  1701 => x"9d0b8814",
  1702 => x"0c900b8c",
  1703 => x"140c8c13",
  1704 => x"0870812a",
  1705 => x"81065654",
  1706 => x"74f4388c",
  1707 => x"13085280",
  1708 => x"c50b8814",
  1709 => x"0c80d00b",
  1710 => x"8c140c8c",
  1711 => x"13087081",
  1712 => x"2a810656",
  1713 => x"5474f438",
  1714 => x"8c130852",
  1715 => x"81ec0b88",
  1716 => x"140c8190",
  1717 => x"0b8c140c",
  1718 => x"8c130870",
  1719 => x"812a8106",
  1720 => x"565474f4",
  1721 => x"388c1308",
  1722 => x"52a10b88",
  1723 => x"140c900b",
  1724 => x"8c140c8c",
  1725 => x"13087081",
  1726 => x"2a810656",
  1727 => x"5474f438",
  1728 => x"8c130852",
  1729 => x"890b8814",
  1730 => x"0c80d00b",
  1731 => x"8c140c8c",
  1732 => x"13087081",
  1733 => x"2a810656",
  1734 => x"5474f438",
  1735 => x"8c130852",
  1736 => x"81ec0b88",
  1737 => x"140c8190",
  1738 => x"0b8c140c",
  1739 => x"8c130870",
  1740 => x"812a8106",
  1741 => x"565474f4",
  1742 => x"388c1308",
  1743 => x"52b30b88",
  1744 => x"140c900b",
  1745 => x"8c140c8c",
  1746 => x"13087081",
  1747 => x"2a810656",
  1748 => x"5474f438",
  1749 => x"8c130852",
  1750 => x"880b8814",
  1751 => x"0c80d00b",
  1752 => x"8c140c8c",
  1753 => x"13087081",
  1754 => x"2a810656",
  1755 => x"5474f438",
  1756 => x"8c130852",
  1757 => x"81ec0b88",
  1758 => x"140c8190",
  1759 => x"0b8c140c",
  1760 => x"8c130870",
  1761 => x"812a8106",
  1762 => x"565474f4",
  1763 => x"388c1308",
  1764 => x"52b40b88",
  1765 => x"140c900b",
  1766 => x"8c140c8c",
  1767 => x"13087081",
  1768 => x"2a810656",
  1769 => x"5474f438",
  1770 => x"8c130852",
  1771 => x"960b8814",
  1772 => x"0c80d00b",
  1773 => x"8c140c8c",
  1774 => x"13087081",
  1775 => x"2a810656",
  1776 => x"5474f438",
  1777 => x"8c130852",
  1778 => x"81ec0b88",
  1779 => x"140c8190",
  1780 => x"0b8c140c",
  1781 => x"8c130870",
  1782 => x"812a8106",
  1783 => x"565474f4",
  1784 => x"388c1308",
  1785 => x"52b60b88",
  1786 => x"140c900b",
  1787 => x"8c140c8c",
  1788 => x"13087081",
  1789 => x"2a810656",
  1790 => x"5474f438",
  1791 => x"8c130852",
  1792 => x"80e00b88",
  1793 => x"140c80d0",
  1794 => x"0b8c140c",
  1795 => x"8c130870",
  1796 => x"812a8106",
  1797 => x"565474f4",
  1798 => x"388c1308",
  1799 => x"5281ec0b",
  1800 => x"88140c81",
  1801 => x"900b8c14",
  1802 => x"0c8c1308",
  1803 => x"70812a81",
  1804 => x"06565474",
  1805 => x"f4388c13",
  1806 => x"085280c9",
  1807 => x"0b88140c",
  1808 => x"900b8c14",
  1809 => x"0c8c1308",
  1810 => x"70812a81",
  1811 => x"06565474",
  1812 => x"f4388c13",
  1813 => x"085281c0",
  1814 => x"0b88140c",
  1815 => x"80d00b8c",
  1816 => x"140c8c13",
  1817 => x"0870812a",
  1818 => x"81065654",
  1819 => x"74f4388c",
  1820 => x"130852f9",
  1821 => x"cc39ff3d",
  1822 => x"0d028f05",
  1823 => x"3380f0d4",
  1824 => x"0852710c",
  1825 => x"800b800c",
  1826 => x"833d0d04",
  1827 => x"ff3d0d02",
  1828 => x"8f053351",
  1829 => x"818acc08",
  1830 => x"52712d80",
  1831 => x"0881ff06",
  1832 => x"800c833d",
  1833 => x"0d04fe3d",
  1834 => x"0d747033",
  1835 => x"53537180",
  1836 => x"2e933881",
  1837 => x"13725281",
  1838 => x"8acc0853",
  1839 => x"53712d72",
  1840 => x"335271ef",
  1841 => x"38843d0d",
  1842 => x"04f43d0d",
  1843 => x"7f028405",
  1844 => x"bb053355",
  1845 => x"57880b8c",
  1846 => x"3d5a5a89",
  1847 => x"5380edf8",
  1848 => x"5278518a",
  1849 => x"b33f737a",
  1850 => x"2e80fa38",
  1851 => x"79567390",
  1852 => x"2e80e738",
  1853 => x"02a70558",
  1854 => x"768f0654",
  1855 => x"738926bf",
  1856 => x"387518b0",
  1857 => x"15555573",
  1858 => x"75347684",
  1859 => x"2aff1770",
  1860 => x"81ff0658",
  1861 => x"555775e0",
  1862 => x"38791955",
  1863 => x"75753478",
  1864 => x"70335555",
  1865 => x"73802e93",
  1866 => x"38811574",
  1867 => x"52818acc",
  1868 => x"08575575",
  1869 => x"2d743354",
  1870 => x"73ef388e",
  1871 => x"3d0d0475",
  1872 => x"18b71555",
  1873 => x"55737534",
  1874 => x"76842aff",
  1875 => x"177081ff",
  1876 => x"06585557",
  1877 => x"75ffa138",
  1878 => x"c0398470",
  1879 => x"575a02a7",
  1880 => x"0558ff94",
  1881 => x"39827057",
  1882 => x"5af439f2",
  1883 => x"3d0d608c",
  1884 => x"3d705b5b",
  1885 => x"53807356",
  1886 => x"57767324",
  1887 => x"81803878",
  1888 => x"17548a52",
  1889 => x"745184e2",
  1890 => x"3f8008b0",
  1891 => x"05537274",
  1892 => x"34811757",
  1893 => x"8a527451",
  1894 => x"84ab3f80",
  1895 => x"08558008",
  1896 => x"de388008",
  1897 => x"779f2a18",
  1898 => x"70812c5a",
  1899 => x"56568078",
  1900 => x"259e3878",
  1901 => x"17ff0555",
  1902 => x"75197033",
  1903 => x"55537433",
  1904 => x"73347375",
  1905 => x"348116ff",
  1906 => x"16565677",
  1907 => x"7624e938",
  1908 => x"76195680",
  1909 => x"76347681",
  1910 => x"ff067a70",
  1911 => x"33555654",
  1912 => x"72802e93",
  1913 => x"38811573",
  1914 => x"52818acc",
  1915 => x"08585576",
  1916 => x"2d743353",
  1917 => x"72ef3873",
  1918 => x"800c903d",
  1919 => x"0d04ad7a",
  1920 => x"3402a905",
  1921 => x"73307119",
  1922 => x"5656598a",
  1923 => x"52745183",
  1924 => x"d93f8008",
  1925 => x"b0055372",
  1926 => x"74348117",
  1927 => x"578a5274",
  1928 => x"5183a23f",
  1929 => x"80085580",
  1930 => x"08fed438",
  1931 => x"fef439fd",
  1932 => x"3d0d80f0",
  1933 => x"cc0876b2",
  1934 => x"e4299412",
  1935 => x"0c54850b",
  1936 => x"98150c98",
  1937 => x"14087081",
  1938 => x"06515372",
  1939 => x"f638853d",
  1940 => x"0d04803d",
  1941 => x"0d80f0cc",
  1942 => x"0851870b",
  1943 => x"84120cff",
  1944 => x"0bb4120c",
  1945 => x"a70bb812",
  1946 => x"0c87e80b",
  1947 => x"a4120ca7",
  1948 => x"0ba8120c",
  1949 => x"b2e40b94",
  1950 => x"120c870b",
  1951 => x"98120c82",
  1952 => x"3d0d0480",
  1953 => x"3d0d80f0",
  1954 => x"d00851b8",
  1955 => x"0b8c120c",
  1956 => x"830b8812",
  1957 => x"0c823d0d",
  1958 => x"04803d0d",
  1959 => x"80f0d008",
  1960 => x"84110881",
  1961 => x"06800c51",
  1962 => x"823d0d04",
  1963 => x"ff3d0d80",
  1964 => x"f0d00852",
  1965 => x"84120870",
  1966 => x"81065151",
  1967 => x"70802ef4",
  1968 => x"38710870",
  1969 => x"81ff0680",
  1970 => x"0c51833d",
  1971 => x"0d04fe3d",
  1972 => x"0d029305",
  1973 => x"3353728a",
  1974 => x"2e9c3880",
  1975 => x"f0d00852",
  1976 => x"84120870",
  1977 => x"892a7081",
  1978 => x"06515151",
  1979 => x"70f23872",
  1980 => x"720c843d",
  1981 => x"0d0480f0",
  1982 => x"d0085284",
  1983 => x"12087089",
  1984 => x"2a708106",
  1985 => x"51515170",
  1986 => x"f2388d72",
  1987 => x"0c841208",
  1988 => x"70892a70",
  1989 => x"81065151",
  1990 => x"5170c538",
  1991 => x"d239803d",
  1992 => x"0d80f0c4",
  1993 => x"0851800b",
  1994 => x"84120c83",
  1995 => x"fe800b88",
  1996 => x"120c800b",
  1997 => x"818ad034",
  1998 => x"800b818a",
  1999 => x"d434823d",
  2000 => x"0d04fa3d",
  2001 => x"0d02a305",
  2002 => x"3380f0c4",
  2003 => x"08818ad0",
  2004 => x"337081ff",
  2005 => x"06701010",
  2006 => x"11818ad4",
  2007 => x"337081ff",
  2008 => x"06729029",
  2009 => x"1170882b",
  2010 => x"7807770c",
  2011 => x"535b5b55",
  2012 => x"55595454",
  2013 => x"738a2e98",
  2014 => x"387480cf",
  2015 => x"2e923873",
  2016 => x"8c2ea438",
  2017 => x"81165372",
  2018 => x"818ad434",
  2019 => x"883d0d04",
  2020 => x"71a326a3",
  2021 => x"38811752",
  2022 => x"71818ad0",
  2023 => x"34800b81",
  2024 => x"8ad43488",
  2025 => x"3d0d0480",
  2026 => x"5271882b",
  2027 => x"730c8112",
  2028 => x"52979072",
  2029 => x"26f33880",
  2030 => x"0b818ad0",
  2031 => x"34800b81",
  2032 => x"8ad434df",
  2033 => x"398c0802",
  2034 => x"8c0cfd3d",
  2035 => x"0d80538c",
  2036 => x"088c0508",
  2037 => x"528c0888",
  2038 => x"05085182",
  2039 => x"de3f8008",
  2040 => x"70800c54",
  2041 => x"853d0d8c",
  2042 => x"0c048c08",
  2043 => x"028c0cfd",
  2044 => x"3d0d8153",
  2045 => x"8c088c05",
  2046 => x"08528c08",
  2047 => x"88050851",
  2048 => x"82b93f80",
  2049 => x"0870800c",
  2050 => x"54853d0d",
  2051 => x"8c0c048c",
  2052 => x"08028c0c",
  2053 => x"f93d0d80",
  2054 => x"0b8c08fc",
  2055 => x"050c8c08",
  2056 => x"88050880",
  2057 => x"25ab388c",
  2058 => x"08880508",
  2059 => x"308c0888",
  2060 => x"050c800b",
  2061 => x"8c08f405",
  2062 => x"0c8c08fc",
  2063 => x"05088838",
  2064 => x"810b8c08",
  2065 => x"f4050c8c",
  2066 => x"08f40508",
  2067 => x"8c08fc05",
  2068 => x"0c8c088c",
  2069 => x"05088025",
  2070 => x"ab388c08",
  2071 => x"8c050830",
  2072 => x"8c088c05",
  2073 => x"0c800b8c",
  2074 => x"08f0050c",
  2075 => x"8c08fc05",
  2076 => x"08883881",
  2077 => x"0b8c08f0",
  2078 => x"050c8c08",
  2079 => x"f005088c",
  2080 => x"08fc050c",
  2081 => x"80538c08",
  2082 => x"8c050852",
  2083 => x"8c088805",
  2084 => x"085181a7",
  2085 => x"3f800870",
  2086 => x"8c08f805",
  2087 => x"0c548c08",
  2088 => x"fc050880",
  2089 => x"2e8c388c",
  2090 => x"08f80508",
  2091 => x"308c08f8",
  2092 => x"050c8c08",
  2093 => x"f8050870",
  2094 => x"800c5489",
  2095 => x"3d0d8c0c",
  2096 => x"048c0802",
  2097 => x"8c0cfb3d",
  2098 => x"0d800b8c",
  2099 => x"08fc050c",
  2100 => x"8c088805",
  2101 => x"08802593",
  2102 => x"388c0888",
  2103 => x"0508308c",
  2104 => x"0888050c",
  2105 => x"810b8c08",
  2106 => x"fc050c8c",
  2107 => x"088c0508",
  2108 => x"80258c38",
  2109 => x"8c088c05",
  2110 => x"08308c08",
  2111 => x"8c050c81",
  2112 => x"538c088c",
  2113 => x"0508528c",
  2114 => x"08880508",
  2115 => x"51ad3f80",
  2116 => x"08708c08",
  2117 => x"f8050c54",
  2118 => x"8c08fc05",
  2119 => x"08802e8c",
  2120 => x"388c08f8",
  2121 => x"0508308c",
  2122 => x"08f8050c",
  2123 => x"8c08f805",
  2124 => x"0870800c",
  2125 => x"54873d0d",
  2126 => x"8c0c048c",
  2127 => x"08028c0c",
  2128 => x"fd3d0d81",
  2129 => x"0b8c08fc",
  2130 => x"050c800b",
  2131 => x"8c08f805",
  2132 => x"0c8c088c",
  2133 => x"05088c08",
  2134 => x"88050827",
  2135 => x"ac388c08",
  2136 => x"fc050880",
  2137 => x"2ea33880",
  2138 => x"0b8c088c",
  2139 => x"05082499",
  2140 => x"388c088c",
  2141 => x"0508108c",
  2142 => x"088c050c",
  2143 => x"8c08fc05",
  2144 => x"08108c08",
  2145 => x"fc050cc9",
  2146 => x"398c08fc",
  2147 => x"0508802e",
  2148 => x"80c9388c",
  2149 => x"088c0508",
  2150 => x"8c088805",
  2151 => x"0826a138",
  2152 => x"8c088805",
  2153 => x"088c088c",
  2154 => x"0508318c",
  2155 => x"0888050c",
  2156 => x"8c08f805",
  2157 => x"088c08fc",
  2158 => x"0508078c",
  2159 => x"08f8050c",
  2160 => x"8c08fc05",
  2161 => x"08812a8c",
  2162 => x"08fc050c",
  2163 => x"8c088c05",
  2164 => x"08812a8c",
  2165 => x"088c050c",
  2166 => x"ffaf398c",
  2167 => x"08900508",
  2168 => x"802e8f38",
  2169 => x"8c088805",
  2170 => x"08708c08",
  2171 => x"f4050c51",
  2172 => x"8d398c08",
  2173 => x"f8050870",
  2174 => x"8c08f405",
  2175 => x"0c518c08",
  2176 => x"f4050880",
  2177 => x"0c853d0d",
  2178 => x"8c0c0480",
  2179 => x"3d0d8651",
  2180 => x"84963f81",
  2181 => x"519f873f",
  2182 => x"fc3d0d76",
  2183 => x"70797b55",
  2184 => x"5555558f",
  2185 => x"72278c38",
  2186 => x"72750783",
  2187 => x"06517080",
  2188 => x"2ea738ff",
  2189 => x"125271ff",
  2190 => x"2e983872",
  2191 => x"70810554",
  2192 => x"33747081",
  2193 => x"055634ff",
  2194 => x"125271ff",
  2195 => x"2e098106",
  2196 => x"ea387480",
  2197 => x"0c863d0d",
  2198 => x"04745172",
  2199 => x"70840554",
  2200 => x"08717084",
  2201 => x"05530c72",
  2202 => x"70840554",
  2203 => x"08717084",
  2204 => x"05530c72",
  2205 => x"70840554",
  2206 => x"08717084",
  2207 => x"05530c72",
  2208 => x"70840554",
  2209 => x"08717084",
  2210 => x"05530cf0",
  2211 => x"1252718f",
  2212 => x"26c93883",
  2213 => x"72279538",
  2214 => x"72708405",
  2215 => x"54087170",
  2216 => x"8405530c",
  2217 => x"fc125271",
  2218 => x"8326ed38",
  2219 => x"7054ff83",
  2220 => x"39fd3d0d",
  2221 => x"755384d8",
  2222 => x"1308802e",
  2223 => x"8a388053",
  2224 => x"72800c85",
  2225 => x"3d0d0481",
  2226 => x"80527251",
  2227 => x"8a883f80",
  2228 => x"0884d814",
  2229 => x"0cff5380",
  2230 => x"08802ee4",
  2231 => x"38800854",
  2232 => x"9f538074",
  2233 => x"70840556",
  2234 => x"0cff1353",
  2235 => x"807324ce",
  2236 => x"38807470",
  2237 => x"8405560c",
  2238 => x"ff135372",
  2239 => x"8025e338",
  2240 => x"ffbc39fd",
  2241 => x"3d0d7577",
  2242 => x"55539f74",
  2243 => x"278d3896",
  2244 => x"730cff52",
  2245 => x"71800c85",
  2246 => x"3d0d0484",
  2247 => x"d8130852",
  2248 => x"71802e93",
  2249 => x"38731010",
  2250 => x"12700879",
  2251 => x"720c5152",
  2252 => x"71800c85",
  2253 => x"3d0d0472",
  2254 => x"51fef63f",
  2255 => x"ff528008",
  2256 => x"d33884d8",
  2257 => x"13087410",
  2258 => x"10117008",
  2259 => x"7a720c51",
  2260 => x"5152dd39",
  2261 => x"f93d0d79",
  2262 => x"7b585676",
  2263 => x"9f2680e8",
  2264 => x"3884d816",
  2265 => x"08547380",
  2266 => x"2eaa3876",
  2267 => x"10101470",
  2268 => x"08555573",
  2269 => x"802eba38",
  2270 => x"80587381",
  2271 => x"2e8f3873",
  2272 => x"ff2ea338",
  2273 => x"80750c76",
  2274 => x"51732d80",
  2275 => x"5877800c",
  2276 => x"893d0d04",
  2277 => x"7551fe99",
  2278 => x"3fff5880",
  2279 => x"08ef3884",
  2280 => x"d8160854",
  2281 => x"c6399676",
  2282 => x"0c810b80",
  2283 => x"0c893d0d",
  2284 => x"04755181",
  2285 => x"ed3f7653",
  2286 => x"80085275",
  2287 => x"5181ad3f",
  2288 => x"8008800c",
  2289 => x"893d0d04",
  2290 => x"96760cff",
  2291 => x"0b800c89",
  2292 => x"3d0d04fc",
  2293 => x"3d0d7678",
  2294 => x"5653ff54",
  2295 => x"749f26b1",
  2296 => x"3884d813",
  2297 => x"08527180",
  2298 => x"2eae3874",
  2299 => x"10101270",
  2300 => x"08535381",
  2301 => x"5471802e",
  2302 => x"98388254",
  2303 => x"71ff2e91",
  2304 => x"38835471",
  2305 => x"812e8a38",
  2306 => x"80730c74",
  2307 => x"51712d80",
  2308 => x"5473800c",
  2309 => x"863d0d04",
  2310 => x"7251fd95",
  2311 => x"3f8008f1",
  2312 => x"3884d813",
  2313 => x"0852c439",
  2314 => x"ff3d0d73",
  2315 => x"5280f0d8",
  2316 => x"0851fea0",
  2317 => x"3f833d0d",
  2318 => x"04fe3d0d",
  2319 => x"75537452",
  2320 => x"80f0d808",
  2321 => x"51fdbc3f",
  2322 => x"843d0d04",
  2323 => x"803d0d80",
  2324 => x"f0d80851",
  2325 => x"fcdb3f82",
  2326 => x"3d0d04ff",
  2327 => x"3d0d7352",
  2328 => x"80f0d808",
  2329 => x"51feec3f",
  2330 => x"833d0d04",
  2331 => x"fc3d0d80",
  2332 => x"0b818ae0",
  2333 => x"0c785277",
  2334 => x"5199973f",
  2335 => x"80085480",
  2336 => x"08ff2e88",
  2337 => x"3873800c",
  2338 => x"863d0d04",
  2339 => x"818ae008",
  2340 => x"5574802e",
  2341 => x"f0387675",
  2342 => x"710c5373",
  2343 => x"800c863d",
  2344 => x"0d0498e9",
  2345 => x"3f04fc3d",
  2346 => x"0d767079",
  2347 => x"70730783",
  2348 => x"06545454",
  2349 => x"557080c3",
  2350 => x"38717008",
  2351 => x"700970f7",
  2352 => x"fbfdff13",
  2353 => x"0670f884",
  2354 => x"82818006",
  2355 => x"51515353",
  2356 => x"5470a638",
  2357 => x"84147274",
  2358 => x"70840556",
  2359 => x"0c700870",
  2360 => x"0970f7fb",
  2361 => x"fdff1306",
  2362 => x"70f88482",
  2363 => x"81800651",
  2364 => x"51535354",
  2365 => x"70802edc",
  2366 => x"38735271",
  2367 => x"70810553",
  2368 => x"33517073",
  2369 => x"70810555",
  2370 => x"3470f038",
  2371 => x"74800c86",
  2372 => x"3d0d04fd",
  2373 => x"3d0d7570",
  2374 => x"71830653",
  2375 => x"555270b8",
  2376 => x"38717008",
  2377 => x"7009f7fb",
  2378 => x"fdff1206",
  2379 => x"70f88482",
  2380 => x"81800651",
  2381 => x"51525370",
  2382 => x"9d388413",
  2383 => x"70087009",
  2384 => x"f7fbfdff",
  2385 => x"120670f8",
  2386 => x"84828180",
  2387 => x"06515152",
  2388 => x"5370802e",
  2389 => x"e5387252",
  2390 => x"71335170",
  2391 => x"802e8a38",
  2392 => x"81127033",
  2393 => x"525270f8",
  2394 => x"38717431",
  2395 => x"800c853d",
  2396 => x"0d04fa3d",
  2397 => x"0d787a7c",
  2398 => x"70545555",
  2399 => x"5272802e",
  2400 => x"80d93871",
  2401 => x"74078306",
  2402 => x"5170802e",
  2403 => x"80d438ff",
  2404 => x"135372ff",
  2405 => x"2eb13871",
  2406 => x"33743356",
  2407 => x"5174712e",
  2408 => x"098106a9",
  2409 => x"3872802e",
  2410 => x"81873870",
  2411 => x"81ff0651",
  2412 => x"70802e80",
  2413 => x"fc388112",
  2414 => x"8115ff15",
  2415 => x"55555272",
  2416 => x"ff2e0981",
  2417 => x"06d13871",
  2418 => x"33743356",
  2419 => x"517081ff",
  2420 => x"067581ff",
  2421 => x"06717131",
  2422 => x"51525270",
  2423 => x"800c883d",
  2424 => x"0d047174",
  2425 => x"57558373",
  2426 => x"27883871",
  2427 => x"0874082e",
  2428 => x"88387476",
  2429 => x"5552ff97",
  2430 => x"39fc1353",
  2431 => x"72802eb1",
  2432 => x"38740870",
  2433 => x"09f7fbfd",
  2434 => x"ff120670",
  2435 => x"f8848281",
  2436 => x"80065151",
  2437 => x"51709a38",
  2438 => x"84158417",
  2439 => x"57558373",
  2440 => x"27d03874",
  2441 => x"0876082e",
  2442 => x"d0387476",
  2443 => x"5552fedf",
  2444 => x"39800b80",
  2445 => x"0c883d0d",
  2446 => x"04f33d0d",
  2447 => x"60626472",
  2448 => x"5a5a5d5d",
  2449 => x"805e7670",
  2450 => x"81055833",
  2451 => x"80ee8511",
  2452 => x"3370832a",
  2453 => x"70810651",
  2454 => x"55555672",
  2455 => x"e93875ad",
  2456 => x"2e81ff38",
  2457 => x"75ab2e81",
  2458 => x"fb387730",
  2459 => x"70790780",
  2460 => x"25799032",
  2461 => x"70307072",
  2462 => x"07802573",
  2463 => x"07535757",
  2464 => x"51537280",
  2465 => x"2e873875",
  2466 => x"b02e81e2",
  2467 => x"38778a38",
  2468 => x"885875b0",
  2469 => x"2e83388a",
  2470 => x"587752ff",
  2471 => x"51f2a63f",
  2472 => x"80087853",
  2473 => x"5aff51f2",
  2474 => x"c13f8008",
  2475 => x"5b80705a",
  2476 => x"5580ee85",
  2477 => x"16337082",
  2478 => x"2a708106",
  2479 => x"51545472",
  2480 => x"802e80c1",
  2481 => x"38d01656",
  2482 => x"75782580",
  2483 => x"d7388079",
  2484 => x"24757b26",
  2485 => x"07537293",
  2486 => x"38747a2e",
  2487 => x"80eb387a",
  2488 => x"762580ed",
  2489 => x"3872802e",
  2490 => x"80e738ff",
  2491 => x"77708105",
  2492 => x"59335759",
  2493 => x"80ee8516",
  2494 => x"3370822a",
  2495 => x"70810651",
  2496 => x"545472c1",
  2497 => x"38738306",
  2498 => x"5372802e",
  2499 => x"97387381",
  2500 => x"06c91755",
  2501 => x"53728538",
  2502 => x"ffa91654",
  2503 => x"73567776",
  2504 => x"24ffab38",
  2505 => x"80792481",
  2506 => x"89387d80",
  2507 => x"2e843874",
  2508 => x"30557b80",
  2509 => x"2e8c38ff",
  2510 => x"17537883",
  2511 => x"387c5372",
  2512 => x"7c0c7480",
  2513 => x"0c8f3d0d",
  2514 => x"04815375",
  2515 => x"7b24ff95",
  2516 => x"38817579",
  2517 => x"29177870",
  2518 => x"81055a33",
  2519 => x"585659ff",
  2520 => x"9339815e",
  2521 => x"76708105",
  2522 => x"583356fd",
  2523 => x"fd398077",
  2524 => x"33545472",
  2525 => x"80f82e80",
  2526 => x"c3387280",
  2527 => x"d8327030",
  2528 => x"70802576",
  2529 => x"07515153",
  2530 => x"72802efe",
  2531 => x"80388117",
  2532 => x"33821858",
  2533 => x"56907053",
  2534 => x"58ff51f0",
  2535 => x"a83f8008",
  2536 => x"78535aff",
  2537 => x"51f0c33f",
  2538 => x"80085b80",
  2539 => x"705a55fe",
  2540 => x"8039ff60",
  2541 => x"5455a273",
  2542 => x"0cfef739",
  2543 => x"8154ffba",
  2544 => x"39fd3d0d",
  2545 => x"77547653",
  2546 => x"755280f0",
  2547 => x"d80851fc",
  2548 => x"e83f853d",
  2549 => x"0d04f33d",
  2550 => x"0d7f618b",
  2551 => x"1170f806",
  2552 => x"5c55555e",
  2553 => x"72962683",
  2554 => x"38905980",
  2555 => x"7924747a",
  2556 => x"26075380",
  2557 => x"5472742e",
  2558 => x"09810680",
  2559 => x"cb387d51",
  2560 => x"8bca3f78",
  2561 => x"83f72680",
  2562 => x"c6387883",
  2563 => x"2a701010",
  2564 => x"1080f894",
  2565 => x"058c1108",
  2566 => x"59595a76",
  2567 => x"782e83b0",
  2568 => x"38841708",
  2569 => x"fc06568c",
  2570 => x"17088818",
  2571 => x"08718c12",
  2572 => x"0c88120c",
  2573 => x"58751784",
  2574 => x"11088107",
  2575 => x"84120c53",
  2576 => x"7d518b89",
  2577 => x"3f881754",
  2578 => x"73800c8f",
  2579 => x"3d0d0478",
  2580 => x"892a7983",
  2581 => x"2a5b5372",
  2582 => x"802ebf38",
  2583 => x"78862ab8",
  2584 => x"055a8473",
  2585 => x"27b43880",
  2586 => x"db135a94",
  2587 => x"7327ab38",
  2588 => x"788c2a80",
  2589 => x"ee055a80",
  2590 => x"d473279e",
  2591 => x"38788f2a",
  2592 => x"80f7055a",
  2593 => x"82d47327",
  2594 => x"91387892",
  2595 => x"2a80fc05",
  2596 => x"5a8ad473",
  2597 => x"27843880",
  2598 => x"fe5a7910",
  2599 => x"101080f8",
  2600 => x"94058c11",
  2601 => x"08585576",
  2602 => x"752ea338",
  2603 => x"841708fc",
  2604 => x"06707a31",
  2605 => x"5556738f",
  2606 => x"2488d538",
  2607 => x"738025fe",
  2608 => x"e6388c17",
  2609 => x"08577675",
  2610 => x"2e098106",
  2611 => x"df38811a",
  2612 => x"5a80f8a4",
  2613 => x"08577680",
  2614 => x"f89c2e82",
  2615 => x"c0388417",
  2616 => x"08fc0670",
  2617 => x"7a315556",
  2618 => x"738f2481",
  2619 => x"f93880f8",
  2620 => x"9c0b80f8",
  2621 => x"a80c80f8",
  2622 => x"9c0b80f8",
  2623 => x"a40c7380",
  2624 => x"25feb238",
  2625 => x"83ff7627",
  2626 => x"83df3875",
  2627 => x"892a7683",
  2628 => x"2a555372",
  2629 => x"802ebf38",
  2630 => x"75862ab8",
  2631 => x"05548473",
  2632 => x"27b43880",
  2633 => x"db135494",
  2634 => x"7327ab38",
  2635 => x"758c2a80",
  2636 => x"ee055480",
  2637 => x"d473279e",
  2638 => x"38758f2a",
  2639 => x"80f70554",
  2640 => x"82d47327",
  2641 => x"91387592",
  2642 => x"2a80fc05",
  2643 => x"548ad473",
  2644 => x"27843880",
  2645 => x"fe547310",
  2646 => x"101080f8",
  2647 => x"94058811",
  2648 => x"08565874",
  2649 => x"782e86cf",
  2650 => x"38841508",
  2651 => x"fc065375",
  2652 => x"73278d38",
  2653 => x"88150855",
  2654 => x"74782e09",
  2655 => x"8106ea38",
  2656 => x"8c150880",
  2657 => x"f8940b84",
  2658 => x"0508718c",
  2659 => x"1a0c7688",
  2660 => x"1a0c7888",
  2661 => x"130c788c",
  2662 => x"180c5d58",
  2663 => x"7953807a",
  2664 => x"2483e638",
  2665 => x"72822c81",
  2666 => x"712b5c53",
  2667 => x"7a7c2681",
  2668 => x"98387b7b",
  2669 => x"06537282",
  2670 => x"f13879fc",
  2671 => x"0684055a",
  2672 => x"7a10707d",
  2673 => x"06545b72",
  2674 => x"82e03884",
  2675 => x"1a5af139",
  2676 => x"88178c11",
  2677 => x"08585876",
  2678 => x"782e0981",
  2679 => x"06fcc238",
  2680 => x"821a5afd",
  2681 => x"ec397817",
  2682 => x"79810784",
  2683 => x"190c7080",
  2684 => x"f8a80c70",
  2685 => x"80f8a40c",
  2686 => x"80f89c0b",
  2687 => x"8c120c8c",
  2688 => x"11088812",
  2689 => x"0c748107",
  2690 => x"84120c74",
  2691 => x"1175710c",
  2692 => x"51537d51",
  2693 => x"87b73f88",
  2694 => x"1754fcac",
  2695 => x"3980f894",
  2696 => x"0b840508",
  2697 => x"7a545c79",
  2698 => x"8025fef8",
  2699 => x"3882da39",
  2700 => x"7a097c06",
  2701 => x"7080f894",
  2702 => x"0b84050c",
  2703 => x"5c7a105b",
  2704 => x"7a7c2685",
  2705 => x"387a85b8",
  2706 => x"3880f894",
  2707 => x"0b880508",
  2708 => x"70841208",
  2709 => x"fc06707c",
  2710 => x"317c7226",
  2711 => x"8f722507",
  2712 => x"57575c5d",
  2713 => x"5572802e",
  2714 => x"80db3879",
  2715 => x"7a1680f8",
  2716 => x"8c081b90",
  2717 => x"115a5557",
  2718 => x"5b80f888",
  2719 => x"08ff2e88",
  2720 => x"38a08f13",
  2721 => x"e0800657",
  2722 => x"76527d51",
  2723 => x"86c03f80",
  2724 => x"08548008",
  2725 => x"ff2e9038",
  2726 => x"80087627",
  2727 => x"82993874",
  2728 => x"80f8942e",
  2729 => x"82913880",
  2730 => x"f8940b88",
  2731 => x"05085584",
  2732 => x"1508fc06",
  2733 => x"707a317a",
  2734 => x"72268f72",
  2735 => x"25075255",
  2736 => x"537283e6",
  2737 => x"38747981",
  2738 => x"0784170c",
  2739 => x"79167080",
  2740 => x"f8940b88",
  2741 => x"050c7581",
  2742 => x"0784120c",
  2743 => x"547e5257",
  2744 => x"85eb3f88",
  2745 => x"1754fae0",
  2746 => x"3975832a",
  2747 => x"70545480",
  2748 => x"7424819b",
  2749 => x"3872822c",
  2750 => x"81712b80",
  2751 => x"f8980807",
  2752 => x"7080f894",
  2753 => x"0b84050c",
  2754 => x"75101010",
  2755 => x"80f89405",
  2756 => x"88110858",
  2757 => x"5a5d5377",
  2758 => x"8c180c74",
  2759 => x"88180c76",
  2760 => x"88190c76",
  2761 => x"8c160cfc",
  2762 => x"f339797a",
  2763 => x"10101080",
  2764 => x"f8940570",
  2765 => x"57595d8c",
  2766 => x"15085776",
  2767 => x"752ea338",
  2768 => x"841708fc",
  2769 => x"06707a31",
  2770 => x"5556738f",
  2771 => x"2483ca38",
  2772 => x"73802584",
  2773 => x"81388c17",
  2774 => x"08577675",
  2775 => x"2e098106",
  2776 => x"df388815",
  2777 => x"811b7083",
  2778 => x"06555b55",
  2779 => x"72c9387c",
  2780 => x"83065372",
  2781 => x"802efdb8",
  2782 => x"38ff1df8",
  2783 => x"19595d88",
  2784 => x"1808782e",
  2785 => x"ea38fdb5",
  2786 => x"39831a53",
  2787 => x"fc963983",
  2788 => x"1470822c",
  2789 => x"81712b80",
  2790 => x"f8980807",
  2791 => x"7080f894",
  2792 => x"0b84050c",
  2793 => x"76101010",
  2794 => x"80f89405",
  2795 => x"88110859",
  2796 => x"5b5e5153",
  2797 => x"fee13980",
  2798 => x"f7d80817",
  2799 => x"58800876",
  2800 => x"2e818d38",
  2801 => x"80f88808",
  2802 => x"ff2e83ec",
  2803 => x"38737631",
  2804 => x"1880f7d8",
  2805 => x"0c738706",
  2806 => x"70575372",
  2807 => x"802e8838",
  2808 => x"88733170",
  2809 => x"15555676",
  2810 => x"149fff06",
  2811 => x"a0807131",
  2812 => x"1770547f",
  2813 => x"53575383",
  2814 => x"d53f8008",
  2815 => x"538008ff",
  2816 => x"2e81a038",
  2817 => x"80f7d808",
  2818 => x"167080f7",
  2819 => x"d80c7475",
  2820 => x"80f8940b",
  2821 => x"88050c74",
  2822 => x"76311870",
  2823 => x"81075155",
  2824 => x"56587b80",
  2825 => x"f8942e83",
  2826 => x"9c38798f",
  2827 => x"2682cb38",
  2828 => x"810b8415",
  2829 => x"0c841508",
  2830 => x"fc06707a",
  2831 => x"317a7226",
  2832 => x"8f722507",
  2833 => x"52555372",
  2834 => x"802efcf9",
  2835 => x"3880db39",
  2836 => x"80089fff",
  2837 => x"065372fe",
  2838 => x"eb387780",
  2839 => x"f7d80c80",
  2840 => x"f8940b88",
  2841 => x"05087b18",
  2842 => x"81078412",
  2843 => x"0c5580f8",
  2844 => x"84087827",
  2845 => x"86387780",
  2846 => x"f8840c80",
  2847 => x"f8800878",
  2848 => x"27fcac38",
  2849 => x"7780f880",
  2850 => x"0c841508",
  2851 => x"fc06707a",
  2852 => x"317a7226",
  2853 => x"8f722507",
  2854 => x"52555372",
  2855 => x"802efca5",
  2856 => x"38883980",
  2857 => x"745456fe",
  2858 => x"db397d51",
  2859 => x"829f3f80",
  2860 => x"0b800c8f",
  2861 => x"3d0d0473",
  2862 => x"53807424",
  2863 => x"a9387282",
  2864 => x"2c81712b",
  2865 => x"80f89808",
  2866 => x"077080f8",
  2867 => x"940b8405",
  2868 => x"0c5d5377",
  2869 => x"8c180c74",
  2870 => x"88180c76",
  2871 => x"88190c76",
  2872 => x"8c160cf9",
  2873 => x"b7398314",
  2874 => x"70822c81",
  2875 => x"712b80f8",
  2876 => x"98080770",
  2877 => x"80f8940b",
  2878 => x"84050c5e",
  2879 => x"5153d439",
  2880 => x"7b7b0653",
  2881 => x"72fca338",
  2882 => x"841a7b10",
  2883 => x"5c5af139",
  2884 => x"ff1a8111",
  2885 => x"515af7b9",
  2886 => x"39781779",
  2887 => x"81078419",
  2888 => x"0c8c1808",
  2889 => x"88190871",
  2890 => x"8c120c88",
  2891 => x"120c5970",
  2892 => x"80f8a80c",
  2893 => x"7080f8a4",
  2894 => x"0c80f89c",
  2895 => x"0b8c120c",
  2896 => x"8c110888",
  2897 => x"120c7481",
  2898 => x"0784120c",
  2899 => x"74117571",
  2900 => x"0c5153f9",
  2901 => x"bd397517",
  2902 => x"84110881",
  2903 => x"0784120c",
  2904 => x"538c1708",
  2905 => x"88180871",
  2906 => x"8c120c88",
  2907 => x"120c587d",
  2908 => x"5180da3f",
  2909 => x"881754f5",
  2910 => x"cf397284",
  2911 => x"150cf41a",
  2912 => x"f8067084",
  2913 => x"1e088106",
  2914 => x"07841e0c",
  2915 => x"701d545b",
  2916 => x"850b8414",
  2917 => x"0c850b88",
  2918 => x"140c8f7b",
  2919 => x"27fdcf38",
  2920 => x"881c527d",
  2921 => x"5182903f",
  2922 => x"80f8940b",
  2923 => x"88050880",
  2924 => x"f7d80859",
  2925 => x"55fdb739",
  2926 => x"7780f7d8",
  2927 => x"0c7380f8",
  2928 => x"880cfc91",
  2929 => x"39728415",
  2930 => x"0cfda339",
  2931 => x"0404fd3d",
  2932 => x"0d800b81",
  2933 => x"8ae00c76",
  2934 => x"5186cc3f",
  2935 => x"80085380",
  2936 => x"08ff2e88",
  2937 => x"3872800c",
  2938 => x"853d0d04",
  2939 => x"818ae008",
  2940 => x"5473802e",
  2941 => x"f0387574",
  2942 => x"710c5272",
  2943 => x"800c853d",
  2944 => x"0d04fb3d",
  2945 => x"0d777052",
  2946 => x"56c23f80",
  2947 => x"f8940b88",
  2948 => x"05088411",
  2949 => x"08fc0670",
  2950 => x"7b319fef",
  2951 => x"05e08006",
  2952 => x"e0800556",
  2953 => x"5653a080",
  2954 => x"74249438",
  2955 => x"80527551",
  2956 => x"ff9c3f80",
  2957 => x"f89c0815",
  2958 => x"53728008",
  2959 => x"2e8f3875",
  2960 => x"51ff8a3f",
  2961 => x"80537280",
  2962 => x"0c873d0d",
  2963 => x"04733052",
  2964 => x"7551fefa",
  2965 => x"3f8008ff",
  2966 => x"2ea83880",
  2967 => x"f8940b88",
  2968 => x"05087575",
  2969 => x"31810784",
  2970 => x"120c5380",
  2971 => x"f7d80874",
  2972 => x"3180f7d8",
  2973 => x"0c7551fe",
  2974 => x"d43f810b",
  2975 => x"800c873d",
  2976 => x"0d048052",
  2977 => x"7551fec6",
  2978 => x"3f80f894",
  2979 => x"0b880508",
  2980 => x"80087131",
  2981 => x"56538f75",
  2982 => x"25ffa438",
  2983 => x"800880f8",
  2984 => x"88083180",
  2985 => x"f7d80c74",
  2986 => x"81078414",
  2987 => x"0c7551fe",
  2988 => x"9c3f8053",
  2989 => x"ff9039f6",
  2990 => x"3d0d7c7e",
  2991 => x"545b7280",
  2992 => x"2e828338",
  2993 => x"7a51fe84",
  2994 => x"3ff81384",
  2995 => x"110870fe",
  2996 => x"06701384",
  2997 => x"1108fc06",
  2998 => x"5d585954",
  2999 => x"5880f89c",
  3000 => x"08752e82",
  3001 => x"de387884",
  3002 => x"160c8073",
  3003 => x"8106545a",
  3004 => x"727a2e81",
  3005 => x"d5387815",
  3006 => x"84110881",
  3007 => x"06515372",
  3008 => x"a0387817",
  3009 => x"577981e6",
  3010 => x"38881508",
  3011 => x"537280f8",
  3012 => x"9c2e82f9",
  3013 => x"388c1508",
  3014 => x"708c150c",
  3015 => x"7388120c",
  3016 => x"56768107",
  3017 => x"84190c76",
  3018 => x"1877710c",
  3019 => x"53798191",
  3020 => x"3883ff77",
  3021 => x"2781c838",
  3022 => x"76892a77",
  3023 => x"832a5653",
  3024 => x"72802ebf",
  3025 => x"3876862a",
  3026 => x"b8055584",
  3027 => x"7327b438",
  3028 => x"80db1355",
  3029 => x"947327ab",
  3030 => x"38768c2a",
  3031 => x"80ee0555",
  3032 => x"80d47327",
  3033 => x"9e38768f",
  3034 => x"2a80f705",
  3035 => x"5582d473",
  3036 => x"27913876",
  3037 => x"922a80fc",
  3038 => x"05558ad4",
  3039 => x"73278438",
  3040 => x"80fe5574",
  3041 => x"10101080",
  3042 => x"f8940588",
  3043 => x"11085556",
  3044 => x"73762e82",
  3045 => x"b3388414",
  3046 => x"08fc0653",
  3047 => x"7673278d",
  3048 => x"38881408",
  3049 => x"5473762e",
  3050 => x"098106ea",
  3051 => x"388c1408",
  3052 => x"708c1a0c",
  3053 => x"74881a0c",
  3054 => x"7888120c",
  3055 => x"56778c15",
  3056 => x"0c7a51fc",
  3057 => x"883f8c3d",
  3058 => x"0d047708",
  3059 => x"78713159",
  3060 => x"77058819",
  3061 => x"08545772",
  3062 => x"80f89c2e",
  3063 => x"80e0388c",
  3064 => x"1808708c",
  3065 => x"150c7388",
  3066 => x"120c56fe",
  3067 => x"89398815",
  3068 => x"088c1608",
  3069 => x"708c130c",
  3070 => x"5788170c",
  3071 => x"fea33976",
  3072 => x"832a7054",
  3073 => x"55807524",
  3074 => x"81983872",
  3075 => x"822c8171",
  3076 => x"2b80f898",
  3077 => x"080780f8",
  3078 => x"940b8405",
  3079 => x"0c537410",
  3080 => x"101080f8",
  3081 => x"94058811",
  3082 => x"08555675",
  3083 => x"8c190c73",
  3084 => x"88190c77",
  3085 => x"88170c77",
  3086 => x"8c150cff",
  3087 => x"8439815a",
  3088 => x"fdb43978",
  3089 => x"17738106",
  3090 => x"54577298",
  3091 => x"38770878",
  3092 => x"71315977",
  3093 => x"058c1908",
  3094 => x"881a0871",
  3095 => x"8c120c88",
  3096 => x"120c5757",
  3097 => x"76810784",
  3098 => x"190c7780",
  3099 => x"f8940b88",
  3100 => x"050c80f8",
  3101 => x"90087726",
  3102 => x"fec73880",
  3103 => x"f88c0852",
  3104 => x"7a51fafe",
  3105 => x"3f7a51fa",
  3106 => x"c43ffeba",
  3107 => x"3981788c",
  3108 => x"150c7888",
  3109 => x"150c738c",
  3110 => x"1a0c7388",
  3111 => x"1a0c5afd",
  3112 => x"80398315",
  3113 => x"70822c81",
  3114 => x"712b80f8",
  3115 => x"98080780",
  3116 => x"f8940b84",
  3117 => x"050c5153",
  3118 => x"74101010",
  3119 => x"80f89405",
  3120 => x"88110855",
  3121 => x"56fee439",
  3122 => x"74538075",
  3123 => x"24a73872",
  3124 => x"822c8171",
  3125 => x"2b80f898",
  3126 => x"080780f8",
  3127 => x"940b8405",
  3128 => x"0c53758c",
  3129 => x"190c7388",
  3130 => x"190c7788",
  3131 => x"170c778c",
  3132 => x"150cfdcd",
  3133 => x"39831570",
  3134 => x"822c8171",
  3135 => x"2b80f898",
  3136 => x"080780f8",
  3137 => x"940b8405",
  3138 => x"0c5153d6",
  3139 => x"39810b80",
  3140 => x"0c04803d",
  3141 => x"0d72812e",
  3142 => x"8938800b",
  3143 => x"800c823d",
  3144 => x"0d047351",
  3145 => x"80f83ffe",
  3146 => x"3d0d818a",
  3147 => x"d8085170",
  3148 => x"8a38818a",
  3149 => x"e470818a",
  3150 => x"d80c5170",
  3151 => x"75125252",
  3152 => x"ff537087",
  3153 => x"fb808026",
  3154 => x"88387081",
  3155 => x"8ad80c71",
  3156 => x"5372800c",
  3157 => x"843d0d04",
  3158 => x"fd3d0d80",
  3159 => x"0b80f0ac",
  3160 => x"08545472",
  3161 => x"812e9c38",
  3162 => x"73818adc",
  3163 => x"0cffa6b3",
  3164 => x"3fffa58c",
  3165 => x"3f81809c",
  3166 => x"528151cf",
  3167 => x"943f8008",
  3168 => x"51a23f72",
  3169 => x"818adc0c",
  3170 => x"ffa6983f",
  3171 => x"ffa4f13f",
  3172 => x"81809c52",
  3173 => x"8151cef9",
  3174 => x"3f800851",
  3175 => x"873f00ff",
  3176 => x"3900ff39",
  3177 => x"f73d0d7b",
  3178 => x"80f0d808",
  3179 => x"82c81108",
  3180 => x"5a545a77",
  3181 => x"802e80da",
  3182 => x"38818818",
  3183 => x"841908ff",
  3184 => x"0581712b",
  3185 => x"59555980",
  3186 => x"742480ea",
  3187 => x"38807424",
  3188 => x"b5387382",
  3189 => x"2b781188",
  3190 => x"05565681",
  3191 => x"80190877",
  3192 => x"06537280",
  3193 => x"2eb63878",
  3194 => x"16700853",
  3195 => x"53795174",
  3196 => x"0853722d",
  3197 => x"ff14fc17",
  3198 => x"fc177981",
  3199 => x"2c5a5757",
  3200 => x"54738025",
  3201 => x"d6387708",
  3202 => x"5877ffad",
  3203 => x"3880f0d8",
  3204 => x"0853bc13",
  3205 => x"08a53879",
  3206 => x"51ff833f",
  3207 => x"74085372",
  3208 => x"2dff14fc",
  3209 => x"17fc1779",
  3210 => x"812c5a57",
  3211 => x"57547380",
  3212 => x"25ffa838",
  3213 => x"d1398057",
  3214 => x"ff933972",
  3215 => x"51bc1308",
  3216 => x"53722d79",
  3217 => x"51fed73f",
  3218 => x"ff3d0d81",
  3219 => x"80a40bfc",
  3220 => x"05700852",
  3221 => x"5270ff2e",
  3222 => x"9138702d",
  3223 => x"fc127008",
  3224 => x"525270ff",
  3225 => x"2e098106",
  3226 => x"f138833d",
  3227 => x"0d0404ff",
  3228 => x"a59e3f04",
  3229 => x"00000040",
  3230 => x"68656c70",
  3231 => x"00000000",
  3232 => x"3e200000",
  3233 => x"636f6d6d",
  3234 => x"616e6420",
  3235 => x"6e6f7420",
  3236 => x"666f756e",
  3237 => x"642e0a00",
  3238 => x"73757070",
  3239 => x"6f727465",
  3240 => x"6420636f",
  3241 => x"6d6d616e",
  3242 => x"64733a0a",
  3243 => x"0a000000",
  3244 => x"202d2000",
  3245 => x"62706d00",
  3246 => x"73686f77",
  3247 => x"2042504d",
  3248 => x"20726567",
  3249 => x"69737465",
  3250 => x"72730000",
  3251 => x"63686563",
  3252 => x"6b000000",
  3253 => x"63686563",
  3254 => x"6b204932",
  3255 => x"43206164",
  3256 => x"64726573",
  3257 => x"73000000",
  3258 => x"65646964",
  3259 => x"00000000",
  3260 => x"72656164",
  3261 => x"20454449",
  3262 => x"44206469",
  3263 => x"73706c61",
  3264 => x"79206461",
  3265 => x"74610000",
  3266 => x"63726561",
  3267 => x"64000000",
  3268 => x"72656164",
  3269 => x"20636872",
  3270 => x"6f6e7465",
  3271 => x"6c207265",
  3272 => x"67697374",
  3273 => x"65727300",
  3274 => x"63696e69",
  3275 => x"74000000",
  3276 => x"696e6974",
  3277 => x"20636872",
  3278 => x"6f6e7465",
  3279 => x"6c207265",
  3280 => x"67697374",
  3281 => x"65727300",
  3282 => x"63777269",
  3283 => x"74650000",
  3284 => x"77726974",
  3285 => x"65206368",
  3286 => x"726f6e74",
  3287 => x"656c2072",
  3288 => x"65676973",
  3289 => x"74657220",
  3290 => x"3c726567",
  3291 => x"3e203c76",
  3292 => x"616c7565",
  3293 => x"3e000000",
  3294 => x"6d656d00",
  3295 => x"616c6961",
  3296 => x"7320666f",
  3297 => x"72207800",
  3298 => x"776d656d",
  3299 => x"00000000",
  3300 => x"77726974",
  3301 => x"6520776f",
  3302 => x"72640000",
  3303 => x"6558616d",
  3304 => x"696e6520",
  3305 => x"6d656d6f",
  3306 => x"72790000",
  3307 => x"636c6561",
  3308 => x"72000000",
  3309 => x"636c6561",
  3310 => x"72207363",
  3311 => x"7265656e",
  3312 => x"00000000",
  3313 => x"71756974",
  3314 => x"00000000",
  3315 => x"30780000",
  3316 => x"0a307800",
  3317 => x"203a2000",
  3318 => x"69326320",
  3319 => x"4456490a",
  3320 => x"00000000",
  3321 => x"69326320",
  3322 => x"464d430a",
  3323 => x"00000000",
  3324 => x"69326320",
  3325 => x"61646472",
  3326 => x"6573733a",
  3327 => x"20307800",
  3328 => x"2020202d",
  3329 => x"2d3e2020",
  3330 => x"2041434b",
  3331 => x"0a000000",
  3332 => x"72656164",
  3333 => x"20454449",
  3334 => x"44206461",
  3335 => x"74612028",
  3336 => x"00000000",
  3337 => x"20627974",
  3338 => x"65732920",
  3339 => x"66726f6d",
  3340 => x"20493243",
  3341 => x"2d616464",
  3342 => x"72657373",
  3343 => x"20307800",
  3344 => x"0a0a0000",
  3345 => x"6368726f",
  3346 => x"6e74656c",
  3347 => x"20726567",
  3348 => x"20307800",
  3349 => x"3a203078",
  3350 => x"00000000",
  3351 => x"206e6163",
  3352 => x"6b000000",
  3353 => x"76616c75",
  3354 => x"653a2030",
  3355 => x"78000000",
  3356 => x"6572726f",
  3357 => x"7220286e",
  3358 => x"61636b29",
  3359 => x"00000000",
  3360 => x"6265616d",
  3361 => x"20706f73",
  3362 => x"6974696f",
  3363 => x"6e206d6f",
  3364 => x"6e69746f",
  3365 => x"72207265",
  3366 => x"67697374",
  3367 => x"65727300",
  3368 => x"0a202020",
  3369 => x"20202020",
  3370 => x"20202020",
  3371 => x"20202020",
  3372 => x"20202020",
  3373 => x"20202020",
  3374 => x"20636861",
  3375 => x"6e6e656c",
  3376 => x"20302020",
  3377 => x"20636861",
  3378 => x"6e6e656c",
  3379 => x"20312020",
  3380 => x"20636861",
  3381 => x"6e6e656c",
  3382 => x"20322020",
  3383 => x"20636861",
  3384 => x"6e6e656c",
  3385 => x"20330000",
  3386 => x"0a202020",
  3387 => x"20202020",
  3388 => x"20202020",
  3389 => x"20202020",
  3390 => x"20202020",
  3391 => x"20202020",
  3392 => x"202d2d2d",
  3393 => x"2d20686f",
  3394 => x"72697a6f",
  3395 => x"6e74616c",
  3396 => x"202d2d2d",
  3397 => x"2d2d2020",
  3398 => x"202d2d2d",
  3399 => x"2d2d2d20",
  3400 => x"76657274",
  3401 => x"6963616c",
  3402 => x"202d2d2d",
  3403 => x"2d2d0000",
  3404 => x"0a736361",
  3405 => x"6c657220",
  3406 => x"76616c75",
  3407 => x"65732020",
  3408 => x"20202020",
  3409 => x"20202020",
  3410 => x"20000000",
  3411 => x"0a6e6f69",
  3412 => x"73652063",
  3413 => x"6f6d7065",
  3414 => x"6e736174",
  3415 => x"696f6e20",
  3416 => x"20202020",
  3417 => x"20000000",
  3418 => x"0a6d6561",
  3419 => x"73757265",
  3420 => x"6d656e74",
  3421 => x"20202020",
  3422 => x"20202020",
  3423 => x"20202020",
  3424 => x"20000000",
  3425 => x"0a73756d",
  3426 => x"20636861",
  3427 => x"6e6e656c",
  3428 => x"2020203a",
  3429 => x"20000000",
  3430 => x"0a706f73",
  3431 => x"6974696f",
  3432 => x"6e20636f",
  3433 => x"6d707574",
  3434 => x"6174696f",
  3435 => x"6e000000",
  3436 => x"0a202073",
  3437 => x"63616c65",
  3438 => x"72207661",
  3439 => x"6c756573",
  3440 => x"20202020",
  3441 => x"20202020",
  3442 => x"20000000",
  3443 => x"0a20206f",
  3444 => x"66667365",
  3445 => x"74202020",
  3446 => x"20202020",
  3447 => x"20202020",
  3448 => x"20202020",
  3449 => x"20000000",
  3450 => x"0a6f7574",
  3451 => x"70757420",
  3452 => x"73656c65",
  3453 => x"6374203a",
  3454 => x"20000000",
  3455 => x"6368616e",
  3456 => x"6e656c20",
  3457 => x"30000000",
  3458 => x"76657274",
  3459 => x"6963616c",
  3460 => x"00000000",
  3461 => x"686f7269",
  3462 => x"7a6f6e74",
  3463 => x"616c0000",
  3464 => x"73756d00",
  3465 => x"6368616e",
  3466 => x"6e656c20",
  3467 => x"33000000",
  3468 => x"6368616e",
  3469 => x"6e656c20",
  3470 => x"32000000",
  3471 => x"6368616e",
  3472 => x"6e656c20",
  3473 => x"31000000",
  3474 => x"6265616d",
  3475 => x"20706f73",
  3476 => x"6974696f",
  3477 => x"6e206d6f",
  3478 => x"6e69746f",
  3479 => x"72000000",
  3480 => x"20286f6e",
  3481 => x"2073696d",
  3482 => x"290a0000",
  3483 => x"0a636f6d",
  3484 => x"70696c65",
  3485 => x"643a204d",
  3486 => x"61792020",
  3487 => x"32203230",
  3488 => x"31312020",
  3489 => x"31313a34",
  3490 => x"303a3339",
  3491 => x"00000000",
  3492 => x"0a737973",
  3493 => x"74656d20",
  3494 => x"636c6f63",
  3495 => x"6b3a2000",
  3496 => x"204d487a",
  3497 => x"0a000000",
  3498 => x"44454255",
  3499 => x"47204d4f",
  3500 => x"4445204f",
  3501 => x"4e0a0000",
  3502 => x"000018cb",
  3503 => x"00001908",
  3504 => x"000018ff",
  3505 => x"000018f6",
  3506 => x"000018ed",
  3507 => x"000018e4",
  3508 => x"000018db",
  3509 => x"30622020",
  3510 => x"20202020",
  3511 => x"20202020",
  3512 => x"20202020",
  3513 => x"20202020",
  3514 => x"20202020",
  3515 => x"20202020",
  3516 => x"20202020",
  3517 => x"20200000",
  3518 => x"20202020",
  3519 => x"20202020",
  3520 => x"00000000",
  3521 => x"00202020",
  3522 => x"20202020",
  3523 => x"20202828",
  3524 => x"28282820",
  3525 => x"20202020",
  3526 => x"20202020",
  3527 => x"20202020",
  3528 => x"20202020",
  3529 => x"20881010",
  3530 => x"10101010",
  3531 => x"10101010",
  3532 => x"10101010",
  3533 => x"10040404",
  3534 => x"04040404",
  3535 => x"04040410",
  3536 => x"10101010",
  3537 => x"10104141",
  3538 => x"41414141",
  3539 => x"01010101",
  3540 => x"01010101",
  3541 => x"01010101",
  3542 => x"01010101",
  3543 => x"01010101",
  3544 => x"10101010",
  3545 => x"10104242",
  3546 => x"42424242",
  3547 => x"02020202",
  3548 => x"02020202",
  3549 => x"02020202",
  3550 => x"02020202",
  3551 => x"02020202",
  3552 => x"10101010",
  3553 => x"20000000",
  3554 => x"00000000",
  3555 => x"00000000",
  3556 => x"00000000",
  3557 => x"00000000",
  3558 => x"00000000",
  3559 => x"00000000",
  3560 => x"00000000",
  3561 => x"00000000",
  3562 => x"00000000",
  3563 => x"00000000",
  3564 => x"00000000",
  3565 => x"00000000",
  3566 => x"00000000",
  3567 => x"00000000",
  3568 => x"00000000",
  3569 => x"00000000",
  3570 => x"00000000",
  3571 => x"00000000",
  3572 => x"00000000",
  3573 => x"00000000",
  3574 => x"00000000",
  3575 => x"00000000",
  3576 => x"00000000",
  3577 => x"00000000",
  3578 => x"00000000",
  3579 => x"00000000",
  3580 => x"00000000",
  3581 => x"00000000",
  3582 => x"00000000",
  3583 => x"00000000",
  3584 => x"00000000",
  3585 => x"00000000",
  3586 => x"43000000",
  3587 => x"64756d6d",
  3588 => x"792e6578",
  3589 => x"65000000",
  3590 => x"00ffffff",
  3591 => x"ff00ffff",
  3592 => x"ffff00ff",
  3593 => x"ffffff00",
  3594 => x"00000000",
  3595 => x"00000000",
  3596 => x"00000000",
  3597 => x"0000402c",
  3598 => x"80000a00",
  3599 => x"80000700",
  3600 => x"80000800",
  3601 => x"80000600",
  3602 => x"80000400",
  3603 => x"80000200",
  3604 => x"80000100",
  3605 => x"80000000",
  3606 => x"0000385c",
  3607 => x"00000000",
  3608 => x"00003ac4",
  3609 => x"00003b20",
  3610 => x"00003b7c",
  3611 => x"00000000",
  3612 => x"00000000",
  3613 => x"00000000",
  3614 => x"00000000",
  3615 => x"00000000",
  3616 => x"00000000",
  3617 => x"00000000",
  3618 => x"00000000",
  3619 => x"00000000",
  3620 => x"00003808",
  3621 => x"00000000",
  3622 => x"00000000",
  3623 => x"00000000",
  3624 => x"00000000",
  3625 => x"00000000",
  3626 => x"00000000",
  3627 => x"00000000",
  3628 => x"00000000",
  3629 => x"00000000",
  3630 => x"00000000",
  3631 => x"00000000",
  3632 => x"00000000",
  3633 => x"00000000",
  3634 => x"00000000",
  3635 => x"00000000",
  3636 => x"00000000",
  3637 => x"00000000",
  3638 => x"00000000",
  3639 => x"00000000",
  3640 => x"00000000",
  3641 => x"00000000",
  3642 => x"00000000",
  3643 => x"00000000",
  3644 => x"00000000",
  3645 => x"00000000",
  3646 => x"00000000",
  3647 => x"00000000",
  3648 => x"00000000",
  3649 => x"00000001",
  3650 => x"330eabcd",
  3651 => x"1234e66d",
  3652 => x"deec0005",
  3653 => x"000b0000",
  3654 => x"00000000",
  3655 => x"00000000",
  3656 => x"00000000",
  3657 => x"00000000",
  3658 => x"00000000",
  3659 => x"00000000",
  3660 => x"00000000",
  3661 => x"00000000",
  3662 => x"00000000",
  3663 => x"00000000",
  3664 => x"00000000",
  3665 => x"00000000",
  3666 => x"00000000",
  3667 => x"00000000",
  3668 => x"00000000",
  3669 => x"00000000",
  3670 => x"00000000",
  3671 => x"00000000",
  3672 => x"00000000",
  3673 => x"00000000",
  3674 => x"00000000",
  3675 => x"00000000",
  3676 => x"00000000",
  3677 => x"00000000",
  3678 => x"00000000",
  3679 => x"00000000",
  3680 => x"00000000",
  3681 => x"00000000",
  3682 => x"00000000",
  3683 => x"00000000",
  3684 => x"00000000",
  3685 => x"00000000",
  3686 => x"00000000",
  3687 => x"00000000",
  3688 => x"00000000",
  3689 => x"00000000",
  3690 => x"00000000",
  3691 => x"00000000",
  3692 => x"00000000",
  3693 => x"00000000",
  3694 => x"00000000",
  3695 => x"00000000",
  3696 => x"00000000",
  3697 => x"00000000",
  3698 => x"00000000",
  3699 => x"00000000",
  3700 => x"00000000",
  3701 => x"00000000",
  3702 => x"00000000",
  3703 => x"00000000",
  3704 => x"00000000",
  3705 => x"00000000",
  3706 => x"00000000",
  3707 => x"00000000",
  3708 => x"00000000",
  3709 => x"00000000",
  3710 => x"00000000",
  3711 => x"00000000",
  3712 => x"00000000",
  3713 => x"00000000",
  3714 => x"00000000",
  3715 => x"00000000",
  3716 => x"00000000",
  3717 => x"00000000",
  3718 => x"00000000",
  3719 => x"00000000",
  3720 => x"00000000",
  3721 => x"00000000",
  3722 => x"00000000",
  3723 => x"00000000",
  3724 => x"00000000",
  3725 => x"00000000",
  3726 => x"00000000",
  3727 => x"00000000",
  3728 => x"00000000",
  3729 => x"00000000",
  3730 => x"00000000",
  3731 => x"00000000",
  3732 => x"00000000",
  3733 => x"00000000",
  3734 => x"00000000",
  3735 => x"00000000",
  3736 => x"00000000",
  3737 => x"00000000",
  3738 => x"00000000",
  3739 => x"00000000",
  3740 => x"00000000",
  3741 => x"00000000",
  3742 => x"00000000",
  3743 => x"00000000",
  3744 => x"00000000",
  3745 => x"00000000",
  3746 => x"00000000",
  3747 => x"00000000",
  3748 => x"00000000",
  3749 => x"00000000",
  3750 => x"00000000",
  3751 => x"00000000",
  3752 => x"00000000",
  3753 => x"00000000",
  3754 => x"00000000",
  3755 => x"00000000",
  3756 => x"00000000",
  3757 => x"00000000",
  3758 => x"00000000",
  3759 => x"00000000",
  3760 => x"00000000",
  3761 => x"00000000",
  3762 => x"00000000",
  3763 => x"00000000",
  3764 => x"00000000",
  3765 => x"00000000",
  3766 => x"00000000",
  3767 => x"00000000",
  3768 => x"00000000",
  3769 => x"00000000",
  3770 => x"00000000",
  3771 => x"00000000",
  3772 => x"00000000",
  3773 => x"00000000",
  3774 => x"00000000",
  3775 => x"00000000",
  3776 => x"00000000",
  3777 => x"00000000",
  3778 => x"00000000",
  3779 => x"00000000",
  3780 => x"00000000",
  3781 => x"00000000",
  3782 => x"00000000",
  3783 => x"00000000",
  3784 => x"00000000",
  3785 => x"00000000",
  3786 => x"00000000",
  3787 => x"00000000",
  3788 => x"00000000",
  3789 => x"00000000",
  3790 => x"00000000",
  3791 => x"00000000",
  3792 => x"00000000",
  3793 => x"00000000",
  3794 => x"00000000",
  3795 => x"00000000",
  3796 => x"00000000",
  3797 => x"00000000",
  3798 => x"00000000",
  3799 => x"00000000",
  3800 => x"00000000",
  3801 => x"00000000",
  3802 => x"00000000",
  3803 => x"00000000",
  3804 => x"00000000",
  3805 => x"00000000",
  3806 => x"00000000",
  3807 => x"00000000",
  3808 => x"00000000",
  3809 => x"00000000",
  3810 => x"00000000",
  3811 => x"00000000",
  3812 => x"00000000",
  3813 => x"00000000",
  3814 => x"00000000",
  3815 => x"00000000",
  3816 => x"00000000",
  3817 => x"00000000",
  3818 => x"00000000",
  3819 => x"00000000",
  3820 => x"00000000",
  3821 => x"00000000",
  3822 => x"00000000",
  3823 => x"00000000",
  3824 => x"00000000",
  3825 => x"00000000",
  3826 => x"00000000",
  3827 => x"00000000",
  3828 => x"00000000",
  3829 => x"00000000",
  3830 => x"00000000",
  3831 => x"00000000",
  3832 => x"00000000",
  3833 => x"00000000",
  3834 => x"00000000",
  3835 => x"00000000",
  3836 => x"00000000",
  3837 => x"00000000",
  3838 => x"00000000",
  3839 => x"00000000",
  3840 => x"00000000",
  3841 => x"00000000",
  3842 => x"ffffffff",
  3843 => x"00000000",
  3844 => x"00020000",
  3845 => x"00000000",
  3846 => x"00000000",
  3847 => x"00003c14",
  3848 => x"00003c14",
  3849 => x"00003c1c",
  3850 => x"00003c1c",
  3851 => x"00003c24",
  3852 => x"00003c24",
  3853 => x"00003c2c",
  3854 => x"00003c2c",
  3855 => x"00003c34",
  3856 => x"00003c34",
  3857 => x"00003c3c",
  3858 => x"00003c3c",
  3859 => x"00003c44",
  3860 => x"00003c44",
  3861 => x"00003c4c",
  3862 => x"00003c4c",
  3863 => x"00003c54",
  3864 => x"00003c54",
  3865 => x"00003c5c",
  3866 => x"00003c5c",
  3867 => x"00003c64",
  3868 => x"00003c64",
  3869 => x"00003c6c",
  3870 => x"00003c6c",
  3871 => x"00003c74",
  3872 => x"00003c74",
  3873 => x"00003c7c",
  3874 => x"00003c7c",
  3875 => x"00003c84",
  3876 => x"00003c84",
  3877 => x"00003c8c",
  3878 => x"00003c8c",
  3879 => x"00003c94",
  3880 => x"00003c94",
  3881 => x"00003c9c",
  3882 => x"00003c9c",
  3883 => x"00003ca4",
  3884 => x"00003ca4",
  3885 => x"00003cac",
  3886 => x"00003cac",
  3887 => x"00003cb4",
  3888 => x"00003cb4",
  3889 => x"00003cbc",
  3890 => x"00003cbc",
  3891 => x"00003cc4",
  3892 => x"00003cc4",
  3893 => x"00003ccc",
  3894 => x"00003ccc",
  3895 => x"00003cd4",
  3896 => x"00003cd4",
  3897 => x"00003cdc",
  3898 => x"00003cdc",
  3899 => x"00003ce4",
  3900 => x"00003ce4",
  3901 => x"00003cec",
  3902 => x"00003cec",
  3903 => x"00003cf4",
  3904 => x"00003cf4",
  3905 => x"00003cfc",
  3906 => x"00003cfc",
  3907 => x"00003d04",
  3908 => x"00003d04",
  3909 => x"00003d0c",
  3910 => x"00003d0c",
  3911 => x"00003d14",
  3912 => x"00003d14",
  3913 => x"00003d1c",
  3914 => x"00003d1c",
  3915 => x"00003d24",
  3916 => x"00003d24",
  3917 => x"00003d2c",
  3918 => x"00003d2c",
  3919 => x"00003d34",
  3920 => x"00003d34",
  3921 => x"00003d3c",
  3922 => x"00003d3c",
  3923 => x"00003d44",
  3924 => x"00003d44",
  3925 => x"00003d4c",
  3926 => x"00003d4c",
  3927 => x"00003d54",
  3928 => x"00003d54",
  3929 => x"00003d5c",
  3930 => x"00003d5c",
  3931 => x"00003d64",
  3932 => x"00003d64",
  3933 => x"00003d6c",
  3934 => x"00003d6c",
  3935 => x"00003d74",
  3936 => x"00003d74",
  3937 => x"00003d7c",
  3938 => x"00003d7c",
  3939 => x"00003d84",
  3940 => x"00003d84",
  3941 => x"00003d8c",
  3942 => x"00003d8c",
  3943 => x"00003d94",
  3944 => x"00003d94",
  3945 => x"00003d9c",
  3946 => x"00003d9c",
  3947 => x"00003da4",
  3948 => x"00003da4",
  3949 => x"00003dac",
  3950 => x"00003dac",
  3951 => x"00003db4",
  3952 => x"00003db4",
  3953 => x"00003dbc",
  3954 => x"00003dbc",
  3955 => x"00003dc4",
  3956 => x"00003dc4",
  3957 => x"00003dcc",
  3958 => x"00003dcc",
  3959 => x"00003dd4",
  3960 => x"00003dd4",
  3961 => x"00003ddc",
  3962 => x"00003ddc",
  3963 => x"00003de4",
  3964 => x"00003de4",
  3965 => x"00003dec",
  3966 => x"00003dec",
  3967 => x"00003df4",
  3968 => x"00003df4",
  3969 => x"00003dfc",
  3970 => x"00003dfc",
  3971 => x"00003e04",
  3972 => x"00003e04",
  3973 => x"00003e0c",
  3974 => x"00003e0c",
  3975 => x"00003e14",
  3976 => x"00003e14",
  3977 => x"00003e1c",
  3978 => x"00003e1c",
  3979 => x"00003e24",
  3980 => x"00003e24",
  3981 => x"00003e2c",
  3982 => x"00003e2c",
  3983 => x"00003e34",
  3984 => x"00003e34",
  3985 => x"00003e3c",
  3986 => x"00003e3c",
  3987 => x"00003e44",
  3988 => x"00003e44",
  3989 => x"00003e4c",
  3990 => x"00003e4c",
  3991 => x"00003e54",
  3992 => x"00003e54",
  3993 => x"00003e5c",
  3994 => x"00003e5c",
  3995 => x"00003e64",
  3996 => x"00003e64",
  3997 => x"00003e6c",
  3998 => x"00003e6c",
  3999 => x"00003e74",
  4000 => x"00003e74",
  4001 => x"00003e7c",
  4002 => x"00003e7c",
  4003 => x"00003e84",
  4004 => x"00003e84",
  4005 => x"00003e8c",
  4006 => x"00003e8c",
  4007 => x"00003e94",
  4008 => x"00003e94",
  4009 => x"00003e9c",
  4010 => x"00003e9c",
  4011 => x"00003ea4",
  4012 => x"00003ea4",
  4013 => x"00003eac",
  4014 => x"00003eac",
  4015 => x"00003eb4",
  4016 => x"00003eb4",
  4017 => x"00003ebc",
  4018 => x"00003ebc",
  4019 => x"00003ec4",
  4020 => x"00003ec4",
  4021 => x"00003ecc",
  4022 => x"00003ecc",
  4023 => x"00003ed4",
  4024 => x"00003ed4",
  4025 => x"00003edc",
  4026 => x"00003edc",
  4027 => x"00003ee4",
  4028 => x"00003ee4",
  4029 => x"00003eec",
  4030 => x"00003eec",
  4031 => x"00003ef4",
  4032 => x"00003ef4",
  4033 => x"00003efc",
  4034 => x"00003efc",
  4035 => x"00003f04",
  4036 => x"00003f04",
  4037 => x"00003f0c",
  4038 => x"00003f0c",
  4039 => x"00003f14",
  4040 => x"00003f14",
  4041 => x"00003f1c",
  4042 => x"00003f1c",
  4043 => x"00003f24",
  4044 => x"00003f24",
  4045 => x"00003f2c",
  4046 => x"00003f2c",
  4047 => x"00003f34",
  4048 => x"00003f34",
  4049 => x"00003f3c",
  4050 => x"00003f3c",
  4051 => x"00003f44",
  4052 => x"00003f44",
  4053 => x"00003f4c",
  4054 => x"00003f4c",
  4055 => x"00003f54",
  4056 => x"00003f54",
  4057 => x"00003f5c",
  4058 => x"00003f5c",
  4059 => x"00003f64",
  4060 => x"00003f64",
  4061 => x"00003f6c",
  4062 => x"00003f6c",
  4063 => x"00003f74",
  4064 => x"00003f74",
  4065 => x"00003f7c",
  4066 => x"00003f7c",
  4067 => x"00003f84",
  4068 => x"00003f84",
  4069 => x"00003f8c",
  4070 => x"00003f8c",
  4071 => x"00003f94",
  4072 => x"00003f94",
  4073 => x"00003f9c",
  4074 => x"00003f9c",
  4075 => x"00003fa4",
  4076 => x"00003fa4",
  4077 => x"00003fac",
  4078 => x"00003fac",
  4079 => x"00003fb4",
  4080 => x"00003fb4",
  4081 => x"00003fbc",
  4082 => x"00003fbc",
  4083 => x"00003fc4",
  4084 => x"00003fc4",
  4085 => x"00003fcc",
  4086 => x"00003fcc",
  4087 => x"00003fd4",
  4088 => x"00003fd4",
  4089 => x"00003fdc",
  4090 => x"00003fdc",
  4091 => x"00003fe4",
  4092 => x"00003fe4",
  4093 => x"00003fec",
  4094 => x"00003fec",
  4095 => x"00003ff4",
  4096 => x"00003ff4",
  4097 => x"00003ffc",
  4098 => x"00003ffc",
  4099 => x"00004004",
  4100 => x"00004004",
  4101 => x"0000400c",
  4102 => x"0000400c",
  4103 => x"0000380c",
  4104 => x"ffffffff",
  4105 => x"00000000",
  4106 => x"ffffffff",
  4107 => x"00000000",
  4108 => x"00000000",
	others => x"aaaaaaaa" -- mask for mem check
	--others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
