--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:    11:47:36 03/22/05
-- Design Name:    
-- Module Name:    mem_sys - behave
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description:
--
-- Dependencies:
-- 				  
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;
library zylin;
use zylin.zpu_config.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


signal	low				: std_logic;
signal	high				: std_logic;
signal  re : std_logic;
																		 
begin

	high <= '1';
	low <= '0';
	re <= '1';


   ZPU_RAM0 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"01A100E100010001003600770002006D000F0000000F06AD000302940008003C",
      INIT_01 => X"7D4000000741F68100C800030000377935990003000300030003002A00150001",
      INIT_02 => X"0007584101010C3D55555555370000000092800000001490000000066A594EBB",
      INIT_03 => X"0009015555932D564C093A4024055555564CB555593C1569EA90C00000007000",
      INIT_04 => X"BF8AA55961BE2A956586C40A4CB00932C00024A80000024C9569C893C0024E90",
      INIT_05 => X"18A1251E2A956586F8AA55961BF8AA55961BE2A956586FE2A956586F8AA55961",
      INIT_06 => X"51349D53764E258A2043E21BE5645DE5C4FC00E0100430C140E4665595558750",
      INIT_07 => X"47B1656A855555D435575A815D077558E475559E755715A1C364945042425555",
      INIT_08 => X"5555F123348C17657C405070D5E745A518B58DD5555F55551D5506F00D707B15",
      INIT_09 => X"C141C74DD5137120D51C0715094CC4F01006A8131DD91531B913118944815155",
      INIT_0A => X"5E559655003D3549550D458C5994A04D476568D05B0F45451D143E53D0F2CD6B",
      INIT_0B => X"4D1E1C5D3474C5C5A1E1C5D34787171C44DC7844D3451D37974D164DD55DD555",
      INIT_0C => X"2074532E4C3A5074DE129D074D1137134477D546C01D374DD348774DE15D3717",
      INIT_0D => X"875650117671948CB05545A5A2615074889149341D04D4956F843575543E1A19",
      INIT_0E => X"F804036D9753106651D5140E6905C158D8979404C7459123540DD9955A43F563",
      INIT_0F => X"7958D037C3557056405549520F96E88622775767141BA3755D1418E1BE234480",
      INIT_10 => X"294A1C405ACCC3705D5599D55037776149584D8F98F98F98FDD00D904D205421",
      INIT_11 => X"74710D5C26798346751441DD555BE179544D8F98F98F98FDD00D910DC3D357C3",
      INIT_12 => X"605D5570051840119D04C0DC3755B61D7951D9A9522D995D51D5BB106B90F7C0",
      INIT_13 => X"D81BC3646611D695A02D1A9419695D695422C40110C0F85D6F899E4D0D555BC3",
      INIT_14 => X"28531104D5F01EDD204141807555735D38346423303676407555545F6B945696",
      INIT_15 => X"5212D7645155503146685C599546660676E81041C85D570DCE1B07116F116021",
      INIT_16 => X"5F9D03530F840406A5725910604E420D910DD521D6170F9AF0F940D91836445D",
      INIT_17 => X"83E03E03C03414D5D5F5D9BE7550DD55775514A145E5405657024C3664F3059C",
      INIT_18 => X"444C7584143756C431049D594DC444FD19CE181427555124440155503F58E14D",
      INIT_19 => X"D54521B201810644D895159C568F40C6C85503E135203FCF555151102C7343CC",
      INIT_1A => X"5A95904431351D93820C4D1AA2C7FD0CD95555311185802971639A1755607515",
      INIT_1B => X"E7D41815C826057201815C826057201815C806057209815C82741C75D1BF4336",
      INIT_1C => X"41BD443664E14155000C4191440445305B46A8D40443A3E115495503116861C3",
      INIT_1D => X"A1520F9C10F850FC18DB80D4777F1D5757195241D35F9754D755DD35F40D9D99",
      INIT_1E => X"65E6A10F206870F0557411545536F0D5FA1765C8D5443E658956E52727558D14",
      INIT_1F => X"DDD2151D31A956A0400F03FC754175510FD4A34252E0DC4076A5EC66A10FB312",
      INIT_20 => X"77C1676610FBD310C3C3CC76F05C9FF20755DC17ECE5451D3472D9D215D34C40",
      INIT_21 => X"55556189C508B6C3F0F0FF1D9F4561676610F207A5EF52D7957CC0F8800F7726",
      INIT_22 => X"8890203480C224080B251D4352F126920C8CF13E00C15A16445A44DA4F105554",
      INIT_23 => X"0F203CF4495240B82923890203080E20B8809249524080C2C0B490210C803203",
      INIT_24 => X"854F25C74C20400C1030000B24838A6F858A08E24080F2823890203C80D203C8",
      INIT_25 => X"00000C000000001F75D5D74FC0000000000000003FFFFFFFEAAA95438104DA47",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000154000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(1 downto 0),      -- Port A 2-bit Data Output
      DOB => memBRead(1 downto 0),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(1 downto 0),      -- Port A 2-bit Data Input
      DIB => memBWrite(1 downto 0),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => low,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM1 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"01510111000100020061006B0000004000100002001005510001059A00360064",
      INIT_01 => X"40300000064005640380001E0001543802180002000200010002000500110005",
      INIT_02 => X"000653709D19C24E555555552400000000920000000024000000000162843876",
      INIT_03 => X"0000CC55555DC1557EC5DC00033155555577055555D315607655000000007000",
      INIT_04 => X"74818211417206084505C705770000F940000398000001765560745D30017700",
      INIT_05 => X"165081C206084505C8182114174818211417206084505D206084505C81821141",
      INIT_06 => X"51200592163801450816D095E0044564ADB5C58C82606080118051A1162881C8",
      INIT_07 => X"550175554516163566505D44014118AA4818516C185014519662131830201616",
      INIT_08 => X"96140906D01981608AF43685992015DA5245D45628675859062835B511755017",
      INIT_09 => X"6000B8F861B22CE39C0EC602ED202FC596B59458405845C55118595694001162",
      INIT_0A => X"55A58300016D31668D5941040556516111611710005B4D4545716E190280595B",
      INIT_0B => X"C968C00BA5BE80B2C68C00B65A3002C1BC8BA32CBE70C3EA02C9CAC89C59458A",
      INIT_0C => X"0B1A0D6164EC408F8A047008D9CB622E2D19546CB32362C8BE8312FACC4BA202",
      INIT_0D => X"4455CCCC1601143B2E45916976DC147401104104059F14685B456418596D1171",
      INIT_0E => X"B4B55655D7453C5DA01654441070416015693378C475DC495A0458256156D15F",
      INIT_0F => X"468751645665865943F040105B8164446641416011165018A11454D15D007415",
      INIT_10 => X"8175134656FB96434615446289641B554684057595597595D066598611165695",
      INIT_11 => X"18A6599B55F856501AD764059656556684017495497495C066598559C91D555D",
      INIT_12 => X"5346166005EB404406411356518A35554684656685DD4686446112185F85B684",
      INIT_13 => X"D555D6601585546854151468D5568546895EB4044115B4595F454E12599655D6",
      INIT_14 => X"335D511B5557C55D467C504218A4E119C7135101456604AE1A05A1555F861668",
      INIT_15 => X"91101161116169E0F5D448156855955595171C7110462859E41D55815FD556C1",
      INIT_16 => X"153011465B440F059A495550560474598A50591544045B8105B8459841662905",
      INIT_17 => X"16E16C16C16514546104654E051C0615418A9450651A1155A1B165662D1D417D",
      INIT_18 => X"700111F690095D6159A445904D270024D7D3C3B711855915976D62896C56D165",
      INIT_19 => X"62A10F7C5B0C0557D468857E5149D00170C316D15CCD6EC558AD0441D72116D2",
      INIT_1A => X"97681F4400824581000023D4516DE3E2517161920D8D38057557861185921514",
      INIT_1B => X"E152154484F551212D544846551210954484D551212154484515A45C3B78F895",
      INIT_1C => X"457E256626804961925697473A0E2C44D0F51470F47849C431468400D048CD56",
      INIT_1D => X"51105B8C05B445B315555C05417946285153C440619C2166018A4619C8598151",
      INIT_1E => X"4595955BA2EA0761584405655975B59920519556E9056E0566859A4581645C14",
      INIT_1F => X"9055965A909455530D5B16F1185118A55B15520D55159076C55AF455155B50B6",
      INIT_20 => X"8085515155B6E90616D6E0146830806841851156724A0EC620DD04559653A415",
      INIT_21 => X"75858C001F40514145B5B40507C305515155BA2D93E496D5695545B4605B9418",
      INIT_22 => X"0810203080F20408032DA18003C200E266D1C15050400CF788038803844E58A1",
      INIT_23 => X"0F203CCF4CF040B12103010203480F208C80A24CF04080D0C03C1023BC82F203",
      INIT_24 => X"0600F6CFD04155043040000C38832340070840C04080F2103010203C803203C8",
      INIT_25 => X"0A000C00000020061C7185CFEAAAAAAAAAAAAAAA95555555555555540B080387",
      INIT_26 => X"0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A",
      INIT_27 => X"313A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A",
      INIT_28 => X"00000000000000000000000000000000000000000001F0000000000000030000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(3 downto 2),      -- Port A 2-bit Data Output
      DOB => memBRead(3 downto 2),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(3 downto 2),      -- Port A 2-bit Data Input
      DIB => memBWrite(3 downto 2),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM2 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"0008000800000000000000010001002A000200000002000800000080000800C6",
      INIT_01 => X"023AAAAAA028A040002A0000000002B000000000000000000000000000080000",
      INIT_02 => X"AAA00B000020000C0000000002AAAAAAAA082AAAAAAA828AAAAAAAA008223032",
      INIT_03 => X"AAA8CC000000E0000CC00E2AA33000000003800000030008300C2AAAAAAA3AAA",
      INIT_04 => X"3C2828002830A0A000A0C020038AA8F02AAAA302AAAAA8000008300032A8038A",
      INIT_05 => X"820800C0A0A000A0C282800283C2828002830A0A000A0F0A0A000A0C28280028",
      INIT_06 => X"00000C00303000208600C841C0008C028AB00806C170000010000C0080002A30",
      INIT_07 => X"8AB83808200000C000020C2000023002A830001E300380080002A00230100000",
      INIT_08 => X"0000C00C00322300330800E0008020C088C0E280000B0003CC0020F08038AB83",
      INIT_09 => X"40001DA0C0200401080400000CD880A23C00C23008C00A3B20303010102C8000",
      INIT_0A => X"0000002AEC0C70000A0093220A8008C0230028EE00032A008CA00C230004F00B",
      INIT_0B => X"9030420240C820130704202C1C108041C900C10A2CD04E0C00B34C80380E4000",
      INIT_0C => X"8E32028C080030DA0244070DA342C0BC26AA40880A36C0A020D1008304020040",
      INIT_0D => X"20A0303230280000AC0020A828028A20220000000C2080000B200030000C82C2",
      INIT_0E => X"323200204380C300000080880B80A80B83008D037820E3A00008C0400000C203",
      INIT_0F => X"00004800400008012C2000000300820808A323008D800A30008083C81C801000",
      INIT_10 => X"8030808000C0002F8C0008C0000230000002200882883881C8CB0002FA000000",
      INIT_11 => X"3080000A8030002A3220A08C0002800002200882883881C8CB000200C1200170",
      INIT_12 => X"2F8C000AB0282A0A8CAFA006230000040008C8300080100408C08A820B003028",
      INIT_13 => X"0002C0020208400002C8C1020800040002C282A0A800320003203C02000000C0",
      INIT_14 => X"28002208005C2A840002A08A3009090828820E0900000A823200200507004300",
      INIT_15 => X"0880A3000000020F00420E030000A080A0208208828C00000821810007080322",
      INIT_16 => X"85002D080320300040088382000800000008C080E0AA0300E030A0000000008C",
      INIT_17 => X"80C00C00C0010088C088C83C00028C002300800820000200013834000010B03C",
      INIT_18 => X"0A20108A00290E4080038C088C00A20081C12810A30000E0A0A000000C02C804",
      INIT_19 => X"C000020C0223C020C300000C002300C20882C0C813280FEF0008C0A8280900C0",
      INIT_1A => X"8200000030428C0E008C100108E0CC084020000ABA882800380702E300026028",
      INIT_1B => X"C0CE4280A240A02890280A240A02890280A200A02880280A2230228824330210",
      INIT_1C => X"081C8000008000008C00C204DC280368800042CE0002C1C0A0000383A00E0280",
      INIT_1D => X"0880030E803200308281822223088C00020082C0C08C630003008C08CA000000",
      INIT_1E => X"00206003248C882E00238008023030008EB33021D0D00C002020400323020E80",
      INIT_1F => X"08CA008A00888008AE0300F230223002030008AE02A00808A040812060030823",
      INIT_20 => X"88B0060A0032E00880C0C8322821A22AA3020D83B00D808C182E28CA00878020",
      INIT_21 => X"20000C003280A28E2030320C8B8220060A003248C6EA80C3003820302403026A",
      INIT_22 => X"C2BA0AAC2AA0AE82A93AAEABA2A0B110EAAFA3EFEE8ABBAAC2C442444F300000",
      INIT_23 => X"A90AA4BABAAAE82F04946BA0AAC2AA0AC82AE0BAAAE82AB24E5ABA09E42B90AA",
      INIT_24 => X"AA8FAAAAACFBBEE8BED8AAA9EC0AEEBECAC1251AE82A905946BA0AA42AA0AA42",
      INIT_25 => X"FAA00C000000700562A2FC8FC00000000000000000000000000000000E02C44E",
      INIT_26 => X"FAA5500FFAA5500FFAA5500FFAA5500FFAA5500FFAA5500FFAA5500FFAA5500F",
      INIT_27 => X"0D25500FFAA5500FFAA5500FFAA5500FFAA5500FFAA5500FFAA5500FFAA5500F",
      INIT_28 => X"0000000000000000000000000000000000000000000080000000000000020000",
      INIT_29 => X"00000000000000000CF000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(5 downto 4),      -- Port A 2-bit Data Output
      DOB => memBRead(5 downto 4),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(5 downto 4),      -- Port A 2-bit Data Input
      DIB => memBWrite(5 downto 4),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM3 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"00040044000000020008000200020115000500020005000400020000000C0089",
      INIT_01 => X"2975555550165082031500000000017218820002000200020002002000040000",
      INIT_02 => X"5550070B0150281C000000008155555555849555555561555555555404117230",
      INIT_03 => X"5555EE000000D8000CE00D9557B8000000036000000B80053000555555553555",
      INIT_04 => X"31141484143450521050E090036555F0955557015555540000053200B9540365",
      INIT_05 => X"4305181450521050D1414841431141484143450521050C450521050D14148414",
      INIT_06 => X"088A0C0830B088305988C583C9824C914136660AEABA8A2AAA2A08084081160A",
      INIT_07 => X"1544300C14808010800A0C1694A932055632082D3208420448095991A8684080",
      INIT_08 => X"008210800A02130B030A8092006990C04620C540821702028C8290F568315443",
      INIT_09 => X"9AB92A20C8084AAB01A820AB082640D53AA081A164C265B750A1702032124808",
      INIT_0A => X"08016955148DF82021207E5595420685930996D9952351204C588C926A2FC00B",
      INIT_0B => X"20E9A590C3A2192A9E9A590C3A6964A7A312A6830CEBA08A6433AA21310CA020",
      INIT_0C => X"6E31A15036890AA312FD78AA33A084ACBE61820106E8843108A6A4229A90C4A4",
      INIT_0D => X"11510AC9309402005C20185021614512190A28A28CF042020F108232008C45C4",
      INIT_0E => X"31214814832100080940422454855404420142448520CC9E00A4C2C40808D90B",
      INIT_0F => X"20268482C800150257062188232541244453130942420532044203C43C593612",
      INIT_10 => X"7830466802C008134C8064C8208132082025942102102103D4C6202525980008",
      INIT_11 => X"3241200540B2481531105A4C0002082025942102102103D4C6202520FB5002B0",
      INIT_12 => X"134C801D711635AD4C525809932060882024C4202648202924C855430F223516",
      INIT_13 => X"8282C80B91A8820265040201042028202691635AD44231040B103C99200003C8",
      INIT_14 => X"9600999400AC154C98015A653207468C14C808871080914131A01A0A0F24C301",
      INIT_15 => X"044853098808030C00C111820210C16080C44104654C8220949E86A80B240B19",
      INIT_16 => X"4B46A224231280A0801E421B0AA401202064C048D1552324123252026480814C",
      INIT_17 => X"48E88E88E8828204C864C42C90814C8053204205108099080A743C809070883D",
      INIT_18 => X"0596A8858AA60CAA58004C066C60594203DB16B053201012505808208D03C468",
      INIT_19 => X"C818807D4458A0C2C202603D081702E6862888C460988FDF02089AD4164688C6",
      INIT_1A => X"420200A2B99B4C29286E640205F1CC088844081F49601684300F25132009D084",
      INIT_1B => X"C9C2831215A0C4856831215A0C4856831215A0C485683121593251515C730222",
      INIT_1C => X"203D4080904A20086864E4682C918096010081C30A0292C6442020EBD9160148",
      INIT_1D => X"0548232D623112344203115113204C82084015E8C94D930063204C94D5202448",
      INIT_1E => X"1080842348196501021064050170B2005553108554208C902010C06313012D42",
      INIT_1F => X"04C500542A464205692388F93219320523420569084206041080560084234606",
      INIT_20 => X"660408084234C2A548C8D63106851905632142433C9D654C965D54C5005B0A92",
      INIT_21 => X"00201E21706259615232358C576854080842348195C541C3003112361A235591",
      INIT_22 => X"005000100050140005055541515105505555514554414515441544554002020A",
      INIT_23 => X"0500145455514015051545000140050014001055514000514054500114005001",
      INIT_24 => X"4545554554515544005000055401555541414551400050515450001400500140",
      INIT_25 => X"FFF00C000000501394E93A4FC000000000000000000000000000000005041545",
      INIT_26 => X"FFFFFFFAAAAAAAA5555555500000000FFFFFFFFAAAAAAAA5555555500000000F",
      INIT_27 => X"093FFFFAAAAAAAA5555555500000000FFFFFFFFAAAAAAAA5555555500000000F",
      INIT_28 => X"0000000000000000000000000000000000000000000070000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(7 downto 6),      -- Port A 2-bit Data Output
      DOB => memBRead(7 downto 6),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(7 downto 6),      -- Port A 2-bit Data Input
      DIB => memBWrite(7 downto 6),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM4 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"02550195000200030077007600030359001E0003001C09DD000307EA00000064",
      INIT_01 => X"706555555755A365027600130001222837780003000300030003001600120005",
      INIT_02 => X"555709831042087800000000D355555554DA5555555536355555554D5AA46DF7",
      INIT_03 => X"5541AA00002A2800AC82A25506A8000000A8A00002A200018329555555559555",
      INIT_04 => X"A6956586F8AA55961BE2AAACA89541B85555060D555554AAC001822A2154A895",
      INIT_05 => X"15564C3A55961BE2A956586F8A6956586F8AA55961BE29A55961BE2A956586F8",
      INIT_06 => X"C4DD0F9C3E254D554C5A94D4A3500F07C1D00B5C330CF3C3F3CC5544DD52494A",
      INIT_07 => X"E1B5D755571D97818E76755CE71835646436755036461D5558E13248A5555D99",
      INIT_08 => X"DD953042010B03E0024CD486B931E7579D27491D5550765A0D55154409D21B5D",
      INIT_09 => X"4424F150D91D3714CDB070020425D4601515551100F8018994D19555114041D5",
      INIT_0A => X"75543554959F55D556679190489D554403E0072C4060DE140F41BA11D6E44451",
      INIT_0B => X"6845704D611544DC545704D5111C1371144C1DC79E5C71E113697174D0747754",
      INIT_0C => X"38344823553107174E413471697193C477905D84C7455344DE19D378574D9313",
      INIT_0D => X"55DD48483E1B310505675CCD58860351454104100F441D5552558C3655B95098",
      INIT_0E => X"65111AF8DD1AD055541D1D54F08F41D115509285CE0754B47450F82DDB5B6556",
      INIT_0F => X"D550499F18E4B076DA4214846A8499649843C3E382555435685D9495496C3106",
      INIT_10 => X"4DD55C3555001BD40D9110D5558C3701D5515951951D5114D0D2678221658145",
      INIT_11 => X"340D6B9445289AC434711C0F9F15CDD5515951951D5114D0D2678267C4950175",
      INIT_12 => X"F40D912D604235CD0D221D444356E005D550D1555381555500D97D875686A420",
      INIT_13 => X"80549BE357DF5D553D7DD55A1DD555D557D4336CD746A5475E5D6A216391175A",
      INIT_14 => X"010501F5405D40C8D5940C1435580D3849CE5740B18E1910340745C556881D5B",
      INIT_15 => X"9B4603E049D9C0084555521555D5710555774D34040D536B8421F9D453441141",
      INIT_16 => X"041175106E554455555F9551036500638510F943D169668356285678818E340F",
      INIT_17 => X"D8F98F98F98FDD00D920DD6A08440D9103545D563755637555C621AE0505C164",
      INIT_18 => X"1157D3918169757BC8590F9710611503950440C103644653210DD555BE179544",
      INIT_19 => X"D54C433594B0854455550145755140154527D89514BD8B95754C1CD64F0D1906",
      INIT_1A => X"5551405045830F8D75D16D155464110C4D99D918486C8049DD528503667CD750",
      INIT_1B => X"A3429553102554C409553102554C409553102554C4095531003C972139044313",
      INIT_1C => X"D151519E005111D94414170D204D0484CA4555500503216C59D5301C3526441B",
      INIT_1D => X"57046685066556A495D5DD4103D10D51773591C0DE4C83E503570DE4CD6B889D",
      INIT_1E => X"1775776F4CCF97A4766261D877D536396DC347407021AA255525558D03E7055D",
      INIT_1F => X"30F31DBD15BBDD56706F9BF83648357C6F5D547377B6FD0855545F35776F3A33",
      INIT_20 => X"8837575776B0C15859D9843C816FE39A4366411D28401C0D41F3E0FB1D9F4566",
      INIT_21 => X"07670D146590C32F1676610FF31267545776B40CCCCFC89D59D5A6E8DC6F2CDF",
      INIT_22 => X"CC30300C00300C000C320499A95208E1C4535A2755E92DCB882389238A427556",
      INIT_23 => X"000002951C50C080313003030BC02D003400811C50C002CB87E43003F803E300",
      INIT_24 => X"5841550C544F955C0740000C380831B1C14C8C00C0C023330030300800D00000",
      INIT_25 => X"FFF00C000000F01400FFEAB3C0000000000000003FFFFFFFEAAA9543850823A8",
      INIT_26 => X"555555555555555555555555555555500000000000000000000000000000000F",
      INIT_27 => X"3A3FFFFFFFFFFFFFFFFFFFFFFFFFFFFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA5",
      INIT_28 => X"00000000000000000000000000000000000000000000B0000000000000020000",
      INIT_29 => X"00000000000000000CE000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(9 downto 8),      -- Port A 2-bit Data Output
      DOB => memBRead(9 downto 8),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(9 downto 8),      -- Port A 2-bit Data Input
      DIB => memBWrite(9 downto 8),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM5 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"0028016800040002006B00A40002002500150002001500200002078500620060",
      INIT_01 => X"090555555A16501F0555001E00011554543400020002000200020008001C0004",
      INIT_02 => X"555A082282D08E55000000009355555555841555555561455555555058510938",
      INIT_03 => X"5564320000C598030D3C595590C80000031660000C58C0246FC1555555550555",
      INIT_04 => X"12084505C8182114172040DF165564345555903D55555715C0246FC58D571655",
      INIT_05 => X"96296A48211417206084505C81A084505C8182114172058211417206084505C8",
      INIT_06 => X"E18B5B896D1CD962A7546A5450CF5B71580861C4E138618E91B8586205916041",
      INIT_07 => X"17146758A54584656E0B18A04CF16646C1660945661A862854D183703F0F0588",
      INIT_08 => X"0582C0F063C156D030459915F861A18480718705961516185996751FBC617146",
      INIT_09 => X"378E9CA59823E272012C64BB400C144101558A49B5B4BD50710945615F380059",
      INIT_0A => X"1852855419554461645F509EE3462926D6D2F546F1595CCC5B756511B2343155",
      INIT_0B => X"B7702AFAD5CB6C8B1702AFAD9C0AB629CBD9C4BA28082E8CBEA02C8E801A1166",
      INIT_0C => X"0166AC531C4502C8D941902C80263E735D40066BA5723A8DA8CCBEA322DAFEBE",
      INIT_0D => X"A01240416D1107E5A19151016694527B3730C30C5B44061651A15D6601668510",
      INIT_0E => X"DA01D4D9861C12585D05065D2811A8519615D0104661940514C5B41453955451",
      INIT_0F => X"6168095D15E114149C58BE2F5542950D5956D6D080162966440614694692E3C5",
      INIT_10 => X"40628441544996DA5988A599654D643461695D65165D65D45596534A07012D74",
      INIT_11 => X"668D5784B55457D16459CA5B8496B061695D65165D65D4559653465304D4BC14",
      INIT_12 => X"CA5985D59F72958459207121566453606155996169016161A5985D5559451715",
      INIT_13 => X"4D5555D195940616913116116061606165B7295844555A2759A175215B85D555",
      INIT_14 => X"70B417352F056B6A715694656668C4C6756858D0D14D121D66E164A05D440611",
      INIT_15 => X"80ACD6D20058E080458A141616C58D8595B41041C55991577DC058B25D774D57",
      INIT_16 => X"A01F145855A314C58515165132DC89574495B80B0855514715545534054D025B",
      INIT_17 => X"17495497495C066598559D45356659889666462941859D185867416D14046975",
      INIT_18 => X"99524CDD7720192513505B84634995CA1454710996622409D9C0596565546840",
      INIT_19 => X"996DF895A74805A21616894518A86430CC0D5568440545001645484671C4D444",
      INIT_1A => X"561B22C94D195B472D1345162807D10000A4582043DF16F464514116627A61A5",
      INIT_1B => X"5100966998A59A662966998A59A662966998A59A66296699896E9892E1FC400C",
      INIT_1C => X"6545195D1AC85458697806A50148143DF1458A102C00D046646190140D247717",
      INIT_1D => X"280F5144451A15D51616D05456C1599118412815927256E196655927215B4460",
      INIT_1E => X"11858751486456951621685817855578511641A9DF0165016105845C16E02E06",
      INIT_1F => X"35B8051B0CB846294559D7456619664659462A441B75B441C587E5058759A619",
      INIT_20 => X"641759587598E0C15454556E8BAA56A5566140865C12B2596B3255B40507C305",
      INIT_21 => X"C1632BBD073618665515155B50B647595875948676CA8846106405D4D05DA420",
      INIT_22 => X"C030003C40F10C040D284715799040C1155498499FE9FDA30103010304C41658",
      INIT_23 => X"0D1036025D60C0F617D18300080422103440125D60C0420B00C4301190424003",
      INIT_24 => X"D0456C31905419FC4108000C300999F50245F460C000C14D1830003040D10344",
      INIT_25 => X"AAA00C000000002AAA555573EAAAAAAAAAAAAAAA955555555555555407010320",
      INIT_26 => X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA",
      INIT_27 => X"003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
      INIT_28 => X"0000000000000000000000000000000000000000000060000000000000020000",
      INIT_29 => X"00000000000000000CE000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(11 downto 10),      -- Port A 2-bit Data Output
      DOB => memBRead(11 downto 10),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(11 downto 10),      -- Port A 2-bit Data Input
      DIB => memBWrite(11 downto 10),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM6 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"00000000000000000001000200000000000200000002008800000300000000B0",
      INIT_01 => X"202000000800080A010000000000080202B20000000000000000000200000000",
      INIT_02 => X"0008A20300A00C02AAAAAAAA0B00000000020000000000000000000002002830",
      INIT_03 => X"0000B8AAAAC002AB2CBC000002E2AAAAAB000AAAAC0EEA800FC8000000000000",
      INIT_04 => X"84A000A0C2828002830A22CF000000B00000023C00000300EA800FC0EC030000",
      INIT_05 => X"000003028002830A0A000A0C284A000A0C2828002830A328002830A0A000A0C2",
      INIT_06 => X"3C0003000CA33000040300400B38030004028238020082002600000C8C080000",
      INIT_07 => X"8A08CB00028C0A803C31300EA08000208000200800208C0003C8380232828C02",
      INIT_08 => X"8C000B04881380C8800F0400B03803020093020C000A30280000202224C0A08C",
      INIT_09 => X"003914C000B6C0E02C000003000820C882A00080003200900D800800B802D8C0",
      INIT_0A => X"30003002B808C8C004033000800C020000C802409E0608CE03080080A00C0302",
      INIT_0B => X"C0D00083034C08010D100830340028034CB3403C3000030420C004DA00322302",
      INIT_0C => X"E0002A07384C004DB0C22004D00B6894C2820CAE22D364D8304820C120932820",
      INIT_0D => X"00E002C00C811C0028A3282C08228A2400CB2CB203C08C0000002C0008000200",
      INIT_0E => X"000E80CACC0B80002A0C0C80280088C20008800A22B32C0E30803220CB808800",
      INIT_0F => X"C002283E00C289320830C830042028000200C0C8200000002A8C80000022BC30",
      INIT_10 => X"88C0020880BB82C800080000003C02F8C0000C08408008008002032202088038",
      INIT_11 => X"022C0B02300202C0000020030A00B8C0000C0840800800800203220B08800010",
      INIT_12 => X"C8000A04800A12240020200280022F80C000000001080000200000010020A080",
      INIT_13 => X"BE8081C90A260C0010BA8008A8C000C00100A122401000030C0030880F0A0080",
      INIT_14 => X"0A00822000040020688002080028208008480200401C8A80002302800C200C08",
      INIT_15 => X"00A000C8D8C0C0800000028000E00C20200082082000080B202050200E020802",
      INIT_16 => X"000218020C02208000050088F8834C0F2A20300FB400002380C20072201CA803",
      INIT_17 => X"00882883881C8CB000200C008880000800028C00230002300003203C81004038",
      INIT_18 => X"000008428210320A080A03020820002200880A80000202B92028C00028000022",
      INIT_19 => X"00890210803420210000280A30001020B8C8C200000C1800302F82430A2083B2",
      INIT_1A => X"0000D0B68823032CC0A208000200000C20A8C0E000830008C800228000B06320",
      INIT_1B => X"0820808E8CA023A12808E84A023A12808E84A023A12808E8480C0B8AE0040304",
      INIT_1C => X"C808003C8233A0C00C30080800009008320000000B83A00828C0082808800001",
      INIT_1D => X"00B00820E0C000A08080022200C6000A322860C0083880C000020083800F2028",
      INIT_1E => X"E320230E188022AA300E24C13380203035000332ED0C20800080020E80C03C8C",
      INIT_1F => X"70320C8A08388C003602C18800000022028C00363330F3888002A2E0230A2220",
      INIT_20 => X"2263020230E1E0880182800C92308AAA0000384C8C202300C23220320C8B8220",
      INIT_21 => X"E303800A0100820A0060A003082303020230E18800DAB48C08C8B0E0C80202AA",
      INIT_22 => X"4AAA2AA4AAA2AA8AAB2AEEEAE2A12512CFEFA2FAAA8F2AA2C59444944F803000",
      INIT_23 => X"A32A8CAAABAAA8EF04892AA3AC4AB02AD0AAC2ABAAA8AB12CF7EAA2B4CA932AA",
      INIT_24 => X"AE8EEAAFA8FBFAA8AE94AAAAAC8FABAA8A81224AA8EA305892AA3A8CAAB2A8CA",
      INIT_25 => X"00000C000000100000000033C00000000000000000000000000000000A04944E",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"1500000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"00000000000000000000000000000000000000000000A0000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(13 downto 12),      -- Port A 2-bit Data Output
      DOB => memBRead(13 downto 12),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(13 downto 12),      -- Port A 2-bit Data Input
      DIB => memBWrite(13 downto 12),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM7 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"028200020002000000020081000001800000000000000A4600000320002A00CA",
      INIT_01 => X"905000000C800680020000080000444101710000000000000000001100000002",
      INIT_02 => X"000C51A6981A9A015555555587000000002140000000081000000006010850B2",
      INIT_03 => X"0001745555E001579D7E000005D15555578005555E0DD5410FE400000000A000",
      INIT_04 => X"4C521050D1414841434519CF80000172000005BC00000380D5410FE0DC038000",
      INIT_05 => X"00800311484143450521050D148521050D1414841434521484143450521050D1",
      INIT_06 => X"B21023208C60000808020082040823582DA15A0A0A828A202A0202024C040620",
      INIT_07 => X"5454C702054C25583CB23201564080111480B02080B14C8202C4451530504C29",
      INIT_08 => X"4C2CD70F843F88C6782C0E40B2442321A663258C008530942000508418C9454C",
      INIT_09 => X"90332AA202A8C4867C420A02E68152956550205C02310276425C64087C4124C0",
      INIT_0A => X"320900014031E4C8090F7980048C817008C409D4390C4DAD23442049465EBE08",
      INIT_0B => X"A6EA40229BAA42128EA40229BA900843AA22A93A69924E9A08A64AA22E319301",
      INIT_0C => X"1080551FB198A8AA21E92A8AA64A88A82A6D8C6B22EA88A329A508A694328808",
      INIT_0D => X"091921E08C46AC38145316580551649C4024924923E24C8008083C80A4202506",
      INIT_0E => X"809103D78C9C4802118C8C50462554C94085486515E31E1D32123198C7831708",
      INIT_0F => X"C805903D82C942314421C0700C1514904108C8C518408080114C42002005E000",
      INIT_10 => X"64C82514423FC3D4202E1200002C8134C8000C048048048202080B1484546834",
      INIT_11 => X"81380F25708102D882181023258074C8000C048048048202080B140BA642AAA2",
      INIT_12 => X"D42025987905A11A208844A948010368C80200080368080812025822081080C0",
      INIT_13 => X"0D4202C615198C803475408494C808C802D05A11A220C0A30C0830540B258202",
      INIT_14 => X"45A24450AAA8001ED44005148016322E0482011A9C2C554C8013056A0C128C84",
      INIT_15 => X"267108C424C2CAA22020854080D02C10102165961120040B501AB6060C09A404",
      INIT_16 => X"2A80668308085210208B405C3410A90B1512326F49010C17408110F1542C5423",
      INIT_17 => X"42102102103D4C6202520C204660202E08014C80932001320243982C52A28031",
      INIT_18 => X"800422C160763185560523251E58003082160568080B914B1814C00020820259",
      INIT_19 => X"00470222620A101A808054213206208A2193C202621C225A301FD1A305320225",
      INIT_1A => X"408028096013231C01580480818028AE6674C292201F5104C60814480A709312",
      INIT_1B => X"05A8405D4A5017529405D4A5017529405D4A5017529405D4A48D445D900A2B99",
      INIT_1C => X"C421882C5F0098C24E6697488A6D6201F520208A80EBD91434C81A9690E40082",
      INIT_1D => X"81700C11108080C14040851988D92005316491C20534C8C808012053440F1254",
      INIT_1E => X"1310130866891415309108C2332080B255482315568030580850212D48C9BC4C",
      INIT_1F => X"B2358C41A1714C810908C22080848011084C81093370B4E690215110130841A2",
      INIT_20 => X"119301013086DA150202108D206544150809068C5E980520407852358C576850",
      INIT_21 => X"D30B40018241451440808423460613010130866895E50E4C84C54086C6085545",
      INIT_22 => X"4410101440510404051545555151455155455154554145554515451540283001",
      INIT_23 => X"0510145455504015151141010144051054405055504040514154101054415101",
      INIT_24 => X"5445551554515554415400041401555541454450404051511410101440510144",
      INIT_25 => X"55500C000000D00000000033C000000000000000000000000000000005051544",
      INIT_26 => X"5555555555555555555555555555555555555555555555555555555555555555",
      INIT_27 => X"1515555555555555555555555555555555555555555555555555555555555555",
      INIT_28 => X"00000000000000000000000000000000000000000000E0000000000000010000",
      INIT_29 => X"00000000000000000CD000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(15 downto 14),      -- Port A 2-bit Data Output
      DOB => memBRead(15 downto 14),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(15 downto 14),      -- Port A 2-bit Data Input
      DIB => memBWrite(15 downto 14),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM8 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"015502550005000300F6005200030357002A0003002A066500030BDD001C000F",
      INIT_01 => X"793000000D4EC7C70123002F0001191522250003000300030003003D00060009",
      INIT_02 => X"000D601010C040A555555554DA00000001DCC000000077600000001645953DFD",
      INIT_03 => X"0024C9555693855A7CB92A00932555555A4E15556932D564899E00000000A000",
      INIT_04 => X"5D961BE2A956586F8AA567064E0024F0000093A4000002405564CB932C024A80",
      INIT_05 => X"5D510E56586F8AA55961BE2A955961BE2A956586F8AA566586F8AA55961BE2A9",
      INIT_06 => X"A2CD6E8D995445D50415505D54486DAC86F2014401004100D90F76420F951317",
      INIT_07 => X"1510D0756C0F85016A08356D69D1AE7545BE09D1BE090D551595211564540F86",
      INIT_08 => X"0F805644C511DB9595044165E874C364C783450F96543E146F9B074370D9510D",
      INIT_09 => X"D0059716B8C5137DC0372001534D13641227546416A51443126409D9590120F9",
      INIT_0A => X"36560854A95A40D9CF52944C950D51909A94912C5C5517E569C5555639E4D274",
      INIT_0B => X"1C5D34787171C74DC5D34787174D1531714974D1874D34571E113716083403E4",
      INIT_0C => X"11BC45059E74587172579D87113C5A54D9100D71F15C56148574D215D3785A1E",
      INIT_0D => X"57101951A951691C0443C079D85206791520820865500D917555498E15555D43",
      INIT_0E => X"5643D4020DC94C76460F0D54FD2FB0F89D9E0713B48365143E566570FDD56475",
      INIT_0F => X"D9515D4955A1203DB50398E455555344471A9996A41D51BE6B0D1D51D5B6B105",
      INIT_10 => X"10D5514C5D3FD4116B8D1639C1459E40D9C401D0DD3DD2DD36BE5659440CD400",
      INIT_11 => X"9F7C5E85475555A1AF08416284DD00D9F401D01D31D21D36BE56595B07104410",
      INIT_12 => X"016B86C4001110346B344830DAE76470D916F1D9C089D9C816783811755571F1",
      INIT_13 => X"905DD595B4040D9C0A341D9FD0D9C0D98D1111034FC55553757DD5545E865D17",
      INIT_14 => X"11907484261415500C0179A5BE6373A31C467445C5596D8D8C03C3F0755C0D9D",
      INIT_15 => X"83E4589420F845D51755749D9C37408777410410826F9657E7434002771C0034",
      INIT_16 => X"354053475556521764441D2BC0A4815E5456A851083F555955557525B559536A",
      INIT_17 => X"951951D5114D0D2678263DD55BD1678D58E60D5903659436431C1549535241DD",
      INIT_18 => X"44003B04E4403403010B6681900440719D0110345BE343C85440F9715CDD5515",
      INIT_19 => X"7986431374C5975D9D99B9D835502D49FC805555310551403E56034C107395E0",
      INIT_1A => X"9D9120C85C8066553413241D5C5014B168B0F8D350CD1D40D275549BE1100366",
      INIT_1B => X"54B49D071CE741C739D071CE741C739D071C2741C739D071CD815C8654051858",
      INIT_1C => X"D1D145596B4080F8C1518D8456E6310CD53754060C2C353430D91D85BC110115",
      INIT_1D => X"5264555525557571DDDD84001BD76B9437189636B0241BA01AE46B024D525D40",
      INIT_1E => X"0377485474C5E3903E3400F03FC755E86D59C3478B415575D96767055BA26C0D",
      INIT_1F => X"E6A10F207A310D5D0455154D8E21AE7F540D550437D5EC0C6767EA6748574D31",
      INIT_20 => X"EF2D7675C576C499D515DDAD233DBA2F18E0360D814C1E67410C66A10FB31265",
      INIT_21 => X"03E10116505841CC7565776BFB332B767485444C49EF430D90DD1554E856A57E",
      INIT_22 => X"060010B042F18004022C024D1C0C8C024C88055CCD9726B03330313015D43E70",
      INIT_23 => X"2E10B94C860800712F77200103040C105040C086080040C8029A0013B84AE10B",
      INIT_24 => X"7D02A0C02689FCD84294002EC00712EB68CBDDC80042C2F7720010B040210B84",
      INIT_25 => X"00008C00000000000000003CC0000000000000003FFFFFFFEAAA954349323032",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000C20000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(17 downto 16),      -- Port A 2-bit Data Output
      DOB => memBRead(17 downto 16),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(17 downto 16),      -- Port A 2-bit Data Input
      DIB => memBWrite(17 downto 16),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM9 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"009600160000000600E4009200060557000C0006000C02960006039300FA003A",
      INIT_01 => X"B5D000000581E4BC081000060000110A155A0006000600060006004200740002",
      INIT_02 => X"000959D19C274612555555558600000001AD000000006B60000000120541D009",
      INIT_03 => X"00176555560F45581050E6005D955555583D155560F955579000000000002000",
      INIT_04 => X"811417206084505C818201B03D00174C00005DC0000000331557D00F94003980",
      INIT_05 => X"05904844505C8182114172060811417206084505C818204505C8182114172060",
      INIT_06 => X"00B95D4956847059025610062B41597E299E04403812086A800816305B801AB3",
      INIT_07 => X"16159116405B452D7501664AC09D5E01854D00657D01599654685565C7F75B44",
      INIT_08 => X"5B405444511054691C433355D45496618696555B86456D155784919B25916159",
      INIT_09 => X"970A02C57472B208C4E68B5073F10827B8D166E7551A574890E7B45841D905B8",
      INIT_0A => X"6608B8000D640598E4514E75D5599B9D54695D15555904C55955628C08C3901A",
      INIT_0B => X"C00B65A3002C1BE880B25A3002E96FA02CB02E9C30CB670268CB22CAE16696E1",
      INIT_0C => X"356F85644232302C85304B02CBE7201284D6591C100B20C8302FA0CCBEB32C68",
      INIT_0D => X"5A1BF03D468501103796DC24564AC421C50C30C3550C59841859454D1161632D",
      INIT_0E => X"85D4D448590820161C5B595667C5A5B00581FCE8121643C16C95DA45B0D65418",
      INIT_0F => X"985951471451596F6CB8120458A153154515546A2F45996E0059061061011525",
      INIT_10 => X"659969F546555451534615B81D455DA5981400574554574665B551AAF5F542E5",
      INIT_11 => X"6E55514D618A545D4CF26151450565984400574554574665B151AA555CD50306",
      INIT_12 => X"615B4500879C03135F4F516357E04A6598053058E04058E495F4D4C818A5A16D",
      INIT_13 => X"2B06D5689712598E0D3485815598E5986439C031312585AA184862965D454615",
      INIT_14 => X"5C56557980C2D511356D69554E245A019110147CD1668D555F16CD6E18AD5981",
      INIT_15 => X"4547156A05B44C709165B5058C4155014151861854578151255C0A1E1890E155",
      INIT_16 => X"2C2148055859485162900507A804095DA5159403033C58A4458A051A45469451",
      INIT_17 => X"D65165D65D4559653465B062850D534657E159901662056619D03156BAC41061",
      INIT_18 => X"B40CA027558966CDB0B5594581EB405406459A4355D1A9405265B84963061695",
      INIT_19 => X"B88C400052E3616445894869665813035A621616A3C160716E0031309D5A160E",
      INIT_1A => X"85810003DF1055A137F7C24592C0B0534655B4753E2568459918A017D1809655",
      INIT_1B => X"2ABF45A916115A458456916115A458456916D15A4584569161554844B32CD4D2",
      INIT_1C => X"90665146A34835B4405B2243F45997E25841667C00140D3415982F3F5F100D16",
      INIT_1D => X"914458A14585B58D0505057316525381649A743537DD175394E25B7DD251A445",
      INIT_1E => X"564156596A42E5216D10D5B16F1195145157D6798BF562805801602E55501859",
      INIT_1F => X"55955BA2D8F159910159565D4D217E105A5995016785D8328160E61156594E90",
      INIT_20 => X"ED891416A5952D91D6561D652197FA6617D2065983117557579455155B50B645",
      INIT_21 => X"96D1C15CCF5965D07595875966192514156597A438065D59859925A5D55A7182",
      INIT_22 => X"86601098427198040F00102D2065F4638C0066147C25890194D197D1A48D6E32",
      INIT_23 => X"2F10BD01DBE980D133F4660103040C10F04001DBE98040CF435E60123048C109",
      INIT_24 => X"41CC71F0461277C043200020184454DCA90C7D198042D31F466010B440F10BC4",
      INIT_25 => X"00000C00000000000000003CEAAAAAAAAAAAAAAA95555555555555540D14D180",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000B70000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(19 downto 18),      -- Port A 2-bit Data Output
      DOB => memBRead(19 downto 18),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(19 downto 18),      -- Port A 2-bit Data Input
      DIB => memBWrite(19 downto 18),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM10 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"00000000000200000042000800000003000A0000000A00000000038300200000",
      INIT_01 => X"300AAAAAA020C232008800040000088008000000000000000000000800020000",
      INIT_02 => X"AAA00002000008000000000000AAAAAAA8042AAAAAAA010AAAAAAA8020080088",
      INIT_03 => X"AA800000008F00020208C0AA00000000023C000008F00000088CAAAAAAAA0AAA",
      INIT_04 => X"0002830A0A000A0C282820323C2A800CAAAA00E2AAAAAA330000C88F02AA302A",
      INIT_05 => X"8C0800000A0C2828002830A0A0002830A0A000A0C2828000A0C2828002830A0A",
      INIT_06 => X"00300020200000C0A1000A0C000002088CA200005C130CB400003000030080C3",
      INIT_07 => X"020002302E0320083088002282802C00880C88C83C880000C000083000800320",
      INIT_08 => X"0322C80CE030C20033203A80C2CB0000E00022030A800C830F0A2321A0082000",
      INIT_09 => X"020C00407253203845C00010EF0EF6002003008C60406000008C08C000200030",
      INIT_0A => X"000003AAA80820008C020809000002318101802138028CC00E20000838403030",
      INIT_0B => X"4202C0C108040C8010241C108090720804C0093413A20D00B042004C0C0000C0",
      INIT_0C => X"802D008C8E130004D020800042893401283000252C01344D1008344020C13030",
      INIT_0D => X"008A4000100000328380C228C82C20A028000000063200023000082C800000C0",
      INIT_0E => X"02A8408800BCD830040300828028A0328C009022AA0000000EA0800030C08030",
      INIT_0F => X"00A0000A0008280C031A0E8000000B8020C18000808C083C0A000C08C0A20800",
      INIT_10 => X"000000808C9540880F24C0F0A0183C8000A2A0C78C78C68C90B000080080A800",
      INIT_11 => X"0C100020230080883C080804208C8000A2A0C78C78C68C90B00008020822A882",
      INIT_12 => X"880720A2880288820F00008800C0A800008070C0C0A8C0C140320BE030002868",
      INIT_13 => X"A00C000080A0000C0A120C004000C000880028882000002E3028C0000C208C00",
      INIT_14 => X"02A03008AA200022008010800C001222002A3008243000041C40D082300C0002",
      INIT_15 => X"20808202003208CF6300308C0EA32823032C208220030202210210BA32028B30",
      INIT_16 => X"08D080B10000B62300200C028200260C0080C20B80FF0000000030003800020C",
      INIT_17 => X"C084080080080020322030C02A200B2401C0000880028000200AA000258210C8",
      INIT_18 => X"82A22200A08000200A0A0820C2282A1A8CA0000800C90280080030A00B8C0000",
      INIT_19 => X"7038030C21E023288C0238C80023663238A100000C2002080C000822021200A2",
      INIT_1A => X"8C0C088083000C003020CD8C08382EA2083032C0008420000A3000C0C8000020",
      INIT_1B => X"00F08C08A0A3022828C08A0A3022828C08A023022828C08A08280A2C0D0B6882",
      INIT_1C => X"00C800000108003200820121208428084F63002088280880B000FC0A230B8800",
      INIT_1D => X"088000002000300C8C0CB208838A0300000AA21072EA030B82C00F2EA2000820",
      INIT_1E => X"802328022802E2A80C8AE0300F2320023A02C0294F080038C023003C03080E00",
      INIT_1F => X"206003248E340008E002008C3C903C08020008E00380E000E30008A328021E00",
      INIT_20 => X"ECAA3232802208C0C0808C386200BAA2C3C8E20012002B0B0281206003082300",
      INIT_21 => X"00C82C04338C00893020230E2220EA32328022800A22AC00000AA020E00200AA",
      INIT_22 => X"8BAA2AC8AB22EA8AAA3AAAABAEF12242EAEEFAAAEAEAB9EB858904893FB00C38",
      INIT_23 => X"B62ADAAFAAAEA88604013AA2AD8AB62AA8AAA3AAAEA8AB6ECAA3AA299CAE72AC",
      INIT_24 => X"FA8BABAAF8BEAEACBAC0AABBF88B3FAB8FC1804EA8AB706013AA2ADCAA22AD8A",
      INIT_25 => X"00000C00000000000000003CC00000000000000000000000000000000B05893B",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"00000000000000000000000000000000000000000002C0000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(21 downto 20),      -- Port A 2-bit Data Output
      DOB => memBRead(21 downto 20),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(21 downto 20),      -- Port A 2-bit Data Input
      DIB => memBWrite(21 downto 20),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM11 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"010002800005000000C1008400000003002100000021040000000B0B00000080",
      INIT_01 => X"300555555818C13E024600280002446044400000000000000000001400210008",
      INIT_02 => X"5558001502C05488000000002055555554085555555502055555554490240A60",
      INIT_03 => X"55400000005F20014925C05500000000017C800005F080001652555555554555",
      INIT_04 => X"284143450521050D141494397C95402E555500D95555557B8000D65F09557015",
      INIT_05 => X"4C06A011050D1414841434505284143450521050D1414A1050D1414841434505",
      INIT_06 => X"08300810202228C05A80858C82220C544955A62AAEABAEBA2AA230A8232640C7",
      INIT_07 => X"81820930112311843064801515403C98683C64CC3C642000820254B002222311",
      INIT_08 => X"2319C42EE8BAC200709BF860C11608091088112325648C440F25531652041820",
      INIT_09 => X"0AAA64A0B1AA88B6AE80A0F9CB0D89600123002ED080D0A1082E04C2601C8232",
      INIT_0A => X"80B1F855540592024B086067802000BB42034297B9016AC008640821B6A83830",
      INIT_0B => X"A590C3A6964A7A3129083A696430E8864AA6423AE830CEA4A9A084AA0C8048C8",
      INIT_0C => X"402E609E6DA6824AA1855024A08AA99B160820AA6292A9AA6A4229A908A6A9E9",
      INIT_0D => X"0155C680202440B64308D144C55D125014820820088920293200203C44080420",
      INIT_0E => X"21158224204A263099232052441402364C257115550828288DD0801236C05232",
      INIT_0F => X"025008204204448D20BD0F420204075350030300404C042C95208C84C8591480",
      INIT_10 => X"120000824C6A82140F18C0B258202D42025358CF4CF4CF4C70F6080202425682",
      INIT_11 => X"2D2E0814132042102D960C0C114C42025358CF4CF4CF4C70F608020811195469",
      INIT_12 => X"140F1159658164C80B60264402C9144202E0B8C2CA74C2C6C0F140DA32001498",
      INIT_13 => X"508C820240D8202CA5A58C268202C2024698164C8BB0201D3214C8120C114C82",
      INIT_14 => X"41582246551A8099826834902C91209986B53201DC3018282FC8F041320C2024",
      INIT_15 => X"14404302823121C09300314C2D531653231C1041590B25085301B0E5318547A2",
      INIT_16 => X"812A614202024993081A8C9343921D0C01408167603C02062020808004200508",
      INIT_17 => X"C048048048202080B140B8C815580B1803C9200648096080914544201F19B8C4",
      INIT_18 => X"635309A05A60803045A50814A916352D4C51801602C6196216023258074C8000",
      INIT_19 => X"B2642B997AD453154C2904C48011F864F8BA80800C1809048C988C8B81208071",
      INIT_1A => X"4C2886A01F5A0808B007D24C040A0258047231C180889E2205320603C46A4810",
      INIT_1B => X"80704C945513251544C945513251544C945513251544C9455031215D42809601",
      INIT_1C => X"08C528201A2E02316950461B05582C08889300706A9690E6B2029C005E94E8C0",
      INIT_1D => X"044202085020302C4C8C718442140B248247C1B0F4D18206C3C90B4D15080612",
      INIT_1E => X"4813140150A9C5588C5692388F9310815542C81567040804C25309BC02058D20",
      INIT_1F => X"80842348197820041901405C3C782C95012004188320C6849309555314016C2A",
      INIT_20 => X"CC55313140158184C0404C219A25715003C510202846A50F6A46008423460610",
      INIT_21 => X"08C41C890A4D24963010130841A215313140150A91905D2022045012D6015414",
      INIT_22 => X"4050001400501400051411551455445144445554554505515511551140808CB4",
      INIT_23 => X"0500154555414015155545000500140050004155414001414154500154015001",
      INIT_24 => X"5545515054551554015400055445555541451551400051455450001400500140",
      INIT_25 => X"00000C00000000000000003CC000000000000000000000000000000001151151",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000300000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(23 downto 22),      -- Port A 2-bit Data Output
      DOB => memBRead(23 downto 22),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(23 downto 22),      -- Port A 2-bit Data Input
      DIB => memBWrite(23 downto 22),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM12 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"039A019A000D000B001200DA0007023A001E000F001E0FDA000F0BD9003C00CC",
      INIT_01 => X"B69555554C5750DF077600150001D65619160003000B0003000B007E00620009",
      INIT_02 => X"554C39042084105A00000001DD55555555D955555555769555555565615EB5BE",
      INIT_03 => X"554AAC0000192000620183552AB000000064800001B8800A0819555555549555",
      INIT_04 => X"686F8AA55961BE2A9565862064954A8855552A255555506A800A481B855060D5",
      INIT_05 => X"0F947491BE2A956586F8AA559686F8AA55961BE2A9565A1BE2A956586F8AA559",
      INIT_06 => X"55E4555D553130F9471D940D531356044986430CC330E31F333C3E346A848391",
      INIT_07 => X"35D6B03E5162555DD551BE454D416A32594950D1695D6F969D55D0B050106257",
      INIT_08 => X"6A55650674135555948D2557551899E1D319DC6686C599575286C34146735D6B",
      INIT_09 => X"0B511375E55C5CCB20300054564209022543E5E74557415004E410F8141746E8",
      INIT_0A => X"AE0A5E5545D396F84475FC1100639791155105719777D7445735D550CB8C5434",
      INIT_0B => X"704D5111C1371164C4DA119C13584551371134971C79E5D3C571D371018C5BA1",
      INIT_0C => X"994753E402D391371FF80D1371A5C46D51346795104DC671DD378774DE15C546",
      INIT_0D => X"5B5A9011555CD497541A5760FB60D8541C4D34D354C86B843665D9495DD99522",
      INIT_0E => X"64695D546782203E03646F924107E6D50F86A6360919C905A7E55556E49D9436",
      INIT_0F => X"B8440DDE1D5511B9048D4B53755C343160951559A40F957A056F0D90D94114C7",
      INIT_10 => X"D679D4140D155DD85255D5E851D14116B87360F80F80F00D0537757F43D40796",
      INIT_11 => X"7410755803559DF9600C1C55540FD6387360F80F80F00D0534757C75D144000D",
      INIT_12 => X"D8525415078455CE5804350557A1910638D530F845D0F840E5651B0C35474055",
      INIT_13 => X"450D5D5551C06F8451150F8B46F8467840C8455CEC0766083640D5A775540D9D",
      INIT_14 => X"C435C39600054001D41427915A29110183343D0001D5B8055FDAF500354C6B86",
      INIT_15 => X"5E50155F46A5765083E7050F8583D043C3C4D34D43568A75400001C83704D943",
      INIT_16 => X"092310E176738BC3E0850F1317C143755645556B5856754057556754DDD55B55",
      INIT_17 => X"1D05D35D25D36BE56595F0D52318565417A1679C5AE171AE108065D5B81070DC",
      INIT_18 => X"137710413751AC75D19455584241371D0D284586159535150C16284DD40D9740",
      INIT_19 => X"68B51C594F5503C60F85C0DDBE728B201C6CDD960905D341AA04DCE847119D04",
      INIT_1A => X"0F8C5FD0CDD555441033720F9048321F20C6655390C4D1167C355C5495C159F5",
      INIT_1B => X"54650F25F943C97E50F25F943C97E50F25F943C97E50F25F99553100D20C86C8",
      INIT_1C => X"B0D3CDD5C10D16651A0001CA4C27190C4C83E467FD85FC2686B8D90E8F841C1D",
      INIT_1D => X"9B517557476727680F0FB03495F05689BECE30C59D995556D6A05DD991756036",
      INIT_1E => X"9AC3CC76F058CBDDA96706F9BF837755E8D719DE3645D500F8C3E26C15549C6B",
      INIT_1F => X"75776F40CEB46F9098761DF5694D6A1D776B9C198FF7418483E18F83EC767C15",
      INIT_20 => X"CF6C3C3EC76E0CC7DD9D71515318703B9794416707741951E1AF35776F3A3327",
      INIT_21 => X"1995184149CDC7DFA76748564D310C3C3CC76F45BAFA416F86F01755E5775604",
      INIT_22 => X"C13000BC02E04C002D999D80225BDDC38B0652041E3E0C672F772F7700859A10",
      INIT_23 => X"3900D6125104C0BE1369130006001000D000C25104C001872DE13009E407500B",
      INIT_24 => X"9B24DA1D155701E2091800057049300F44449A44C003B116913000DC02D00F40",
      INIT_25 => X"00000C00000000000000003F00000000000000003FFFFFFFEAAA954314EF7729",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"00000000000000000000000000000000000000000002B0000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(25 downto 24),      -- Port A 2-bit Data Output
      DOB => memBRead(25 downto 24),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(25 downto 24),      -- Port A 2-bit Data Input
      DIB => memBWrite(25 downto 24),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM13 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"048000800000000200D00184000A017000000002000011200002000000180188",
      INIT_01 => X"7C5555555854138606440000000108641104000E0006000A0002005000C00000",
      INIT_02 => X"5558042D08A0B41A00000001AD555555549155555555E41555555541A0206648",
      INIT_03 => X"55715C000240F00919240F55C57000000903C000243480300640555555555555",
      INIT_04 => X"405C8182114172060845114903D571635555C5955555590C80300643455903D5",
      INIT_05 => X"5B801D017206084505C818211405C8182114172060845017206084505C818211",
      INIT_06 => X"CF9158A961AC95B82D05825991BD5A818146BA784E178E05EE196D1F5140921C",
      INIT_07 => X"B005756E115DA14862955E25811175003146959146905384061691264ACA55A0",
      INIT_08 => X"59A42C80120D1614043907018A5255D15255DD5D458556865145564855BB005F",
      INIT_09 => X"01CCB2259A0B2392C28EB25C2C44439D7556E1C065846DC42FC145B4B017F5D4",
      INIT_0A => X"5D045055085455F440192D596B5B87059615B7094314F0445810596FD2990D67",
      INIT_0B => X"2AFAD9C0AB629CBFAFADDC0ABEB572DBE2CBEB0208A280BA712A3A2C017F5451",
      INIT_0C => X"11556380E4B31F22CC8459F22A00B2C9AD2F53440AC8B22C8BAA332CA8CCB170",
      INIT_0D => X"20521D116161320750D75445BA63043113F3CF3C5A8353456600614680580100",
      INIT_0E => X"61C0465D5B55056D2C59536A410615565B4484160756D1354445850590451166",
      INIT_0F => X"34540464C6282165840F2FC01644185361165611845B8175155F598598574301",
      INIT_10 => X"95B81610590006D555A145D454614515B44D55B85B05B059451518414910F155",
      INIT_11 => X"754218A4566586A15676D758A25B95745945B85B05B05945151841195403B8C5",
      INIT_12 => X"D551A2D57526556851549CC515512185746555B44C55B454651AD2896651552D",
      INIT_13 => X"8559861581715344E5155B4405F4557449226556808162B96615991018A25946",
      INIT_14 => X"26810900EE302D971042C7156514441D7E116C47006114D165575485665C5744",
      INIT_15 => X"A0C05611F51A011016E3015B4416DC56D6D50410605144194847857167575649",
      INIT_16 => X"8501D75816390056D02C5B13154B001851558A06B000164401658184C0614458",
      INIT_17 => X"0574554574665B151AA515999DD755A194515B8256D1855D195248612057559C",
      INIT_18 => X"294541ADD1C95F545C0658A6DD729444592D35B5D46841BCF6D5145056598440",
      INIT_19 => X"149C18D3853DD6ED5B46C5954E2306988017058001305075452D168064440507",
      INIT_1A => X"5B45DE3E255C5866C889405B844000F7C4859A19500318D5F56654D4686755D5",
      INIT_1B => X"94C55B661556D98555B661556D98555B661556D98555B6615966998090003DF1",
      INIT_1C => X"3592E46160BFE5DAB10482E8425701001416E005E33F6F15057471E127141505",
      INIT_1D => X"80C9165B516301415B5B0701161251457D340D55D4531628D7525D4509184AA5",
      INIT_1E => X"16D6E0146835CA997694559D7456518A815556F59C405905B416D01856291657",
      INIT_1F => X"8587514864C4538C5A1605E146B57504145784994C01A31416D14956D0141E0C",
      INIT_20 => X"CD516D6D0145C6464505A965E90EB3E9566B0C5F1536A2596A25058759A61921",
      INIT_21 => X"5468563D4019C7D5514156594E90616D6E0146C37529415345B4115925148658",
      INIT_22 => X"01C0003000C07000268DD053D75C7D13203354162007003471F473F46485451C",
      INIT_23 => X"020009137507003F200E1C000C003400D00003750700030D29C1C00BC00F0003",
      INIT_24 => X"CC244C4D1D8522020A340015444E300FD448038700000200E1C0000002D00080",
      INIT_25 => X"00000C00000000000000003F2AAAAAAAAAAAAAAA95555555555555541931F475",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000300000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(27 downto 26),      -- Port A 2-bit Data Output
      DOB => memBRead(27 downto 26),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(27 downto 26),      -- Port A 2-bit Data Input
      DIB => memBWrite(27 downto 26),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM14 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"000A000A00020008000A0002000400B2000A0008000A008A000C000A00100010",
      INIT_01 => X"3C00000002000B2100020000000000020882000C000800000004000A00060002",
      INIT_02 => X"0002800A00C02800AAAAAAA80400000003080000000042000000000008082020",
      INIT_03 => X"00300EAAA808FAA00C008F00C03AAAAAA023EAAA80B02AB22008000000000000",
      INIT_04 => X"2A0C2828002830A0A000802023C0303B0000C0000000002E2AB2200B000023C0",
      INIT_05 => X"0302A00830A0A000A0C2828002A0C2828002830A0A000A830A0A000A0C282800",
      INIT_06 => X"322C0000000F2030098C00000AC20218800000408020003A00A00C9008220000",
      INIT_07 => X"3000B00C08080028C0002C008CC030B82000000000000B0A0C00001031310403",
      INIT_08 => X"080003203C800000000302230088C3CB2C00CF0420E030020020000200F3000F",
      INIT_09 => X"0284200000013410000200FB000402024000C082C002C087A08260320D0F0002",
      INIT_0A => X"1C88F20068CB00320032CA23C00F020B000B0203C230201A00B0C00610320001",
      INIT_0B => X"00830340024034CA0830340020C0D302C0420C0001C30028D0036C04002D0108",
      INIT_0C => X"CC390F8224230200473B002007401083A38D0B0080801204828C120B304810D1",
      INIT_0D => X"2B020380000CCE810202820030002ACC0B082082000003200008C80000C02802",
      INIT_0E => X"004C8C800F22000C8E0E072BB02AA0A003228022B000F80018400000228C0000",
      INIT_0F => X"7202A8CC8C002008E004CD363022A22F0A808008200300308807000000200D83",
      INIT_10 => X"4070A00200000C00000240C208C0188072012030030030004022302201020A80",
      INIT_11 => X"3802300200028CA00A8A040000030032012030030030004022302232C0A80B28",
      INIT_12 => X"000000000880004802201A200008A820F24020320800321260002A2000232800",
      INIT_13 => X"A0008C000C4A0B208080032230B210720008000488830208000000823000008C",
      INIT_14 => X"0008812A02CA808202280340308C0A8280900FC200C08BE03940902800240B22",
      INIT_15 => X"0234800B00400A0000C3A0032000C200C0C820820A0022322904885000800281",
      INIT_16 => X"2209082030310040C888038181680230000000030082302223002302E8C00200",
      INIT_17 => X"0C78C78C68C90B0000802000A02800020008070001C8203C880808C0A0281003",
      INIT_18 => X"A121A82029842D1002A00002420A1204002880CA000088080A004208C8000A2A",
      INIT_19 => X"0233E882882000C80320E0080C0E0A284C208C024008C0AC10800488800A8C00",
      INIT_1A => X"032E0CC0840800023421000303022020C080C00080C20BA070002200000E03C0",
      INIT_1B => X"0B000302E000C0B800302E000C0B800302E000C0B800302E0808E84000880830",
      INIT_1C => X"B002E8C088442000220300C83023800C1400C300CC0A33000032C00B0700280C",
      INIT_1D => X"003630032303A32803032088808800201CC82C30E08A000243080E0882302220",
      INIT_1E => X"82C0C8322820D2881003602C1880230035C081C88008C0A032C0C80E00000C0B",
      INIT_1F => X"20230E18800B030389304CE000303088320703880C23280000C88880C8322E08",
      INIT_20 => X"DE080C0C8320883A8C8CA008A00036AA8300AE0F0221300E1312E0230A2220E3",
      INIT_21 => X"03000BCE003CC3C2A32328021E00880C0C83228208AAA00720B0E32A223212A9",
      INIT_22 => X"0ABA2A90AA42AE8AB02AAEFA8AC18042EFAACFBAAB4AAEAB060104013F402082",
      INIT_23 => X"AC2AB3AAAEEAE8940911ABA2AB8AAE2AB8AAE2AEEAE8AAE84B2ABA2DB0A6C2A9",
      INIT_24 => X"AB4EAAEAB2AAAAB4BA84AAAAB08BAAAA2A42C46AE8AAD0B11ABA2AB4AB42AB0A",
      INIT_25 => X"00000C00000000000000003F000000000000000000000000000000002E06012A",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000170000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(29 downto 28),      -- Port A 2-bit Data Output
      DOB => memBRead(29 downto 28),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(29 downto 28),      -- Port A 2-bit Data Input
      DIB => memBWrite(29 downto 28),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
   ZPU_RAM15 : RAMB16_S2_S2
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"0", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"0", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      INIT_00 => X"012501250005000C00850021000C04790015000800150445000C06A500A20022",
      INIT_01 => X"3E0000000102861A0021001A000062014461000800080008000C000500090005",
      INIT_02 => X"00016181A9A606405555555408000000020400000000C1800000002406860012",
      INIT_03 => X"00380D555416F5504C816F00E0355555505BD555417215799015000000000000",
      INIT_04 => X"150D141484143450521044505BC038370000E0000000005D1579901720005BC0",
      INIT_05 => X"232560943450521050D141484150D1414841434505210543450521050D141484",
      INIT_06 => X"00220200080CA232424C242006C10156652140C2A0A8208A00A08C600C152802",
      INIT_07 => X"7960B48C94080954C8002C90603830464420020820060B290C804A2B0A8A0808",
      INIT_08 => X"0801A099B260808262038663204603C45802DC0C111020210811482500B7960F",
      INIT_09 => X"B21A08408092A834489A08F2B02D6019E008C8D9C021C81E70D9D231028F00C1",
      INIT_0A => X"3C65F50054C400B126310D53AA0B236700872053A93255150278C00D7442A482",
      INIT_0B => X"40229BA900843AA20229BA9008A6EA90C4A08A6493A69908EA4E884AE83E0304",
      INIT_0C => X"083213991D0B0084AC3620084E992813008A0B666021294A508A694329A528EA",
      INIT_0D => X"941900480802026609C30522351855428704104100200F1080A4C42028C29489",
      INIT_0E => X"09924C500B55848C49080F5E48945081231541904403C48021D020A0854C8880",
      INIT_0F => X"F11354CE4C829821D2282A093015515E4540408412232430540F202202542263",
      INIT_10 => X"C0B252C920AA8C820809A0C114C82140F11A123A23A23A20A08132192B490540",
      INIT_11 => X"31A9320188014C4821458A02082340F11A123A23A23A20A08132193189540F14",
      INIT_12 => X"82080840056000820852B53082055430F180823121423135908045108013168C",
      INIT_13 => X"50204C8060860B121484231580B130B12056000826630914809200493208204C",
      INIT_14 => X"60147B5503C56A444956B3C8304DAD4164688CA9A8C840D832822238801B0B15",
      INIT_15 => X"050A408700809D8A08CB58231148D108C8D65965050811315FBC68B48264017B",
      INIT_16 => X"3987081A30B361C8C641238A42DC6932092020630669301593001321D4C82502",
      INIT_17 => X"8CF4CF4CF4C70F60802082005016080982040F2403C4582C4D2424C852942208",
      INIT_18 => X"5A12D4581F1C3F2241500201C105A1AA20896085820254018580C114C4202535",
      INIT_19 => X"81709601658808D02311D2042C992E2EAE684C29A084C9682040482661AD4CA0",
      INIT_1A => X"231F1CC0888102070A2228232621A807D66080894AE65C90B4801182024003D0",
      INIT_1B => X"060023511408D445023511408D445023511408D4450235114405D4AA486A01F5",
      INIT_1C => X"F208D4C846C8108005EA29C4245760AE6A08CA81CC005E9120F1C00A4B12968C",
      INIT_1D => X"26093003130B531623235855404608102D249870C644408183040C6451321180",
      INIT_1E => X"42C8D6310685E5402010908C22081320554202D55024C0523108C58D80818C0F",
      INIT_1F => X"1013086689640B2442308CC820343062310B24402E93142648C56148D6315DA1",
      INIT_20 => X"ED148C8D631068854C4C500542A579414301690F86B5240C527110130841A213",
      INIT_21 => X"82028B29217CE3C1531314016C2A548C8D6310685441680F10F6131181315052",
      INIT_22 => X"4150005401505400051555515555155155055515155504555455555540A03041",
      INIT_23 => X"1100451145454055115515000500140050004145454001414151500144051005",
      INIT_24 => X"5544555515551154011400155405100554441545400111055150004400500440",
      INIT_25 => X"00000C00000000000000003F0000000000000000000000000000000015545555",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000300000000000000000000",
      INIT_29 => X"00000000000000000CC000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => memARead(31 downto 30),      -- Port A 2-bit Data Output
      DOB => memBRead(31 downto 30),      -- Port B 2-bit Data Output
      ADDRA => memAAddr(14 downto 2),  -- Port A 13-bit Address Input
      ADDRB => memBAddr(14 downto 2),  -- Port B 13-bit Address Input
      CLKA => clk,    -- Port A Clock
      CLKB => clk,    -- Port B Clock
      DIA => memAWrite(31 downto 30),      -- Port A 2-bit Data Input
      DIB => memBWrite(31 downto 30),      -- Port B 2-bit Data Input
      ENA => re,      -- Port A RAM Enable Input
      ENB => high,     -- PortB RAM Enable Input
      SSRA => low,    -- Port A Synchronous Set/Reset Input
      SSRB => low,    -- Port B Synchronous Set/Reset Input
      WEA => memAWriteEnable,      -- Port A Write Enable Input
      WEB => memBWriteEnable       -- Port B Write Enable Input
   );
end dualport_ram_arch;
