library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity DualPortRAM is
   generic(
      WORD_SIZE    : integer:=32;  -- Word Size 16/32
      BYTE_BITS    : integer:=2;   -- Bits used to address bytes
      BRAM_W       : integer:=15); -- Address Width
   port(
      clk_i     : in  std_logic;
      -- Port A
      a_we_i    : in  std_logic;
      a_addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      a_write_i : in  unsigned(WORD_SIZE-1 downto 0);
      a_read_o  : out unsigned(WORD_SIZE-1 downto 0);
      -- Port B
      b_we_i    : in  std_logic;
      b_addr_i  : in  unsigned(BRAM_W-1 downto BYTE_BITS);
      b_write_i : in  unsigned(WORD_SIZE-1 downto 0);
      b_read_o  : out unsigned(WORD_SIZE-1 downto 0));
end entity DualPortRAM;

architecture DualPort_Arch of DualPortRAM is
   type ram_type is array(natural range 0 to ((2**BRAM_W)/4)-1) of unsigned(WORD_SIZE-1 downto 0);

   shared variable ram : ram_type:=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80cd800c",
     3 => x"3a0b0b80",
     4 => x"c58f0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80c5d62d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80cc",
   162 => x"ec738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8b",
   171 => x"8a2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8c",
   179 => x"bc2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80ccfc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82c73f80",
   257 => x"c4913f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"fe3d0d0b",
   281 => x"0b80dce8",
   282 => x"08538413",
   283 => x"0870882a",
   284 => x"70810651",
   285 => x"52527080",
   286 => x"2ef03871",
   287 => x"81ff0680",
   288 => x"0c843d0d",
   289 => x"04ff3d0d",
   290 => x"0b0b80dc",
   291 => x"e8085271",
   292 => x"0870882a",
   293 => x"81327081",
   294 => x"06515151",
   295 => x"70f13873",
   296 => x"720c833d",
   297 => x"0d0480cc",
   298 => x"fc08802e",
   299 => x"a43880cd",
   300 => x"8008822e",
   301 => x"bd388380",
   302 => x"800b0b0b",
   303 => x"80dce80c",
   304 => x"82a0800b",
   305 => x"80dcec0c",
   306 => x"8290800b",
   307 => x"80dcf00c",
   308 => x"04f88080",
   309 => x"80a40b0b",
   310 => x"0b80dce8",
   311 => x"0cf88080",
   312 => x"82800b80",
   313 => x"dcec0cf8",
   314 => x"80808480",
   315 => x"0b80dcf0",
   316 => x"0c0480c0",
   317 => x"a8808c0b",
   318 => x"0b0b80dc",
   319 => x"e80c80c0",
   320 => x"a880940b",
   321 => x"80dcec0c",
   322 => x"0b0b80cc",
   323 => x"c40b80dc",
   324 => x"f00c04ff",
   325 => x"3d0d80dc",
   326 => x"f4335170",
   327 => x"a73880cd",
   328 => x"88087008",
   329 => x"52527080",
   330 => x"2e943884",
   331 => x"1280cd88",
   332 => x"0c702d80",
   333 => x"cd880870",
   334 => x"08525270",
   335 => x"ee38810b",
   336 => x"80dcf434",
   337 => x"833d0d04",
   338 => x"04803d0d",
   339 => x"0b0b80dc",
   340 => x"e408802e",
   341 => x"8e380b0b",
   342 => x"0b0b800b",
   343 => x"802e0981",
   344 => x"06853882",
   345 => x"3d0d040b",
   346 => x"0b80dce4",
   347 => x"510b0b0b",
   348 => x"f58e3f82",
   349 => x"3d0d0404",
   350 => x"803d0d80",
   351 => x"ccc85185",
   352 => x"de3f800b",
   353 => x"800c823d",
   354 => x"0d048c08",
   355 => x"028c0cf9",
   356 => x"3d0d800b",
   357 => x"8c08fc05",
   358 => x"0c8c0888",
   359 => x"05088025",
   360 => x"ab388c08",
   361 => x"88050830",
   362 => x"8c088805",
   363 => x"0c800b8c",
   364 => x"08f4050c",
   365 => x"8c08fc05",
   366 => x"08883881",
   367 => x"0b8c08f4",
   368 => x"050c8c08",
   369 => x"f405088c",
   370 => x"08fc050c",
   371 => x"8c088c05",
   372 => x"088025ab",
   373 => x"388c088c",
   374 => x"0508308c",
   375 => x"088c050c",
   376 => x"800b8c08",
   377 => x"f0050c8c",
   378 => x"08fc0508",
   379 => x"8838810b",
   380 => x"8c08f005",
   381 => x"0c8c08f0",
   382 => x"05088c08",
   383 => x"fc050c80",
   384 => x"538c088c",
   385 => x"0508528c",
   386 => x"08880508",
   387 => x"5181a73f",
   388 => x"8008708c",
   389 => x"08f8050c",
   390 => x"548c08fc",
   391 => x"0508802e",
   392 => x"8c388c08",
   393 => x"f8050830",
   394 => x"8c08f805",
   395 => x"0c8c08f8",
   396 => x"05087080",
   397 => x"0c54893d",
   398 => x"0d8c0c04",
   399 => x"8c08028c",
   400 => x"0cfb3d0d",
   401 => x"800b8c08",
   402 => x"fc050c8c",
   403 => x"08880508",
   404 => x"80259338",
   405 => x"8c088805",
   406 => x"08308c08",
   407 => x"88050c81",
   408 => x"0b8c08fc",
   409 => x"050c8c08",
   410 => x"8c050880",
   411 => x"258c388c",
   412 => x"088c0508",
   413 => x"308c088c",
   414 => x"050c8153",
   415 => x"8c088c05",
   416 => x"08528c08",
   417 => x"88050851",
   418 => x"ad3f8008",
   419 => x"708c08f8",
   420 => x"050c548c",
   421 => x"08fc0508",
   422 => x"802e8c38",
   423 => x"8c08f805",
   424 => x"08308c08",
   425 => x"f8050c8c",
   426 => x"08f80508",
   427 => x"70800c54",
   428 => x"873d0d8c",
   429 => x"0c048c08",
   430 => x"028c0cfd",
   431 => x"3d0d810b",
   432 => x"8c08fc05",
   433 => x"0c800b8c",
   434 => x"08f8050c",
   435 => x"8c088c05",
   436 => x"088c0888",
   437 => x"050827ac",
   438 => x"388c08fc",
   439 => x"0508802e",
   440 => x"a338800b",
   441 => x"8c088c05",
   442 => x"08249938",
   443 => x"8c088c05",
   444 => x"08108c08",
   445 => x"8c050c8c",
   446 => x"08fc0508",
   447 => x"108c08fc",
   448 => x"050cc939",
   449 => x"8c08fc05",
   450 => x"08802e80",
   451 => x"c9388c08",
   452 => x"8c05088c",
   453 => x"08880508",
   454 => x"26a1388c",
   455 => x"08880508",
   456 => x"8c088c05",
   457 => x"08318c08",
   458 => x"88050c8c",
   459 => x"08f80508",
   460 => x"8c08fc05",
   461 => x"08078c08",
   462 => x"f8050c8c",
   463 => x"08fc0508",
   464 => x"812a8c08",
   465 => x"fc050c8c",
   466 => x"088c0508",
   467 => x"812a8c08",
   468 => x"8c050cff",
   469 => x"af398c08",
   470 => x"90050880",
   471 => x"2e8f388c",
   472 => x"08880508",
   473 => x"708c08f4",
   474 => x"050c518d",
   475 => x"398c08f8",
   476 => x"0508708c",
   477 => x"08f4050c",
   478 => x"518c08f4",
   479 => x"0508800c",
   480 => x"853d0d8c",
   481 => x"0c04fc3d",
   482 => x"0d767079",
   483 => x"7b555555",
   484 => x"558f7227",
   485 => x"8c387275",
   486 => x"07830651",
   487 => x"70802ea7",
   488 => x"38ff1252",
   489 => x"71ff2e98",
   490 => x"38727081",
   491 => x"05543374",
   492 => x"70810556",
   493 => x"34ff1252",
   494 => x"71ff2e09",
   495 => x"8106ea38",
   496 => x"74800c86",
   497 => x"3d0d0474",
   498 => x"51727084",
   499 => x"05540871",
   500 => x"70840553",
   501 => x"0c727084",
   502 => x"05540871",
   503 => x"70840553",
   504 => x"0c727084",
   505 => x"05540871",
   506 => x"70840553",
   507 => x"0c727084",
   508 => x"05540871",
   509 => x"70840553",
   510 => x"0cf01252",
   511 => x"718f26c9",
   512 => x"38837227",
   513 => x"95387270",
   514 => x"84055408",
   515 => x"71708405",
   516 => x"530cfc12",
   517 => x"52718326",
   518 => x"ed387054",
   519 => x"ff8339f7",
   520 => x"3d0d7c70",
   521 => x"525380c8",
   522 => x"3f725480",
   523 => x"085580cc",
   524 => x"d8568157",
   525 => x"80088105",
   526 => x"5a8b3de4",
   527 => x"11595382",
   528 => x"59f41352",
   529 => x"7b881108",
   530 => x"52538183",
   531 => x"3f800830",
   532 => x"70800807",
   533 => x"9f2c8a07",
   534 => x"800c538b",
   535 => x"3d0d04ff",
   536 => x"3d0d7352",
   537 => x"80cd8c08",
   538 => x"51ffb43f",
   539 => x"833d0d04",
   540 => x"fd3d0d75",
   541 => x"70718306",
   542 => x"53555270",
   543 => x"b8387170",
   544 => x"087009f7",
   545 => x"fbfdff12",
   546 => x"0670f884",
   547 => x"82818006",
   548 => x"51515253",
   549 => x"709d3884",
   550 => x"13700870",
   551 => x"09f7fbfd",
   552 => x"ff120670",
   553 => x"f8848281",
   554 => x"80065151",
   555 => x"52537080",
   556 => x"2ee53872",
   557 => x"52713351",
   558 => x"70802e8a",
   559 => x"38811270",
   560 => x"33525270",
   561 => x"f8387174",
   562 => x"31800c85",
   563 => x"3d0d04f2",
   564 => x"3d0d6062",
   565 => x"88110870",
   566 => x"57575f5a",
   567 => x"74802e81",
   568 => x"90388c1a",
   569 => x"2270832a",
   570 => x"81327081",
   571 => x"06515558",
   572 => x"73863890",
   573 => x"1a089138",
   574 => x"795190a2",
   575 => x"3fff5480",
   576 => x"0880ee38",
   577 => x"8c1a2258",
   578 => x"7d085780",
   579 => x"7883ffff",
   580 => x"06700a10",
   581 => x"0a708106",
   582 => x"51565755",
   583 => x"73752e80",
   584 => x"d7387490",
   585 => x"38760884",
   586 => x"18088819",
   587 => x"59565974",
   588 => x"802ef238",
   589 => x"74548880",
   590 => x"75278438",
   591 => x"88805473",
   592 => x"5378529c",
   593 => x"1a0851a4",
   594 => x"1a085473",
   595 => x"2d800b80",
   596 => x"082582e6",
   597 => x"38800819",
   598 => x"75800831",
   599 => x"7f880508",
   600 => x"80083170",
   601 => x"6188050c",
   602 => x"56565973",
   603 => x"ffb43880",
   604 => x"5473800c",
   605 => x"903d0d04",
   606 => x"75813270",
   607 => x"81067641",
   608 => x"51547380",
   609 => x"2e81c138",
   610 => x"74903876",
   611 => x"08841808",
   612 => x"88195956",
   613 => x"5974802e",
   614 => x"f238881a",
   615 => x"087883ff",
   616 => x"ff067089",
   617 => x"2a708106",
   618 => x"51565956",
   619 => x"73802e82",
   620 => x"fa387575",
   621 => x"278d3877",
   622 => x"872a7081",
   623 => x"06515473",
   624 => x"82b53874",
   625 => x"76278338",
   626 => x"74567553",
   627 => x"78527908",
   628 => x"5185823f",
   629 => x"881a0876",
   630 => x"31881b0c",
   631 => x"7908167a",
   632 => x"0c745675",
   633 => x"19757731",
   634 => x"7f880508",
   635 => x"78317061",
   636 => x"88050c56",
   637 => x"56597380",
   638 => x"2efef438",
   639 => x"8c1a2258",
   640 => x"ff863977",
   641 => x"78547953",
   642 => x"7b525684",
   643 => x"c83f881a",
   644 => x"08783188",
   645 => x"1b0c7908",
   646 => x"187a0c7c",
   647 => x"76315d7c",
   648 => x"8e387951",
   649 => x"8fdc3f80",
   650 => x"08818f38",
   651 => x"80085f75",
   652 => x"19757731",
   653 => x"7f880508",
   654 => x"78317061",
   655 => x"88050c56",
   656 => x"56597380",
   657 => x"2efea838",
   658 => x"74818338",
   659 => x"76088418",
   660 => x"08881959",
   661 => x"56597480",
   662 => x"2ef23874",
   663 => x"538a5278",
   664 => x"5182d33f",
   665 => x"80087931",
   666 => x"81055d80",
   667 => x"08843881",
   668 => x"155d815f",
   669 => x"7c58747d",
   670 => x"27833874",
   671 => x"58941a08",
   672 => x"881b0811",
   673 => x"575c807a",
   674 => x"085c5490",
   675 => x"1a087b27",
   676 => x"83388154",
   677 => x"75782584",
   678 => x"3873ba38",
   679 => x"7b7824fe",
   680 => x"e2387b53",
   681 => x"78529c1a",
   682 => x"0851a41a",
   683 => x"0854732d",
   684 => x"80085680",
   685 => x"088024fe",
   686 => x"e2388c1a",
   687 => x"2280c007",
   688 => x"54738c1b",
   689 => x"23ff5473",
   690 => x"800c903d",
   691 => x"0d047eff",
   692 => x"a338ff87",
   693 => x"39755378",
   694 => x"527a5182",
   695 => x"f83f7908",
   696 => x"167a0c79",
   697 => x"518e9b3f",
   698 => x"8008cf38",
   699 => x"7c76315d",
   700 => x"7cfebc38",
   701 => x"feac3990",
   702 => x"1a087a08",
   703 => x"71317611",
   704 => x"70565a57",
   705 => x"5280cd8c",
   706 => x"0851848c",
   707 => x"3f800880",
   708 => x"2effa738",
   709 => x"8008901b",
   710 => x"0c800816",
   711 => x"7a0c7794",
   712 => x"1b0c7488",
   713 => x"1b0c7456",
   714 => x"fd993979",
   715 => x"0858901a",
   716 => x"08782783",
   717 => x"38815475",
   718 => x"75278438",
   719 => x"73b33894",
   720 => x"1a085675",
   721 => x"752680d3",
   722 => x"38755378",
   723 => x"529c1a08",
   724 => x"51a41a08",
   725 => x"54732d80",
   726 => x"08568008",
   727 => x"8024fd83",
   728 => x"388c1a22",
   729 => x"80c00754",
   730 => x"738c1b23",
   731 => x"ff54fed7",
   732 => x"39755378",
   733 => x"52775181",
   734 => x"dc3f7908",
   735 => x"167a0c79",
   736 => x"518cff3f",
   737 => x"8008802e",
   738 => x"fcd9388c",
   739 => x"1a2280c0",
   740 => x"0754738c",
   741 => x"1b23ff54",
   742 => x"fead3974",
   743 => x"75547953",
   744 => x"78525681",
   745 => x"b03f881a",
   746 => x"08753188",
   747 => x"1b0c7908",
   748 => x"157a0cfc",
   749 => x"ae39fa3d",
   750 => x"0d7a7902",
   751 => x"8805a705",
   752 => x"33565253",
   753 => x"8373278a",
   754 => x"38708306",
   755 => x"5271802e",
   756 => x"a838ff13",
   757 => x"5372ff2e",
   758 => x"97387033",
   759 => x"5273722e",
   760 => x"91388111",
   761 => x"ff145451",
   762 => x"72ff2e09",
   763 => x"8106eb38",
   764 => x"80517080",
   765 => x"0c883d0d",
   766 => x"04707257",
   767 => x"55835175",
   768 => x"82802914",
   769 => x"ff125256",
   770 => x"708025f3",
   771 => x"38837327",
   772 => x"bf387408",
   773 => x"76327009",
   774 => x"f7fbfdff",
   775 => x"120670f8",
   776 => x"84828180",
   777 => x"06515151",
   778 => x"70802e99",
   779 => x"38745180",
   780 => x"52703357",
   781 => x"73772eff",
   782 => x"b9388111",
   783 => x"81135351",
   784 => x"837227ed",
   785 => x"38fc1384",
   786 => x"16565372",
   787 => x"8326c338",
   788 => x"7451fefe",
   789 => x"39fa3d0d",
   790 => x"787a7c72",
   791 => x"72725757",
   792 => x"57595656",
   793 => x"747627b2",
   794 => x"38761551",
   795 => x"757127aa",
   796 => x"38707717",
   797 => x"ff145455",
   798 => x"5371ff2e",
   799 => x"9638ff14",
   800 => x"ff145454",
   801 => x"72337434",
   802 => x"ff125271",
   803 => x"ff2e0981",
   804 => x"06ec3875",
   805 => x"800c883d",
   806 => x"0d04768f",
   807 => x"269738ff",
   808 => x"125271ff",
   809 => x"2eed3872",
   810 => x"70810554",
   811 => x"33747081",
   812 => x"055634eb",
   813 => x"39747607",
   814 => x"83065170",
   815 => x"e2387575",
   816 => x"54517270",
   817 => x"84055408",
   818 => x"71708405",
   819 => x"530c7270",
   820 => x"84055408",
   821 => x"71708405",
   822 => x"530c7270",
   823 => x"84055408",
   824 => x"71708405",
   825 => x"530c7270",
   826 => x"84055408",
   827 => x"71708405",
   828 => x"530cf012",
   829 => x"52718f26",
   830 => x"c9388372",
   831 => x"27953872",
   832 => x"70840554",
   833 => x"08717084",
   834 => x"05530cfc",
   835 => x"12527183",
   836 => x"26ed3870",
   837 => x"54ff8839",
   838 => x"ef3d0d63",
   839 => x"6567405d",
   840 => x"427b802e",
   841 => x"84fa3861",
   842 => x"51a5b63f",
   843 => x"f81c7084",
   844 => x"120870fc",
   845 => x"0670628b",
   846 => x"0570f806",
   847 => x"4159455b",
   848 => x"5c415796",
   849 => x"742782c3",
   850 => x"38807b24",
   851 => x"7e7c2607",
   852 => x"59805478",
   853 => x"742e0981",
   854 => x"0682a938",
   855 => x"777b2581",
   856 => x"fc387717",
   857 => x"80d4c80b",
   858 => x"8805085e",
   859 => x"567c762e",
   860 => x"84bd3884",
   861 => x"160870fe",
   862 => x"06178411",
   863 => x"08810651",
   864 => x"55557382",
   865 => x"8b3874fc",
   866 => x"06597c76",
   867 => x"2e84dd38",
   868 => x"77195f7e",
   869 => x"7b2581fd",
   870 => x"38798106",
   871 => x"547382bf",
   872 => x"38767708",
   873 => x"31841108",
   874 => x"fc06565a",
   875 => x"75802e91",
   876 => x"387c762e",
   877 => x"84ea3874",
   878 => x"19185978",
   879 => x"7b258489",
   880 => x"3879802e",
   881 => x"82993877",
   882 => x"15567a76",
   883 => x"24829038",
   884 => x"8c1a0888",
   885 => x"1b08718c",
   886 => x"120c8812",
   887 => x"0c557976",
   888 => x"59578817",
   889 => x"61fc0557",
   890 => x"5975a426",
   891 => x"85ef387b",
   892 => x"79555593",
   893 => x"762780c9",
   894 => x"387b7084",
   895 => x"055d087c",
   896 => x"56790c74",
   897 => x"70840556",
   898 => x"088c180c",
   899 => x"9017549b",
   900 => x"7627ae38",
   901 => x"74708405",
   902 => x"5608740c",
   903 => x"74708405",
   904 => x"56089418",
   905 => x"0c981754",
   906 => x"a3762795",
   907 => x"38747084",
   908 => x"05560874",
   909 => x"0c747084",
   910 => x"0556089c",
   911 => x"180ca017",
   912 => x"54747084",
   913 => x"05560874",
   914 => x"70840556",
   915 => x"0c747084",
   916 => x"05560874",
   917 => x"70840556",
   918 => x"0c740874",
   919 => x"0c777b31",
   920 => x"56758f26",
   921 => x"80c93884",
   922 => x"17088106",
   923 => x"78078418",
   924 => x"0c771784",
   925 => x"11088107",
   926 => x"84120c54",
   927 => x"6151a2e2",
   928 => x"3f881754",
   929 => x"73800c93",
   930 => x"3d0d0490",
   931 => x"5bfdba39",
   932 => x"7856fe85",
   933 => x"398c1608",
   934 => x"88170871",
   935 => x"8c120c88",
   936 => x"120c557e",
   937 => x"707c3157",
   938 => x"588f7627",
   939 => x"ffb9387a",
   940 => x"17841808",
   941 => x"81067c07",
   942 => x"84190c76",
   943 => x"81078412",
   944 => x"0c761184",
   945 => x"11088107",
   946 => x"84120c55",
   947 => x"88055261",
   948 => x"518cf73f",
   949 => x"6151a28a",
   950 => x"3f881754",
   951 => x"ffa6397d",
   952 => x"52615194",
   953 => x"f73f8008",
   954 => x"59800880",
   955 => x"2e81a338",
   956 => x"8008f805",
   957 => x"60840508",
   958 => x"fe066105",
   959 => x"55577674",
   960 => x"2e83e638",
   961 => x"fc185675",
   962 => x"a42681aa",
   963 => x"387b8008",
   964 => x"55559376",
   965 => x"2780d838",
   966 => x"74708405",
   967 => x"56088008",
   968 => x"70840580",
   969 => x"0c0c8008",
   970 => x"75708405",
   971 => x"57087170",
   972 => x"8405530c",
   973 => x"549b7627",
   974 => x"b6387470",
   975 => x"84055608",
   976 => x"74708405",
   977 => x"560c7470",
   978 => x"84055608",
   979 => x"74708405",
   980 => x"560ca376",
   981 => x"27993874",
   982 => x"70840556",
   983 => x"08747084",
   984 => x"05560c74",
   985 => x"70840556",
   986 => x"08747084",
   987 => x"05560c74",
   988 => x"70840556",
   989 => x"08747084",
   990 => x"05560c74",
   991 => x"70840556",
   992 => x"08747084",
   993 => x"05560c74",
   994 => x"08740c7b",
   995 => x"5261518b",
   996 => x"b93f6151",
   997 => x"a0cc3f78",
   998 => x"5473800c",
   999 => x"933d0d04",
  1000 => x"7d526151",
  1001 => x"93b63f80",
  1002 => x"08800c93",
  1003 => x"3d0d0484",
  1004 => x"160855fb",
  1005 => x"d1397553",
  1006 => x"7b528008",
  1007 => x"51efc73f",
  1008 => x"7b526151",
  1009 => x"8b843fca",
  1010 => x"398c1608",
  1011 => x"88170871",
  1012 => x"8c120c88",
  1013 => x"120c558c",
  1014 => x"1a08881b",
  1015 => x"08718c12",
  1016 => x"0c88120c",
  1017 => x"55797959",
  1018 => x"57fbf739",
  1019 => x"7719901c",
  1020 => x"55557375",
  1021 => x"24fba238",
  1022 => x"7a177080",
  1023 => x"d4c80b88",
  1024 => x"050c757c",
  1025 => x"31810784",
  1026 => x"120c5d84",
  1027 => x"17088106",
  1028 => x"7b078418",
  1029 => x"0c61519f",
  1030 => x"c93f8817",
  1031 => x"54fce539",
  1032 => x"74191890",
  1033 => x"1c555d73",
  1034 => x"7d24fb95",
  1035 => x"388c1a08",
  1036 => x"881b0871",
  1037 => x"8c120c88",
  1038 => x"120c5588",
  1039 => x"1a61fc05",
  1040 => x"575975a4",
  1041 => x"2681ae38",
  1042 => x"7b795555",
  1043 => x"93762780",
  1044 => x"c9387b70",
  1045 => x"84055d08",
  1046 => x"7c56790c",
  1047 => x"74708405",
  1048 => x"56088c1b",
  1049 => x"0c901a54",
  1050 => x"9b7627ae",
  1051 => x"38747084",
  1052 => x"05560874",
  1053 => x"0c747084",
  1054 => x"05560894",
  1055 => x"1b0c981a",
  1056 => x"54a37627",
  1057 => x"95387470",
  1058 => x"84055608",
  1059 => x"740c7470",
  1060 => x"84055608",
  1061 => x"9c1b0ca0",
  1062 => x"1a547470",
  1063 => x"84055608",
  1064 => x"74708405",
  1065 => x"560c7470",
  1066 => x"84055608",
  1067 => x"74708405",
  1068 => x"560c7408",
  1069 => x"740c7a1a",
  1070 => x"7080d4c8",
  1071 => x"0b88050c",
  1072 => x"7d7c3181",
  1073 => x"0784120c",
  1074 => x"54841a08",
  1075 => x"81067b07",
  1076 => x"841b0c61",
  1077 => x"519e8b3f",
  1078 => x"7854fdbd",
  1079 => x"3975537b",
  1080 => x"527851ed",
  1081 => x"a13ffaf5",
  1082 => x"39841708",
  1083 => x"fc061860",
  1084 => x"5858fae9",
  1085 => x"3975537b",
  1086 => x"527851ed",
  1087 => x"893f7a1a",
  1088 => x"7080d4c8",
  1089 => x"0b88050c",
  1090 => x"7d7c3181",
  1091 => x"0784120c",
  1092 => x"54841a08",
  1093 => x"81067b07",
  1094 => x"841b0cff",
  1095 => x"b639fa3d",
  1096 => x"0d7880cd",
  1097 => x"8c085455",
  1098 => x"b8130880",
  1099 => x"2e81b638",
  1100 => x"8c152270",
  1101 => x"83ffff06",
  1102 => x"70832a81",
  1103 => x"32708106",
  1104 => x"51555556",
  1105 => x"72802e80",
  1106 => x"dc387384",
  1107 => x"2a813281",
  1108 => x"0657ff53",
  1109 => x"7680f738",
  1110 => x"73822a70",
  1111 => x"81065153",
  1112 => x"72802eb9",
  1113 => x"38b01508",
  1114 => x"5473802e",
  1115 => x"9c3880c0",
  1116 => x"15537373",
  1117 => x"2e8f3873",
  1118 => x"5280cd8c",
  1119 => x"085187ca",
  1120 => x"3f8c1522",
  1121 => x"5676b016",
  1122 => x"0c75db06",
  1123 => x"53728c16",
  1124 => x"23800b84",
  1125 => x"160c9015",
  1126 => x"08750c72",
  1127 => x"56758807",
  1128 => x"53728c16",
  1129 => x"23901508",
  1130 => x"802e80c1",
  1131 => x"388c1522",
  1132 => x"70810655",
  1133 => x"53739e38",
  1134 => x"720a100a",
  1135 => x"70810651",
  1136 => x"53728538",
  1137 => x"94150854",
  1138 => x"7388160c",
  1139 => x"80537280",
  1140 => x"0c883d0d",
  1141 => x"04800b88",
  1142 => x"160c9415",
  1143 => x"08309816",
  1144 => x"0c8053ea",
  1145 => x"39725182",
  1146 => x"fb3ffec4",
  1147 => x"3974518c",
  1148 => x"e83f8c15",
  1149 => x"22708106",
  1150 => x"55537380",
  1151 => x"2effb938",
  1152 => x"d439f83d",
  1153 => x"0d7a5877",
  1154 => x"802e8199",
  1155 => x"3880cd8c",
  1156 => x"0854b814",
  1157 => x"08802e80",
  1158 => x"ed388c18",
  1159 => x"2270902b",
  1160 => x"70902c70",
  1161 => x"832a8132",
  1162 => x"81065c51",
  1163 => x"57547880",
  1164 => x"cd389018",
  1165 => x"08577680",
  1166 => x"2e80c338",
  1167 => x"77087731",
  1168 => x"77790c76",
  1169 => x"83067a58",
  1170 => x"55557385",
  1171 => x"38941808",
  1172 => x"56758819",
  1173 => x"0c807525",
  1174 => x"a5387453",
  1175 => x"76529c18",
  1176 => x"0851a418",
  1177 => x"0854732d",
  1178 => x"800b8008",
  1179 => x"2580c938",
  1180 => x"80081775",
  1181 => x"80083156",
  1182 => x"57748024",
  1183 => x"dd38800b",
  1184 => x"800c8a3d",
  1185 => x"0d047351",
  1186 => x"81da3f8c",
  1187 => x"18227090",
  1188 => x"2b70902c",
  1189 => x"70832a81",
  1190 => x"3281065c",
  1191 => x"51575478",
  1192 => x"dd38ff8e",
  1193 => x"39a48252",
  1194 => x"80cd8c08",
  1195 => x"5189f13f",
  1196 => x"8008800c",
  1197 => x"8a3d0d04",
  1198 => x"8c182280",
  1199 => x"c0075473",
  1200 => x"8c1923ff",
  1201 => x"0b800c8a",
  1202 => x"3d0d0480",
  1203 => x"3d0d7251",
  1204 => x"80710c80",
  1205 => x"0b84120c",
  1206 => x"800b8812",
  1207 => x"0c028e05",
  1208 => x"228c1223",
  1209 => x"02920522",
  1210 => x"8e122380",
  1211 => x"0b90120c",
  1212 => x"800b9412",
  1213 => x"0c800b98",
  1214 => x"120c709c",
  1215 => x"120c80c0",
  1216 => x"970ba012",
  1217 => x"0c80c0e3",
  1218 => x"0ba4120c",
  1219 => x"80c1df0b",
  1220 => x"a8120c80",
  1221 => x"c2b00bac",
  1222 => x"120c823d",
  1223 => x"0d04fa3d",
  1224 => x"0d797080",
  1225 => x"dc298c11",
  1226 => x"547a5356",
  1227 => x"578cad3f",
  1228 => x"80088008",
  1229 => x"55568008",
  1230 => x"802ea238",
  1231 => x"80088c05",
  1232 => x"54800b80",
  1233 => x"080c7680",
  1234 => x"0884050c",
  1235 => x"73800888",
  1236 => x"050c7453",
  1237 => x"80527351",
  1238 => x"97f83f75",
  1239 => x"5473800c",
  1240 => x"883d0d04",
  1241 => x"fc3d0d76",
  1242 => x"a8f70bbc",
  1243 => x"120c5581",
  1244 => x"0bb8160c",
  1245 => x"800b84dc",
  1246 => x"160c830b",
  1247 => x"84e0160c",
  1248 => x"84e81584",
  1249 => x"e4160c74",
  1250 => x"54805384",
  1251 => x"52841508",
  1252 => x"51feb83f",
  1253 => x"74548153",
  1254 => x"89528815",
  1255 => x"0851feab",
  1256 => x"3f745482",
  1257 => x"538a528c",
  1258 => x"150851fe",
  1259 => x"9e3f863d",
  1260 => x"0d04f93d",
  1261 => x"0d7980cd",
  1262 => x"8c085457",
  1263 => x"b8130880",
  1264 => x"2e80c838",
  1265 => x"84dc1356",
  1266 => x"88160884",
  1267 => x"1708ff05",
  1268 => x"55558074",
  1269 => x"249f388c",
  1270 => x"15227090",
  1271 => x"2b70902c",
  1272 => x"51545872",
  1273 => x"802e80ca",
  1274 => x"3880dc15",
  1275 => x"ff155555",
  1276 => x"738025e3",
  1277 => x"38750853",
  1278 => x"72802e9f",
  1279 => x"38725688",
  1280 => x"16088417",
  1281 => x"08ff0555",
  1282 => x"55c83972",
  1283 => x"51fed53f",
  1284 => x"80cd8c08",
  1285 => x"84dc0556",
  1286 => x"ffae3984",
  1287 => x"527651fd",
  1288 => x"fd3f8008",
  1289 => x"760c8008",
  1290 => x"802e80c0",
  1291 => x"38800856",
  1292 => x"ce39810b",
  1293 => x"8c162372",
  1294 => x"750c7288",
  1295 => x"160c7284",
  1296 => x"160c7290",
  1297 => x"160c7294",
  1298 => x"160c7298",
  1299 => x"160cff0b",
  1300 => x"8e162372",
  1301 => x"b0160c72",
  1302 => x"b4160c72",
  1303 => x"80c4160c",
  1304 => x"7280c816",
  1305 => x"0c74800c",
  1306 => x"893d0d04",
  1307 => x"8c770c80",
  1308 => x"0b800c89",
  1309 => x"3d0d04ff",
  1310 => x"3d0da482",
  1311 => x"52735186",
  1312 => x"9f3f833d",
  1313 => x"0d04803d",
  1314 => x"0d80cd8c",
  1315 => x"0851e83f",
  1316 => x"823d0d04",
  1317 => x"fb3d0d77",
  1318 => x"70525696",
  1319 => x"c43f80d4",
  1320 => x"c80b8805",
  1321 => x"08841108",
  1322 => x"fc06707b",
  1323 => x"319fef05",
  1324 => x"e08006e0",
  1325 => x"80055656",
  1326 => x"53a08074",
  1327 => x"24943880",
  1328 => x"52755196",
  1329 => x"9e3f80d4",
  1330 => x"d0081553",
  1331 => x"7280082e",
  1332 => x"8f387551",
  1333 => x"968c3f80",
  1334 => x"5372800c",
  1335 => x"873d0d04",
  1336 => x"73305275",
  1337 => x"5195fc3f",
  1338 => x"8008ff2e",
  1339 => x"a83880d4",
  1340 => x"c80b8805",
  1341 => x"08757531",
  1342 => x"81078412",
  1343 => x"0c5380d4",
  1344 => x"8c087431",
  1345 => x"80d48c0c",
  1346 => x"755195d6",
  1347 => x"3f810b80",
  1348 => x"0c873d0d",
  1349 => x"04805275",
  1350 => x"5195c83f",
  1351 => x"80d4c80b",
  1352 => x"88050880",
  1353 => x"08713156",
  1354 => x"538f7525",
  1355 => x"ffa43880",
  1356 => x"0880d4bc",
  1357 => x"083180d4",
  1358 => x"8c0c7481",
  1359 => x"0784140c",
  1360 => x"7551959e",
  1361 => x"3f8053ff",
  1362 => x"9039f63d",
  1363 => x"0d7c7e54",
  1364 => x"5b72802e",
  1365 => x"8283387a",
  1366 => x"5195863f",
  1367 => x"f8138411",
  1368 => x"0870fe06",
  1369 => x"70138411",
  1370 => x"08fc065d",
  1371 => x"58595458",
  1372 => x"80d4d008",
  1373 => x"752e82de",
  1374 => x"38788416",
  1375 => x"0c807381",
  1376 => x"06545a72",
  1377 => x"7a2e81d5",
  1378 => x"38781584",
  1379 => x"11088106",
  1380 => x"515372a0",
  1381 => x"38781757",
  1382 => x"7981e638",
  1383 => x"88150853",
  1384 => x"7280d4d0",
  1385 => x"2e82f938",
  1386 => x"8c150870",
  1387 => x"8c150c73",
  1388 => x"88120c56",
  1389 => x"76810784",
  1390 => x"190c7618",
  1391 => x"77710c53",
  1392 => x"79819138",
  1393 => x"83ff7727",
  1394 => x"81c83876",
  1395 => x"892a7783",
  1396 => x"2a565372",
  1397 => x"802ebf38",
  1398 => x"76862ab8",
  1399 => x"05558473",
  1400 => x"27b43880",
  1401 => x"db135594",
  1402 => x"7327ab38",
  1403 => x"768c2a80",
  1404 => x"ee055580",
  1405 => x"d473279e",
  1406 => x"38768f2a",
  1407 => x"80f70555",
  1408 => x"82d47327",
  1409 => x"91387692",
  1410 => x"2a80fc05",
  1411 => x"558ad473",
  1412 => x"27843880",
  1413 => x"fe557410",
  1414 => x"101080d4",
  1415 => x"c8058811",
  1416 => x"08555673",
  1417 => x"762e82b3",
  1418 => x"38841408",
  1419 => x"fc065376",
  1420 => x"73278d38",
  1421 => x"88140854",
  1422 => x"73762e09",
  1423 => x"8106ea38",
  1424 => x"8c140870",
  1425 => x"8c1a0c74",
  1426 => x"881a0c78",
  1427 => x"88120c56",
  1428 => x"778c150c",
  1429 => x"7a51938a",
  1430 => x"3f8c3d0d",
  1431 => x"04770878",
  1432 => x"71315977",
  1433 => x"05881908",
  1434 => x"54577280",
  1435 => x"d4d02e80",
  1436 => x"e0388c18",
  1437 => x"08708c15",
  1438 => x"0c738812",
  1439 => x"0c56fe89",
  1440 => x"39881508",
  1441 => x"8c160870",
  1442 => x"8c130c57",
  1443 => x"88170cfe",
  1444 => x"a3397683",
  1445 => x"2a705455",
  1446 => x"80752481",
  1447 => x"98387282",
  1448 => x"2c81712b",
  1449 => x"80d4cc08",
  1450 => x"0780d4c8",
  1451 => x"0b84050c",
  1452 => x"53741010",
  1453 => x"1080d4c8",
  1454 => x"05881108",
  1455 => x"5556758c",
  1456 => x"190c7388",
  1457 => x"190c7788",
  1458 => x"170c778c",
  1459 => x"150cff84",
  1460 => x"39815afd",
  1461 => x"b4397817",
  1462 => x"73810654",
  1463 => x"57729838",
  1464 => x"77087871",
  1465 => x"31597705",
  1466 => x"8c190888",
  1467 => x"1a08718c",
  1468 => x"120c8812",
  1469 => x"0c575776",
  1470 => x"81078419",
  1471 => x"0c7780d4",
  1472 => x"c80b8805",
  1473 => x"0c80d4c4",
  1474 => x"087726fe",
  1475 => x"c73880d4",
  1476 => x"c008527a",
  1477 => x"51fafd3f",
  1478 => x"7a5191c6",
  1479 => x"3ffeba39",
  1480 => x"81788c15",
  1481 => x"0c788815",
  1482 => x"0c738c1a",
  1483 => x"0c73881a",
  1484 => x"0c5afd80",
  1485 => x"39831570",
  1486 => x"822c8171",
  1487 => x"2b80d4cc",
  1488 => x"080780d4",
  1489 => x"c80b8405",
  1490 => x"0c515374",
  1491 => x"10101080",
  1492 => x"d4c80588",
  1493 => x"11085556",
  1494 => x"fee43974",
  1495 => x"53807524",
  1496 => x"a7387282",
  1497 => x"2c81712b",
  1498 => x"80d4cc08",
  1499 => x"0780d4c8",
  1500 => x"0b84050c",
  1501 => x"53758c19",
  1502 => x"0c738819",
  1503 => x"0c778817",
  1504 => x"0c778c15",
  1505 => x"0cfdcd39",
  1506 => x"83157082",
  1507 => x"2c81712b",
  1508 => x"80d4cc08",
  1509 => x"0780d4c8",
  1510 => x"0b84050c",
  1511 => x"5153d639",
  1512 => x"f93d0d79",
  1513 => x"7b585380",
  1514 => x"0b80cd8c",
  1515 => x"08535672",
  1516 => x"722e80c0",
  1517 => x"3884dc13",
  1518 => x"5574762e",
  1519 => x"b7388815",
  1520 => x"08841608",
  1521 => x"ff055454",
  1522 => x"8073249d",
  1523 => x"388c1422",
  1524 => x"70902b70",
  1525 => x"902c5153",
  1526 => x"587180d8",
  1527 => x"3880dc14",
  1528 => x"ff145454",
  1529 => x"728025e5",
  1530 => x"38740855",
  1531 => x"74d03880",
  1532 => x"cd8c0852",
  1533 => x"84dc1255",
  1534 => x"74802eb1",
  1535 => x"38881508",
  1536 => x"841608ff",
  1537 => x"05545480",
  1538 => x"73249c38",
  1539 => x"8c142270",
  1540 => x"902b7090",
  1541 => x"2c515358",
  1542 => x"71ad3880",
  1543 => x"dc14ff14",
  1544 => x"54547280",
  1545 => x"25e63874",
  1546 => x"085574d1",
  1547 => x"3875800c",
  1548 => x"893d0d04",
  1549 => x"7351762d",
  1550 => x"75800807",
  1551 => x"80dc15ff",
  1552 => x"15555556",
  1553 => x"ff9e3973",
  1554 => x"51762d75",
  1555 => x"80080780",
  1556 => x"dc15ff15",
  1557 => x"555556ca",
  1558 => x"39ea3d0d",
  1559 => x"688c1122",
  1560 => x"700a100a",
  1561 => x"81065758",
  1562 => x"567480e4",
  1563 => x"388e1622",
  1564 => x"70902b70",
  1565 => x"902c5155",
  1566 => x"58807424",
  1567 => x"b138983d",
  1568 => x"c4055373",
  1569 => x"5280cd8c",
  1570 => x"085192ac",
  1571 => x"3f800b80",
  1572 => x"08249738",
  1573 => x"7983e080",
  1574 => x"06547380",
  1575 => x"c0802e81",
  1576 => x"8f387382",
  1577 => x"80802e81",
  1578 => x"91388c16",
  1579 => x"22577690",
  1580 => x"80075473",
  1581 => x"8c172388",
  1582 => x"805280cd",
  1583 => x"8c085181",
  1584 => x"9b3f8008",
  1585 => x"9d388c16",
  1586 => x"22820754",
  1587 => x"738c1723",
  1588 => x"80c31670",
  1589 => x"770c9017",
  1590 => x"0c810b94",
  1591 => x"170c983d",
  1592 => x"0d0480cd",
  1593 => x"8c08a8f7",
  1594 => x"0bbc120c",
  1595 => x"548c1622",
  1596 => x"81800754",
  1597 => x"738c1723",
  1598 => x"8008760c",
  1599 => x"80089017",
  1600 => x"0c88800b",
  1601 => x"94170c74",
  1602 => x"802ed338",
  1603 => x"8e162270",
  1604 => x"902b7090",
  1605 => x"2c535558",
  1606 => x"98a23f80",
  1607 => x"08802eff",
  1608 => x"bd388c16",
  1609 => x"22810754",
  1610 => x"738c1723",
  1611 => x"983d0d04",
  1612 => x"810b8c17",
  1613 => x"225855fe",
  1614 => x"f539a816",
  1615 => x"0880c1df",
  1616 => x"2e098106",
  1617 => x"fee4388c",
  1618 => x"16228880",
  1619 => x"0754738c",
  1620 => x"17238880",
  1621 => x"0b80cc17",
  1622 => x"0cfedc39",
  1623 => x"f33d0d7f",
  1624 => x"618b1170",
  1625 => x"f8065c55",
  1626 => x"555e7296",
  1627 => x"26833890",
  1628 => x"59807924",
  1629 => x"747a2607",
  1630 => x"53805472",
  1631 => x"742e0981",
  1632 => x"0680cb38",
  1633 => x"7d518cd9",
  1634 => x"3f7883f7",
  1635 => x"2680c638",
  1636 => x"78832a70",
  1637 => x"10101080",
  1638 => x"d4c8058c",
  1639 => x"11085959",
  1640 => x"5a76782e",
  1641 => x"83b03884",
  1642 => x"1708fc06",
  1643 => x"568c1708",
  1644 => x"88180871",
  1645 => x"8c120c88",
  1646 => x"120c5875",
  1647 => x"17841108",
  1648 => x"81078412",
  1649 => x"0c537d51",
  1650 => x"8c983f88",
  1651 => x"17547380",
  1652 => x"0c8f3d0d",
  1653 => x"0478892a",
  1654 => x"79832a5b",
  1655 => x"5372802e",
  1656 => x"bf387886",
  1657 => x"2ab8055a",
  1658 => x"847327b4",
  1659 => x"3880db13",
  1660 => x"5a947327",
  1661 => x"ab38788c",
  1662 => x"2a80ee05",
  1663 => x"5a80d473",
  1664 => x"279e3878",
  1665 => x"8f2a80f7",
  1666 => x"055a82d4",
  1667 => x"73279138",
  1668 => x"78922a80",
  1669 => x"fc055a8a",
  1670 => x"d4732784",
  1671 => x"3880fe5a",
  1672 => x"79101010",
  1673 => x"80d4c805",
  1674 => x"8c110858",
  1675 => x"5576752e",
  1676 => x"a3388417",
  1677 => x"08fc0670",
  1678 => x"7a315556",
  1679 => x"738f2488",
  1680 => x"d5387380",
  1681 => x"25fee638",
  1682 => x"8c170857",
  1683 => x"76752e09",
  1684 => x"8106df38",
  1685 => x"811a5a80",
  1686 => x"d4d80857",
  1687 => x"7680d4d0",
  1688 => x"2e82c038",
  1689 => x"841708fc",
  1690 => x"06707a31",
  1691 => x"5556738f",
  1692 => x"2481f938",
  1693 => x"80d4d00b",
  1694 => x"80d4dc0c",
  1695 => x"80d4d00b",
  1696 => x"80d4d80c",
  1697 => x"738025fe",
  1698 => x"b23883ff",
  1699 => x"762783df",
  1700 => x"3875892a",
  1701 => x"76832a55",
  1702 => x"5372802e",
  1703 => x"bf387586",
  1704 => x"2ab80554",
  1705 => x"847327b4",
  1706 => x"3880db13",
  1707 => x"54947327",
  1708 => x"ab38758c",
  1709 => x"2a80ee05",
  1710 => x"5480d473",
  1711 => x"279e3875",
  1712 => x"8f2a80f7",
  1713 => x"055482d4",
  1714 => x"73279138",
  1715 => x"75922a80",
  1716 => x"fc05548a",
  1717 => x"d4732784",
  1718 => x"3880fe54",
  1719 => x"73101010",
  1720 => x"80d4c805",
  1721 => x"88110856",
  1722 => x"5874782e",
  1723 => x"86cf3884",
  1724 => x"1508fc06",
  1725 => x"53757327",
  1726 => x"8d388815",
  1727 => x"08557478",
  1728 => x"2e098106",
  1729 => x"ea388c15",
  1730 => x"0880d4c8",
  1731 => x"0b840508",
  1732 => x"718c1a0c",
  1733 => x"76881a0c",
  1734 => x"7888130c",
  1735 => x"788c180c",
  1736 => x"5d587953",
  1737 => x"807a2483",
  1738 => x"e6387282",
  1739 => x"2c81712b",
  1740 => x"5c537a7c",
  1741 => x"26819838",
  1742 => x"7b7b0653",
  1743 => x"7282f138",
  1744 => x"79fc0684",
  1745 => x"055a7a10",
  1746 => x"707d0654",
  1747 => x"5b7282e0",
  1748 => x"38841a5a",
  1749 => x"f1398817",
  1750 => x"8c110858",
  1751 => x"5876782e",
  1752 => x"098106fc",
  1753 => x"c238821a",
  1754 => x"5afdec39",
  1755 => x"78177981",
  1756 => x"0784190c",
  1757 => x"7080d4dc",
  1758 => x"0c7080d4",
  1759 => x"d80c80d4",
  1760 => x"d00b8c12",
  1761 => x"0c8c1108",
  1762 => x"88120c74",
  1763 => x"81078412",
  1764 => x"0c741175",
  1765 => x"710c5153",
  1766 => x"7d5188c6",
  1767 => x"3f881754",
  1768 => x"fcac3980",
  1769 => x"d4c80b84",
  1770 => x"05087a54",
  1771 => x"5c798025",
  1772 => x"fef83882",
  1773 => x"da397a09",
  1774 => x"7c067080",
  1775 => x"d4c80b84",
  1776 => x"050c5c7a",
  1777 => x"105b7a7c",
  1778 => x"2685387a",
  1779 => x"85b83880",
  1780 => x"d4c80b88",
  1781 => x"05087084",
  1782 => x"1208fc06",
  1783 => x"707c317c",
  1784 => x"72268f72",
  1785 => x"25075757",
  1786 => x"5c5d5572",
  1787 => x"802e80db",
  1788 => x"38797a16",
  1789 => x"80d4c008",
  1790 => x"1b90115a",
  1791 => x"55575b80",
  1792 => x"d4bc08ff",
  1793 => x"2e8838a0",
  1794 => x"8f13e080",
  1795 => x"06577652",
  1796 => x"7d5187cf",
  1797 => x"3f800854",
  1798 => x"8008ff2e",
  1799 => x"90388008",
  1800 => x"76278299",
  1801 => x"387480d4",
  1802 => x"c82e8291",
  1803 => x"3880d4c8",
  1804 => x"0b880508",
  1805 => x"55841508",
  1806 => x"fc06707a",
  1807 => x"317a7226",
  1808 => x"8f722507",
  1809 => x"52555372",
  1810 => x"83e63874",
  1811 => x"79810784",
  1812 => x"170c7916",
  1813 => x"7080d4c8",
  1814 => x"0b88050c",
  1815 => x"75810784",
  1816 => x"120c547e",
  1817 => x"525786fa",
  1818 => x"3f881754",
  1819 => x"fae03975",
  1820 => x"832a7054",
  1821 => x"54807424",
  1822 => x"819b3872",
  1823 => x"822c8171",
  1824 => x"2b80d4cc",
  1825 => x"08077080",
  1826 => x"d4c80b84",
  1827 => x"050c7510",
  1828 => x"101080d4",
  1829 => x"c8058811",
  1830 => x"08585a5d",
  1831 => x"53778c18",
  1832 => x"0c748818",
  1833 => x"0c768819",
  1834 => x"0c768c16",
  1835 => x"0cfcf339",
  1836 => x"797a1010",
  1837 => x"1080d4c8",
  1838 => x"05705759",
  1839 => x"5d8c1508",
  1840 => x"5776752e",
  1841 => x"a3388417",
  1842 => x"08fc0670",
  1843 => x"7a315556",
  1844 => x"738f2483",
  1845 => x"ca387380",
  1846 => x"25848138",
  1847 => x"8c170857",
  1848 => x"76752e09",
  1849 => x"8106df38",
  1850 => x"8815811b",
  1851 => x"70830655",
  1852 => x"5b5572c9",
  1853 => x"387c8306",
  1854 => x"5372802e",
  1855 => x"fdb838ff",
  1856 => x"1df81959",
  1857 => x"5d881808",
  1858 => x"782eea38",
  1859 => x"fdb53983",
  1860 => x"1a53fc96",
  1861 => x"39831470",
  1862 => x"822c8171",
  1863 => x"2b80d4cc",
  1864 => x"08077080",
  1865 => x"d4c80b84",
  1866 => x"050c7610",
  1867 => x"101080d4",
  1868 => x"c8058811",
  1869 => x"08595b5e",
  1870 => x"5153fee1",
  1871 => x"3980d48c",
  1872 => x"08175880",
  1873 => x"08762e81",
  1874 => x"8d3880d4",
  1875 => x"bc08ff2e",
  1876 => x"83ec3873",
  1877 => x"76311880",
  1878 => x"d48c0c73",
  1879 => x"87067057",
  1880 => x"5372802e",
  1881 => x"88388873",
  1882 => x"31701555",
  1883 => x"5676149f",
  1884 => x"ff06a080",
  1885 => x"71311770",
  1886 => x"547f5357",
  1887 => x"5384e43f",
  1888 => x"80085380",
  1889 => x"08ff2e81",
  1890 => x"a03880d4",
  1891 => x"8c081670",
  1892 => x"80d48c0c",
  1893 => x"747580d4",
  1894 => x"c80b8805",
  1895 => x"0c747631",
  1896 => x"18708107",
  1897 => x"51555658",
  1898 => x"7b80d4c8",
  1899 => x"2e839c38",
  1900 => x"798f2682",
  1901 => x"cb38810b",
  1902 => x"84150c84",
  1903 => x"1508fc06",
  1904 => x"707a317a",
  1905 => x"72268f72",
  1906 => x"25075255",
  1907 => x"5372802e",
  1908 => x"fcf93880",
  1909 => x"db398008",
  1910 => x"9fff0653",
  1911 => x"72feeb38",
  1912 => x"7780d48c",
  1913 => x"0c80d4c8",
  1914 => x"0b880508",
  1915 => x"7b188107",
  1916 => x"84120c55",
  1917 => x"80d4b808",
  1918 => x"78278638",
  1919 => x"7780d4b8",
  1920 => x"0c80d4b4",
  1921 => x"087827fc",
  1922 => x"ac387780",
  1923 => x"d4b40c84",
  1924 => x"1508fc06",
  1925 => x"707a317a",
  1926 => x"72268f72",
  1927 => x"25075255",
  1928 => x"5372802e",
  1929 => x"fca53888",
  1930 => x"39807454",
  1931 => x"56fedb39",
  1932 => x"7d5183ae",
  1933 => x"3f800b80",
  1934 => x"0c8f3d0d",
  1935 => x"04735380",
  1936 => x"7424a938",
  1937 => x"72822c81",
  1938 => x"712b80d4",
  1939 => x"cc080770",
  1940 => x"80d4c80b",
  1941 => x"84050c5d",
  1942 => x"53778c18",
  1943 => x"0c748818",
  1944 => x"0c768819",
  1945 => x"0c768c16",
  1946 => x"0cf9b739",
  1947 => x"83147082",
  1948 => x"2c81712b",
  1949 => x"80d4cc08",
  1950 => x"077080d4",
  1951 => x"c80b8405",
  1952 => x"0c5e5153",
  1953 => x"d4397b7b",
  1954 => x"065372fc",
  1955 => x"a338841a",
  1956 => x"7b105c5a",
  1957 => x"f139ff1a",
  1958 => x"8111515a",
  1959 => x"f7b93978",
  1960 => x"17798107",
  1961 => x"84190c8c",
  1962 => x"18088819",
  1963 => x"08718c12",
  1964 => x"0c88120c",
  1965 => x"597080d4",
  1966 => x"dc0c7080",
  1967 => x"d4d80c80",
  1968 => x"d4d00b8c",
  1969 => x"120c8c11",
  1970 => x"0888120c",
  1971 => x"74810784",
  1972 => x"120c7411",
  1973 => x"75710c51",
  1974 => x"53f9bd39",
  1975 => x"75178411",
  1976 => x"08810784",
  1977 => x"120c538c",
  1978 => x"17088818",
  1979 => x"08718c12",
  1980 => x"0c88120c",
  1981 => x"587d5181",
  1982 => x"e93f8817",
  1983 => x"54f5cf39",
  1984 => x"7284150c",
  1985 => x"f41af806",
  1986 => x"70841e08",
  1987 => x"81060784",
  1988 => x"1e0c701d",
  1989 => x"545b850b",
  1990 => x"84140c85",
  1991 => x"0b88140c",
  1992 => x"8f7b27fd",
  1993 => x"cf38881c",
  1994 => x"527d51ec",
  1995 => x"9d3f80d4",
  1996 => x"c80b8805",
  1997 => x"0880d48c",
  1998 => x"085955fd",
  1999 => x"b7397780",
  2000 => x"d48c0c73",
  2001 => x"80d4bc0c",
  2002 => x"fc913972",
  2003 => x"84150cfd",
  2004 => x"a339fc3d",
  2005 => x"0d767971",
  2006 => x"028c059f",
  2007 => x"05335755",
  2008 => x"53558372",
  2009 => x"278a3874",
  2010 => x"83065170",
  2011 => x"802ea238",
  2012 => x"ff125271",
  2013 => x"ff2e9338",
  2014 => x"73737081",
  2015 => x"055534ff",
  2016 => x"125271ff",
  2017 => x"2e098106",
  2018 => x"ef387480",
  2019 => x"0c863d0d",
  2020 => x"04747488",
  2021 => x"2b750770",
  2022 => x"71902b07",
  2023 => x"5154518f",
  2024 => x"7227a538",
  2025 => x"72717084",
  2026 => x"05530c72",
  2027 => x"71708405",
  2028 => x"530c7271",
  2029 => x"70840553",
  2030 => x"0c727170",
  2031 => x"8405530c",
  2032 => x"f0125271",
  2033 => x"8f26dd38",
  2034 => x"83722790",
  2035 => x"38727170",
  2036 => x"8405530c",
  2037 => x"fc125271",
  2038 => x"8326f238",
  2039 => x"7053ff90",
  2040 => x"390404fd",
  2041 => x"3d0d800b",
  2042 => x"80dd800c",
  2043 => x"765184ee",
  2044 => x"3f800853",
  2045 => x"8008ff2e",
  2046 => x"88387280",
  2047 => x"0c853d0d",
  2048 => x"0480dd80",
  2049 => x"08547380",
  2050 => x"2ef03875",
  2051 => x"74710c52",
  2052 => x"72800c85",
  2053 => x"3d0d04f9",
  2054 => x"3d0d797c",
  2055 => x"557b548e",
  2056 => x"11227090",
  2057 => x"2b70902c",
  2058 => x"555780cd",
  2059 => x"8c085358",
  2060 => x"5683f33f",
  2061 => x"80085780",
  2062 => x"0b800824",
  2063 => x"933880d0",
  2064 => x"16088008",
  2065 => x"0580d017",
  2066 => x"0c76800c",
  2067 => x"893d0d04",
  2068 => x"8c162283",
  2069 => x"dfff0655",
  2070 => x"748c1723",
  2071 => x"76800c89",
  2072 => x"3d0d04fa",
  2073 => x"3d0d788c",
  2074 => x"11227088",
  2075 => x"2a708106",
  2076 => x"51575856",
  2077 => x"74a9388c",
  2078 => x"162283df",
  2079 => x"ff065574",
  2080 => x"8c17237a",
  2081 => x"5479538e",
  2082 => x"16227090",
  2083 => x"2b70902c",
  2084 => x"545680cd",
  2085 => x"8c085256",
  2086 => x"81b23f88",
  2087 => x"3d0d0482",
  2088 => x"5480538e",
  2089 => x"16227090",
  2090 => x"2b70902c",
  2091 => x"545680cd",
  2092 => x"8c085257",
  2093 => x"82b83f8c",
  2094 => x"162283df",
  2095 => x"ff065574",
  2096 => x"8c17237a",
  2097 => x"5479538e",
  2098 => x"16227090",
  2099 => x"2b70902c",
  2100 => x"545680cd",
  2101 => x"8c085256",
  2102 => x"80f23f88",
  2103 => x"3d0d04f9",
  2104 => x"3d0d797c",
  2105 => x"557b548e",
  2106 => x"11227090",
  2107 => x"2b70902c",
  2108 => x"555780cd",
  2109 => x"8c085358",
  2110 => x"5681f33f",
  2111 => x"80085780",
  2112 => x"08ff2e99",
  2113 => x"388c1622",
  2114 => x"a0800755",
  2115 => x"748c1723",
  2116 => x"800880d0",
  2117 => x"170c7680",
  2118 => x"0c893d0d",
  2119 => x"048c1622",
  2120 => x"83dfff06",
  2121 => x"55748c17",
  2122 => x"2376800c",
  2123 => x"893d0d04",
  2124 => x"fe3d0d74",
  2125 => x"8e112270",
  2126 => x"902b7090",
  2127 => x"2c555151",
  2128 => x"5380cd8c",
  2129 => x"0851bd3f",
  2130 => x"843d0d04",
  2131 => x"fb3d0d80",
  2132 => x"0b80dd80",
  2133 => x"0c7a5379",
  2134 => x"52785182",
  2135 => x"fc3f8008",
  2136 => x"558008ff",
  2137 => x"2e883874",
  2138 => x"800c873d",
  2139 => x"0d0480dd",
  2140 => x"80085675",
  2141 => x"802ef038",
  2142 => x"7776710c",
  2143 => x"5474800c",
  2144 => x"873d0d04",
  2145 => x"fd3d0d80",
  2146 => x"0b80dd80",
  2147 => x"0c765184",
  2148 => x"c63f8008",
  2149 => x"538008ff",
  2150 => x"2e883872",
  2151 => x"800c853d",
  2152 => x"0d0480dd",
  2153 => x"80085473",
  2154 => x"802ef038",
  2155 => x"7574710c",
  2156 => x"5272800c",
  2157 => x"853d0d04",
  2158 => x"fc3d0d80",
  2159 => x"0b80dd80",
  2160 => x"0c785277",
  2161 => x"5186ac3f",
  2162 => x"80085480",
  2163 => x"08ff2e88",
  2164 => x"3873800c",
  2165 => x"863d0d04",
  2166 => x"80dd8008",
  2167 => x"5574802e",
  2168 => x"f0387675",
  2169 => x"710c5373",
  2170 => x"800c863d",
  2171 => x"0d04fb3d",
  2172 => x"0d800b80",
  2173 => x"dd800c7a",
  2174 => x"53795278",
  2175 => x"5184893f",
  2176 => x"80085580",
  2177 => x"08ff2e88",
  2178 => x"3874800c",
  2179 => x"873d0d04",
  2180 => x"80dd8008",
  2181 => x"5675802e",
  2182 => x"f0387776",
  2183 => x"710c5474",
  2184 => x"800c873d",
  2185 => x"0d04fb3d",
  2186 => x"0d800b80",
  2187 => x"dd800c7a",
  2188 => x"53795278",
  2189 => x"5182963f",
  2190 => x"80085580",
  2191 => x"08ff2e88",
  2192 => x"3874800c",
  2193 => x"873d0d04",
  2194 => x"80dd8008",
  2195 => x"5675802e",
  2196 => x"f0387776",
  2197 => x"710c5474",
  2198 => x"800c873d",
  2199 => x"0d04fe3d",
  2200 => x"0d80dcf8",
  2201 => x"0851708a",
  2202 => x"3880dd84",
  2203 => x"7080dcf8",
  2204 => x"0c517075",
  2205 => x"125252ff",
  2206 => x"537087fb",
  2207 => x"80802688",
  2208 => x"387080dc",
  2209 => x"f80c7153",
  2210 => x"72800c84",
  2211 => x"3d0d04fd",
  2212 => x"3d0d800b",
  2213 => x"80cd8008",
  2214 => x"54547281",
  2215 => x"2e9b3873",
  2216 => x"80dcfc0c",
  2217 => x"c4803fc2",
  2218 => x"d73f80dc",
  2219 => x"d0528151",
  2220 => x"c5c63f80",
  2221 => x"085185bb",
  2222 => x"3f7280dc",
  2223 => x"fc0cc3e6",
  2224 => x"3fc2bd3f",
  2225 => x"80dcd052",
  2226 => x"8151c5ac",
  2227 => x"3f800851",
  2228 => x"85a13f00",
  2229 => x"ff3900ff",
  2230 => x"39f53d0d",
  2231 => x"7e6080dc",
  2232 => x"fc08705b",
  2233 => x"585b5b75",
  2234 => x"80c23877",
  2235 => x"7a25a138",
  2236 => x"771b7033",
  2237 => x"7081ff06",
  2238 => x"58585975",
  2239 => x"8a2e9838",
  2240 => x"7681ff06",
  2241 => x"51c2fe3f",
  2242 => x"81185879",
  2243 => x"7824e138",
  2244 => x"79800c8d",
  2245 => x"3d0d048d",
  2246 => x"51c2ea3f",
  2247 => x"78337081",
  2248 => x"ff065257",
  2249 => x"c2df3f81",
  2250 => x"1858e039",
  2251 => x"79557a54",
  2252 => x"7d538552",
  2253 => x"8d3dfc05",
  2254 => x"51c2873f",
  2255 => x"80085684",
  2256 => x"ab3f7b80",
  2257 => x"080c7580",
  2258 => x"0c8d3d0d",
  2259 => x"04f63d0d",
  2260 => x"7d7f80dc",
  2261 => x"fc08705b",
  2262 => x"585a5a75",
  2263 => x"80c13877",
  2264 => x"7925b338",
  2265 => x"c1fa3f80",
  2266 => x"0881ff06",
  2267 => x"708d3270",
  2268 => x"30709f2a",
  2269 => x"51515757",
  2270 => x"768a2e80",
  2271 => x"c3387580",
  2272 => x"2ebe3877",
  2273 => x"1a567676",
  2274 => x"347651c1",
  2275 => x"f83f8118",
  2276 => x"58787824",
  2277 => x"cf387756",
  2278 => x"75800c8c",
  2279 => x"3d0d0478",
  2280 => x"5579547c",
  2281 => x"5384528c",
  2282 => x"3dfc0551",
  2283 => x"c1943f80",
  2284 => x"085683b8",
  2285 => x"3f7a8008",
  2286 => x"0c75800c",
  2287 => x"8c3d0d04",
  2288 => x"771a568a",
  2289 => x"76348118",
  2290 => x"588d51c1",
  2291 => x"b83f8a51",
  2292 => x"c1b33f77",
  2293 => x"56c239fb",
  2294 => x"3d0d80dc",
  2295 => x"fc087056",
  2296 => x"54738838",
  2297 => x"74800c87",
  2298 => x"3d0d0477",
  2299 => x"53835287",
  2300 => x"3dfc0551",
  2301 => x"c0cc3f80",
  2302 => x"085482f0",
  2303 => x"3f758008",
  2304 => x"0c73800c",
  2305 => x"873d0d04",
  2306 => x"fa3d0d80",
  2307 => x"dcfc0880",
  2308 => x"2ea2387a",
  2309 => x"55795478",
  2310 => x"53865288",
  2311 => x"3dfc0551",
  2312 => x"c0a03f80",
  2313 => x"085682c4",
  2314 => x"3f768008",
  2315 => x"0c75800c",
  2316 => x"883d0d04",
  2317 => x"82b63f9d",
  2318 => x"0b80080c",
  2319 => x"ff0b800c",
  2320 => x"883d0d04",
  2321 => x"fb3d0d77",
  2322 => x"79565680",
  2323 => x"70545473",
  2324 => x"75259f38",
  2325 => x"74101010",
  2326 => x"f8055272",
  2327 => x"16703370",
  2328 => x"742b7607",
  2329 => x"8116f816",
  2330 => x"56565651",
  2331 => x"51747324",
  2332 => x"ea387380",
  2333 => x"0c873d0d",
  2334 => x"04fc3d0d",
  2335 => x"76785555",
  2336 => x"bc538052",
  2337 => x"7351f5ca",
  2338 => x"3f845274",
  2339 => x"51ffb53f",
  2340 => x"80087423",
  2341 => x"84528415",
  2342 => x"51ffa93f",
  2343 => x"80088215",
  2344 => x"23845288",
  2345 => x"1551ff9c",
  2346 => x"3f800884",
  2347 => x"150c8452",
  2348 => x"8c1551ff",
  2349 => x"8f3f8008",
  2350 => x"88152384",
  2351 => x"52901551",
  2352 => x"ff823f80",
  2353 => x"088a1523",
  2354 => x"84529415",
  2355 => x"51fef53f",
  2356 => x"80088c15",
  2357 => x"23845298",
  2358 => x"1551fee8",
  2359 => x"3f80088e",
  2360 => x"15238852",
  2361 => x"9c1551fe",
  2362 => x"db3f8008",
  2363 => x"90150c86",
  2364 => x"3d0d04e9",
  2365 => x"3d0d6a80",
  2366 => x"dcfc0857",
  2367 => x"57759338",
  2368 => x"80c0800b",
  2369 => x"84180c75",
  2370 => x"ac180c75",
  2371 => x"800c993d",
  2372 => x"0d04893d",
  2373 => x"70556a54",
  2374 => x"558a5299",
  2375 => x"3dffbc05",
  2376 => x"51ffbe9e",
  2377 => x"3f800877",
  2378 => x"53755256",
  2379 => x"fecb3fbc",
  2380 => x"3f778008",
  2381 => x"0c75800c",
  2382 => x"993d0d04",
  2383 => x"fc3d0d81",
  2384 => x"5480dcfc",
  2385 => x"08883873",
  2386 => x"800c863d",
  2387 => x"0d047653",
  2388 => x"97b95286",
  2389 => x"3dfc0551",
  2390 => x"ffbde73f",
  2391 => x"8008548c",
  2392 => x"3f748008",
  2393 => x"0c73800c",
  2394 => x"863d0d04",
  2395 => x"80cd8c08",
  2396 => x"800c04f7",
  2397 => x"3d0d7b80",
  2398 => x"cd8c0882",
  2399 => x"c811085a",
  2400 => x"545a7780",
  2401 => x"2e80da38",
  2402 => x"81881884",
  2403 => x"1908ff05",
  2404 => x"81712b59",
  2405 => x"55598074",
  2406 => x"2480ea38",
  2407 => x"807424b5",
  2408 => x"3873822b",
  2409 => x"78118805",
  2410 => x"56568180",
  2411 => x"19087706",
  2412 => x"5372802e",
  2413 => x"b6387816",
  2414 => x"70085353",
  2415 => x"79517408",
  2416 => x"53722dff",
  2417 => x"14fc17fc",
  2418 => x"1779812c",
  2419 => x"5a575754",
  2420 => x"738025d6",
  2421 => x"38770858",
  2422 => x"77ffad38",
  2423 => x"80cd8c08",
  2424 => x"53bc1308",
  2425 => x"a5387951",
  2426 => x"f9e93f74",
  2427 => x"0853722d",
  2428 => x"ff14fc17",
  2429 => x"fc177981",
  2430 => x"2c5a5757",
  2431 => x"54738025",
  2432 => x"ffa838d1",
  2433 => x"398057ff",
  2434 => x"93397251",
  2435 => x"bc130853",
  2436 => x"722d7951",
  2437 => x"f9bd3fff",
  2438 => x"3d0d80dc",
  2439 => x"d80bfc05",
  2440 => x"70085252",
  2441 => x"70ff2e91",
  2442 => x"38702dfc",
  2443 => x"12700852",
  2444 => x"5270ff2e",
  2445 => x"098106f1",
  2446 => x"38833d0d",
  2447 => x"0404ffbd",
  2448 => x"d23f0400",
  2449 => x"00000040",
  2450 => x"48656c6c",
  2451 => x"6f20776f",
  2452 => x"726c6421",
  2453 => x"00000000",
  2454 => x"0a000000",
  2455 => x"43000000",
  2456 => x"64756d6d",
  2457 => x"792e6578",
  2458 => x"65000000",
  2459 => x"00ffffff",
  2460 => x"ff00ffff",
  2461 => x"ffff00ff",
  2462 => x"ffffff00",
  2463 => x"00000000",
  2464 => x"00000000",
  2465 => x"00000000",
  2466 => x"00002e60",
  2467 => x"00002690",
  2468 => x"00000000",
  2469 => x"000028f8",
  2470 => x"00002954",
  2471 => x"000029b0",
  2472 => x"00000000",
  2473 => x"00000000",
  2474 => x"00000000",
  2475 => x"00000000",
  2476 => x"00000000",
  2477 => x"00000000",
  2478 => x"00000000",
  2479 => x"00000000",
  2480 => x"00000000",
  2481 => x"0000265c",
  2482 => x"00000000",
  2483 => x"00000000",
  2484 => x"00000000",
  2485 => x"00000000",
  2486 => x"00000000",
  2487 => x"00000000",
  2488 => x"00000000",
  2489 => x"00000000",
  2490 => x"00000000",
  2491 => x"00000000",
  2492 => x"00000000",
  2493 => x"00000000",
  2494 => x"00000000",
  2495 => x"00000000",
  2496 => x"00000000",
  2497 => x"00000000",
  2498 => x"00000000",
  2499 => x"00000000",
  2500 => x"00000000",
  2501 => x"00000000",
  2502 => x"00000000",
  2503 => x"00000000",
  2504 => x"00000000",
  2505 => x"00000000",
  2506 => x"00000000",
  2507 => x"00000000",
  2508 => x"00000000",
  2509 => x"00000000",
  2510 => x"00000001",
  2511 => x"330eabcd",
  2512 => x"1234e66d",
  2513 => x"deec0005",
  2514 => x"000b0000",
  2515 => x"00000000",
  2516 => x"00000000",
  2517 => x"00000000",
  2518 => x"00000000",
  2519 => x"00000000",
  2520 => x"00000000",
  2521 => x"00000000",
  2522 => x"00000000",
  2523 => x"00000000",
  2524 => x"00000000",
  2525 => x"00000000",
  2526 => x"00000000",
  2527 => x"00000000",
  2528 => x"00000000",
  2529 => x"00000000",
  2530 => x"00000000",
  2531 => x"00000000",
  2532 => x"00000000",
  2533 => x"00000000",
  2534 => x"00000000",
  2535 => x"00000000",
  2536 => x"00000000",
  2537 => x"00000000",
  2538 => x"00000000",
  2539 => x"00000000",
  2540 => x"00000000",
  2541 => x"00000000",
  2542 => x"00000000",
  2543 => x"00000000",
  2544 => x"00000000",
  2545 => x"00000000",
  2546 => x"00000000",
  2547 => x"00000000",
  2548 => x"00000000",
  2549 => x"00000000",
  2550 => x"00000000",
  2551 => x"00000000",
  2552 => x"00000000",
  2553 => x"00000000",
  2554 => x"00000000",
  2555 => x"00000000",
  2556 => x"00000000",
  2557 => x"00000000",
  2558 => x"00000000",
  2559 => x"00000000",
  2560 => x"00000000",
  2561 => x"00000000",
  2562 => x"00000000",
  2563 => x"00000000",
  2564 => x"00000000",
  2565 => x"00000000",
  2566 => x"00000000",
  2567 => x"00000000",
  2568 => x"00000000",
  2569 => x"00000000",
  2570 => x"00000000",
  2571 => x"00000000",
  2572 => x"00000000",
  2573 => x"00000000",
  2574 => x"00000000",
  2575 => x"00000000",
  2576 => x"00000000",
  2577 => x"00000000",
  2578 => x"00000000",
  2579 => x"00000000",
  2580 => x"00000000",
  2581 => x"00000000",
  2582 => x"00000000",
  2583 => x"00000000",
  2584 => x"00000000",
  2585 => x"00000000",
  2586 => x"00000000",
  2587 => x"00000000",
  2588 => x"00000000",
  2589 => x"00000000",
  2590 => x"00000000",
  2591 => x"00000000",
  2592 => x"00000000",
  2593 => x"00000000",
  2594 => x"00000000",
  2595 => x"00000000",
  2596 => x"00000000",
  2597 => x"00000000",
  2598 => x"00000000",
  2599 => x"00000000",
  2600 => x"00000000",
  2601 => x"00000000",
  2602 => x"00000000",
  2603 => x"00000000",
  2604 => x"00000000",
  2605 => x"00000000",
  2606 => x"00000000",
  2607 => x"00000000",
  2608 => x"00000000",
  2609 => x"00000000",
  2610 => x"00000000",
  2611 => x"00000000",
  2612 => x"00000000",
  2613 => x"00000000",
  2614 => x"00000000",
  2615 => x"00000000",
  2616 => x"00000000",
  2617 => x"00000000",
  2618 => x"00000000",
  2619 => x"00000000",
  2620 => x"00000000",
  2621 => x"00000000",
  2622 => x"00000000",
  2623 => x"00000000",
  2624 => x"00000000",
  2625 => x"00000000",
  2626 => x"00000000",
  2627 => x"00000000",
  2628 => x"00000000",
  2629 => x"00000000",
  2630 => x"00000000",
  2631 => x"00000000",
  2632 => x"00000000",
  2633 => x"00000000",
  2634 => x"00000000",
  2635 => x"00000000",
  2636 => x"00000000",
  2637 => x"00000000",
  2638 => x"00000000",
  2639 => x"00000000",
  2640 => x"00000000",
  2641 => x"00000000",
  2642 => x"00000000",
  2643 => x"00000000",
  2644 => x"00000000",
  2645 => x"00000000",
  2646 => x"00000000",
  2647 => x"00000000",
  2648 => x"00000000",
  2649 => x"00000000",
  2650 => x"00000000",
  2651 => x"00000000",
  2652 => x"00000000",
  2653 => x"00000000",
  2654 => x"00000000",
  2655 => x"00000000",
  2656 => x"00000000",
  2657 => x"00000000",
  2658 => x"00000000",
  2659 => x"00000000",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000000",
  2683 => x"00000000",
  2684 => x"00000000",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"ffffffff",
  2704 => x"00000000",
  2705 => x"00020000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00002a48",
  2709 => x"00002a48",
  2710 => x"00002a50",
  2711 => x"00002a50",
  2712 => x"00002a58",
  2713 => x"00002a58",
  2714 => x"00002a60",
  2715 => x"00002a60",
  2716 => x"00002a68",
  2717 => x"00002a68",
  2718 => x"00002a70",
  2719 => x"00002a70",
  2720 => x"00002a78",
  2721 => x"00002a78",
  2722 => x"00002a80",
  2723 => x"00002a80",
  2724 => x"00002a88",
  2725 => x"00002a88",
  2726 => x"00002a90",
  2727 => x"00002a90",
  2728 => x"00002a98",
  2729 => x"00002a98",
  2730 => x"00002aa0",
  2731 => x"00002aa0",
  2732 => x"00002aa8",
  2733 => x"00002aa8",
  2734 => x"00002ab0",
  2735 => x"00002ab0",
  2736 => x"00002ab8",
  2737 => x"00002ab8",
  2738 => x"00002ac0",
  2739 => x"00002ac0",
  2740 => x"00002ac8",
  2741 => x"00002ac8",
  2742 => x"00002ad0",
  2743 => x"00002ad0",
  2744 => x"00002ad8",
  2745 => x"00002ad8",
  2746 => x"00002ae0",
  2747 => x"00002ae0",
  2748 => x"00002ae8",
  2749 => x"00002ae8",
  2750 => x"00002af0",
  2751 => x"00002af0",
  2752 => x"00002af8",
  2753 => x"00002af8",
  2754 => x"00002b00",
  2755 => x"00002b00",
  2756 => x"00002b08",
  2757 => x"00002b08",
  2758 => x"00002b10",
  2759 => x"00002b10",
  2760 => x"00002b18",
  2761 => x"00002b18",
  2762 => x"00002b20",
  2763 => x"00002b20",
  2764 => x"00002b28",
  2765 => x"00002b28",
  2766 => x"00002b30",
  2767 => x"00002b30",
  2768 => x"00002b38",
  2769 => x"00002b38",
  2770 => x"00002b40",
  2771 => x"00002b40",
  2772 => x"00002b48",
  2773 => x"00002b48",
  2774 => x"00002b50",
  2775 => x"00002b50",
  2776 => x"00002b58",
  2777 => x"00002b58",
  2778 => x"00002b60",
  2779 => x"00002b60",
  2780 => x"00002b68",
  2781 => x"00002b68",
  2782 => x"00002b70",
  2783 => x"00002b70",
  2784 => x"00002b78",
  2785 => x"00002b78",
  2786 => x"00002b80",
  2787 => x"00002b80",
  2788 => x"00002b88",
  2789 => x"00002b88",
  2790 => x"00002b90",
  2791 => x"00002b90",
  2792 => x"00002b98",
  2793 => x"00002b98",
  2794 => x"00002ba0",
  2795 => x"00002ba0",
  2796 => x"00002ba8",
  2797 => x"00002ba8",
  2798 => x"00002bb0",
  2799 => x"00002bb0",
  2800 => x"00002bb8",
  2801 => x"00002bb8",
  2802 => x"00002bc0",
  2803 => x"00002bc0",
  2804 => x"00002bc8",
  2805 => x"00002bc8",
  2806 => x"00002bd0",
  2807 => x"00002bd0",
  2808 => x"00002bd8",
  2809 => x"00002bd8",
  2810 => x"00002be0",
  2811 => x"00002be0",
  2812 => x"00002be8",
  2813 => x"00002be8",
  2814 => x"00002bf0",
  2815 => x"00002bf0",
  2816 => x"00002bf8",
  2817 => x"00002bf8",
  2818 => x"00002c00",
  2819 => x"00002c00",
  2820 => x"00002c08",
  2821 => x"00002c08",
  2822 => x"00002c10",
  2823 => x"00002c10",
  2824 => x"00002c18",
  2825 => x"00002c18",
  2826 => x"00002c20",
  2827 => x"00002c20",
  2828 => x"00002c28",
  2829 => x"00002c28",
  2830 => x"00002c30",
  2831 => x"00002c30",
  2832 => x"00002c38",
  2833 => x"00002c38",
  2834 => x"00002c40",
  2835 => x"00002c40",
  2836 => x"00002c48",
  2837 => x"00002c48",
  2838 => x"00002c50",
  2839 => x"00002c50",
  2840 => x"00002c58",
  2841 => x"00002c58",
  2842 => x"00002c60",
  2843 => x"00002c60",
  2844 => x"00002c68",
  2845 => x"00002c68",
  2846 => x"00002c70",
  2847 => x"00002c70",
  2848 => x"00002c78",
  2849 => x"00002c78",
  2850 => x"00002c80",
  2851 => x"00002c80",
  2852 => x"00002c88",
  2853 => x"00002c88",
  2854 => x"00002c90",
  2855 => x"00002c90",
  2856 => x"00002c98",
  2857 => x"00002c98",
  2858 => x"00002ca0",
  2859 => x"00002ca0",
  2860 => x"00002ca8",
  2861 => x"00002ca8",
  2862 => x"00002cb0",
  2863 => x"00002cb0",
  2864 => x"00002cb8",
  2865 => x"00002cb8",
  2866 => x"00002cc0",
  2867 => x"00002cc0",
  2868 => x"00002cc8",
  2869 => x"00002cc8",
  2870 => x"00002cd0",
  2871 => x"00002cd0",
  2872 => x"00002cd8",
  2873 => x"00002cd8",
  2874 => x"00002ce0",
  2875 => x"00002ce0",
  2876 => x"00002ce8",
  2877 => x"00002ce8",
  2878 => x"00002cf0",
  2879 => x"00002cf0",
  2880 => x"00002cf8",
  2881 => x"00002cf8",
  2882 => x"00002d00",
  2883 => x"00002d00",
  2884 => x"00002d08",
  2885 => x"00002d08",
  2886 => x"00002d10",
  2887 => x"00002d10",
  2888 => x"00002d18",
  2889 => x"00002d18",
  2890 => x"00002d20",
  2891 => x"00002d20",
  2892 => x"00002d28",
  2893 => x"00002d28",
  2894 => x"00002d30",
  2895 => x"00002d30",
  2896 => x"00002d38",
  2897 => x"00002d38",
  2898 => x"00002d40",
  2899 => x"00002d40",
  2900 => x"00002d48",
  2901 => x"00002d48",
  2902 => x"00002d50",
  2903 => x"00002d50",
  2904 => x"00002d58",
  2905 => x"00002d58",
  2906 => x"00002d60",
  2907 => x"00002d60",
  2908 => x"00002d68",
  2909 => x"00002d68",
  2910 => x"00002d70",
  2911 => x"00002d70",
  2912 => x"00002d78",
  2913 => x"00002d78",
  2914 => x"00002d80",
  2915 => x"00002d80",
  2916 => x"00002d88",
  2917 => x"00002d88",
  2918 => x"00002d90",
  2919 => x"00002d90",
  2920 => x"00002d98",
  2921 => x"00002d98",
  2922 => x"00002da0",
  2923 => x"00002da0",
  2924 => x"00002da8",
  2925 => x"00002da8",
  2926 => x"00002db0",
  2927 => x"00002db0",
  2928 => x"00002db8",
  2929 => x"00002db8",
  2930 => x"00002dc0",
  2931 => x"00002dc0",
  2932 => x"00002dc8",
  2933 => x"00002dc8",
  2934 => x"00002dd0",
  2935 => x"00002dd0",
  2936 => x"00002dd8",
  2937 => x"00002dd8",
  2938 => x"00002de0",
  2939 => x"00002de0",
  2940 => x"00002de8",
  2941 => x"00002de8",
  2942 => x"00002df0",
  2943 => x"00002df0",
  2944 => x"00002df8",
  2945 => x"00002df8",
  2946 => x"00002e00",
  2947 => x"00002e00",
  2948 => x"00002e08",
  2949 => x"00002e08",
  2950 => x"00002e10",
  2951 => x"00002e10",
  2952 => x"00002e18",
  2953 => x"00002e18",
  2954 => x"00002e20",
  2955 => x"00002e20",
  2956 => x"00002e28",
  2957 => x"00002e28",
  2958 => x"00002e30",
  2959 => x"00002e30",
  2960 => x"00002e38",
  2961 => x"00002e38",
  2962 => x"00002e40",
  2963 => x"00002e40",
  2964 => x"00002660",
  2965 => x"ffffffff",
  2966 => x"00000000",
  2967 => x"ffffffff",
  2968 => x"00000000",
  2969 => x"00000000",

others => x"00000000"
);
begin
   do_port_a:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         if (a_we_i='1') and (b_we_i='1') and (a_addr_i=b_addr_i) and (a_write_i/=b_write_i) then
            report "DualPortRAM write collision" severity failure;
         end if;
         iaddr:=to_integer(a_addr_i);
         if a_we_i='1' then
            ram(iaddr):=a_write_i;
            a_read_o <= a_write_i;
         else
            a_read_o <= ram(iaddr);
         end if;
      end if;
   end process do_port_a;

   do_port_b:
   process (clk_i)
      variable iaddr : integer;
   begin
      if rising_edge(clk_i) then
         iaddr:=to_integer(b_addr_i);
         if b_we_i='1' then
            ram(iaddr):=b_write_i;
            b_read_o <= b_write_i;
         else
            b_read_o <= ram(iaddr);
         end if;
      end if;
   end process do_port_b;
end architecture DualPort_Arch; -- Entity: DualPortRAM
