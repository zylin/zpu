-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80e6840c",
     3 => x"3a0b0b80",
     4 => x"d5a20400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80d5eb2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80e5",
   162 => x"f0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80d0",
   171 => x"8d2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80d1",
   179 => x"bf2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80e6800c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"cf8c3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80e68008",
   281 => x"802ea438",
   282 => x"80e68408",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80ed",
   286 => x"c00c82a0",
   287 => x"800b80ed",
   288 => x"c40c8290",
   289 => x"800b80ed",
   290 => x"c80c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"edc00cf8",
   294 => x"80808280",
   295 => x"0b80edc4",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"edc80c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80edc00c",
   302 => x"80c0a880",
   303 => x"940b80ed",
   304 => x"c40c0b0b",
   305 => x"80d7c00b",
   306 => x"80edc80c",
   307 => x"04ff3d0d",
   308 => x"80edcc33",
   309 => x"5170a738",
   310 => x"80e68c08",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"e68c0c70",
   315 => x"2d80e68c",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80ed",
   319 => x"cc34833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80edbc08",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"edbc510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404fb3d",
   333 => x"0d775680",
   334 => x"55747627",
   335 => x"81993880",
   336 => x"e6a00854",
   337 => x"bfa9bc0b",
   338 => x"94150c85",
   339 => x"0b98150c",
   340 => x"98140870",
   341 => x"81065153",
   342 => x"72f638bf",
   343 => x"a9bc0b94",
   344 => x"150c850b",
   345 => x"98150c98",
   346 => x"14087081",
   347 => x"06515372",
   348 => x"f638bfa9",
   349 => x"bc0b9415",
   350 => x"0c850b98",
   351 => x"150c9814",
   352 => x"08708106",
   353 => x"515372f6",
   354 => x"38bfa9bc",
   355 => x"0b94150c",
   356 => x"850b9815",
   357 => x"0c981408",
   358 => x"70810651",
   359 => x"5372f638",
   360 => x"bfa9bc0b",
   361 => x"94150c85",
   362 => x"0b98150c",
   363 => x"98140870",
   364 => x"81065153",
   365 => x"72f638bf",
   366 => x"a9bc0b94",
   367 => x"150c850b",
   368 => x"98150c98",
   369 => x"14087081",
   370 => x"06515372",
   371 => x"f6388115",
   372 => x"55757526",
   373 => x"feee3887",
   374 => x"3d0d0480",
   375 => x"3d0d80e6",
   376 => x"a0085187",
   377 => x"0b84120c",
   378 => x"823d0d04",
   379 => x"f83d0d7a",
   380 => x"7c595380",
   381 => x"73565776",
   382 => x"732480de",
   383 => x"38771754",
   384 => x"8a527451",
   385 => x"80c3e13f",
   386 => x"8008b005",
   387 => x"53727434",
   388 => x"8117578a",
   389 => x"52745180",
   390 => x"c3a93f80",
   391 => x"08558008",
   392 => x"dc388008",
   393 => x"779f2a18",
   394 => x"70812c5b",
   395 => x"56568079",
   396 => x"259e3877",
   397 => x"17ff0555",
   398 => x"75187033",
   399 => x"55537433",
   400 => x"73347375",
   401 => x"348116ff",
   402 => x"16565678",
   403 => x"7624e938",
   404 => x"76185680",
   405 => x"76348a3d",
   406 => x"0d04ad78",
   407 => x"7081055a",
   408 => x"34723078",
   409 => x"1855558a",
   410 => x"52745180",
   411 => x"c2fa3f80",
   412 => x"08b00553",
   413 => x"72743481",
   414 => x"17578a52",
   415 => x"745180c2",
   416 => x"c23f8008",
   417 => x"558008fe",
   418 => x"f438ff96",
   419 => x"39f93d0d",
   420 => x"79707133",
   421 => x"7081ff06",
   422 => x"54555555",
   423 => x"70802eb1",
   424 => x"3880e6a4",
   425 => x"08527281",
   426 => x"ff068115",
   427 => x"5553728a",
   428 => x"2e80f538",
   429 => x"84120870",
   430 => x"822a8106",
   431 => x"52577080",
   432 => x"2ef23872",
   433 => x"720c7333",
   434 => x"7081ff06",
   435 => x"595377d6",
   436 => x"38747533",
   437 => x"52567080",
   438 => x"2e80c938",
   439 => x"7080e69c",
   440 => x"08595381",
   441 => x"1680edd4",
   442 => x"337081ff",
   443 => x"06701010",
   444 => x"1180edd8",
   445 => x"337081ff",
   446 => x"06729029",
   447 => x"1170882b",
   448 => x"7a077f0c",
   449 => x"53595954",
   450 => x"54585672",
   451 => x"8a2ebe38",
   452 => x"7380cf2e",
   453 => x"b8388115",
   454 => x"537280ed",
   455 => x"d8347533",
   456 => x"5372c038",
   457 => x"893d0d04",
   458 => x"84120870",
   459 => x"822a8106",
   460 => x"57587580",
   461 => x"2ef2388d",
   462 => x"720c8412",
   463 => x"0870822a",
   464 => x"81065257",
   465 => x"70802efe",
   466 => x"eb38fef7",
   467 => x"3971a326",
   468 => x"99388117",
   469 => x"527180ed",
   470 => x"d434800b",
   471 => x"80edd834",
   472 => x"75335372",
   473 => x"fefd38ff",
   474 => x"bb39800b",
   475 => x"80edd434",
   476 => x"800b80ed",
   477 => x"d834e939",
   478 => x"fd3d0d80",
   479 => x"e6980854",
   480 => x"80d50b84",
   481 => x"150c80e6",
   482 => x"a4085284",
   483 => x"12088106",
   484 => x"5170802e",
   485 => x"f6387108",
   486 => x"7081ff06",
   487 => x"f6115254",
   488 => x"5170ae26",
   489 => x"8c387010",
   490 => x"1080e3f0",
   491 => x"05517008",
   492 => x"04841208",
   493 => x"70822a70",
   494 => x"81065151",
   495 => x"5170802e",
   496 => x"f038ab72",
   497 => x"0c728a2e",
   498 => x"aa388412",
   499 => x"0870822a",
   500 => x"70810651",
   501 => x"51517080",
   502 => x"2ef03872",
   503 => x"720c8412",
   504 => x"0870822a",
   505 => x"81065153",
   506 => x"72802ef2",
   507 => x"38ad720c",
   508 => x"ff993984",
   509 => x"12087082",
   510 => x"2a708106",
   511 => x"51515170",
   512 => x"802ef038",
   513 => x"8d720c84",
   514 => x"12087082",
   515 => x"2a708106",
   516 => x"51515170",
   517 => x"802effb2",
   518 => x"38c13981",
   519 => x"ff0b8415",
   520 => x"0cfee839",
   521 => x"80ff0b84",
   522 => x"150cfedf",
   523 => x"39bf0b84",
   524 => x"150cfed7",
   525 => x"399f0b84",
   526 => x"150cfecf",
   527 => x"398f0b84",
   528 => x"150cfec7",
   529 => x"39870b84",
   530 => x"150cfebf",
   531 => x"39830b84",
   532 => x"150cfeb7",
   533 => x"39810b84",
   534 => x"150cfeaf",
   535 => x"39800b84",
   536 => x"150cfea7",
   537 => x"39d73d0d",
   538 => x"80e69c08",
   539 => x"55800b84",
   540 => x"160cfe80",
   541 => x"0a0b8816",
   542 => x"0c800b80",
   543 => x"edd43480",
   544 => x"0b80edd8",
   545 => x"34a63d70",
   546 => x"5380e694",
   547 => x"088c1108",
   548 => x"53555bfa",
   549 => x"d73f80da",
   550 => x"ec0b80da",
   551 => x"ec33555a",
   552 => x"73802e80",
   553 => x"cc3880e6",
   554 => x"9c087457",
   555 => x"5c811a80",
   556 => x"edd43370",
   557 => x"81ff0670",
   558 => x"10101180",
   559 => x"edd83370",
   560 => x"81ff0672",
   561 => x"90291170",
   562 => x"882b7d07",
   563 => x"630c445c",
   564 => x"5c42575a",
   565 => x"5a758a2e",
   566 => x"87bd3876",
   567 => x"80cf2e87",
   568 => x"b6388118",
   569 => x"577680ed",
   570 => x"d8347933",
   571 => x"5675ffbd",
   572 => x"387a7b33",
   573 => x"555a7380",
   574 => x"2e80cc38",
   575 => x"80e69c08",
   576 => x"74575b81",
   577 => x"1a80edd4",
   578 => x"337081ff",
   579 => x"06701010",
   580 => x"1180edd8",
   581 => x"337081ff",
   582 => x"06729029",
   583 => x"1170882b",
   584 => x"7d07620c",
   585 => x"465c5c44",
   586 => x"575a5a75",
   587 => x"8a2e8785",
   588 => x"387680cf",
   589 => x"2e86fe38",
   590 => x"81185978",
   591 => x"80edd834",
   592 => x"79335675",
   593 => x"ffbd3880",
   594 => x"db840b80",
   595 => x"db843355",
   596 => x"5a73802e",
   597 => x"80cc3880",
   598 => x"e69c0874",
   599 => x"575b811a",
   600 => x"80edd433",
   601 => x"7081ff06",
   602 => x"70101011",
   603 => x"80edd833",
   604 => x"7081ff06",
   605 => x"72902911",
   606 => x"70882b7d",
   607 => x"07620c49",
   608 => x"5c5c5757",
   609 => x"5a5a758a",
   610 => x"2e85ee38",
   611 => x"7680cf2e",
   612 => x"85e73881",
   613 => x"185d7c80",
   614 => x"edd83479",
   615 => x"335675ff",
   616 => x"bd3880e6",
   617 => x"94087008",
   618 => x"a53d5b57",
   619 => x"5a8b5380",
   620 => x"d7c45278",
   621 => x"5180c0d1",
   622 => x"3f820284",
   623 => x"05818905",
   624 => x"5957758f",
   625 => x"06547389",
   626 => x"26859238",
   627 => x"7618b015",
   628 => x"55557375",
   629 => x"3475842a",
   630 => x"ff187081",
   631 => x"ff06595c",
   632 => x"5676df38",
   633 => x"78793355",
   634 => x"5a73802e",
   635 => x"80cc3880",
   636 => x"e69c0874",
   637 => x"575b811a",
   638 => x"80edd433",
   639 => x"7081ff06",
   640 => x"70101011",
   641 => x"80edd833",
   642 => x"7081ff06",
   643 => x"72902911",
   644 => x"70882b7d",
   645 => x"07620c45",
   646 => x"5c5c5f57",
   647 => x"5a5a758a",
   648 => x"2e87f338",
   649 => x"7680cf2e",
   650 => x"87ec3881",
   651 => x"18577680",
   652 => x"edd83479",
   653 => x"335675ff",
   654 => x"bd3880db",
   655 => x"900b80db",
   656 => x"9033555a",
   657 => x"73802e80",
   658 => x"cc3880e6",
   659 => x"9c087457",
   660 => x"5b811a80",
   661 => x"edd43370",
   662 => x"81ff0670",
   663 => x"10101180",
   664 => x"edd83370",
   665 => x"81ff0672",
   666 => x"90291170",
   667 => x"882b7d07",
   668 => x"620c475c",
   669 => x"5c45575a",
   670 => x"5a758a2e",
   671 => x"87b63876",
   672 => x"80cf2e87",
   673 => x"af388118",
   674 => x"597880ed",
   675 => x"d8347933",
   676 => x"5675ffbd",
   677 => x"38805f89",
   678 => x"0a5cac3d",
   679 => x"087f2e09",
   680 => x"810687ca",
   681 => x"387ea13d",
   682 => x"02880580",
   683 => x"fd054041",
   684 => x"5d7cbf06",
   685 => x"436285d4",
   686 => x"3880dae4",
   687 => x"0b80dae4",
   688 => x"33555a73",
   689 => x"802e80cc",
   690 => x"3880e69c",
   691 => x"0874575b",
   692 => x"811a80ed",
   693 => x"d4337081",
   694 => x"ff067010",
   695 => x"101180ed",
   696 => x"d8337081",
   697 => x"ff067290",
   698 => x"29117088",
   699 => x"2b7d0762",
   700 => x"0c475c5c",
   701 => x"45575a5a",
   702 => x"758a2e84",
   703 => x"8a387680",
   704 => x"cf2e8483",
   705 => x"38811856",
   706 => x"7580edd8",
   707 => x"34793356",
   708 => x"75ffbd38",
   709 => x"7b568b53",
   710 => x"80d7c452",
   711 => x"7f51bde9",
   712 => x"3f885775",
   713 => x"8f065473",
   714 => x"892683d2",
   715 => x"38761eb0",
   716 => x"15555573",
   717 => x"75347584",
   718 => x"2aff1870",
   719 => x"81ff0659",
   720 => x"5b5676df",
   721 => x"387f6033",
   722 => x"555a7380",
   723 => x"2e85bf38",
   724 => x"80e69c08",
   725 => x"74575b81",
   726 => x"1a80edd4",
   727 => x"337081ff",
   728 => x"06701010",
   729 => x"1180edd8",
   730 => x"337081ff",
   731 => x"06729029",
   732 => x"1170882b",
   733 => x"7d07620c",
   734 => x"5a5c5c44",
   735 => x"575a5a75",
   736 => x"8a2e83bf",
   737 => x"387680cf",
   738 => x"2e83b838",
   739 => x"81185978",
   740 => x"80edd834",
   741 => x"79335675",
   742 => x"ffbd3880",
   743 => x"db940b80",
   744 => x"db943355",
   745 => x"5a73802e",
   746 => x"80c73873",
   747 => x"56811a80",
   748 => x"edd43370",
   749 => x"81ff0670",
   750 => x"10101180",
   751 => x"edd83370",
   752 => x"81ff0672",
   753 => x"90291170",
   754 => x"882b7d07",
   755 => x"620c495c",
   756 => x"5c57575a",
   757 => x"5a758a2e",
   758 => x"82cb3876",
   759 => x"80cf2e82",
   760 => x"c4388118",
   761 => x"557480ed",
   762 => x"d8347933",
   763 => x"5675ffbd",
   764 => x"387b087c",
   765 => x"32703071",
   766 => x"07709f2a",
   767 => x"7081ff06",
   768 => x"b0117081",
   769 => x"ff0680ed",
   770 => x"d4337081",
   771 => x"ff067010",
   772 => x"101180ed",
   773 => x"d8337081",
   774 => x"ff067290",
   775 => x"29117088",
   776 => x"2b770767",
   777 => x"0c4e5859",
   778 => x"5c535f46",
   779 => x"5a52595b",
   780 => x"58608a2e",
   781 => x"83a43876",
   782 => x"80cf2e83",
   783 => x"9d388118",
   784 => x"416080ed",
   785 => x"d834791f",
   786 => x"841d811f",
   787 => x"5f5d5f8f",
   788 => x"ff7d27fc",
   789 => x"dc387e80",
   790 => x"0cab3d0d",
   791 => x"047618b7",
   792 => x"15555573",
   793 => x"75347584",
   794 => x"2aff1870",
   795 => x"81ff0659",
   796 => x"5c5676fa",
   797 => x"cd38faec",
   798 => x"3974a326",
   799 => x"80f13881",
   800 => x"19557480",
   801 => x"edd43480",
   802 => x"0b80edd8",
   803 => x"34793356",
   804 => x"75f9cb38",
   805 => x"fa8c3974",
   806 => x"a32680c4",
   807 => x"38811956",
   808 => x"7580edd4",
   809 => x"34800b80",
   810 => x"edd83479",
   811 => x"335675f7",
   812 => x"fc38f8bd",
   813 => x"3974a326",
   814 => x"99388119",
   815 => x"587780ed",
   816 => x"d434800b",
   817 => x"80edd834",
   818 => x"79335675",
   819 => x"f8b538f8",
   820 => x"f639800b",
   821 => x"80edd434",
   822 => x"800b80ed",
   823 => x"d834e939",
   824 => x"800b80ed",
   825 => x"d434800b",
   826 => x"80edd834",
   827 => x"ffbd3980",
   828 => x"0b80edd4",
   829 => x"34800b80",
   830 => x"edd834ff",
   831 => x"9039761e",
   832 => x"b7155555",
   833 => x"fcad3974",
   834 => x"a32680f1",
   835 => x"38811955",
   836 => x"7480edd4",
   837 => x"34800b80",
   838 => x"edd83479",
   839 => x"335675fb",
   840 => x"af38fbf0",
   841 => x"3974a326",
   842 => x"80c43881",
   843 => x"19587780",
   844 => x"edd43480",
   845 => x"0b80edd8",
   846 => x"34793356",
   847 => x"75fcee38",
   848 => x"fdaf3974",
   849 => x"a3269938",
   850 => x"81195776",
   851 => x"80edd434",
   852 => x"800b80ed",
   853 => x"d8347933",
   854 => x"5675fbfb",
   855 => x"38fcbc39",
   856 => x"800b80ed",
   857 => x"d434800b",
   858 => x"80edd834",
   859 => x"e939800b",
   860 => x"80edd434",
   861 => x"800b80ed",
   862 => x"d834ffbd",
   863 => x"39800b80",
   864 => x"edd43480",
   865 => x"0b80edd8",
   866 => x"34ff9039",
   867 => x"80e69c08",
   868 => x"7c087d32",
   869 => x"70307107",
   870 => x"709f2a70",
   871 => x"81ff06b0",
   872 => x"117081ff",
   873 => x"0680edd4",
   874 => x"337081ff",
   875 => x"06701010",
   876 => x"1180edd8",
   877 => x"337081ff",
   878 => x"06729029",
   879 => x"1170882b",
   880 => x"77077d0c",
   881 => x"4f58595d",
   882 => x"5340475b",
   883 => x"525a5c59",
   884 => x"5b608a2e",
   885 => x"098106fc",
   886 => x"de3875a3",
   887 => x"26a23881",
   888 => x"195b7a80",
   889 => x"edd43480",
   890 => x"0b80edd8",
   891 => x"34791f84",
   892 => x"1d811f5f",
   893 => x"5d5f8fff",
   894 => x"7d27f9b5",
   895 => x"38fcd739",
   896 => x"800b80ed",
   897 => x"d434800b",
   898 => x"80edd834",
   899 => x"e03980e6",
   900 => x"9c085bfb",
   901 => x"863974a3",
   902 => x"2680c438",
   903 => x"81195675",
   904 => x"80edd434",
   905 => x"800b80ed",
   906 => x"d8347933",
   907 => x"5675f7c6",
   908 => x"38f88739",
   909 => x"74a32699",
   910 => x"38811958",
   911 => x"7780edd4",
   912 => x"34800b80",
   913 => x"edd83479",
   914 => x"335675f8",
   915 => x"8438f8c5",
   916 => x"39800b80",
   917 => x"edd43480",
   918 => x"0b80edd8",
   919 => x"34e93980",
   920 => x"0b80edd4",
   921 => x"34800b80",
   922 => x"edd834ff",
   923 => x"bd397b7f",
   924 => x"9f3d028c",
   925 => x"0580f105",
   926 => x"983d0294",
   927 => x"0580cd05",
   928 => x"45424543",
   929 => x"445d80da",
   930 => x"e40b80da",
   931 => x"e433555a",
   932 => x"73802e80",
   933 => x"cc3880e6",
   934 => x"9c087457",
   935 => x"5b811a80",
   936 => x"edd43370",
   937 => x"81ff0670",
   938 => x"10101180",
   939 => x"edd83370",
   940 => x"81ff0672",
   941 => x"90291170",
   942 => x"882b7d07",
   943 => x"620c5a5c",
   944 => x"5c5f575a",
   945 => x"5a758a2e",
   946 => x"84833876",
   947 => x"80cf2e83",
   948 => x"fc388118",
   949 => x"577680ed",
   950 => x"d8347933",
   951 => x"5675ffbd",
   952 => x"387c568b",
   953 => x"5380d7c4",
   954 => x"526051b6",
   955 => x"9c3f8857",
   956 => x"758f0654",
   957 => x"73892683",
   958 => x"cb386117",
   959 => x"b0155555",
   960 => x"73753475",
   961 => x"842aff18",
   962 => x"7081ff06",
   963 => x"595b5676",
   964 => x"df386061",
   965 => x"33555a73",
   966 => x"802e84e3",
   967 => x"3880e69c",
   968 => x"0874575b",
   969 => x"811a80ed",
   970 => x"d4337081",
   971 => x"ff067010",
   972 => x"101180ed",
   973 => x"d8337081",
   974 => x"ff067290",
   975 => x"29117088",
   976 => x"2b7d0762",
   977 => x"0c425c5c",
   978 => x"57575a5a",
   979 => x"758a2e83",
   980 => x"9a387680",
   981 => x"cf2e8393",
   982 => x"38811859",
   983 => x"7880edd8",
   984 => x"34793356",
   985 => x"75ffbd38",
   986 => x"80edd433",
   987 => x"7081ff06",
   988 => x"70101011",
   989 => x"80edd833",
   990 => x"7081ff06",
   991 => x"72902911",
   992 => x"70882ba0",
   993 => x"07610c41",
   994 => x"595a5657",
   995 => x"587480cf",
   996 => x"2e84a038",
   997 => x"81175675",
   998 => x"80edd834",
   999 => x"7c087058",
  1000 => x"5ca35380",
  1001 => x"d7d0527d",
  1002 => x"51b4de3f",
  1003 => x"a0567f16",
  1004 => x"77b106b0",
  1005 => x"07565974",
  1006 => x"7934760a",
  1007 => x"100aff17",
  1008 => x"7081ff06",
  1009 => x"58595775",
  1010 => x"e5387d7e",
  1011 => x"33555a73",
  1012 => x"802e8488",
  1013 => x"3880e69c",
  1014 => x"0874575b",
  1015 => x"811a80ed",
  1016 => x"d4337081",
  1017 => x"ff067010",
  1018 => x"101180ed",
  1019 => x"d8337081",
  1020 => x"ff067290",
  1021 => x"29117088",
  1022 => x"2b7d0762",
  1023 => x"0c535c5c",
  1024 => x"57575a5a",
  1025 => x"758a2e82",
  1026 => x"80387680",
  1027 => x"cf2e81f9",
  1028 => x"38811856",
  1029 => x"7580edd8",
  1030 => x"34793356",
  1031 => x"75ffbd38",
  1032 => x"80edd433",
  1033 => x"7081ff06",
  1034 => x"70101011",
  1035 => x"80edd833",
  1036 => x"7081ff06",
  1037 => x"72902911",
  1038 => x"70882ba0",
  1039 => x"07610c5a",
  1040 => x"5e5a5657",
  1041 => x"587980cf",
  1042 => x"2e83c538",
  1043 => x"81175877",
  1044 => x"80edd834",
  1045 => x"7c7c2e83",
  1046 => x"d43880db",
  1047 => x"980b80db",
  1048 => x"9833555a",
  1049 => x"73802e80",
  1050 => x"c7387356",
  1051 => x"811a80ed",
  1052 => x"d4337081",
  1053 => x"ff067010",
  1054 => x"101180ed",
  1055 => x"d8337081",
  1056 => x"ff067290",
  1057 => x"29117088",
  1058 => x"2b7d0762",
  1059 => x"0c425c5c",
  1060 => x"57575a5a",
  1061 => x"758a2e81",
  1062 => x"8d387680",
  1063 => x"cf2e8186",
  1064 => x"38811857",
  1065 => x"7680edd8",
  1066 => x"34793356",
  1067 => x"75ffbd38",
  1068 => x"841d6381",
  1069 => x"05445d9f",
  1070 => x"6327fbca",
  1071 => x"387e800c",
  1072 => x"ab3d0d04",
  1073 => x"6117b715",
  1074 => x"5555fcb4",
  1075 => x"3974a326",
  1076 => x"81803881",
  1077 => x"19567580",
  1078 => x"edd43480",
  1079 => x"0b80edd8",
  1080 => x"34793356",
  1081 => x"75fbb638",
  1082 => x"fbf73974",
  1083 => x"a32680f1",
  1084 => x"38811958",
  1085 => x"7780edd4",
  1086 => x"34800b80",
  1087 => x"edd83479",
  1088 => x"335675fc",
  1089 => x"9f38fce0",
  1090 => x"3974a326",
  1091 => x"b7388119",
  1092 => x"577680ed",
  1093 => x"d434800b",
  1094 => x"80edd834",
  1095 => x"79335675",
  1096 => x"fdba38fd",
  1097 => x"fb3974a3",
  1098 => x"2680c538",
  1099 => x"81195574",
  1100 => x"80edd434",
  1101 => x"800b80ed",
  1102 => x"d8347933",
  1103 => x"5675feac",
  1104 => x"38feed39",
  1105 => x"800b80ed",
  1106 => x"d434800b",
  1107 => x"80edd834",
  1108 => x"cb39800b",
  1109 => x"80edd434",
  1110 => x"800b80ed",
  1111 => x"d834ff81",
  1112 => x"39800b80",
  1113 => x"edd43480",
  1114 => x"0b80edd8",
  1115 => x"34ff9039",
  1116 => x"800b80ed",
  1117 => x"d434800b",
  1118 => x"80edd834",
  1119 => x"ffbc3980",
  1120 => x"e69c0880",
  1121 => x"edd43370",
  1122 => x"81ff0670",
  1123 => x"10101180",
  1124 => x"edd83370",
  1125 => x"81ff0672",
  1126 => x"90291170",
  1127 => x"882ba007",
  1128 => x"770c425a",
  1129 => x"5b575859",
  1130 => x"5b7480cf",
  1131 => x"2e098106",
  1132 => x"fbe23875",
  1133 => x"a32682b8",
  1134 => x"3881185b",
  1135 => x"7a80edd4",
  1136 => x"34800b80",
  1137 => x"edd8347c",
  1138 => x"0870585c",
  1139 => x"a35380d7",
  1140 => x"d0527d51",
  1141 => x"b0b33fa0",
  1142 => x"56fbd339",
  1143 => x"80e69c08",
  1144 => x"80edd433",
  1145 => x"7081ff06",
  1146 => x"70101011",
  1147 => x"80edd833",
  1148 => x"7081ff06",
  1149 => x"72902911",
  1150 => x"70882ba0",
  1151 => x"07770c5b",
  1152 => x"5f5b5758",
  1153 => x"595b7980",
  1154 => x"cf2e0981",
  1155 => x"06fcbd38",
  1156 => x"75a32681",
  1157 => x"cc388118",
  1158 => x"577680ed",
  1159 => x"d434800b",
  1160 => x"80edd834",
  1161 => x"7c7c2e09",
  1162 => x"8106fcae",
  1163 => x"3880dba0",
  1164 => x"0b80dba0",
  1165 => x"33555a73",
  1166 => x"802efcf4",
  1167 => x"3873811b",
  1168 => x"80edd433",
  1169 => x"7081ff06",
  1170 => x"70101011",
  1171 => x"80edd833",
  1172 => x"7081ff06",
  1173 => x"72902911",
  1174 => x"70882b78",
  1175 => x"07630c5b",
  1176 => x"5d5d4058",
  1177 => x"5b5b5675",
  1178 => x"8a2e80ca",
  1179 => x"387680cf",
  1180 => x"2e80c338",
  1181 => x"81185978",
  1182 => x"80edd834",
  1183 => x"79335675",
  1184 => x"802efcac",
  1185 => x"38811a80",
  1186 => x"edd43370",
  1187 => x"81ff0670",
  1188 => x"10101180",
  1189 => x"edd83370",
  1190 => x"81ff0672",
  1191 => x"90291170",
  1192 => x"882b7d07",
  1193 => x"620c5a5c",
  1194 => x"5c5f575a",
  1195 => x"5a758a2e",
  1196 => x"098106ff",
  1197 => x"b83874a3",
  1198 => x"26993881",
  1199 => x"19567580",
  1200 => x"edd43480",
  1201 => x"0b80edd8",
  1202 => x"34793356",
  1203 => x"75ffb638",
  1204 => x"fbde3980",
  1205 => x"0b80edd4",
  1206 => x"34800b80",
  1207 => x"edd834e9",
  1208 => x"39800b80",
  1209 => x"edd43480",
  1210 => x"0b80edd8",
  1211 => x"34feb539",
  1212 => x"800b80ed",
  1213 => x"d434800b",
  1214 => x"80edd834",
  1215 => x"fdc939d9",
  1216 => x"3d0d80db",
  1217 => x"a851e785",
  1218 => x"3f80e690",
  1219 => x"08700880",
  1220 => x"dbb8535d",
  1221 => x"55e6f63f",
  1222 => x"a63d7053",
  1223 => x"7c81ffff",
  1224 => x"06525de5",
  1225 => x"c73f7c51",
  1226 => x"e6e33f80",
  1227 => x"dbcc51e6",
  1228 => x"dc3f7b8f",
  1229 => x"2a8106a4",
  1230 => x"3d5a568b",
  1231 => x"5380d7c4",
  1232 => x"527851ad",
  1233 => x"c43f8202",
  1234 => x"84058189",
  1235 => x"05595775",
  1236 => x"8f065473",
  1237 => x"892689b3",
  1238 => x"387618b0",
  1239 => x"15555573",
  1240 => x"75347584",
  1241 => x"2aff1870",
  1242 => x"81ff0659",
  1243 => x"5b5676df",
  1244 => x"38787933",
  1245 => x"55577380",
  1246 => x"2ea93873",
  1247 => x"80e6a408",
  1248 => x"56568117",
  1249 => x"57758a2e",
  1250 => x"899d3884",
  1251 => x"15087082",
  1252 => x"2a81065b",
  1253 => x"5b79802e",
  1254 => x"f2387575",
  1255 => x"0c763356",
  1256 => x"75e03878",
  1257 => x"7933555a",
  1258 => x"73802e80",
  1259 => x"cc387380",
  1260 => x"e69c085c",
  1261 => x"56811a80",
  1262 => x"edd43370",
  1263 => x"81ff0670",
  1264 => x"10101180",
  1265 => x"edd83370",
  1266 => x"81ff0672",
  1267 => x"90291170",
  1268 => x"882b7d07",
  1269 => x"620c535c",
  1270 => x"5c57575a",
  1271 => x"5a758a2e",
  1272 => x"89863876",
  1273 => x"80cf2e88",
  1274 => x"ff388118",
  1275 => x"577680ed",
  1276 => x"d8347933",
  1277 => x"5675ffbd",
  1278 => x"3880dbe0",
  1279 => x"51e58e3f",
  1280 => x"7b902a81",
  1281 => x"06a13d5a",
  1282 => x"568b5380",
  1283 => x"d7c45278",
  1284 => x"51abf63f",
  1285 => x"82028405",
  1286 => x"80fd0559",
  1287 => x"57758f06",
  1288 => x"54738926",
  1289 => x"88a63876",
  1290 => x"18b01555",
  1291 => x"55737534",
  1292 => x"75842aff",
  1293 => x"187081ff",
  1294 => x"06595656",
  1295 => x"76df3878",
  1296 => x"79335557",
  1297 => x"73802ea9",
  1298 => x"3880e6a4",
  1299 => x"08745755",
  1300 => x"81175775",
  1301 => x"8a2e88bb",
  1302 => x"38841508",
  1303 => x"70822a81",
  1304 => x"06555873",
  1305 => x"802ef238",
  1306 => x"75750c76",
  1307 => x"335675e0",
  1308 => x"38787933",
  1309 => x"555a7380",
  1310 => x"2e80cc38",
  1311 => x"80e69c08",
  1312 => x"74575b81",
  1313 => x"1a80edd4",
  1314 => x"337081ff",
  1315 => x"06701010",
  1316 => x"1180edd8",
  1317 => x"337081ff",
  1318 => x"06729029",
  1319 => x"1170882b",
  1320 => x"7d07620c",
  1321 => x"535c5c57",
  1322 => x"575a5a75",
  1323 => x"8a2e93a1",
  1324 => x"387680cf",
  1325 => x"2e939a38",
  1326 => x"81185776",
  1327 => x"80edd834",
  1328 => x"79335675",
  1329 => x"ffbd3880",
  1330 => x"dbf451e3",
  1331 => x"c03f7b95",
  1332 => x"2a830654",
  1333 => x"73812e94",
  1334 => x"fa388174",
  1335 => x"2694ea38",
  1336 => x"73822e94",
  1337 => x"f8387383",
  1338 => x"2e88e138",
  1339 => x"80dc8851",
  1340 => x"e39b3f7c",
  1341 => x"527b972a",
  1342 => x"87068305",
  1343 => x"81712b52",
  1344 => x"5ae1e93f",
  1345 => x"7c51e385",
  1346 => x"3f80dc9c",
  1347 => x"51e2fe3f",
  1348 => x"80dca451",
  1349 => x"e2f73f7c",
  1350 => x"527b9a2a",
  1351 => x"81068105",
  1352 => x"51e1c93f",
  1353 => x"7c51e2e5",
  1354 => x"3f80dcb8",
  1355 => x"51e2de3f",
  1356 => x"7c527b9b",
  1357 => x"2a870683",
  1358 => x"0551e1b0",
  1359 => x"3f7c51e2",
  1360 => x"cc3f80dc",
  1361 => x"cc51e2c5",
  1362 => x"3f7c527b",
  1363 => x"9e2a8207",
  1364 => x"51e1993f",
  1365 => x"7c51e2b5",
  1366 => x"3f80dce0",
  1367 => x"51e2ae3f",
  1368 => x"7b9f2a9e",
  1369 => x"3d5a568b",
  1370 => x"5380d7c4",
  1371 => x"527851a9",
  1372 => x"983f8202",
  1373 => x"840580f1",
  1374 => x"05595775",
  1375 => x"8f065473",
  1376 => x"892690f6",
  1377 => x"387618b0",
  1378 => x"15555573",
  1379 => x"75347584",
  1380 => x"2aff1870",
  1381 => x"81ff0659",
  1382 => x"5d5676df",
  1383 => x"38787933",
  1384 => x"55577380",
  1385 => x"2ea93880",
  1386 => x"e6a40874",
  1387 => x"57558117",
  1388 => x"57758a2e",
  1389 => x"86823884",
  1390 => x"15087082",
  1391 => x"2a810659",
  1392 => x"5477802e",
  1393 => x"f2387575",
  1394 => x"0c763356",
  1395 => x"75e03878",
  1396 => x"7933555a",
  1397 => x"73802e80",
  1398 => x"cc3880e6",
  1399 => x"9c087457",
  1400 => x"5b811a80",
  1401 => x"edd43370",
  1402 => x"81ff0670",
  1403 => x"10101180",
  1404 => x"edd83370",
  1405 => x"81ff0672",
  1406 => x"90291170",
  1407 => x"882b7d07",
  1408 => x"620c5a5c",
  1409 => x"5c5f575a",
  1410 => x"5a758a2e",
  1411 => x"90e13876",
  1412 => x"80cf2e90",
  1413 => x"da388118",
  1414 => x"577680ed",
  1415 => x"d8347933",
  1416 => x"5675ffbd",
  1417 => x"3880e690",
  1418 => x"08841108",
  1419 => x"80dcf453",
  1420 => x"5658e0d9",
  1421 => x"3f7c5274",
  1422 => x"9fff0651",
  1423 => x"dfae3f7c",
  1424 => x"51e0ca3f",
  1425 => x"80dd8851",
  1426 => x"e0c33f7c",
  1427 => x"52748c2a",
  1428 => x"87068305",
  1429 => x"81712b52",
  1430 => x"5bdf913f",
  1431 => x"7c51e0ad",
  1432 => x"3f748f2a",
  1433 => x"810680dd",
  1434 => x"9c525ce0",
  1435 => x"a03f7b9b",
  1436 => x"3d5a568b",
  1437 => x"5380d7c4",
  1438 => x"527851a7",
  1439 => x"8c3f8202",
  1440 => x"840580e5",
  1441 => x"05595775",
  1442 => x"8f065473",
  1443 => x"89268efc",
  1444 => x"387618b0",
  1445 => x"15555573",
  1446 => x"75347584",
  1447 => x"2aff1870",
  1448 => x"81ff0659",
  1449 => x"555676df",
  1450 => x"38787933",
  1451 => x"55577380",
  1452 => x"2ea93880",
  1453 => x"e6a40874",
  1454 => x"57558117",
  1455 => x"57758a2e",
  1456 => x"849b3884",
  1457 => x"15087082",
  1458 => x"2a810655",
  1459 => x"5a73802e",
  1460 => x"f2387575",
  1461 => x"0c763356",
  1462 => x"75e03878",
  1463 => x"7933555a",
  1464 => x"73802e80",
  1465 => x"cc3880e6",
  1466 => x"9c087457",
  1467 => x"5b811a80",
  1468 => x"edd43370",
  1469 => x"81ff0670",
  1470 => x"10101180",
  1471 => x"edd83370",
  1472 => x"81ff0672",
  1473 => x"90291170",
  1474 => x"882b7d07",
  1475 => x"620c535c",
  1476 => x"5c57575a",
  1477 => x"5a758a2e",
  1478 => x"8e993876",
  1479 => x"80cf2e8e",
  1480 => x"92388118",
  1481 => x"577680ed",
  1482 => x"d8347933",
  1483 => x"5675ffbd",
  1484 => x"387b83f3",
  1485 => x"3880e690",
  1486 => x"08901108",
  1487 => x"80ddb053",
  1488 => x"5856dec9",
  1489 => x"3f768f3d",
  1490 => x"5a568b53",
  1491 => x"80d7c452",
  1492 => x"7851a5b5",
  1493 => x"3f880284",
  1494 => x"05b50559",
  1495 => x"57758f06",
  1496 => x"54738926",
  1497 => x"8d9d3876",
  1498 => x"18b01555",
  1499 => x"55737534",
  1500 => x"75842aff",
  1501 => x"187081ff",
  1502 => x"06595c56",
  1503 => x"76df3878",
  1504 => x"79335557",
  1505 => x"73802ea9",
  1506 => x"3880e6a4",
  1507 => x"08745755",
  1508 => x"81175775",
  1509 => x"8a2e82ea",
  1510 => x"38841508",
  1511 => x"70822a81",
  1512 => x"065d5b7b",
  1513 => x"802ef238",
  1514 => x"75750c76",
  1515 => x"335675e0",
  1516 => x"38787933",
  1517 => x"555a7380",
  1518 => x"2e80cc38",
  1519 => x"80e69c08",
  1520 => x"74575b81",
  1521 => x"1a80edd4",
  1522 => x"337081ff",
  1523 => x"06701010",
  1524 => x"1180edd8",
  1525 => x"337081ff",
  1526 => x"06729029",
  1527 => x"1170882b",
  1528 => x"7d07620c",
  1529 => x"425c5c40",
  1530 => x"575a5a75",
  1531 => x"8a2e8ca5",
  1532 => x"387680cf",
  1533 => x"2e8c9e38",
  1534 => x"81185978",
  1535 => x"80edd834",
  1536 => x"79335675",
  1537 => x"ffbd38a9",
  1538 => x"3d0d0476",
  1539 => x"18b71555",
  1540 => x"55737534",
  1541 => x"75842aff",
  1542 => x"187081ff",
  1543 => x"06595b56",
  1544 => x"76f6ac38",
  1545 => x"f6cb3984",
  1546 => x"15087082",
  1547 => x"2a810659",
  1548 => x"5477802e",
  1549 => x"f2388d75",
  1550 => x"0c841508",
  1551 => x"70822a81",
  1552 => x"065b5b79",
  1553 => x"802ef6c3",
  1554 => x"38f6cf39",
  1555 => x"7618b715",
  1556 => x"55557375",
  1557 => x"3475842a",
  1558 => x"ff187081",
  1559 => x"ff065956",
  1560 => x"5676f7b9",
  1561 => x"38f7d839",
  1562 => x"74a32699",
  1563 => x"38811956",
  1564 => x"7580edd4",
  1565 => x"34800b80",
  1566 => x"edd83479",
  1567 => x"335675f6",
  1568 => x"b438f6f5",
  1569 => x"39800b80",
  1570 => x"edd43480",
  1571 => x"0b80edd8",
  1572 => x"34e93984",
  1573 => x"15087082",
  1574 => x"2a81065b",
  1575 => x"5b79802e",
  1576 => x"f2388d75",
  1577 => x"0c841508",
  1578 => x"70822a81",
  1579 => x"06555873",
  1580 => x"802ef7a5",
  1581 => x"38f7b139",
  1582 => x"84150870",
  1583 => x"822a8106",
  1584 => x"555a7380",
  1585 => x"2ef2388d",
  1586 => x"750c8415",
  1587 => x"0870822a",
  1588 => x"81065954",
  1589 => x"77802ef9",
  1590 => x"de38f9ea",
  1591 => x"39841508",
  1592 => x"70822a81",
  1593 => x"065c587a",
  1594 => x"802ef238",
  1595 => x"8d750c84",
  1596 => x"15087082",
  1597 => x"2a810655",
  1598 => x"5a73802e",
  1599 => x"fbc538fb",
  1600 => x"d1398415",
  1601 => x"0870822a",
  1602 => x"81065954",
  1603 => x"77802ef2",
  1604 => x"388d750c",
  1605 => x"84150870",
  1606 => x"822a8106",
  1607 => x"5d5b7b80",
  1608 => x"2efcf638",
  1609 => x"fd823980",
  1610 => x"e6900888",
  1611 => x"110880dd",
  1612 => x"c453565c",
  1613 => x"dad73f74",
  1614 => x"87065473",
  1615 => x"862681a5",
  1616 => x"38731010",
  1617 => x"80e5ac05",
  1618 => x"59780804",
  1619 => x"80ddd851",
  1620 => x"dabb3f80",
  1621 => x"dc8851da",
  1622 => x"b43f7c52",
  1623 => x"7b972a87",
  1624 => x"06830581",
  1625 => x"712b525a",
  1626 => x"d9823f7c",
  1627 => x"51da9e3f",
  1628 => x"80dc9c51",
  1629 => x"da973f80",
  1630 => x"dca451da",
  1631 => x"903f7c52",
  1632 => x"7b9a2a81",
  1633 => x"06810551",
  1634 => x"d8e23f7c",
  1635 => x"51d9fe3f",
  1636 => x"80dcb851",
  1637 => x"d9f73f7c",
  1638 => x"527b9b2a",
  1639 => x"87068305",
  1640 => x"51d8c93f",
  1641 => x"7c51d9e5",
  1642 => x"3f80dccc",
  1643 => x"51d9de3f",
  1644 => x"7c527b9e",
  1645 => x"2a820751",
  1646 => x"d8b23f7c",
  1647 => x"51d9ce3f",
  1648 => x"80dce051",
  1649 => x"d9c73f7b",
  1650 => x"9f2a9e3d",
  1651 => x"5a568b53",
  1652 => x"80d7c452",
  1653 => x"7851a0b1",
  1654 => x"3f820284",
  1655 => x"0580f105",
  1656 => x"5957f797",
  1657 => x"3980dde0",
  1658 => x"51d9a23f",
  1659 => x"80dde851",
  1660 => x"d99b3f80",
  1661 => x"ddf051d9",
  1662 => x"943f7483",
  1663 => x"2a830654",
  1664 => x"73812e90",
  1665 => x"e2388174",
  1666 => x"268ae638",
  1667 => x"73822e90",
  1668 => x"ea387383",
  1669 => x"2e90c638",
  1670 => x"80de8451",
  1671 => x"d8ef3f80",
  1672 => x"de8851d8",
  1673 => x"e83f7485",
  1674 => x"2a870654",
  1675 => x"73812e90",
  1676 => x"c0388174",
  1677 => x"268ab038",
  1678 => x"73822e90",
  1679 => x"c8387383",
  1680 => x"2e909038",
  1681 => x"80de9c51",
  1682 => x"d8c33f74",
  1683 => x"902a8706",
  1684 => x"54738526",
  1685 => x"8c387310",
  1686 => x"1080e5c8",
  1687 => x"05547308",
  1688 => x"0480dde0",
  1689 => x"51d8a63f",
  1690 => x"80deb051",
  1691 => x"d89f3f7c",
  1692 => x"5274932a",
  1693 => x"83068207",
  1694 => x"51d6f13f",
  1695 => x"7c51d88d",
  1696 => x"3f80dec4",
  1697 => x"51d8863f",
  1698 => x"7c527494",
  1699 => x"2a8f0651",
  1700 => x"d6da3f7c",
  1701 => x"51d7f63f",
  1702 => x"80ded851",
  1703 => x"d7ef3f7c",
  1704 => x"5274982a",
  1705 => x"81068105",
  1706 => x"51d6c13f",
  1707 => x"7c51d7dd",
  1708 => x"3f80deec",
  1709 => x"51d7d63f",
  1710 => x"7c52749e",
  1711 => x"2a820751",
  1712 => x"d6aa3f7c",
  1713 => x"51d7c63f",
  1714 => x"80df8051",
  1715 => x"d7bf3f74",
  1716 => x"9f2a983d",
  1717 => x"5a568b53",
  1718 => x"80d7c452",
  1719 => x"78519ea9",
  1720 => x"3f820284",
  1721 => x"0580d905",
  1722 => x"5957758f",
  1723 => x"06547389",
  1724 => x"2687d438",
  1725 => x"7618b015",
  1726 => x"55557375",
  1727 => x"3475842a",
  1728 => x"ff187081",
  1729 => x"ff06595e",
  1730 => x"5676df38",
  1731 => x"78793355",
  1732 => x"5773802e",
  1733 => x"a93880e6",
  1734 => x"a4087457",
  1735 => x"55811757",
  1736 => x"758a2e84",
  1737 => x"e6388415",
  1738 => x"0870822a",
  1739 => x"8106555d",
  1740 => x"73802ef2",
  1741 => x"3875750c",
  1742 => x"76335675",
  1743 => x"e0387879",
  1744 => x"33555a73",
  1745 => x"802e80cc",
  1746 => x"3880e69c",
  1747 => x"0874575b",
  1748 => x"811a80ed",
  1749 => x"d4337081",
  1750 => x"ff067010",
  1751 => x"101180ed",
  1752 => x"d8337081",
  1753 => x"ff067290",
  1754 => x"29117088",
  1755 => x"2b7d0762",
  1756 => x"0c425c5c",
  1757 => x"40575a5a",
  1758 => x"758a2e87",
  1759 => x"83387680",
  1760 => x"cf2e86fc",
  1761 => x"38811859",
  1762 => x"7880edd8",
  1763 => x"34793356",
  1764 => x"75ffbd38",
  1765 => x"80e69008",
  1766 => x"94110880",
  1767 => x"df945358",
  1768 => x"56d5ea3f",
  1769 => x"76953d5a",
  1770 => x"568b5380",
  1771 => x"d7c45278",
  1772 => x"519cd63f",
  1773 => x"88028405",
  1774 => x"80cd0559",
  1775 => x"57758f06",
  1776 => x"54738926",
  1777 => x"86933876",
  1778 => x"18b01555",
  1779 => x"55737534",
  1780 => x"75842aff",
  1781 => x"187081ff",
  1782 => x"06595c56",
  1783 => x"76df3878",
  1784 => x"79335557",
  1785 => x"73802ea9",
  1786 => x"3880e6a4",
  1787 => x"08745755",
  1788 => x"81175775",
  1789 => x"8a2e83b8",
  1790 => x"38841508",
  1791 => x"70822a81",
  1792 => x"065d5b7b",
  1793 => x"802ef238",
  1794 => x"75750c76",
  1795 => x"335675e0",
  1796 => x"38787933",
  1797 => x"555a7380",
  1798 => x"2e80cc38",
  1799 => x"80e69c08",
  1800 => x"74575b81",
  1801 => x"1a80edd4",
  1802 => x"337081ff",
  1803 => x"06701010",
  1804 => x"1180edd8",
  1805 => x"337081ff",
  1806 => x"06729029",
  1807 => x"1170882b",
  1808 => x"7d07620c",
  1809 => x"425c5c40",
  1810 => x"575a5a75",
  1811 => x"8a2e8592",
  1812 => x"387680cf",
  1813 => x"2e858b38",
  1814 => x"81185978",
  1815 => x"80edd834",
  1816 => x"79335675",
  1817 => x"ffbd3880",
  1818 => x"e6900898",
  1819 => x"110880df",
  1820 => x"a8535856",
  1821 => x"d4973f76",
  1822 => x"923d5a56",
  1823 => x"8b5380d7",
  1824 => x"c4527851",
  1825 => x"9b833f88",
  1826 => x"02840580",
  1827 => x"c1055957",
  1828 => x"758f0654",
  1829 => x"73892684",
  1830 => x"b7387618",
  1831 => x"b0155555",
  1832 => x"73753475",
  1833 => x"842aff18",
  1834 => x"7081ff06",
  1835 => x"595b5676",
  1836 => x"df387879",
  1837 => x"33555773",
  1838 => x"802ea938",
  1839 => x"80e6a408",
  1840 => x"74575581",
  1841 => x"1757758a",
  1842 => x"2e828a38",
  1843 => x"84150870",
  1844 => x"822a8106",
  1845 => x"5d5a7b80",
  1846 => x"2ef23875",
  1847 => x"750c7633",
  1848 => x"5675e038",
  1849 => x"78793355",
  1850 => x"5a73802e",
  1851 => x"f4c73880",
  1852 => x"e69c0874",
  1853 => x"811c80ed",
  1854 => x"d4337081",
  1855 => x"ff067010",
  1856 => x"101180ed",
  1857 => x"d8337081",
  1858 => x"ff067290",
  1859 => x"29117088",
  1860 => x"2b780779",
  1861 => x"0c445e5e",
  1862 => x"42595c5c",
  1863 => x"575b758a",
  1864 => x"2e80ca38",
  1865 => x"7680cf2e",
  1866 => x"80c33881",
  1867 => x"18597880",
  1868 => x"edd83479",
  1869 => x"33567580",
  1870 => x"2ef3fa38",
  1871 => x"811a80ed",
  1872 => x"d4337081",
  1873 => x"ff067010",
  1874 => x"101180ed",
  1875 => x"d8337081",
  1876 => x"ff067290",
  1877 => x"29117088",
  1878 => x"2b7d0762",
  1879 => x"0c425c5c",
  1880 => x"40575a5a",
  1881 => x"758a2e09",
  1882 => x"8106ffb8",
  1883 => x"3874a326",
  1884 => x"83ab3881",
  1885 => x"19557480",
  1886 => x"edd43480",
  1887 => x"0b80edd8",
  1888 => x"34793356",
  1889 => x"75ffb538",
  1890 => x"f3ab3984",
  1891 => x"15087082",
  1892 => x"2a810659",
  1893 => x"5a77802e",
  1894 => x"f2388d75",
  1895 => x"0c841508",
  1896 => x"70822a81",
  1897 => x"06555d73",
  1898 => x"802efafa",
  1899 => x"38fb8639",
  1900 => x"84150870",
  1901 => x"822a8106",
  1902 => x"59547780",
  1903 => x"2ef2388d",
  1904 => x"750c8415",
  1905 => x"0870822a",
  1906 => x"81065d5b",
  1907 => x"7b802efc",
  1908 => x"a838fcb4",
  1909 => x"39841508",
  1910 => x"70822a81",
  1911 => x"06595477",
  1912 => x"802ef238",
  1913 => x"8d750c84",
  1914 => x"15087082",
  1915 => x"2a81065d",
  1916 => x"5a7b802e",
  1917 => x"fdd638fd",
  1918 => x"e2397618",
  1919 => x"b7155555",
  1920 => x"ef893976",
  1921 => x"18b71555",
  1922 => x"55f2e239",
  1923 => x"7618b715",
  1924 => x"5555f183",
  1925 => x"3974a326",
  1926 => x"819e3881",
  1927 => x"19557480",
  1928 => x"edd43480",
  1929 => x"0b80edd8",
  1930 => x"34793356",
  1931 => x"75f39438",
  1932 => x"f3d53974",
  1933 => x"a32680f1",
  1934 => x"38811956",
  1935 => x"7580edd4",
  1936 => x"34800b80",
  1937 => x"edd83479",
  1938 => x"335675f1",
  1939 => x"a038f1e1",
  1940 => x"3974a326",
  1941 => x"80c43881",
  1942 => x"19567580",
  1943 => x"edd43480",
  1944 => x"0b80edd8",
  1945 => x"34793356",
  1946 => x"75ec9838",
  1947 => x"ecd93974",
  1948 => x"a3269938",
  1949 => x"81195675",
  1950 => x"80edd434",
  1951 => x"800b80ed",
  1952 => x"d8347933",
  1953 => x"5675eed9",
  1954 => x"38ef9a39",
  1955 => x"800b80ed",
  1956 => x"d434800b",
  1957 => x"80edd834",
  1958 => x"e939800b",
  1959 => x"80edd434",
  1960 => x"800b80ed",
  1961 => x"d834ffbd",
  1962 => x"39800b80",
  1963 => x"edd43480",
  1964 => x"0b80edd8",
  1965 => x"34ff9039",
  1966 => x"800b80ed",
  1967 => x"d434800b",
  1968 => x"80edd834",
  1969 => x"fee33976",
  1970 => x"18b71555",
  1971 => x"55f8ab39",
  1972 => x"7618b715",
  1973 => x"5555fbc8",
  1974 => x"397618b7",
  1975 => x"155555f9",
  1976 => x"ec3974a3",
  1977 => x"2680d338",
  1978 => x"81195574",
  1979 => x"80edd434",
  1980 => x"800b80ed",
  1981 => x"d8347933",
  1982 => x"5675faa7",
  1983 => x"38fae839",
  1984 => x"74a326a8",
  1985 => x"38811955",
  1986 => x"7480edd4",
  1987 => x"34800b80",
  1988 => x"edd83479",
  1989 => x"335675f8",
  1990 => x"b738f8f8",
  1991 => x"39800b80",
  1992 => x"edd43480",
  1993 => x"0b80edd8",
  1994 => x"34fcd639",
  1995 => x"800b80ed",
  1996 => x"d434800b",
  1997 => x"80edd834",
  1998 => x"da39800b",
  1999 => x"80edd434",
  2000 => x"800b80ed",
  2001 => x"d834ffae",
  2002 => x"3980dfbc",
  2003 => x"51cebe3f",
  2004 => x"f4813980",
  2005 => x"dfc451ce",
  2006 => x"b43ff3f7",
  2007 => x"3980dfcc",
  2008 => x"51ceaa3f",
  2009 => x"f3ed3980",
  2010 => x"dfd451ce",
  2011 => x"a03ff5d4",
  2012 => x"3980dfdc",
  2013 => x"51ce963f",
  2014 => x"f59e3980",
  2015 => x"dfe051f4",
  2016 => x"e83980df",
  2017 => x"e451f4e1",
  2018 => x"3980dfe8",
  2019 => x"51f4da39",
  2020 => x"80dfec51",
  2021 => x"f4d33980",
  2022 => x"dff051cd",
  2023 => x"f03f80de",
  2024 => x"b051cde9",
  2025 => x"3f7c5274",
  2026 => x"932a8306",
  2027 => x"820751cc",
  2028 => x"bb3f7c51",
  2029 => x"cdd73f80",
  2030 => x"dec451cd",
  2031 => x"d03f7c52",
  2032 => x"74942a8f",
  2033 => x"0651cca4",
  2034 => x"3f7c51cd",
  2035 => x"c03f80de",
  2036 => x"d851cdb9",
  2037 => x"3f7c5274",
  2038 => x"982a8106",
  2039 => x"810551cc",
  2040 => x"8b3f7c51",
  2041 => x"cda73f80",
  2042 => x"deec51cd",
  2043 => x"a03f7c52",
  2044 => x"749e2a82",
  2045 => x"0751cbf4",
  2046 => x"3f7c51cd",
  2047 => x"903f80df",
  2048 => x"8051cd89",
  2049 => x"3f749f2a",
  2050 => x"983d5a56",
  2051 => x"8b5380d7",
  2052 => x"c4527851",
  2053 => x"93f33f82",
  2054 => x"02840580",
  2055 => x"d9055957",
  2056 => x"f5c83980",
  2057 => x"e08051cc",
  2058 => x"e43f80de",
  2059 => x"b051ccdd",
  2060 => x"3f7c5274",
  2061 => x"932a8306",
  2062 => x"820751cb",
  2063 => x"af3f7c51",
  2064 => x"cccb3f80",
  2065 => x"dec451cc",
  2066 => x"c43f7c52",
  2067 => x"74942a8f",
  2068 => x"0651cb98",
  2069 => x"3f7c51cc",
  2070 => x"b43f80de",
  2071 => x"d851ccad",
  2072 => x"3f7c5274",
  2073 => x"982a8106",
  2074 => x"810551ca",
  2075 => x"ff3f7c51",
  2076 => x"cc9b3f80",
  2077 => x"deec51cc",
  2078 => x"943f7c52",
  2079 => x"749e2a82",
  2080 => x"0751cae8",
  2081 => x"3f7c51cc",
  2082 => x"843f80df",
  2083 => x"8051cbfd",
  2084 => x"3f749f2a",
  2085 => x"983d5a56",
  2086 => x"8b5380d7",
  2087 => x"c4527851",
  2088 => x"92e73f82",
  2089 => x"02840580",
  2090 => x"d9055957",
  2091 => x"f4bc3980",
  2092 => x"e08c51cb",
  2093 => x"d83f80de",
  2094 => x"b051cbd1",
  2095 => x"3f7c5274",
  2096 => x"932a8306",
  2097 => x"820751ca",
  2098 => x"a33f7c51",
  2099 => x"cbbf3f80",
  2100 => x"dec451cb",
  2101 => x"b83f7c52",
  2102 => x"74942a8f",
  2103 => x"0651ca8c",
  2104 => x"3f7c51cb",
  2105 => x"a83f80de",
  2106 => x"d851cba1",
  2107 => x"3f7c5274",
  2108 => x"982a8106",
  2109 => x"810551c9",
  2110 => x"f33f7c51",
  2111 => x"cb8f3f80",
  2112 => x"deec51cb",
  2113 => x"883f7c52",
  2114 => x"749e2a82",
  2115 => x"0751c9dc",
  2116 => x"3f7c51ca",
  2117 => x"f83f80df",
  2118 => x"8051caf1",
  2119 => x"3f749f2a",
  2120 => x"983d5a56",
  2121 => x"8b5380d7",
  2122 => x"c4527851",
  2123 => x"91db3f82",
  2124 => x"02840580",
  2125 => x"d9055957",
  2126 => x"f3b03980",
  2127 => x"e09c51ca",
  2128 => x"cc3f80de",
  2129 => x"b051cac5",
  2130 => x"3f7c5274",
  2131 => x"932a8306",
  2132 => x"820751c9",
  2133 => x"973f7c51",
  2134 => x"cab33f80",
  2135 => x"dec451ca",
  2136 => x"ac3f7c52",
  2137 => x"74942a8f",
  2138 => x"0651c980",
  2139 => x"3f7c51ca",
  2140 => x"9c3f80de",
  2141 => x"d851ca95",
  2142 => x"3f7c5274",
  2143 => x"982a8106",
  2144 => x"810551c8",
  2145 => x"e73f7c51",
  2146 => x"ca833f80",
  2147 => x"deec51c9",
  2148 => x"fc3f7c52",
  2149 => x"749e2a82",
  2150 => x"0751c8d0",
  2151 => x"3f7c51c9",
  2152 => x"ec3f80df",
  2153 => x"8051c9e5",
  2154 => x"3f749f2a",
  2155 => x"983d5a56",
  2156 => x"8b5380d7",
  2157 => x"c4527851",
  2158 => x"90cf3f82",
  2159 => x"02840580",
  2160 => x"d9055957",
  2161 => x"f2a43980",
  2162 => x"e0a851c9",
  2163 => x"c03f80de",
  2164 => x"b051c9b9",
  2165 => x"3f7c5274",
  2166 => x"932a8306",
  2167 => x"820751c8",
  2168 => x"8b3f7c51",
  2169 => x"c9a73f80",
  2170 => x"dec451c9",
  2171 => x"a03f7c52",
  2172 => x"74942a8f",
  2173 => x"0651c7f4",
  2174 => x"3f7c51c9",
  2175 => x"903f80de",
  2176 => x"d851c989",
  2177 => x"3f7c5274",
  2178 => x"982a8106",
  2179 => x"810551c7",
  2180 => x"db3f7c51",
  2181 => x"c8f73f80",
  2182 => x"deec51c8",
  2183 => x"f03f7c52",
  2184 => x"749e2a82",
  2185 => x"0751c7c4",
  2186 => x"3f7c51c8",
  2187 => x"e03f80df",
  2188 => x"8051c8d9",
  2189 => x"3f749f2a",
  2190 => x"983d5a56",
  2191 => x"8b5380d7",
  2192 => x"c4527851",
  2193 => x"8fc33f82",
  2194 => x"02840580",
  2195 => x"d9055957",
  2196 => x"f1983980",
  2197 => x"e0b051c8",
  2198 => x"b43fefe8",
  2199 => x"3980e0b4",
  2200 => x"51c8aa3f",
  2201 => x"efb23980",
  2202 => x"e0b851c8",
  2203 => x"a03fefa8",
  2204 => x"3980e0bc",
  2205 => x"51c8963f",
  2206 => x"efca3980",
  2207 => x"e0c451c8",
  2208 => x"8c3fef94",
  2209 => x"3980dfe4",
  2210 => x"51c8823f",
  2211 => x"efb639e9",
  2212 => x"3d0d80e6",
  2213 => x"90088411",
  2214 => x"08709fff",
  2215 => x"06515454",
  2216 => x"8a54bb73",
  2217 => x"2783388f",
  2218 => x"54725287",
  2219 => x"e8518a93",
  2220 => x"3f8008fd",
  2221 => x"05742970",
  2222 => x"83ffff06",
  2223 => x"5b558070",
  2224 => x"5a5ef17e",
  2225 => x"5e5b8f0b",
  2226 => x"80e69408",
  2227 => x"7b305659",
  2228 => x"5c8c1808",
  2229 => x"56737624",
  2230 => x"9638800b",
  2231 => x"84190c77",
  2232 => x"085776ed",
  2233 => x"38770857",
  2234 => x"76802ef3",
  2235 => x"38e33978",
  2236 => x"30790770",
  2237 => x"80257e81",
  2238 => x"32075854",
  2239 => x"76802e81",
  2240 => x"8b388c18",
  2241 => x"0856757a",
  2242 => x"24818138",
  2243 => x"8055890a",
  2244 => x"758fff71",
  2245 => x"27555854",
  2246 => x"74ab3881",
  2247 => x"70740654",
  2248 => x"5672802e",
  2249 => x"a0387453",
  2250 => x"7374082e",
  2251 => x"83387553",
  2252 => x"7281ff06",
  2253 => x"84158119",
  2254 => x"8fff7127",
  2255 => x"56595555",
  2256 => x"74802ed7",
  2257 => x"38747981",
  2258 => x"32545474",
  2259 => x"92388170",
  2260 => x"74065755",
  2261 => x"75802e87",
  2262 => x"38748c19",
  2263 => x"085c5973",
  2264 => x"802e9238",
  2265 => x"81707a06",
  2266 => x"56547480",
  2267 => x"2e873873",
  2268 => x"8c19085d",
  2269 => x"5d800b88",
  2270 => x"190c7708",
  2271 => x"5473feef",
  2272 => x"38770854",
  2273 => x"73802ef2",
  2274 => x"38fee439",
  2275 => x"739f2a53",
  2276 => x"7c802e82",
  2277 => x"b1388170",
  2278 => x"74065b55",
  2279 => x"79802e82",
  2280 => x"a5387b7b",
  2281 => x"31569e76",
  2282 => x"25829f38",
  2283 => x"759f2a16",
  2284 => x"70762c7d",
  2285 => x"7131778c",
  2286 => x"1c087073",
  2287 => x"31535952",
  2288 => x"525f5480",
  2289 => x"74259938",
  2290 => x"ff145480",
  2291 => x"0b84190c",
  2292 => x"77085776",
  2293 => x"ee387708",
  2294 => x"5776802e",
  2295 => x"f338e439",
  2296 => x"800b80e6",
  2297 => x"9c085654",
  2298 => x"73882b75",
  2299 => x"0c811454",
  2300 => x"97907426",
  2301 => x"f338800b",
  2302 => x"80edd434",
  2303 => x"800b80ed",
  2304 => x"d83480da",
  2305 => x"e451c585",
  2306 => x"3f7d802e",
  2307 => x"82e03880",
  2308 => x"e2c051c4",
  2309 => x"f83f80da",
  2310 => x"e451c4f1",
  2311 => x"3f78802e",
  2312 => x"82c53880",
  2313 => x"e2cc51c4",
  2314 => x"e43f80da",
  2315 => x"e451c4dd",
  2316 => x"3f7c802e",
  2317 => x"81a23880",
  2318 => x"e19c51c4",
  2319 => x"d03f80e1",
  2320 => x"a851c4c9",
  2321 => x"3f943d70",
  2322 => x"537b5259",
  2323 => x"c39e3f78",
  2324 => x"51c4ba3f",
  2325 => x"80e1b851",
  2326 => x"c4b33f78",
  2327 => x"527b51c3",
  2328 => x"8b3f7851",
  2329 => x"c4a73f80",
  2330 => x"dae451c4",
  2331 => x"a03f80e1",
  2332 => x"c851c499",
  2333 => x"3f785275",
  2334 => x"51c2f13f",
  2335 => x"7851c48d",
  2336 => x"3f80e2d8",
  2337 => x"51c4863f",
  2338 => x"7852759f",
  2339 => x"2a167081",
  2340 => x"2c525cc2",
  2341 => x"d73f7851",
  2342 => x"c3f33f80",
  2343 => x"dae451c3",
  2344 => x"ec3f80e2",
  2345 => x"8851c3e5",
  2346 => x"3f785280",
  2347 => x"e694088c",
  2348 => x"1108525b",
  2349 => x"c2b63f78",
  2350 => x"51c3d23f",
  2351 => x"7d81ff06",
  2352 => x"800c993d",
  2353 => x"0d047b7b",
  2354 => x"3156a80b",
  2355 => x"8c190870",
  2356 => x"72315256",
  2357 => x"54fdec39",
  2358 => x"80e2a051",
  2359 => x"c3af3f80",
  2360 => x"e1a851c3",
  2361 => x"a83f943d",
  2362 => x"70537b52",
  2363 => x"59c1fd3f",
  2364 => x"7851c399",
  2365 => x"3f80e1b8",
  2366 => x"51c3923f",
  2367 => x"78527b51",
  2368 => x"c1ea3f78",
  2369 => x"51c3863f",
  2370 => x"80dae451",
  2371 => x"c2ff3f80",
  2372 => x"e1c851c2",
  2373 => x"f83f7852",
  2374 => x"7551c1d0",
  2375 => x"3f7851c2",
  2376 => x"ec3f80e2",
  2377 => x"d851c2e5",
  2378 => x"3f785275",
  2379 => x"9f2a1670",
  2380 => x"812c525c",
  2381 => x"c1b63f78",
  2382 => x"51c2d23f",
  2383 => x"80dae451",
  2384 => x"c2cb3f80",
  2385 => x"e28851c2",
  2386 => x"c43f7852",
  2387 => x"80e69408",
  2388 => x"8c110852",
  2389 => x"5bc1953f",
  2390 => x"7851c2b1",
  2391 => x"3f7d81ff",
  2392 => x"06800c99",
  2393 => x"3d0d0480",
  2394 => x"e2e851fd",
  2395 => x"ba3980e2",
  2396 => x"f851fd9f",
  2397 => x"39ea3d0d",
  2398 => x"800b80e6",
  2399 => x"98087008",
  2400 => x"810a0680",
  2401 => x"edd00c57",
  2402 => x"57c0d03f",
  2403 => x"80e6a408",
  2404 => x"54b60b8c",
  2405 => x"150c830b",
  2406 => x"88150c80",
  2407 => x"e69c0877",
  2408 => x"84120c53",
  2409 => x"fe800a0b",
  2410 => x"88140c76",
  2411 => x"80edd434",
  2412 => x"7680edd8",
  2413 => x"3480e690",
  2414 => x"0854fac9",
  2415 => x"8e868c74",
  2416 => x"0c730870",
  2417 => x"842a8106",
  2418 => x"595577f5",
  2419 => x"3880e388",
  2420 => x"51c1ba3f",
  2421 => x"80edd008",
  2422 => x"802e83bc",
  2423 => x"3880e390",
  2424 => x"51c1aa3f",
  2425 => x"80e3a051",
  2426 => x"c1a33f80",
  2427 => x"dab451c1",
  2428 => x"9c3fda8b",
  2429 => x"3f8551ff",
  2430 => x"beb83f89",
  2431 => x"0a5383ff",
  2432 => x"ff547273",
  2433 => x"0c8413ff",
  2434 => x"15555373",
  2435 => x"8025f338",
  2436 => x"f8fd3f80",
  2437 => x"e3c451c0",
  2438 => x"f43f81f9",
  2439 => x"0a537273",
  2440 => x"0cf88013",
  2441 => x"5372890a",
  2442 => x"27f43880",
  2443 => x"56890a55",
  2444 => x"74087532",
  2445 => x"70307072",
  2446 => x"07802578",
  2447 => x"05888018",
  2448 => x"58585454",
  2449 => x"81f90a75",
  2450 => x"27e6388e",
  2451 => x"3d705376",
  2452 => x"5255ffbf",
  2453 => x"973f7451",
  2454 => x"c0b33f80",
  2455 => x"e3d851c0",
  2456 => x"ac3f8551",
  2457 => x"ffbdcb3f",
  2458 => x"800b80e6",
  2459 => x"9c085654",
  2460 => x"73882b75",
  2461 => x"0c811454",
  2462 => x"97907426",
  2463 => x"f338800b",
  2464 => x"80edd434",
  2465 => x"800b80ed",
  2466 => x"d834893d",
  2467 => x"587651c3",
  2468 => x"d43f80e6",
  2469 => x"98087008",
  2470 => x"70872a81",
  2471 => x"06555754",
  2472 => x"72802e8b",
  2473 => x"3880e694",
  2474 => x"0853800b",
  2475 => x"84140c73",
  2476 => x"0870842a",
  2477 => x"81065653",
  2478 => x"74802e8b",
  2479 => x"3880e694",
  2480 => x"0855800b",
  2481 => x"88160c73",
  2482 => x"0870852a",
  2483 => x"81065755",
  2484 => x"75802e81",
  2485 => x"8b3880e6",
  2486 => x"900854fa",
  2487 => x"c98e868c",
  2488 => x"740c7308",
  2489 => x"70842a81",
  2490 => x"06575575",
  2491 => x"f538890a",
  2492 => x"5383ffff",
  2493 => x"5472730c",
  2494 => x"8413ff15",
  2495 => x"55537380",
  2496 => x"25f338f7",
  2497 => x"8a3f80e3",
  2498 => x"c451ffbf",
  2499 => x"803f81f9",
  2500 => x"0a537273",
  2501 => x"0cf88013",
  2502 => x"5372890a",
  2503 => x"27f43880",
  2504 => x"56890a55",
  2505 => x"74087532",
  2506 => x"70307072",
  2507 => x"07802578",
  2508 => x"05888018",
  2509 => x"58585454",
  2510 => x"81f90a75",
  2511 => x"27e63877",
  2512 => x"527551ff",
  2513 => x"bda63f77",
  2514 => x"51ffbec1",
  2515 => x"3f80e3d8",
  2516 => x"51ffbeb9",
  2517 => x"3f8551ff",
  2518 => x"bbd83f80",
  2519 => x"e6980854",
  2520 => x"73087086",
  2521 => x"2a810657",
  2522 => x"5375802e",
  2523 => x"fe9f3880",
  2524 => x"0b80e69c",
  2525 => x"08565473",
  2526 => x"882b750c",
  2527 => x"81145497",
  2528 => x"907426f3",
  2529 => x"38800b80",
  2530 => x"edd43480",
  2531 => x"0b80edd8",
  2532 => x"34768132",
  2533 => x"57fdf639",
  2534 => x"80e3e051",
  2535 => x"ffbdee3f",
  2536 => x"80e3a051",
  2537 => x"ffbde63f",
  2538 => x"80dab451",
  2539 => x"ffbdde3f",
  2540 => x"d6cd3f85",
  2541 => x"51ffbafa",
  2542 => x"3f890a53",
  2543 => x"83ffff54",
  2544 => x"fcc0398c",
  2545 => x"08028c0c",
  2546 => x"fd3d0d80",
  2547 => x"538c088c",
  2548 => x"0508528c",
  2549 => x"08880508",
  2550 => x"5182de3f",
  2551 => x"80087080",
  2552 => x"0c54853d",
  2553 => x"0d8c0c04",
  2554 => x"8c08028c",
  2555 => x"0cfd3d0d",
  2556 => x"81538c08",
  2557 => x"8c050852",
  2558 => x"8c088805",
  2559 => x"085182b9",
  2560 => x"3f800870",
  2561 => x"800c5485",
  2562 => x"3d0d8c0c",
  2563 => x"048c0802",
  2564 => x"8c0cf93d",
  2565 => x"0d800b8c",
  2566 => x"08fc050c",
  2567 => x"8c088805",
  2568 => x"088025ab",
  2569 => x"388c0888",
  2570 => x"0508308c",
  2571 => x"0888050c",
  2572 => x"800b8c08",
  2573 => x"f4050c8c",
  2574 => x"08fc0508",
  2575 => x"8838810b",
  2576 => x"8c08f405",
  2577 => x"0c8c08f4",
  2578 => x"05088c08",
  2579 => x"fc050c8c",
  2580 => x"088c0508",
  2581 => x"8025ab38",
  2582 => x"8c088c05",
  2583 => x"08308c08",
  2584 => x"8c050c80",
  2585 => x"0b8c08f0",
  2586 => x"050c8c08",
  2587 => x"fc050888",
  2588 => x"38810b8c",
  2589 => x"08f0050c",
  2590 => x"8c08f005",
  2591 => x"088c08fc",
  2592 => x"050c8053",
  2593 => x"8c088c05",
  2594 => x"08528c08",
  2595 => x"88050851",
  2596 => x"81a73f80",
  2597 => x"08708c08",
  2598 => x"f8050c54",
  2599 => x"8c08fc05",
  2600 => x"08802e8c",
  2601 => x"388c08f8",
  2602 => x"0508308c",
  2603 => x"08f8050c",
  2604 => x"8c08f805",
  2605 => x"0870800c",
  2606 => x"54893d0d",
  2607 => x"8c0c048c",
  2608 => x"08028c0c",
  2609 => x"fb3d0d80",
  2610 => x"0b8c08fc",
  2611 => x"050c8c08",
  2612 => x"88050880",
  2613 => x"2593388c",
  2614 => x"08880508",
  2615 => x"308c0888",
  2616 => x"050c810b",
  2617 => x"8c08fc05",
  2618 => x"0c8c088c",
  2619 => x"05088025",
  2620 => x"8c388c08",
  2621 => x"8c050830",
  2622 => x"8c088c05",
  2623 => x"0c81538c",
  2624 => x"088c0508",
  2625 => x"528c0888",
  2626 => x"050851ad",
  2627 => x"3f800870",
  2628 => x"8c08f805",
  2629 => x"0c548c08",
  2630 => x"fc050880",
  2631 => x"2e8c388c",
  2632 => x"08f80508",
  2633 => x"308c08f8",
  2634 => x"050c8c08",
  2635 => x"f8050870",
  2636 => x"800c5487",
  2637 => x"3d0d8c0c",
  2638 => x"048c0802",
  2639 => x"8c0cfd3d",
  2640 => x"0d810b8c",
  2641 => x"08fc050c",
  2642 => x"800b8c08",
  2643 => x"f8050c8c",
  2644 => x"088c0508",
  2645 => x"8c088805",
  2646 => x"0827ac38",
  2647 => x"8c08fc05",
  2648 => x"08802ea3",
  2649 => x"38800b8c",
  2650 => x"088c0508",
  2651 => x"2499388c",
  2652 => x"088c0508",
  2653 => x"108c088c",
  2654 => x"050c8c08",
  2655 => x"fc050810",
  2656 => x"8c08fc05",
  2657 => x"0cc9398c",
  2658 => x"08fc0508",
  2659 => x"802e80c9",
  2660 => x"388c088c",
  2661 => x"05088c08",
  2662 => x"88050826",
  2663 => x"a1388c08",
  2664 => x"8805088c",
  2665 => x"088c0508",
  2666 => x"318c0888",
  2667 => x"050c8c08",
  2668 => x"f805088c",
  2669 => x"08fc0508",
  2670 => x"078c08f8",
  2671 => x"050c8c08",
  2672 => x"fc050881",
  2673 => x"2a8c08fc",
  2674 => x"050c8c08",
  2675 => x"8c050881",
  2676 => x"2a8c088c",
  2677 => x"050cffaf",
  2678 => x"398c0890",
  2679 => x"0508802e",
  2680 => x"8f388c08",
  2681 => x"88050870",
  2682 => x"8c08f405",
  2683 => x"0c518d39",
  2684 => x"8c08f805",
  2685 => x"08708c08",
  2686 => x"f4050c51",
  2687 => x"8c08f405",
  2688 => x"08800c85",
  2689 => x"3d0d8c0c",
  2690 => x"04fc3d0d",
  2691 => x"7670797b",
  2692 => x"55555555",
  2693 => x"8f72278c",
  2694 => x"38727507",
  2695 => x"83065170",
  2696 => x"802ea738",
  2697 => x"ff125271",
  2698 => x"ff2e9838",
  2699 => x"72708105",
  2700 => x"54337470",
  2701 => x"81055634",
  2702 => x"ff125271",
  2703 => x"ff2e0981",
  2704 => x"06ea3874",
  2705 => x"800c863d",
  2706 => x"0d047451",
  2707 => x"72708405",
  2708 => x"54087170",
  2709 => x"8405530c",
  2710 => x"72708405",
  2711 => x"54087170",
  2712 => x"8405530c",
  2713 => x"72708405",
  2714 => x"54087170",
  2715 => x"8405530c",
  2716 => x"72708405",
  2717 => x"54087170",
  2718 => x"8405530c",
  2719 => x"f0125271",
  2720 => x"8f26c938",
  2721 => x"83722795",
  2722 => x"38727084",
  2723 => x"05540871",
  2724 => x"70840553",
  2725 => x"0cfc1252",
  2726 => x"718326ed",
  2727 => x"387054ff",
  2728 => x"8339fd3d",
  2729 => x"0d800b80",
  2730 => x"e6840854",
  2731 => x"5472812e",
  2732 => x"9c387380",
  2733 => x"eddc0cff",
  2734 => x"b3a63fff",
  2735 => x"b2c23f80",
  2736 => x"e6a85281",
  2737 => x"51f5ae3f",
  2738 => x"800851a2",
  2739 => x"3f7280ed",
  2740 => x"dc0cffb3",
  2741 => x"8b3fffb2",
  2742 => x"a73f80e6",
  2743 => x"a8528151",
  2744 => x"f5933f80",
  2745 => x"0851873f",
  2746 => x"00ff3900",
  2747 => x"ff39f73d",
  2748 => x"0d7b80e6",
  2749 => x"ac0882c8",
  2750 => x"11085a54",
  2751 => x"5a77802e",
  2752 => x"80da3881",
  2753 => x"88188419",
  2754 => x"08ff0581",
  2755 => x"712b5955",
  2756 => x"59807424",
  2757 => x"80ea3880",
  2758 => x"7424b538",
  2759 => x"73822b78",
  2760 => x"11880556",
  2761 => x"56818019",
  2762 => x"08770653",
  2763 => x"72802eb6",
  2764 => x"38781670",
  2765 => x"08535379",
  2766 => x"51740853",
  2767 => x"722dff14",
  2768 => x"fc17fc17",
  2769 => x"79812c5a",
  2770 => x"57575473",
  2771 => x"8025d638",
  2772 => x"77085877",
  2773 => x"ffad3880",
  2774 => x"e6ac0853",
  2775 => x"bc1308a5",
  2776 => x"387951ff",
  2777 => x"833f7408",
  2778 => x"53722dff",
  2779 => x"14fc17fc",
  2780 => x"1779812c",
  2781 => x"5a575754",
  2782 => x"738025ff",
  2783 => x"a838d139",
  2784 => x"8057ff93",
  2785 => x"397251bc",
  2786 => x"13085372",
  2787 => x"2d7951fe",
  2788 => x"d73fff3d",
  2789 => x"0d80edb0",
  2790 => x"0bfc0570",
  2791 => x"08525270",
  2792 => x"ff2e9138",
  2793 => x"702dfc12",
  2794 => x"70085252",
  2795 => x"70ff2e09",
  2796 => x"8106f138",
  2797 => x"833d0d04",
  2798 => x"04ffb291",
  2799 => x"3f040000",
  2800 => x"00000040",
  2801 => x"30782020",
  2802 => x"20202020",
  2803 => x"20200000",
  2804 => x"30622020",
  2805 => x"20202020",
  2806 => x"20202020",
  2807 => x"20202020",
  2808 => x"20202020",
  2809 => x"20202020",
  2810 => x"20202020",
  2811 => x"20202020",
  2812 => x"20200000",
  2813 => x"0a677265",
  2814 => x"74682072",
  2815 => x"65676973",
  2816 => x"74657273",
  2817 => x"3a000000",
  2818 => x"0a636f6e",
  2819 => x"74726f6c",
  2820 => x"3a202020",
  2821 => x"20202000",
  2822 => x"0a737461",
  2823 => x"7475733a",
  2824 => x"20202020",
  2825 => x"20202000",
  2826 => x"0a6d6163",
  2827 => x"5f6d7362",
  2828 => x"3a202020",
  2829 => x"20202000",
  2830 => x"0a6d6163",
  2831 => x"5f6c7362",
  2832 => x"3a202020",
  2833 => x"20202000",
  2834 => x"0a6d6469",
  2835 => x"6f5f636f",
  2836 => x"6e74726f",
  2837 => x"6c3a2000",
  2838 => x"0a74785f",
  2839 => x"706f696e",
  2840 => x"7465723a",
  2841 => x"20202000",
  2842 => x"0a72785f",
  2843 => x"706f696e",
  2844 => x"7465723a",
  2845 => x"20202000",
  2846 => x"0a656463",
  2847 => x"6c5f6970",
  2848 => x"3a202020",
  2849 => x"20202000",
  2850 => x"0a686173",
  2851 => x"685f6d73",
  2852 => x"623a2020",
  2853 => x"20202000",
  2854 => x"0a686173",
  2855 => x"685f6c73",
  2856 => x"623a2020",
  2857 => x"20202000",
  2858 => x"0a6d6469",
  2859 => x"6f207068",
  2860 => x"79207265",
  2861 => x"67697374",
  2862 => x"65727300",
  2863 => x"0a206d64",
  2864 => x"696f2070",
  2865 => x"68793a20",
  2866 => x"00000000",
  2867 => x"0a202072",
  2868 => x"65673a20",
  2869 => x"00000000",
  2870 => x"2d3e2000",
  2871 => x"0a677265",
  2872 => x"74682d3e",
  2873 => x"636f6e74",
  2874 => x"726f6c20",
  2875 => x"3a000000",
  2876 => x"0a677265",
  2877 => x"74682d3e",
  2878 => x"73746174",
  2879 => x"75732020",
  2880 => x"3a000000",
  2881 => x"0a646573",
  2882 => x"63722d3e",
  2883 => x"636f6e74",
  2884 => x"726f6c20",
  2885 => x"3a000000",
  2886 => x"77726974",
  2887 => x"65206164",
  2888 => x"64726573",
  2889 => x"733a2000",
  2890 => x"20206c65",
  2891 => x"6e677468",
  2892 => x"3a200000",
  2893 => x"0a0a0000",
  2894 => x"72656164",
  2895 => x"20206164",
  2896 => x"64726573",
  2897 => x"733a2000",
  2898 => x"20206578",
  2899 => x"70656374",
  2900 => x"3a200000",
  2901 => x"2020676f",
  2902 => x"743a2000",
  2903 => x"20657272",
  2904 => x"6f720000",
  2905 => x"0a000000",
  2906 => x"206f6b00",
  2907 => x"70686173",
  2908 => x"65207368",
  2909 => x"69667420",
  2910 => x"202d2020",
  2911 => x"76616c75",
  2912 => x"653a2000",
  2913 => x"20207374",
  2914 => x"61747573",
  2915 => x"3a200000",
  2916 => x"20202020",
  2917 => x"20000000",
  2918 => x"4641494c",
  2919 => x"00000000",
  2920 => x"6f6b2020",
  2921 => x"00000000",
  2922 => x"44445220",
  2923 => x"6d656d6f",
  2924 => x"72792069",
  2925 => x"6e666f00",
  2926 => x"0a0a6175",
  2927 => x"746f2074",
  2928 => x"5f524552",
  2929 => x"45534820",
  2930 => x"3a000000",
  2931 => x"0a636c6f",
  2932 => x"636b2065",
  2933 => x"6e61626c",
  2934 => x"6520203a",
  2935 => x"00000000",
  2936 => x"0a696e69",
  2937 => x"74616c69",
  2938 => x"7a652020",
  2939 => x"2020203a",
  2940 => x"00000000",
  2941 => x"0a636f6c",
  2942 => x"756d6e20",
  2943 => x"73697a65",
  2944 => x"2020203a",
  2945 => x"00000000",
  2946 => x"0a62616e",
  2947 => x"6b73697a",
  2948 => x"65202020",
  2949 => x"2020203a",
  2950 => x"00000000",
  2951 => x"4d627974",
  2952 => x"65000000",
  2953 => x"0a745f52",
  2954 => x"43442020",
  2955 => x"20202020",
  2956 => x"2020203a",
  2957 => x"00000000",
  2958 => x"0a745f52",
  2959 => x"46432020",
  2960 => x"20202020",
  2961 => x"2020203a",
  2962 => x"00000000",
  2963 => x"0a745f52",
  2964 => x"50202020",
  2965 => x"20202020",
  2966 => x"2020203a",
  2967 => x"00000000",
  2968 => x"0a726566",
  2969 => x"72657368",
  2970 => x"20656e2e",
  2971 => x"2020203a",
  2972 => x"00000000",
  2973 => x"0a0a4444",
  2974 => x"52206672",
  2975 => x"65717565",
  2976 => x"6e637920",
  2977 => x"3a000000",
  2978 => x"0a444452",
  2979 => x"20646174",
  2980 => x"61207769",
  2981 => x"6474683a",
  2982 => x"00000000",
  2983 => x"0a6d6f62",
  2984 => x"696c6520",
  2985 => x"73757070",
  2986 => x"6f72743a",
  2987 => x"00000000",
  2988 => x"0a0a7374",
  2989 => x"61747573",
  2990 => x"20726561",
  2991 => x"64202020",
  2992 => x"3a000000",
  2993 => x"0a0a7365",
  2994 => x"6c662072",
  2995 => x"65667265",
  2996 => x"73682020",
  2997 => x"3a000000",
  2998 => x"34303639",
  2999 => x"00000000",
  3000 => x"756e6b6e",
  3001 => x"6f776e00",
  3002 => x"20617272",
  3003 => x"61790000",
  3004 => x"0a74656d",
  3005 => x"702d636f",
  3006 => x"6d702072",
  3007 => x"6566723a",
  3008 => x"00000000",
  3009 => x"c2b04300",
  3010 => x"0a647269",
  3011 => x"76652073",
  3012 => x"7472656e",
  3013 => x"6774683a",
  3014 => x"00000000",
  3015 => x"0a706f77",
  3016 => x"65722073",
  3017 => x"6176696e",
  3018 => x"6720203a",
  3019 => x"00000000",
  3020 => x"0a745f58",
  3021 => x"50202020",
  3022 => x"20202020",
  3023 => x"2020203a",
  3024 => x"00000000",
  3025 => x"0a745f58",
  3026 => x"53522020",
  3027 => x"20202020",
  3028 => x"2020203a",
  3029 => x"00000000",
  3030 => x"0a745f43",
  3031 => x"4b452020",
  3032 => x"20202020",
  3033 => x"2020203a",
  3034 => x"00000000",
  3035 => x"0a434153",
  3036 => x"206c6174",
  3037 => x"656e6379",
  3038 => x"2020203a",
  3039 => x"00000000",
  3040 => x"0a6d6f62",
  3041 => x"696c6520",
  3042 => x"656e6162",
  3043 => x"6c65643a",
  3044 => x"00000000",
  3045 => x"0a0a7068",
  3046 => x"7920636f",
  3047 => x"6e666967",
  3048 => x"20302020",
  3049 => x"3a000000",
  3050 => x"0a0a7068",
  3051 => x"7920636f",
  3052 => x"6e666967",
  3053 => x"20312020",
  3054 => x"3a000000",
  3055 => x"20353132",
  3056 => x"00000000",
  3057 => x"31303234",
  3058 => x"00000000",
  3059 => x"32303438",
  3060 => x"00000000",
  3061 => x"66756c6c",
  3062 => x"00000000",
  3063 => x"37300000",
  3064 => x"312f3800",
  3065 => x"312f3400",
  3066 => x"312f3200",
  3067 => x"312f3100",
  3068 => x"64656570",
  3069 => x"20706f77",
  3070 => x"65722064",
  3071 => x"6f776e00",
  3072 => x"636c6f63",
  3073 => x"6b207374",
  3074 => x"6f700000",
  3075 => x"73656c66",
  3076 => x"20726566",
  3077 => x"72657368",
  3078 => x"00000000",
  3079 => x"706f7765",
  3080 => x"7220646f",
  3081 => x"776e0000",
  3082 => x"6e6f6e65",
  3083 => x"00000000",
  3084 => x"332f3400",
  3085 => x"38350000",
  3086 => x"34350000",
  3087 => x"68616c66",
  3088 => x"00000000",
  3089 => x"31350000",
  3090 => x"61646472",
  3091 => x"6573733a",
  3092 => x"20000000",
  3093 => x"20646174",
  3094 => x"613a2000",
  3095 => x"0a0a4443",
  3096 => x"4d207068",
  3097 => x"61736520",
  3098 => x"73686966",
  3099 => x"74207465",
  3100 => x"7374696e",
  3101 => x"67000000",
  3102 => x"0a696e69",
  3103 => x"7469616c",
  3104 => x"3a200000",
  3105 => x"09000000",
  3106 => x"20202020",
  3107 => x"00000000",
  3108 => x"6c6f7720",
  3109 => x"666f756e",
  3110 => x"64000000",
  3111 => x"68696768",
  3112 => x"20666f75",
  3113 => x"6e640000",
  3114 => x"0a6c6f77",
  3115 => x"3a202020",
  3116 => x"20202020",
  3117 => x"20200000",
  3118 => x"0a686967",
  3119 => x"683a2020",
  3120 => x"20202020",
  3121 => x"20200000",
  3122 => x"0a646966",
  3123 => x"663a2020",
  3124 => x"20202020",
  3125 => x"20200000",
  3126 => x"0a6d696e",
  3127 => x"5f657272",
  3128 => x"3a202020",
  3129 => x"20200000",
  3130 => x"0a6d696e",
  3131 => x"5f657272",
  3132 => x"5f706f73",
  3133 => x"3a200000",
  3134 => x"676f206d",
  3135 => x"696e5f65",
  3136 => x"72726f72",
  3137 => x"00000000",
  3138 => x"0a66696e",
  3139 => x"616c3a20",
  3140 => x"20202020",
  3141 => x"20200000",
  3142 => x"676f207a",
  3143 => x"65726f00",
  3144 => x"68696768",
  3145 => x"204e4f54",
  3146 => x"20666f75",
  3147 => x"6e640000",
  3148 => x"6c6f7720",
  3149 => x"4e4f5420",
  3150 => x"666f756e",
  3151 => x"64000000",
  3152 => x"64617461",
  3153 => x"2076616c",
  3154 => x"69640000",
  3155 => x"6c6f7720",
  3156 => x"20666f75",
  3157 => x"6e640000",
  3158 => x"0a646966",
  3159 => x"662f323a",
  3160 => x"20202020",
  3161 => x"20200000",
  3162 => x"6c6f7720",
  3163 => x"204e4f54",
  3164 => x"20666f75",
  3165 => x"6e640000",
  3166 => x"64617461",
  3167 => x"204e4f54",
  3168 => x"2076616c",
  3169 => x"69640000",
  3170 => x"74657374",
  3171 => x"2e632000",
  3172 => x"286f6e20",
  3173 => x"73696d75",
  3174 => x"6c61746f",
  3175 => x"72290a00",
  3176 => x"636f6d70",
  3177 => x"696c6564",
  3178 => x"3a204f63",
  3179 => x"74203237",
  3180 => x"20323031",
  3181 => x"30202031",
  3182 => x"353a3339",
  3183 => x"3a30310a",
  3184 => x"00000000",
  3185 => x"0a0a6d65",
  3186 => x"6d6f7279",
  3187 => x"2073697a",
  3188 => x"65202020",
  3189 => x"3a000000",
  3190 => x"20626c6f",
  3191 => x"636b7300",
  3192 => x"286f6e20",
  3193 => x"68617264",
  3194 => x"77617265",
  3195 => x"290a0000",
  3196 => x"0000078b",
  3197 => x"000007b1",
  3198 => x"000007b1",
  3199 => x"0000078b",
  3200 => x"000007b1",
  3201 => x"000007b1",
  3202 => x"000007b1",
  3203 => x"000007b1",
  3204 => x"000007b1",
  3205 => x"000007b1",
  3206 => x"000007b1",
  3207 => x"000007b1",
  3208 => x"000007b1",
  3209 => x"000007b1",
  3210 => x"000007b1",
  3211 => x"000007b1",
  3212 => x"000007b1",
  3213 => x"000007b1",
  3214 => x"000007b1",
  3215 => x"000007b1",
  3216 => x"000007b1",
  3217 => x"000007b1",
  3218 => x"000007b1",
  3219 => x"000007b1",
  3220 => x"000007b1",
  3221 => x"000007b1",
  3222 => x"000007b1",
  3223 => x"000007b1",
  3224 => x"000007b1",
  3225 => x"000007b1",
  3226 => x"000007b1",
  3227 => x"000007b1",
  3228 => x"000007b1",
  3229 => x"000007b1",
  3230 => x"000007b1",
  3231 => x"000007b1",
  3232 => x"000007b1",
  3233 => x"000007b1",
  3234 => x"0000085d",
  3235 => x"00000855",
  3236 => x"0000084d",
  3237 => x"00000845",
  3238 => x"0000083d",
  3239 => x"00000835",
  3240 => x"0000082d",
  3241 => x"00000824",
  3242 => x"0000081b",
  3243 => x"00001f90",
  3244 => x"00001f89",
  3245 => x"00001f82",
  3246 => x"000019e5",
  3247 => x"000019e5",
  3248 => x"00001f7b",
  3249 => x"00001f7b",
  3250 => x"000021c7",
  3251 => x"0000213b",
  3252 => x"000020af",
  3253 => x"00001a61",
  3254 => x"00002023",
  3255 => x"00001f97",
  3256 => x"64756d6d",
  3257 => x"792e6578",
  3258 => x"65000000",
  3259 => x"43000000",
  3260 => x"00ffffff",
  3261 => x"ff00ffff",
  3262 => x"ffff00ff",
  3263 => x"ffffff00",
  3264 => x"00000000",
  3265 => x"00000000",
  3266 => x"00000000",
  3267 => x"000036b8",
  3268 => x"fff00000",
  3269 => x"80000e00",
  3270 => x"80000800",
  3271 => x"80000600",
  3272 => x"80000200",
  3273 => x"80000100",
  3274 => x"000032e0",
  3275 => x"00003330",
  3276 => x"00000000",
  3277 => x"00003598",
  3278 => x"000035f4",
  3279 => x"00003650",
  3280 => x"00000000",
  3281 => x"00000000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"00000000",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00000000",
  3288 => x"00000000",
  3289 => x"000032ec",
  3290 => x"00000000",
  3291 => x"00000000",
  3292 => x"00000000",
  3293 => x"00000000",
  3294 => x"00000000",
  3295 => x"00000000",
  3296 => x"00000000",
  3297 => x"00000000",
  3298 => x"00000000",
  3299 => x"00000000",
  3300 => x"00000000",
  3301 => x"00000000",
  3302 => x"00000000",
  3303 => x"00000000",
  3304 => x"00000000",
  3305 => x"00000000",
  3306 => x"00000000",
  3307 => x"00000000",
  3308 => x"00000000",
  3309 => x"00000000",
  3310 => x"00000000",
  3311 => x"00000000",
  3312 => x"00000000",
  3313 => x"00000000",
  3314 => x"00000000",
  3315 => x"00000000",
  3316 => x"00000000",
  3317 => x"00000000",
  3318 => x"00000001",
  3319 => x"330eabcd",
  3320 => x"1234e66d",
  3321 => x"deec0005",
  3322 => x"000b0000",
  3323 => x"00000000",
  3324 => x"00000000",
  3325 => x"00000000",
  3326 => x"00000000",
  3327 => x"00000000",
  3328 => x"00000000",
  3329 => x"00000000",
  3330 => x"00000000",
  3331 => x"00000000",
  3332 => x"00000000",
  3333 => x"00000000",
  3334 => x"00000000",
  3335 => x"00000000",
  3336 => x"00000000",
  3337 => x"00000000",
  3338 => x"00000000",
  3339 => x"00000000",
  3340 => x"00000000",
  3341 => x"00000000",
  3342 => x"00000000",
  3343 => x"00000000",
  3344 => x"00000000",
  3345 => x"00000000",
  3346 => x"00000000",
  3347 => x"00000000",
  3348 => x"00000000",
  3349 => x"00000000",
  3350 => x"00000000",
  3351 => x"00000000",
  3352 => x"00000000",
  3353 => x"00000000",
  3354 => x"00000000",
  3355 => x"00000000",
  3356 => x"00000000",
  3357 => x"00000000",
  3358 => x"00000000",
  3359 => x"00000000",
  3360 => x"00000000",
  3361 => x"00000000",
  3362 => x"00000000",
  3363 => x"00000000",
  3364 => x"00000000",
  3365 => x"00000000",
  3366 => x"00000000",
  3367 => x"00000000",
  3368 => x"00000000",
  3369 => x"00000000",
  3370 => x"00000000",
  3371 => x"00000000",
  3372 => x"00000000",
  3373 => x"00000000",
  3374 => x"00000000",
  3375 => x"00000000",
  3376 => x"00000000",
  3377 => x"00000000",
  3378 => x"00000000",
  3379 => x"00000000",
  3380 => x"00000000",
  3381 => x"00000000",
  3382 => x"00000000",
  3383 => x"00000000",
  3384 => x"00000000",
  3385 => x"00000000",
  3386 => x"00000000",
  3387 => x"00000000",
  3388 => x"00000000",
  3389 => x"00000000",
  3390 => x"00000000",
  3391 => x"00000000",
  3392 => x"00000000",
  3393 => x"00000000",
  3394 => x"00000000",
  3395 => x"00000000",
  3396 => x"00000000",
  3397 => x"00000000",
  3398 => x"00000000",
  3399 => x"00000000",
  3400 => x"00000000",
  3401 => x"00000000",
  3402 => x"00000000",
  3403 => x"00000000",
  3404 => x"00000000",
  3405 => x"00000000",
  3406 => x"00000000",
  3407 => x"00000000",
  3408 => x"00000000",
  3409 => x"00000000",
  3410 => x"00000000",
  3411 => x"00000000",
  3412 => x"00000000",
  3413 => x"00000000",
  3414 => x"00000000",
  3415 => x"00000000",
  3416 => x"00000000",
  3417 => x"00000000",
  3418 => x"00000000",
  3419 => x"00000000",
  3420 => x"00000000",
  3421 => x"00000000",
  3422 => x"00000000",
  3423 => x"00000000",
  3424 => x"00000000",
  3425 => x"00000000",
  3426 => x"00000000",
  3427 => x"00000000",
  3428 => x"00000000",
  3429 => x"00000000",
  3430 => x"00000000",
  3431 => x"00000000",
  3432 => x"00000000",
  3433 => x"00000000",
  3434 => x"00000000",
  3435 => x"00000000",
  3436 => x"00000000",
  3437 => x"00000000",
  3438 => x"00000000",
  3439 => x"00000000",
  3440 => x"00000000",
  3441 => x"00000000",
  3442 => x"00000000",
  3443 => x"00000000",
  3444 => x"00000000",
  3445 => x"00000000",
  3446 => x"00000000",
  3447 => x"00000000",
  3448 => x"00000000",
  3449 => x"00000000",
  3450 => x"00000000",
  3451 => x"00000000",
  3452 => x"00000000",
  3453 => x"00000000",
  3454 => x"00000000",
  3455 => x"00000000",
  3456 => x"00000000",
  3457 => x"00000000",
  3458 => x"00000000",
  3459 => x"00000000",
  3460 => x"00000000",
  3461 => x"00000000",
  3462 => x"00000000",
  3463 => x"00000000",
  3464 => x"00000000",
  3465 => x"00000000",
  3466 => x"00000000",
  3467 => x"00000000",
  3468 => x"00000000",
  3469 => x"00000000",
  3470 => x"00000000",
  3471 => x"00000000",
  3472 => x"00000000",
  3473 => x"00000000",
  3474 => x"00000000",
  3475 => x"00000000",
  3476 => x"00000000",
  3477 => x"00000000",
  3478 => x"00000000",
  3479 => x"00000000",
  3480 => x"00000000",
  3481 => x"00000000",
  3482 => x"00000000",
  3483 => x"00000000",
  3484 => x"00000000",
  3485 => x"00000000",
  3486 => x"00000000",
  3487 => x"00000000",
  3488 => x"00000000",
  3489 => x"00000000",
  3490 => x"00000000",
  3491 => x"00000000",
  3492 => x"00000000",
  3493 => x"00000000",
  3494 => x"00000000",
  3495 => x"00000000",
  3496 => x"00000000",
  3497 => x"00000000",
  3498 => x"00000000",
  3499 => x"ffffffff",
  3500 => x"00000000",
  3501 => x"ffffffff",
  3502 => x"00000000",
  3503 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
