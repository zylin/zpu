
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 15;
constant bytes : integer := 17984;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B0BBA";
    when 16#00001# => romdata <= X"F0040000";
    when 16#00002# => romdata <= X"00000000";
    when 16#00003# => romdata <= X"00000000";
    when 16#00004# => romdata <= X"00000000";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"0B0B0BBD";
    when 16#00009# => romdata <= X"D5040000";
    when 16#0000A# => romdata <= X"00000000";
    when 16#0000B# => romdata <= X"00000000";
    when 16#0000C# => romdata <= X"00000000";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B0BBD";
    when 16#00049# => romdata <= X"89040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B0BBCEC";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B80FC";
    when 16#000A2# => romdata <= X"CC738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B0B";
    when 16#000A5# => romdata <= X"BCEF0400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"0B0B0BBD";
    when 16#000A9# => romdata <= X"BD040000";
    when 16#000AA# => romdata <= X"00000000";
    when 16#000AB# => romdata <= X"00000000";
    when 16#000AC# => romdata <= X"00000000";
    when 16#000AD# => romdata <= X"00000000";
    when 16#000AE# => romdata <= X"00000000";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"0B0B0BBD";
    when 16#000B1# => romdata <= X"A5040000";
    when 16#000B2# => romdata <= X"00000000";
    when 16#000B3# => romdata <= X"00000000";
    when 16#000B4# => romdata <= X"00000000";
    when 16#000B5# => romdata <= X"00000000";
    when 16#000B6# => romdata <= X"00000000";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"80FCDC0C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"FF3D0D02";
    when 16#00101# => romdata <= X"8F053351";
    when 16#00102# => romdata <= X"BB893F71";
    when 16#00103# => romdata <= X"B00C833D";
    when 16#00104# => romdata <= X"0D04FD3D";
    when 16#00105# => romdata <= X"0D818CC0";
    when 16#00106# => romdata <= X"0852F881";
    when 16#00107# => romdata <= X"C08E800B";
    when 16#00108# => romdata <= X"80FCE808";
    when 16#00109# => romdata <= X"55537180";
    when 16#0010A# => romdata <= X"2E80F738";
    when 16#0010B# => romdata <= X"7281FF06";
    when 16#0010C# => romdata <= X"84150C80";
    when 16#0010D# => romdata <= X"FCBC3370";
    when 16#0010E# => romdata <= X"81FF0651";
    when 16#0010F# => romdata <= X"5271802E";
    when 16#00110# => romdata <= X"80C23872";
    when 16#00111# => romdata <= X"9F2A7310";
    when 16#00112# => romdata <= X"0753818C";
    when 16#00113# => romdata <= X"C4337081";
    when 16#00114# => romdata <= X"FF065152";
    when 16#00115# => romdata <= X"71802ED4";
    when 16#00116# => romdata <= X"38800B81";
    when 16#00117# => romdata <= X"8CC43494";
    when 16#00118# => romdata <= X"993F80FC";
    when 16#00119# => romdata <= X"B8335473";
    when 16#0011A# => romdata <= X"80E23880";
    when 16#0011B# => romdata <= X"FCE80873";
    when 16#0011C# => romdata <= X"81FF0684";
    when 16#0011D# => romdata <= X"120C80FC";
    when 16#0011E# => romdata <= X"BC337081";
    when 16#0011F# => romdata <= X"FF065153";
    when 16#00120# => romdata <= X"5471C038";
    when 16#00121# => romdata <= X"72812A73";
    when 16#00122# => romdata <= X"9F2B0753";
    when 16#00123# => romdata <= X"FFBC3972";
    when 16#00124# => romdata <= X"812A739F";
    when 16#00125# => romdata <= X"2B075380";
    when 16#00126# => romdata <= X"FD51B8E0";
    when 16#00127# => romdata <= X"3F80FCE8";
    when 16#00128# => romdata <= X"08547281";
    when 16#00129# => romdata <= X"FF068415";
    when 16#0012A# => romdata <= X"0C80FCBC";
    when 16#0012B# => romdata <= X"337081FF";
    when 16#0012C# => romdata <= X"06535471";
    when 16#0012D# => romdata <= X"802ED838";
    when 16#0012E# => romdata <= X"729F2A73";
    when 16#0012F# => romdata <= X"10075380";
    when 16#00130# => romdata <= X"FD51B8B8";
    when 16#00131# => romdata <= X"3F80FCE8";
    when 16#00132# => romdata <= X"0854D739";
    when 16#00133# => romdata <= X"800BB00C";
    when 16#00134# => romdata <= X"853D0D04";
    when 16#00135# => romdata <= X"FB3D0D8A";
    when 16#00136# => romdata <= X"51B4A03F";
    when 16#00137# => romdata <= X"8B823FAC";
    when 16#00138# => romdata <= X"B2530B0B";
    when 16#00139# => romdata <= X"80E69852";
    when 16#0013A# => romdata <= X"0B0B80E6";
    when 16#0013B# => romdata <= X"A8518B83";
    when 16#0013C# => romdata <= X"3FACC953";
    when 16#0013D# => romdata <= X"0B0B80E6";
    when 16#0013E# => romdata <= X"B0520B0B";
    when 16#0013F# => romdata <= X"80E6CC51";
    when 16#00140# => romdata <= X"8AF13F90";
    when 16#00141# => romdata <= X"F4530B0B";
    when 16#00142# => romdata <= X"80E6D452";
    when 16#00143# => romdata <= X"0B0B80E6";
    when 16#00144# => romdata <= X"E4518ADF";
    when 16#00145# => romdata <= X"3FB4DA53";
    when 16#00146# => romdata <= X"0B0B80E6";
    when 16#00147# => romdata <= X"EC520B0B";
    when 16#00148# => romdata <= X"80F2E051";
    when 16#00149# => romdata <= X"8ACD3FB6";
    when 16#0014A# => romdata <= X"C2530B0B";
    when 16#0014B# => romdata <= X"80E78452";
    when 16#0014C# => romdata <= X"0B0B80E6";
    when 16#0014D# => romdata <= X"FC518ABB";
    when 16#0014E# => romdata <= X"3FB8E353";
    when 16#0014F# => romdata <= X"0B0B80E7";
    when 16#00150# => romdata <= X"90520B0B";
    when 16#00151# => romdata <= X"80E7B051";
    when 16#00152# => romdata <= X"8AA93FB9";
    when 16#00153# => romdata <= X"CE530B0B";
    when 16#00154# => romdata <= X"80E7B852";
    when 16#00155# => romdata <= X"0B0B80E7";
    when 16#00156# => romdata <= X"DC518A97";
    when 16#00157# => romdata <= X"3FBA8753";
    when 16#00158# => romdata <= X"0B0B80E7";
    when 16#00159# => romdata <= X"E4520B0B";
    when 16#0015A# => romdata <= X"80E88051";
    when 16#0015B# => romdata <= X"8A853FBA";
    when 16#0015C# => romdata <= X"BD530B0B";
    when 16#0015D# => romdata <= X"80E88852";
    when 16#0015E# => romdata <= X"0B0B80E8";
    when 16#0015F# => romdata <= X"AC5189F3";
    when 16#00160# => romdata <= X"3FB9A353";
    when 16#00161# => romdata <= X"0B0B80E8";
    when 16#00162# => romdata <= X"B4520B0B";
    when 16#00163# => romdata <= X"80E8CC51";
    when 16#00164# => romdata <= X"89E13FB9";
    when 16#00165# => romdata <= X"BC530B0B";
    when 16#00166# => romdata <= X"80E8D452";
    when 16#00167# => romdata <= X"0B0B80E8";
    when 16#00168# => romdata <= X"F05189CF";
    when 16#00169# => romdata <= X"3FB7B853";
    when 16#0016A# => romdata <= X"0B0B80E8";
    when 16#0016B# => romdata <= X"F8520B0B";
    when 16#0016C# => romdata <= X"80E99051";
    when 16#0016D# => romdata <= X"89BD3FB8";
    when 16#0016E# => romdata <= X"8E530B0B";
    when 16#0016F# => romdata <= X"80E99852";
    when 16#00170# => romdata <= X"0B0B80E9";
    when 16#00171# => romdata <= X"B45189AB";
    when 16#00172# => romdata <= X"3F91CD53";
    when 16#00173# => romdata <= X"0B0B80E9";
    when 16#00174# => romdata <= X"BC520B0B";
    when 16#00175# => romdata <= X"80E9D051";
    when 16#00176# => romdata <= X"89993F91";
    when 16#00177# => romdata <= X"8D530B0B";
    when 16#00178# => romdata <= X"80E9D852";
    when 16#00179# => romdata <= X"0B0B80EA";
    when 16#0017A# => romdata <= X"80518987";
    when 16#0017B# => romdata <= X"3FB3BB53";
    when 16#0017C# => romdata <= X"0B0B80EA";
    when 16#0017D# => romdata <= X"88520B0B";
    when 16#0017E# => romdata <= X"80EA9C51";
    when 16#0017F# => romdata <= X"88F53F88";
    when 16#00180# => romdata <= X"92530B0B";
    when 16#00181# => romdata <= X"80EAA452";
    when 16#00182# => romdata <= X"0B0B80EA";
    when 16#00183# => romdata <= X"B45188E3";
    when 16#00184# => romdata <= X"3FA6EB53";
    when 16#00185# => romdata <= X"0B0B80EA";
    when 16#00186# => romdata <= X"B8520B0B";
    when 16#00187# => romdata <= X"80EACC51";
    when 16#00188# => romdata <= X"88D13FA9";
    when 16#00189# => romdata <= X"F3530B0B";
    when 16#0018A# => romdata <= X"80EAD052";
    when 16#0018B# => romdata <= X"0B0B80EA";
    when 16#0018C# => romdata <= X"F85188BF";
    when 16#0018D# => romdata <= X"3FB4AE53";
    when 16#0018E# => romdata <= X"0B0B80EB";
    when 16#0018F# => romdata <= X"80520B0B";
    when 16#00190# => romdata <= X"80EB9051";
    when 16#00191# => romdata <= X"88AD3F92";
    when 16#00192# => romdata <= X"C7530B0B";
    when 16#00193# => romdata <= X"80EB9452";
    when 16#00194# => romdata <= X"0B0B80EB";
    when 16#00195# => romdata <= X"AC51889B";
    when 16#00196# => romdata <= X"3FAAAD53";
    when 16#00197# => romdata <= X"0B0B80EB";
    when 16#00198# => romdata <= X"B4520B0B";
    when 16#00199# => romdata <= X"80EBC051";
    when 16#0019A# => romdata <= X"88893FAB";
    when 16#0019B# => romdata <= X"DC530B0B";
    when 16#0019C# => romdata <= X"80EBC452";
    when 16#0019D# => romdata <= X"0B0B80EB";
    when 16#0019E# => romdata <= X"EC5187F7";
    when 16#0019F# => romdata <= X"3FAAAD53";
    when 16#001A0# => romdata <= X"0B0B80EB";
    when 16#001A1# => romdata <= X"F4520B0B";
    when 16#001A2# => romdata <= X"80EC9451";
    when 16#001A3# => romdata <= X"87E53FAC";
    when 16#001A4# => romdata <= X"A2530B0B";
    when 16#001A5# => romdata <= X"80EC9852";
    when 16#001A6# => romdata <= X"0B0B80EC";
    when 16#001A7# => romdata <= X"A85187D3";
    when 16#001A8# => romdata <= X"3F90C053";
    when 16#001A9# => romdata <= X"0B0B80F6";
    when 16#001AA# => romdata <= X"D8520B0B";
    when 16#001AB# => romdata <= X"80E69051";
    when 16#001AC# => romdata <= X"87C13F8E";
    when 16#001AD# => romdata <= X"A53F8898";
    when 16#001AE# => romdata <= X"3F810B81";
    when 16#001AF# => romdata <= X"A4B43481";
    when 16#001B0# => romdata <= X"8CC43370";
    when 16#001B1# => romdata <= X"81FF0655";
    when 16#001B2# => romdata <= X"557381EA";
    when 16#001B3# => romdata <= X"38B58F3F";
    when 16#001B4# => romdata <= X"B00881D3";
    when 16#001B5# => romdata <= X"3888873F";
    when 16#001B6# => romdata <= X"80FCE808";
    when 16#001B7# => romdata <= X"70087084";
    when 16#001B8# => romdata <= X"2A810651";
    when 16#001B9# => romdata <= X"55567380";
    when 16#001BA# => romdata <= X"2E80F238";
    when 16#001BB# => romdata <= X"F881C08E";
    when 16#001BC# => romdata <= X"8055818C";
    when 16#001BD# => romdata <= X"C008802E";
    when 16#001BE# => romdata <= X"81833874";
    when 16#001BF# => romdata <= X"81FF0684";
    when 16#001C0# => romdata <= X"170C80FC";
    when 16#001C1# => romdata <= X"BC337081";
    when 16#001C2# => romdata <= X"FF065154";
    when 16#001C3# => romdata <= X"73802E80";
    when 16#001C4# => romdata <= X"C138749F";
    when 16#001C5# => romdata <= X"2A751007";
    when 16#001C6# => romdata <= X"55818CC4";
    when 16#001C7# => romdata <= X"337081FF";
    when 16#001C8# => romdata <= X"06515473";
    when 16#001C9# => romdata <= X"802ED438";
    when 16#001CA# => romdata <= X"800B818C";
    when 16#001CB# => romdata <= X"C4348ECA";
    when 16#001CC# => romdata <= X"3F80FCB8";
    when 16#001CD# => romdata <= X"335675A5";
    when 16#001CE# => romdata <= X"3880FCE8";
    when 16#001CF# => romdata <= X"087581FF";
    when 16#001D0# => romdata <= X"0684120C";
    when 16#001D1# => romdata <= X"80FCBC33";
    when 16#001D2# => romdata <= X"7081FF06";
    when 16#001D3# => romdata <= X"51555673";
    when 16#001D4# => romdata <= X"C1387481";
    when 16#001D5# => romdata <= X"2A759F2B";
    when 16#001D6# => romdata <= X"0755FFBD";
    when 16#001D7# => romdata <= X"3981A4B4";
    when 16#001D8# => romdata <= X"335574FE";
    when 16#001D9# => romdata <= X"DA38873D";
    when 16#001DA# => romdata <= X"0D047481";
    when 16#001DB# => romdata <= X"2A759F2B";
    when 16#001DC# => romdata <= X"075580FD";
    when 16#001DD# => romdata <= X"51B3853F";
    when 16#001DE# => romdata <= X"80FCE808";
    when 16#001DF# => romdata <= X"567481FF";
    when 16#001E0# => romdata <= X"0684170C";
    when 16#001E1# => romdata <= X"80FCBC33";
    when 16#001E2# => romdata <= X"7081FF06";
    when 16#001E3# => romdata <= X"57547580";
    when 16#001E4# => romdata <= X"2ED83874";
    when 16#001E5# => romdata <= X"9F2A7510";
    when 16#001E6# => romdata <= X"075580FD";
    when 16#001E7# => romdata <= X"51B2DD3F";
    when 16#001E8# => romdata <= X"80FCE808";
    when 16#001E9# => romdata <= X"56D739B3";
    when 16#001EA# => romdata <= X"C83FB008";
    when 16#001EB# => romdata <= X"81FF0651";
    when 16#001EC# => romdata <= X"879A3FFE";
    when 16#001ED# => romdata <= X"A039800B";
    when 16#001EE# => romdata <= X"818CC434";
    when 16#001EF# => romdata <= X"8DBC3FB3";
    when 16#001F0# => romdata <= X"9D3FB008";
    when 16#001F1# => romdata <= X"802EFE8D";
    when 16#001F2# => romdata <= X"38DD3980";
    when 16#001F3# => romdata <= X"3D0D0B0B";
    when 16#001F4# => romdata <= X"80ECB051";
    when 16#001F5# => romdata <= X"AEBF3F8C";
    when 16#001F6# => romdata <= X"51AEA03F";
    when 16#001F7# => romdata <= X"0B0B80EC";
    when 16#001F8# => romdata <= X"B451AEB1";
    when 16#001F9# => romdata <= X"3F818CC0";
    when 16#001FA# => romdata <= X"08802E8E";
    when 16#001FB# => romdata <= X"380B0B80";
    when 16#001FC# => romdata <= X"ECCC51AE";
    when 16#001FD# => romdata <= X"A03F823D";
    when 16#001FE# => romdata <= X"0D040B0B";
    when 16#001FF# => romdata <= X"80ECD851";
    when 16#00200# => romdata <= X"AE933F81";
    when 16#00201# => romdata <= X"0A51AE8D";
    when 16#00202# => romdata <= X"3F0B0B80";
    when 16#00203# => romdata <= X"ECEC51AE";
    when 16#00204# => romdata <= X"843F0B0B";
    when 16#00205# => romdata <= X"80ED9451";
    when 16#00206# => romdata <= X"ADFB3F80";
    when 16#00207# => romdata <= X"E451AFBF";
    when 16#00208# => romdata <= X"3F0B0B80";
    when 16#00209# => romdata <= X"EDA851AD";
    when 16#0020A# => romdata <= X"EC3F0B0B";
    when 16#0020B# => romdata <= X"80EDB051";
    when 16#0020C# => romdata <= X"ADE33F0B";
    when 16#0020D# => romdata <= X"0B80EDBC";
    when 16#0020E# => romdata <= X"51ADDA3F";
    when 16#0020F# => romdata <= X"823D0D04";
    when 16#00210# => romdata <= X"FF893F8B";
    when 16#00211# => romdata <= X"953F800B";
    when 16#00212# => romdata <= X"B00C04FE";
    when 16#00213# => romdata <= X"3D0D80FC";
    when 16#00214# => romdata <= X"EC089811";
    when 16#00215# => romdata <= X"0870842A";
    when 16#00216# => romdata <= X"70810651";
    when 16#00217# => romdata <= X"53535370";
    when 16#00218# => romdata <= X"802E8D38";
    when 16#00219# => romdata <= X"71EF0698";
    when 16#0021A# => romdata <= X"140C810B";
    when 16#0021B# => romdata <= X"818CC434";
    when 16#0021C# => romdata <= X"843D0D04";
    when 16#0021D# => romdata <= X"803D0D0B";
    when 16#0021E# => romdata <= X"0B80EDC4";
    when 16#0021F# => romdata <= X"51AD963F";
    when 16#00220# => romdata <= X"8A51ACF7";
    when 16#00221# => romdata <= X"3F800BB0";
    when 16#00222# => romdata <= X"0C823D0D";
    when 16#00223# => romdata <= X"04F93D0D";
    when 16#00224# => romdata <= X"81518994";
    when 16#00225# => romdata <= X"3FB00855";
    when 16#00226# => romdata <= X"8251898C";
    when 16#00227# => romdata <= X"3F74B008";
    when 16#00228# => romdata <= X"075399CC";
    when 16#00229# => romdata <= X"57FCE297";
    when 16#0022A# => romdata <= X"F6805872";
    when 16#0022B# => romdata <= X"802E9038";
    when 16#0022C# => romdata <= X"74755457";
    when 16#0022D# => romdata <= X"80548077";
    when 16#0022E# => romdata <= X"0774B008";
    when 16#0022F# => romdata <= X"07595776";
    when 16#00230# => romdata <= X"5177529B";
    when 16#00231# => romdata <= X"FA3F72B0";
    when 16#00232# => romdata <= X"0C893D0D";
    when 16#00233# => romdata <= X"04FB3D0D";
    when 16#00234# => romdata <= X"815187A2";
    when 16#00235# => romdata <= X"3FB00856";
    when 16#00236# => romdata <= X"81538252";
    when 16#00237# => romdata <= X"8051A5A8";
    when 16#00238# => romdata <= X"3F80FCC8";
    when 16#00239# => romdata <= X"08558975";
    when 16#0023A# => romdata <= X"0C80FCE8";
    when 16#0023B# => romdata <= X"08841108";
    when 16#0023C# => romdata <= X"70810A07";
    when 16#0023D# => romdata <= X"84130C55";
    when 16#0023E# => romdata <= X"557551AF";
    when 16#0023F# => romdata <= X"D93F80FC";
    when 16#00240# => romdata <= X"E8088411";
    when 16#00241# => romdata <= X"0870FE0A";
    when 16#00242# => romdata <= X"0684130C";
    when 16#00243# => romdata <= X"55558153";
    when 16#00244# => romdata <= X"82528051";
    when 16#00245# => romdata <= X"A4F23F80";
    when 16#00246# => romdata <= X"FCC80855";
    when 16#00247# => romdata <= X"89750C80";
    when 16#00248# => romdata <= X"FCE80884";
    when 16#00249# => romdata <= X"11087081";
    when 16#0024A# => romdata <= X"0A078413";
    when 16#0024B# => romdata <= X"0C555575";
    when 16#0024C# => romdata <= X"51AFA33F";
    when 16#0024D# => romdata <= X"80FCE808";
    when 16#0024E# => romdata <= X"84110870";
    when 16#0024F# => romdata <= X"FE0A0684";
    when 16#00250# => romdata <= X"130C5555";
    when 16#00251# => romdata <= X"FF9239FE";
    when 16#00252# => romdata <= X"3D0D8151";
    when 16#00253# => romdata <= X"86A83F80";
    when 16#00254# => romdata <= X"FCE80884";
    when 16#00255# => romdata <= X"11087081";
    when 16#00256# => romdata <= X"0A078413";
    when 16#00257# => romdata <= X"0C5353B0";
    when 16#00258# => romdata <= X"0851AEF2";
    when 16#00259# => romdata <= X"3F80FCE8";
    when 16#0025A# => romdata <= X"08841108";
    when 16#0025B# => romdata <= X"70FE0A06";
    when 16#0025C# => romdata <= X"7084140C";
    when 16#0025D# => romdata <= X"B00C5353";
    when 16#0025E# => romdata <= X"843D0D04";
    when 16#0025F# => romdata <= X"FC3D0D80";
    when 16#00260# => romdata <= X"FCE80870";
    when 16#00261# => romdata <= X"08810A06";
    when 16#00262# => romdata <= X"818CC00C";
    when 16#00263# => romdata <= X"54AF913F";
    when 16#00264# => romdata <= X"AFB53F8A";
    when 16#00265# => romdata <= X"C53F938C";
    when 16#00266# => romdata <= X"3F80FCEC";
    when 16#00267# => romdata <= X"08981108";
    when 16#00268# => romdata <= X"70880798";
    when 16#00269# => romdata <= X"130C5555";
    when 16#0026A# => romdata <= X"818CC008";
    when 16#0026B# => romdata <= X"80D53888";
    when 16#0026C# => romdata <= X"800B81A5";
    when 16#0026D# => romdata <= X"900CFC93";
    when 16#0026E# => romdata <= X"3F818CC0";
    when 16#0026F# => romdata <= X"08802E80";
    when 16#00270# => romdata <= X"D3388153";
    when 16#00271# => romdata <= X"82528051";
    when 16#00272# => romdata <= X"A3BE3F80";
    when 16#00273# => romdata <= X"FCC80855";
    when 16#00274# => romdata <= X"89750C80";
    when 16#00275# => romdata <= X"FCE80884";
    when 16#00276# => romdata <= X"11087081";
    when 16#00277# => romdata <= X"0A078413";
    when 16#00278# => romdata <= X"0C555580";
    when 16#00279# => romdata <= X"51ADEF3F";
    when 16#0027A# => romdata <= X"80FCE808";
    when 16#0027B# => romdata <= X"84110870";
    when 16#0027C# => romdata <= X"FE0A0684";
    when 16#0027D# => romdata <= X"130C5555";
    when 16#0027E# => romdata <= X"80FCC808";
    when 16#0027F# => romdata <= X"5580750C";
    when 16#00280# => romdata <= X"B0AB3FBD";
    when 16#00281# => romdata <= X"E50B81A5";
    when 16#00282# => romdata <= X"900CFBBF";
    when 16#00283# => romdata <= X"3F818CC0";
    when 16#00284# => romdata <= X"08FFAF38";
    when 16#00285# => romdata <= X"80C3930B";
    when 16#00286# => romdata <= X"81A5900C";
    when 16#00287# => romdata <= X"F5B63F81";
    when 16#00288# => romdata <= X"53825280";
    when 16#00289# => romdata <= X"51A2E13F";
    when 16#0028A# => romdata <= X"80FCC808";
    when 16#0028B# => romdata <= X"5589750C";
    when 16#0028C# => romdata <= X"80FCE808";
    when 16#0028D# => romdata <= X"84110870";
    when 16#0028E# => romdata <= X"810A0784";
    when 16#0028F# => romdata <= X"130C5555";
    when 16#00290# => romdata <= X"8051AD92";
    when 16#00291# => romdata <= X"3F80FCE8";
    when 16#00292# => romdata <= X"08841108";
    when 16#00293# => romdata <= X"70FE0A06";
    when 16#00294# => romdata <= X"84130C55";
    when 16#00295# => romdata <= X"5580FCC8";
    when 16#00296# => romdata <= X"08558075";
    when 16#00297# => romdata <= X"0CAFCE3F";
    when 16#00298# => romdata <= X"800B81A4";
    when 16#00299# => romdata <= X"AC34800B";
    when 16#0029A# => romdata <= X"81A4A834";
    when 16#0029B# => romdata <= X"800B81A4";
    when 16#0029C# => romdata <= X"B00C04FC";
    when 16#0029D# => romdata <= X"3D0D81A4";
    when 16#0029E# => romdata <= X"A8335372";
    when 16#0029F# => romdata <= X"A72680C5";
    when 16#002A0# => romdata <= X"38765272";
    when 16#002A1# => romdata <= X"10101073";
    when 16#002A2# => romdata <= X"1005818C";
    when 16#002A3# => romdata <= X"C80551B4";
    when 16#002A4# => romdata <= X"B73F7752";
    when 16#002A5# => romdata <= X"81A4A833";
    when 16#002A6# => romdata <= X"70902971";
    when 16#002A7# => romdata <= X"31701010";
    when 16#002A8# => romdata <= X"818FD805";
    when 16#002A9# => romdata <= X"535654B4";
    when 16#002AA# => romdata <= X"9F3F81A4";
    when 16#002AB# => romdata <= X"A8337010";
    when 16#002AC# => romdata <= X"1081A2B8";
    when 16#002AD# => romdata <= X"057A710C";
    when 16#002AE# => romdata <= X"54810553";
    when 16#002AF# => romdata <= X"7281A4A8";
    when 16#002B0# => romdata <= X"34863D0D";
    when 16#002B1# => romdata <= X"0480EDDC";
    when 16#002B2# => romdata <= X"51A8CA3F";
    when 16#002B3# => romdata <= X"863D0D04";
    when 16#002B4# => romdata <= X"803D0D80";
    when 16#002B5# => romdata <= X"EDF851A8";
    when 16#002B6# => romdata <= X"BC3F823D";
    when 16#002B7# => romdata <= X"0D04FE3D";
    when 16#002B8# => romdata <= X"0D81A4B0";
    when 16#002B9# => romdata <= X"08537285";
    when 16#002BA# => romdata <= X"38843D0D";
    when 16#002BB# => romdata <= X"04722DB0";
    when 16#002BC# => romdata <= X"0853800B";
    when 16#002BD# => romdata <= X"81A4B00C";
    when 16#002BE# => romdata <= X"B0088C38";
    when 16#002BF# => romdata <= X"80EDF851";
    when 16#002C0# => romdata <= X"A8933F84";
    when 16#002C1# => romdata <= X"3D0D0480";
    when 16#002C2# => romdata <= X"F9A851A8";
    when 16#002C3# => romdata <= X"883F7283";
    when 16#002C4# => romdata <= X"FFFF26AA";
    when 16#002C5# => romdata <= X"3881FF73";
    when 16#002C6# => romdata <= X"27963872";
    when 16#002C7# => romdata <= X"529051A8";
    when 16#002C8# => romdata <= X"973F8A51";
    when 16#002C9# => romdata <= X"A7D53F80";
    when 16#002CA# => romdata <= X"EDF851A7";
    when 16#002CB# => romdata <= X"E83FD439";
    when 16#002CC# => romdata <= X"72528851";
    when 16#002CD# => romdata <= X"A8823F8A";
    when 16#002CE# => romdata <= X"51A7C03F";
    when 16#002CF# => romdata <= X"EA397252";
    when 16#002D0# => romdata <= X"A051A7F4";
    when 16#002D1# => romdata <= X"3F8A51A7";
    when 16#002D2# => romdata <= X"B23FDC39";
    when 16#002D3# => romdata <= X"FA3D0D02";
    when 16#002D4# => romdata <= X"A3053356";
    when 16#002D5# => romdata <= X"758D2E80";
    when 16#002D6# => romdata <= X"F4387588";
    when 16#002D7# => romdata <= X"32703077";
    when 16#002D8# => romdata <= X"80FF3270";
    when 16#002D9# => romdata <= X"30728025";
    when 16#002DA# => romdata <= X"71802507";
    when 16#002DB# => romdata <= X"54515658";
    when 16#002DC# => romdata <= X"55749538";
    when 16#002DD# => romdata <= X"9F76278C";
    when 16#002DE# => romdata <= X"3881A4AC";
    when 16#002DF# => romdata <= X"335580CE";
    when 16#002E0# => romdata <= X"7527AE38";
    when 16#002E1# => romdata <= X"883D0D04";
    when 16#002E2# => romdata <= X"81A4AC33";
    when 16#002E3# => romdata <= X"5675802E";
    when 16#002E4# => romdata <= X"F3388851";
    when 16#002E5# => romdata <= X"A6E53FA0";
    when 16#002E6# => romdata <= X"51A6E03F";
    when 16#002E7# => romdata <= X"8851A6DB";
    when 16#002E8# => romdata <= X"3F81A4AC";
    when 16#002E9# => romdata <= X"33FF0557";
    when 16#002EA# => romdata <= X"7681A4AC";
    when 16#002EB# => romdata <= X"34883D0D";
    when 16#002EC# => romdata <= X"047551A6";
    when 16#002ED# => romdata <= X"C63F81A4";
    when 16#002EE# => romdata <= X"AC338111";
    when 16#002EF# => romdata <= X"55577381";
    when 16#002F0# => romdata <= X"A4AC3475";
    when 16#002F1# => romdata <= X"81A3D818";
    when 16#002F2# => romdata <= X"34883D0D";
    when 16#002F3# => romdata <= X"048A51A6";
    when 16#002F4# => romdata <= X"AA3F81A4";
    when 16#002F5# => romdata <= X"AC338111";
    when 16#002F6# => romdata <= X"56547481";
    when 16#002F7# => romdata <= X"A4AC3480";
    when 16#002F8# => romdata <= X"0B81A3D8";
    when 16#002F9# => romdata <= X"15348056";
    when 16#002FA# => romdata <= X"800B81A3";
    when 16#002FB# => romdata <= X"D8173356";
    when 16#002FC# => romdata <= X"5474A02E";
    when 16#002FD# => romdata <= X"83388154";
    when 16#002FE# => romdata <= X"74802E90";
    when 16#002FF# => romdata <= X"3873802E";
    when 16#00300# => romdata <= X"8B388116";
    when 16#00301# => romdata <= X"7081FF06";
    when 16#00302# => romdata <= X"5757DD39";
    when 16#00303# => romdata <= X"75802EBF";
    when 16#00304# => romdata <= X"38800B81";
    when 16#00305# => romdata <= X"A4A83355";
    when 16#00306# => romdata <= X"55747427";
    when 16#00307# => romdata <= X"AB387357";
    when 16#00308# => romdata <= X"74101010";
    when 16#00309# => romdata <= X"75100576";
    when 16#0030A# => romdata <= X"5481A3D8";
    when 16#0030B# => romdata <= X"53818CC8";
    when 16#0030C# => romdata <= X"0551B2E0";
    when 16#0030D# => romdata <= X"3FB00880";
    when 16#0030E# => romdata <= X"2EA63881";
    when 16#0030F# => romdata <= X"157081FF";
    when 16#00310# => romdata <= X"06565476";
    when 16#00311# => romdata <= X"7526D938";
    when 16#00312# => romdata <= X"80EDFC51";
    when 16#00313# => romdata <= X"A5C73F80";
    when 16#00314# => romdata <= X"EDF851A5";
    when 16#00315# => romdata <= X"C03F800B";
    when 16#00316# => romdata <= X"81A4AC34";
    when 16#00317# => romdata <= X"883D0D04";
    when 16#00318# => romdata <= X"74101081";
    when 16#00319# => romdata <= X"A2B80570";
    when 16#0031A# => romdata <= X"0881A4B0";
    when 16#0031B# => romdata <= X"0C56800B";
    when 16#0031C# => romdata <= X"81A4AC34";
    when 16#0031D# => romdata <= X"E739F73D";
    when 16#0031E# => romdata <= X"0D02AF05";
    when 16#0031F# => romdata <= X"3359800B";
    when 16#00320# => romdata <= X"81A3D833";
    when 16#00321# => romdata <= X"81A3D859";
    when 16#00322# => romdata <= X"555673A0";
    when 16#00323# => romdata <= X"2E098106";
    when 16#00324# => romdata <= X"96388116";
    when 16#00325# => romdata <= X"7081FF06";
    when 16#00326# => romdata <= X"81A3D811";
    when 16#00327# => romdata <= X"70335359";
    when 16#00328# => romdata <= X"575473A0";
    when 16#00329# => romdata <= X"2EEC3880";
    when 16#0032A# => romdata <= X"58777927";
    when 16#0032B# => romdata <= X"80EA3880";
    when 16#0032C# => romdata <= X"77335654";
    when 16#0032D# => romdata <= X"74742E83";
    when 16#0032E# => romdata <= X"38815474";
    when 16#0032F# => romdata <= X"A02E9A38";
    when 16#00330# => romdata <= X"7380C538";
    when 16#00331# => romdata <= X"74A02E91";
    when 16#00332# => romdata <= X"38811870";
    when 16#00333# => romdata <= X"81FF0659";
    when 16#00334# => romdata <= X"55787826";
    when 16#00335# => romdata <= X"DA3880C0";
    when 16#00336# => romdata <= X"39811670";
    when 16#00337# => romdata <= X"81FF0681";
    when 16#00338# => romdata <= X"A3D81170";
    when 16#00339# => romdata <= X"33575257";
    when 16#0033A# => romdata <= X"5773A02E";
    when 16#0033B# => romdata <= X"098106D9";
    when 16#0033C# => romdata <= X"38811670";
    when 16#0033D# => romdata <= X"81FF0681";
    when 16#0033E# => romdata <= X"A3D81170";
    when 16#0033F# => romdata <= X"33575257";
    when 16#00340# => romdata <= X"5773A02E";
    when 16#00341# => romdata <= X"D438C239";
    when 16#00342# => romdata <= X"81167081";
    when 16#00343# => romdata <= X"FF0681A3";
    when 16#00344# => romdata <= X"D8115957";
    when 16#00345# => romdata <= X"55FF9839";
    when 16#00346# => romdata <= X"80538B3D";
    when 16#00347# => romdata <= X"FC055276";
    when 16#00348# => romdata <= X"51B5B63F";
    when 16#00349# => romdata <= X"8B3D0D04";
    when 16#0034A# => romdata <= X"F73D0D02";
    when 16#0034B# => romdata <= X"AF053359";
    when 16#0034C# => romdata <= X"800B81A3";
    when 16#0034D# => romdata <= X"D83381A3";
    when 16#0034E# => romdata <= X"D8595556";
    when 16#0034F# => romdata <= X"73A02E09";
    when 16#00350# => romdata <= X"81069638";
    when 16#00351# => romdata <= X"81167081";
    when 16#00352# => romdata <= X"FF0681A3";
    when 16#00353# => romdata <= X"D8117033";
    when 16#00354# => romdata <= X"53595754";
    when 16#00355# => romdata <= X"73A02EEC";
    when 16#00356# => romdata <= X"38805877";
    when 16#00357# => romdata <= X"792780EA";
    when 16#00358# => romdata <= X"38807733";
    when 16#00359# => romdata <= X"56547474";
    when 16#0035A# => romdata <= X"2E833881";
    when 16#0035B# => romdata <= X"5474A02E";
    when 16#0035C# => romdata <= X"9A387380";
    when 16#0035D# => romdata <= X"C53874A0";
    when 16#0035E# => romdata <= X"2E913881";
    when 16#0035F# => romdata <= X"187081FF";
    when 16#00360# => romdata <= X"06595578";
    when 16#00361# => romdata <= X"7826DA38";
    when 16#00362# => romdata <= X"80C03981";
    when 16#00363# => romdata <= X"167081FF";
    when 16#00364# => romdata <= X"0681A3D8";
    when 16#00365# => romdata <= X"11703357";
    when 16#00366# => romdata <= X"52575773";
    when 16#00367# => romdata <= X"A02E0981";
    when 16#00368# => romdata <= X"06D93881";
    when 16#00369# => romdata <= X"167081FF";
    when 16#0036A# => romdata <= X"0681A3D8";
    when 16#0036B# => romdata <= X"11703357";
    when 16#0036C# => romdata <= X"52575773";
    when 16#0036D# => romdata <= X"A02ED438";
    when 16#0036E# => romdata <= X"C2398116";
    when 16#0036F# => romdata <= X"7081FF06";
    when 16#00370# => romdata <= X"81A3D811";
    when 16#00371# => romdata <= X"595755FF";
    when 16#00372# => romdata <= X"98399053";
    when 16#00373# => romdata <= X"8B3DFC05";
    when 16#00374# => romdata <= X"527651B7";
    when 16#00375# => romdata <= X"A13F8B3D";
    when 16#00376# => romdata <= X"0D04FC3D";
    when 16#00377# => romdata <= X"0D8A51A2";
    when 16#00378# => romdata <= X"9A3F80EE";
    when 16#00379# => romdata <= X"9051A2AD";
    when 16#0037A# => romdata <= X"3F800B81";
    when 16#0037B# => romdata <= X"A4A83353";
    when 16#0037C# => romdata <= X"53727227";
    when 16#0037D# => romdata <= X"80F53872";
    when 16#0037E# => romdata <= X"10101073";
    when 16#0037F# => romdata <= X"1005818C";
    when 16#00380# => romdata <= X"C8057052";
    when 16#00381# => romdata <= X"54A28E3F";
    when 16#00382# => romdata <= X"72842B70";
    when 16#00383# => romdata <= X"7431822B";
    when 16#00384# => romdata <= X"818FD811";
    when 16#00385# => romdata <= X"33515355";
    when 16#00386# => romdata <= X"71802EB7";
    when 16#00387# => romdata <= X"387351AE";
    when 16#00388# => romdata <= X"943FB008";
    when 16#00389# => romdata <= X"81FF0652";
    when 16#0038A# => romdata <= X"71892693";
    when 16#0038B# => romdata <= X"38A051A1";
    when 16#0038C# => romdata <= X"CA3F8112";
    when 16#0038D# => romdata <= X"7081FF06";
    when 16#0038E# => romdata <= X"53548972";
    when 16#0038F# => romdata <= X"27EF3880";
    when 16#00390# => romdata <= X"EEA851A1";
    when 16#00391# => romdata <= X"D03F7473";
    when 16#00392# => romdata <= X"31822B81";
    when 16#00393# => romdata <= X"8FD80551";
    when 16#00394# => romdata <= X"A1C33F8A";
    when 16#00395# => romdata <= X"51A1A43F";
    when 16#00396# => romdata <= X"81137081";
    when 16#00397# => romdata <= X"FF0681A4";
    when 16#00398# => romdata <= X"A8335454";
    when 16#00399# => romdata <= X"55717326";
    when 16#0039A# => romdata <= X"FF8D388A";
    when 16#0039B# => romdata <= X"51A18C3F";
    when 16#0039C# => romdata <= X"81A4A833";
    when 16#0039D# => romdata <= X"B00C863D";
    when 16#0039E# => romdata <= X"0D04FE3D";
    when 16#0039F# => romdata <= X"0D81A588";
    when 16#003A0# => romdata <= X"22FF0551";
    when 16#003A1# => romdata <= X"7081A588";
    when 16#003A2# => romdata <= X"237083FF";
    when 16#003A3# => romdata <= X"FF065170";
    when 16#003A4# => romdata <= X"80C43881";
    when 16#003A5# => romdata <= X"A58C3351";
    when 16#003A6# => romdata <= X"7081FF2E";
    when 16#003A7# => romdata <= X"B9387010";
    when 16#003A8# => romdata <= X"101081A4";
    when 16#003A9# => romdata <= X"B8055271";
    when 16#003AA# => romdata <= X"3381A58C";
    when 16#003AB# => romdata <= X"34FE7234";
    when 16#003AC# => romdata <= X"81A58C33";
    when 16#003AD# => romdata <= X"70101010";
    when 16#003AE# => romdata <= X"81A4B805";
    when 16#003AF# => romdata <= X"52538211";
    when 16#003B0# => romdata <= X"2281A588";
    when 16#003B1# => romdata <= X"23841208";
    when 16#003B2# => romdata <= X"53722D81";
    when 16#003B3# => romdata <= X"A5882251";
    when 16#003B4# => romdata <= X"70802EFF";
    when 16#003B5# => romdata <= X"BE38843D";
    when 16#003B6# => romdata <= X"0D04FF3D";
    when 16#003B7# => romdata <= X"0D8A5271";
    when 16#003B8# => romdata <= X"10101081";
    when 16#003B9# => romdata <= X"A4B00551";
    when 16#003BA# => romdata <= X"FE7134FF";
    when 16#003BB# => romdata <= X"127081FF";
    when 16#003BC# => romdata <= X"06535171";
    when 16#003BD# => romdata <= X"EA38FF0B";
    when 16#003BE# => romdata <= X"81A58C34";
    when 16#003BF# => romdata <= X"833D0D04";
    when 16#003C0# => romdata <= X"FE3D0D02";
    when 16#003C1# => romdata <= X"93053302";
    when 16#003C2# => romdata <= X"84059705";
    when 16#003C3# => romdata <= X"33545271";
    when 16#003C4# => romdata <= X"842E80D1";
    when 16#003C5# => romdata <= X"38718424";
    when 16#003C6# => romdata <= X"91387181";
    when 16#003C7# => romdata <= X"2EAC3880";
    when 16#003C8# => romdata <= X"EEAC519F";
    when 16#003C9# => romdata <= X"F03F843D";
    when 16#003CA# => romdata <= X"0D047180";
    when 16#003CB# => romdata <= X"D52E0981";
    when 16#003CC# => romdata <= X"06ED3880";
    when 16#003CD# => romdata <= X"EEB8519F";
    when 16#003CE# => romdata <= X"DC3F728C";
    when 16#003CF# => romdata <= X"26B33872";
    when 16#003D0# => romdata <= X"101080F3";
    when 16#003D1# => romdata <= X"AC055271";
    when 16#003D2# => romdata <= X"080480EE";
    when 16#003D3# => romdata <= X"C4519FC5";
    when 16#003D4# => romdata <= X"3FFA1352";
    when 16#003D5# => romdata <= X"7180DB26";
    when 16#003D6# => romdata <= X"98387110";
    when 16#003D7# => romdata <= X"1080F3E0";
    when 16#003D8# => romdata <= X"05527108";
    when 16#003D9# => romdata <= X"0480EED0";
    when 16#003DA# => romdata <= X"519FAA3F";
    when 16#003DB# => romdata <= X"728F2E8C";
    when 16#003DC# => romdata <= X"3880EEDC";
    when 16#003DD# => romdata <= X"519F9E3F";
    when 16#003DE# => romdata <= X"843D0D04";
    when 16#003DF# => romdata <= X"80EEEC51";
    when 16#003E0# => romdata <= X"9F933F84";
    when 16#003E1# => romdata <= X"3D0D0480";
    when 16#003E2# => romdata <= X"EF84519F";
    when 16#003E3# => romdata <= X"883F843D";
    when 16#003E4# => romdata <= X"0D0480EF";
    when 16#003E5# => romdata <= X"94519EFD";
    when 16#003E6# => romdata <= X"3F843D0D";
    when 16#003E7# => romdata <= X"0480EFAC";
    when 16#003E8# => romdata <= X"519EF23F";
    when 16#003E9# => romdata <= X"843D0D04";
    when 16#003EA# => romdata <= X"80EFBC51";
    when 16#003EB# => romdata <= X"9EE73F84";
    when 16#003EC# => romdata <= X"3D0D0480";
    when 16#003ED# => romdata <= X"EFDC519E";
    when 16#003EE# => romdata <= X"DC3F843D";
    when 16#003EF# => romdata <= X"0D0480EF";
    when 16#003F0# => romdata <= X"F8519ED1";
    when 16#003F1# => romdata <= X"3F843D0D";
    when 16#003F2# => romdata <= X"0480F094";
    when 16#003F3# => romdata <= X"519EC63F";
    when 16#003F4# => romdata <= X"843D0D04";
    when 16#003F5# => romdata <= X"80F0A851";
    when 16#003F6# => romdata <= X"9EBB3F84";
    when 16#003F7# => romdata <= X"3D0D0480";
    when 16#003F8# => romdata <= X"F0C4519E";
    when 16#003F9# => romdata <= X"B03F843D";
    when 16#003FA# => romdata <= X"0D0480F0";
    when 16#003FB# => romdata <= X"D4519EA5";
    when 16#003FC# => romdata <= X"3F843D0D";
    when 16#003FD# => romdata <= X"0480F0E4";
    when 16#003FE# => romdata <= X"519E9A3F";
    when 16#003FF# => romdata <= X"843D0D04";
    when 16#00400# => romdata <= X"80F18451";
    when 16#00401# => romdata <= X"9E8F3F84";
    when 16#00402# => romdata <= X"3D0D0480";
    when 16#00403# => romdata <= X"F198519E";
    when 16#00404# => romdata <= X"843F843D";
    when 16#00405# => romdata <= X"0D0480F1";
    when 16#00406# => romdata <= X"B4519DF9";
    when 16#00407# => romdata <= X"3F843D0D";
    when 16#00408# => romdata <= X"0480F1CC";
    when 16#00409# => romdata <= X"519DEE3F";
    when 16#0040A# => romdata <= X"843D0D04";
    when 16#0040B# => romdata <= X"80F1E051";
    when 16#0040C# => romdata <= X"9DE33F84";
    when 16#0040D# => romdata <= X"3D0D0480";
    when 16#0040E# => romdata <= X"F1F0519D";
    when 16#0040F# => romdata <= X"D83F843D";
    when 16#00410# => romdata <= X"0D0480F2";
    when 16#00411# => romdata <= X"84519DCD";
    when 16#00412# => romdata <= X"3F843D0D";
    when 16#00413# => romdata <= X"0480F294";
    when 16#00414# => romdata <= X"519DC23F";
    when 16#00415# => romdata <= X"843D0D04";
    when 16#00416# => romdata <= X"80F2AC51";
    when 16#00417# => romdata <= X"9DB73F84";
    when 16#00418# => romdata <= X"3D0D0480";
    when 16#00419# => romdata <= X"F2C0519D";
    when 16#0041A# => romdata <= X"AC3F843D";
    when 16#0041B# => romdata <= X"0D0480F2";
    when 16#0041C# => romdata <= X"D0519DA1";
    when 16#0041D# => romdata <= X"3F843D0D";
    when 16#0041E# => romdata <= X"04F73D0D";
    when 16#0041F# => romdata <= X"02B30533";
    when 16#00420# => romdata <= X"7C7008C0";
    when 16#00421# => romdata <= X"80800659";
    when 16#00422# => romdata <= X"545A8056";
    when 16#00423# => romdata <= X"75832B77";
    when 16#00424# => romdata <= X"07BFE080";
    when 16#00425# => romdata <= X"07707084";
    when 16#00426# => romdata <= X"05520871";
    when 16#00427# => romdata <= X"088C2ABF";
    when 16#00428# => romdata <= X"FE800679";
    when 16#00429# => romdata <= X"0771982A";
    when 16#0042A# => romdata <= X"728C2A9F";
    when 16#0042B# => romdata <= X"FF067385";
    when 16#0042C# => romdata <= X"2A708F06";
    when 16#0042D# => romdata <= X"759F0656";
    when 16#0042E# => romdata <= X"51585D58";
    when 16#0042F# => romdata <= X"52555874";
    when 16#00430# => romdata <= X"8D388116";
    when 16#00431# => romdata <= X"568F7627";
    when 16#00432# => romdata <= X"C3388B3D";
    when 16#00433# => romdata <= X"0D0480F2";
    when 16#00434# => romdata <= X"E8519CC1";
    when 16#00435# => romdata <= X"3F75519E";
    when 16#00436# => romdata <= X"863F8452";
    when 16#00437# => romdata <= X"B008519F";
    when 16#00438# => romdata <= X"C73F80F2";
    when 16#00439# => romdata <= X"F4519CAD";
    when 16#0043A# => romdata <= X"3F745288";
    when 16#0043B# => romdata <= X"519CC93F";
    when 16#0043C# => romdata <= X"8452B008";
    when 16#0043D# => romdata <= X"519FB13F";
    when 16#0043E# => romdata <= X"80F2FC51";
    when 16#0043F# => romdata <= X"9C973F78";
    when 16#00440# => romdata <= X"5290519C";
    when 16#00441# => romdata <= X"B33F8652";
    when 16#00442# => romdata <= X"B008519F";
    when 16#00443# => romdata <= X"9B3F80F3";
    when 16#00444# => romdata <= X"84519C81";
    when 16#00445# => romdata <= X"3F72519D";
    when 16#00446# => romdata <= X"C63F8452";
    when 16#00447# => romdata <= X"B008519F";
    when 16#00448# => romdata <= X"873F80F3";
    when 16#00449# => romdata <= X"8C519BED";
    when 16#0044A# => romdata <= X"3F73519D";
    when 16#0044B# => romdata <= X"B23F8452";
    when 16#0044C# => romdata <= X"B008519E";
    when 16#0044D# => romdata <= X"F33F80F3";
    when 16#0044E# => romdata <= X"94519BD9";
    when 16#0044F# => romdata <= X"3F7752A0";
    when 16#00450# => romdata <= X"519BF53F";
    when 16#00451# => romdata <= X"8A52B008";
    when 16#00452# => romdata <= X"519EDD3F";
    when 16#00453# => romdata <= X"7992388A";
    when 16#00454# => romdata <= X"519BA83F";
    when 16#00455# => romdata <= X"8116568F";
    when 16#00456# => romdata <= X"7627FEB0";
    when 16#00457# => romdata <= X"38FEEB39";
    when 16#00458# => romdata <= X"7881FF06";
    when 16#00459# => romdata <= X"527451FB";
    when 16#0045A# => romdata <= X"973F8A51";
    when 16#0045B# => romdata <= X"9B8D3FE4";
    when 16#0045C# => romdata <= X"39F83D0D";
    when 16#0045D# => romdata <= X"02AB0533";
    when 16#0045E# => romdata <= X"59805675";
    when 16#0045F# => romdata <= X"852BE090";
    when 16#00460# => romdata <= X"11E08012";
    when 16#00461# => romdata <= X"0870982A";
    when 16#00462# => romdata <= X"718C2A9F";
    when 16#00463# => romdata <= X"FF067285";
    when 16#00464# => romdata <= X"2A708F06";
    when 16#00465# => romdata <= X"749F0655";
    when 16#00466# => romdata <= X"51585B53";
    when 16#00467# => romdata <= X"56595574";
    when 16#00468# => romdata <= X"802E81A1";
    when 16#00469# => romdata <= X"3875BF26";
    when 16#0046A# => romdata <= X"81A93880";
    when 16#0046B# => romdata <= X"F39C519A";
    when 16#0046C# => romdata <= X"E43F7551";
    when 16#0046D# => romdata <= X"9CA93F86";
    when 16#0046E# => romdata <= X"52B00851";
    when 16#0046F# => romdata <= X"9DEA3F80";
    when 16#00470# => romdata <= X"F2F4519A";
    when 16#00471# => romdata <= X"D03F7452";
    when 16#00472# => romdata <= X"88519AEC";
    when 16#00473# => romdata <= X"3F8452B0";
    when 16#00474# => romdata <= X"08519DD4";
    when 16#00475# => romdata <= X"3F80F2FC";
    when 16#00476# => romdata <= X"519ABA3F";
    when 16#00477# => romdata <= X"76529051";
    when 16#00478# => romdata <= X"9AD63F86";
    when 16#00479# => romdata <= X"52B00851";
    when 16#0047A# => romdata <= X"9DBE3F80";
    when 16#0047B# => romdata <= X"F384519A";
    when 16#0047C# => romdata <= X"A43F7251";
    when 16#0047D# => romdata <= X"9BE93F84";
    when 16#0047E# => romdata <= X"52B00851";
    when 16#0047F# => romdata <= X"9DAA3F80";
    when 16#00480# => romdata <= X"F38C519A";
    when 16#00481# => romdata <= X"903F7351";
    when 16#00482# => romdata <= X"9BD53F84";
    when 16#00483# => romdata <= X"52B00851";
    when 16#00484# => romdata <= X"9D963F80";
    when 16#00485# => romdata <= X"F3945199";
    when 16#00486# => romdata <= X"FC3F7708";
    when 16#00487# => romdata <= X"C0808006";
    when 16#00488# => romdata <= X"52A0519A";
    when 16#00489# => romdata <= X"933F8A52";
    when 16#0048A# => romdata <= X"B008519C";
    when 16#0048B# => romdata <= X"FB3F7881";
    when 16#0048C# => romdata <= X"AC388A51";
    when 16#0048D# => romdata <= X"99C53F80";
    when 16#0048E# => romdata <= X"5374812E";
    when 16#0048F# => romdata <= X"81D93876";
    when 16#00490# => romdata <= X"862E81B5";
    when 16#00491# => romdata <= X"38811656";
    when 16#00492# => romdata <= X"80FF7627";
    when 16#00493# => romdata <= X"FEAD388A";
    when 16#00494# => romdata <= X"3D0D0480";
    when 16#00495# => romdata <= X"F3A45199";
    when 16#00496# => romdata <= X"BC3FC016";
    when 16#00497# => romdata <= X"519B803F";
    when 16#00498# => romdata <= X"8652B008";
    when 16#00499# => romdata <= X"519CC13F";
    when 16#0049A# => romdata <= X"80F2F451";
    when 16#0049B# => romdata <= X"99A73F74";
    when 16#0049C# => romdata <= X"52885199";
    when 16#0049D# => romdata <= X"C33F8452";
    when 16#0049E# => romdata <= X"B008519C";
    when 16#0049F# => romdata <= X"AB3F80F2";
    when 16#004A0# => romdata <= X"FC519991";
    when 16#004A1# => romdata <= X"3F765290";
    when 16#004A2# => romdata <= X"5199AD3F";
    when 16#004A3# => romdata <= X"8652B008";
    when 16#004A4# => romdata <= X"519C953F";
    when 16#004A5# => romdata <= X"80F38451";
    when 16#004A6# => romdata <= X"98FB3F72";
    when 16#004A7# => romdata <= X"519AC03F";
    when 16#004A8# => romdata <= X"8452B008";
    when 16#004A9# => romdata <= X"519C813F";
    when 16#004AA# => romdata <= X"80F38C51";
    when 16#004AB# => romdata <= X"98E73F73";
    when 16#004AC# => romdata <= X"519AAC3F";
    when 16#004AD# => romdata <= X"8452B008";
    when 16#004AE# => romdata <= X"519BED3F";
    when 16#004AF# => romdata <= X"80F39451";
    when 16#004B0# => romdata <= X"98D33F77";
    when 16#004B1# => romdata <= X"08C08080";
    when 16#004B2# => romdata <= X"0652A051";
    when 16#004B3# => romdata <= X"98EA3F8A";
    when 16#004B4# => romdata <= X"52B00851";
    when 16#004B5# => romdata <= X"9BD23F78";
    when 16#004B6# => romdata <= X"802EFED6";
    when 16#004B7# => romdata <= X"387681FF";
    when 16#004B8# => romdata <= X"06527451";
    when 16#004B9# => romdata <= X"F89A3F8A";
    when 16#004BA# => romdata <= X"5198903F";
    when 16#004BB# => romdata <= X"80537481";
    when 16#004BC# => romdata <= X"2E098106";
    when 16#004BD# => romdata <= X"FEC9389F";
    when 16#004BE# => romdata <= X"39728106";
    when 16#004BF# => romdata <= X"5776802E";
    when 16#004C0# => romdata <= X"FEC33878";
    when 16#004C1# => romdata <= X"527751FA";
    when 16#004C2# => romdata <= X"F03F8116";
    when 16#004C3# => romdata <= X"5680FF76";
    when 16#004C4# => romdata <= X"27FCE838";
    when 16#004C5# => romdata <= X"FEB93974";
    when 16#004C6# => romdata <= X"5376862E";
    when 16#004C7# => romdata <= X"098106FE";
    when 16#004C8# => romdata <= X"A438D639";
    when 16#004C9# => romdata <= X"803D0D80";
    when 16#004CA# => romdata <= X"FCE40851";
    when 16#004CB# => romdata <= X"B1710C81";
    when 16#004CC# => romdata <= X"800B8412";
    when 16#004CD# => romdata <= X"0C823D0D";
    when 16#004CE# => romdata <= X"04FE3D0D";
    when 16#004CF# => romdata <= X"74028405";
    when 16#004D0# => romdata <= X"97053302";
    when 16#004D1# => romdata <= X"88059B05";
    when 16#004D2# => romdata <= X"3388130C";
    when 16#004D3# => romdata <= X"8C120C53";
    when 16#004D4# => romdata <= X"8C130870";
    when 16#004D5# => romdata <= X"812A8106";
    when 16#004D6# => romdata <= X"515271F4";
    when 16#004D7# => romdata <= X"388C1308";
    when 16#004D8# => romdata <= X"7081FF06";
    when 16#004D9# => romdata <= X"B00C5184";
    when 16#004DA# => romdata <= X"3D0D04FB";
    when 16#004DB# => romdata <= X"3D0D800B";
    when 16#004DC# => romdata <= X"80F6D052";
    when 16#004DD# => romdata <= X"56979E3F";
    when 16#004DE# => romdata <= X"75557410";
    when 16#004DF# => romdata <= X"5381D052";
    when 16#004E0# => romdata <= X"80FCE408";
    when 16#004E1# => romdata <= X"51FFB23F";
    when 16#004E2# => romdata <= X"B008872A";
    when 16#004E3# => romdata <= X"70810651";
    when 16#004E4# => romdata <= X"5473802E";
    when 16#004E5# => romdata <= X"99388115";
    when 16#004E6# => romdata <= X"7081FF06";
    when 16#004E7# => romdata <= X"70982B52";
    when 16#004E8# => romdata <= X"56547380";
    when 16#004E9# => romdata <= X"25D43875";
    when 16#004EA# => romdata <= X"B00C873D";
    when 16#004EB# => romdata <= X"0D0480F6";
    when 16#004EC# => romdata <= X"DC5196E1";
    when 16#004ED# => romdata <= X"3F745288";
    when 16#004EE# => romdata <= X"5196FD3F";
    when 16#004EF# => romdata <= X"80F6E851";
    when 16#004F0# => romdata <= X"96D33F81";
    when 16#004F1# => romdata <= X"167083FF";
    when 16#004F2# => romdata <= X"FF068117";
    when 16#004F3# => romdata <= X"7081FF06";
    when 16#004F4# => romdata <= X"70982B52";
    when 16#004F5# => romdata <= X"58525754";
    when 16#004F6# => romdata <= X"738025FF";
    when 16#004F7# => romdata <= X"9D38C839";
    when 16#004F8# => romdata <= X"F33D0D7F";
    when 16#004F9# => romdata <= X"02840580";
    when 16#004FA# => romdata <= X"C3053302";
    when 16#004FB# => romdata <= X"880580C6";
    when 16#004FC# => romdata <= X"052280F6";
    when 16#004FD# => romdata <= X"F8545B55";
    when 16#004FE# => romdata <= X"58969A3F";
    when 16#004FF# => romdata <= X"785197DF";
    when 16#00500# => romdata <= X"3F80F784";
    when 16#00501# => romdata <= X"51968E3F";
    when 16#00502# => romdata <= X"73528851";
    when 16#00503# => romdata <= X"96AA3F80";
    when 16#00504# => romdata <= X"ECB05196";
    when 16#00505# => romdata <= X"803F8057";
    when 16#00506# => romdata <= X"76792781";
    when 16#00507# => romdata <= X"91387310";
    when 16#00508# => romdata <= X"8E3D5C5A";
    when 16#00509# => romdata <= X"79538190";
    when 16#0050A# => romdata <= X"527751FE";
    when 16#0050B# => romdata <= X"8C3F7688";
    when 16#0050C# => romdata <= X"2A539052";
    when 16#0050D# => romdata <= X"7751FE81";
    when 16#0050E# => romdata <= X"3F7681FF";
    when 16#0050F# => romdata <= X"06539052";
    when 16#00510# => romdata <= X"7751FDF5";
    when 16#00511# => romdata <= X"3F811A53";
    when 16#00512# => romdata <= X"81905277";
    when 16#00513# => romdata <= X"51FDEA3F";
    when 16#00514# => romdata <= X"805380E0";
    when 16#00515# => romdata <= X"527751FD";
    when 16#00516# => romdata <= X"E03FB008";
    when 16#00517# => romdata <= X"872A8106";
    when 16#00518# => romdata <= X"54738A38";
    when 16#00519# => romdata <= X"88180870";
    when 16#0051A# => romdata <= X"81FF065D";
    when 16#0051B# => romdata <= X"567B81FF";
    when 16#0051C# => romdata <= X"0680F9A8";
    when 16#0051D# => romdata <= X"5256959D";
    when 16#0051E# => romdata <= X"3F755288";
    when 16#0051F# => romdata <= X"5195B93F";
    when 16#00520# => romdata <= X"80EED851";
    when 16#00521# => romdata <= X"958F3FE0";
    when 16#00522# => romdata <= X"165480DF";
    when 16#00523# => romdata <= X"7427B638";
    when 16#00524# => romdata <= X"76870670";
    when 16#00525# => romdata <= X"1C5755A0";
    when 16#00526# => romdata <= X"76347487";
    when 16#00527# => romdata <= X"2EB93881";
    when 16#00528# => romdata <= X"177083FF";
    when 16#00529# => romdata <= X"FF065855";
    when 16#0052A# => romdata <= X"787726FE";
    when 16#0052B# => romdata <= X"F73880E0";
    when 16#0052C# => romdata <= X"0B8C190C";
    when 16#0052D# => romdata <= X"8C180870";
    when 16#0052E# => romdata <= X"812A8106";
    when 16#0052F# => romdata <= X"585A76F4";
    when 16#00530# => romdata <= X"388F3D0D";
    when 16#00531# => romdata <= X"04768706";
    when 16#00532# => romdata <= X"701C5555";
    when 16#00533# => romdata <= X"75743474";
    when 16#00534# => romdata <= X"872E0981";
    when 16#00535# => romdata <= X"06C9387A";
    when 16#00536# => romdata <= X"5194BA3F";
    when 16#00537# => romdata <= X"8A51949B";
    when 16#00538# => romdata <= X"3F811770";
    when 16#00539# => romdata <= X"83FFFF06";
    when 16#0053A# => romdata <= X"58557877";
    when 16#0053B# => romdata <= X"26FEB538";
    when 16#0053C# => romdata <= X"FFBC39FB";
    when 16#0053D# => romdata <= X"3D0D8151";
    when 16#0053E# => romdata <= X"EEFC3F82";
    when 16#0053F# => romdata <= X"51F0A93F";
    when 16#00540# => romdata <= X"B00881FF";
    when 16#00541# => romdata <= X"06568351";
    when 16#00542# => romdata <= X"EEEC3FB0";
    when 16#00543# => romdata <= X"0883FFFF";
    when 16#00544# => romdata <= X"0680FCE4";
    when 16#00545# => romdata <= X"08565473";
    when 16#00546# => romdata <= X"84388180";
    when 16#00547# => romdata <= X"54735375";
    when 16#00548# => romdata <= X"527451FD";
    when 16#00549# => romdata <= X"BB3F73B0";
    when 16#0054A# => romdata <= X"0C873D0D";
    when 16#0054B# => romdata <= X"04FB3D0D";
    when 16#0054C# => romdata <= X"8151EFF4";
    when 16#0054D# => romdata <= X"3FB00853";
    when 16#0054E# => romdata <= X"8251EFEC";
    when 16#0054F# => romdata <= X"3FB00856";
    when 16#00550# => romdata <= X"B0088338";
    when 16#00551# => romdata <= X"905672FC";
    when 16#00552# => romdata <= X"06557581";
    when 16#00553# => romdata <= X"2E80F138";
    when 16#00554# => romdata <= X"80547376";
    when 16#00555# => romdata <= X"27AA3873";
    when 16#00556# => romdata <= X"83065372";
    when 16#00557# => romdata <= X"802EAE38";
    when 16#00558# => romdata <= X"80F9A851";
    when 16#00559# => romdata <= X"93AF3F74";
    when 16#0055A# => romdata <= X"70840556";
    when 16#0055B# => romdata <= X"0852A051";
    when 16#0055C# => romdata <= X"93C63FA0";
    when 16#0055D# => romdata <= X"5193843F";
    when 16#0055E# => romdata <= X"81145475";
    when 16#0055F# => romdata <= X"7426D838";
    when 16#00560# => romdata <= X"8A5192F7";
    when 16#00561# => romdata <= X"3F800BB0";
    when 16#00562# => romdata <= X"0C873D0D";
    when 16#00563# => romdata <= X"0480F7A0";
    when 16#00564# => romdata <= X"5193823F";
    when 16#00565# => romdata <= X"7452A051";
    when 16#00566# => romdata <= X"939E3F80";
    when 16#00567# => romdata <= X"F8E85192";
    when 16#00568# => romdata <= X"F43F80F9";
    when 16#00569# => romdata <= X"A85192ED";
    when 16#0056A# => romdata <= X"3F747084";
    when 16#0056B# => romdata <= X"05560852";
    when 16#0056C# => romdata <= X"A0519384";
    when 16#0056D# => romdata <= X"3FA05192";
    when 16#0056E# => romdata <= X"C23F8114";
    when 16#0056F# => romdata <= X"54FFBC39";
    when 16#00570# => romdata <= X"80F9A851";
    when 16#00571# => romdata <= X"92CF3F74";
    when 16#00572# => romdata <= X"0852A051";
    when 16#00573# => romdata <= X"92EA3F8A";
    when 16#00574# => romdata <= X"5192A83F";
    when 16#00575# => romdata <= X"800BB00C";
    when 16#00576# => romdata <= X"873D0D04";
    when 16#00577# => romdata <= X"FC3D0D81";
    when 16#00578# => romdata <= X"51EEC53F";
    when 16#00579# => romdata <= X"B0085282";
    when 16#0057A# => romdata <= X"51ED8B3F";
    when 16#0057B# => romdata <= X"B00881FF";
    when 16#0057C# => romdata <= X"06725653";
    when 16#0057D# => romdata <= X"83547280";
    when 16#0057E# => romdata <= X"2EA13873";
    when 16#0057F# => romdata <= X"51EEA93F";
    when 16#00580# => romdata <= X"81147081";
    when 16#00581# => romdata <= X"FF06FF15";
    when 16#00582# => romdata <= X"7081FF06";
    when 16#00583# => romdata <= X"B0087970";
    when 16#00584# => romdata <= X"84055B0C";
    when 16#00585# => romdata <= X"56525552";
    when 16#00586# => romdata <= X"72E13872";
    when 16#00587# => romdata <= X"B00C863D";
    when 16#00588# => romdata <= X"0D04803D";
    when 16#00589# => romdata <= X"0D8C5191";
    when 16#0058A# => romdata <= X"D23F800B";
    when 16#0058B# => romdata <= X"B00C823D";
    when 16#0058C# => romdata <= X"0D04803D";
    when 16#0058D# => romdata <= X"0D80FCF4";
    when 16#0058E# => romdata <= X"0851F8BB";
    when 16#0058F# => romdata <= X"9586A171";
    when 16#00590# => romdata <= X"0C810BB0";
    when 16#00591# => romdata <= X"0C823D0D";
    when 16#00592# => romdata <= X"04803D0D";
    when 16#00593# => romdata <= X"8151ECA6";
    when 16#00594# => romdata <= X"3FB00881";
    when 16#00595# => romdata <= X"FF0651F6";
    when 16#00596# => romdata <= X"983F800B";
    when 16#00597# => romdata <= X"B00C823D";
    when 16#00598# => romdata <= X"0D04FF3D";
    when 16#00599# => romdata <= X"0D80FCC0";
    when 16#0059A# => romdata <= X"08A01108";
    when 16#0059B# => romdata <= X"7080FF0A";
    when 16#0059C# => romdata <= X"06A0130C";
    when 16#0059D# => romdata <= X"5252BBC8";
    when 16#0059E# => romdata <= X"80800BA0";
    when 16#0059F# => romdata <= X"130C833D";
    when 16#005A0# => romdata <= X"0D04FF3D";
    when 16#005A1# => romdata <= X"0D028F05";
    when 16#005A2# => romdata <= X"3370982B";
    when 16#005A3# => romdata <= X"80FCC008";
    when 16#005A4# => romdata <= X"52B0120C";
    when 16#005A5# => romdata <= X"51833D0D";
    when 16#005A6# => romdata <= X"04FF3D0D";
    when 16#005A7# => romdata <= X"80FCC008";
    when 16#005A8# => romdata <= X"52A41208";
    when 16#005A9# => romdata <= X"70892A70";
    when 16#005AA# => romdata <= X"81065151";
    when 16#005AB# => romdata <= X"5170802E";
    when 16#005AC# => romdata <= X"F038B412";
    when 16#005AD# => romdata <= X"0870902A";
    when 16#005AE# => romdata <= X"B00C5183";
    when 16#005AF# => romdata <= X"3D0D04F8";
    when 16#005B0# => romdata <= X"3D0D7A7C";
    when 16#005B1# => romdata <= X"5755FF9A";
    when 16#005B2# => romdata <= X"3F80FCE8";
    when 16#005B3# => romdata <= X"08841108";
    when 16#005B4# => romdata <= X"82808007";
    when 16#005B5# => romdata <= X"84120C84";
    when 16#005B6# => romdata <= X"1108FDFF";
    when 16#005B7# => romdata <= X"FF068412";
    when 16#005B8# => romdata <= X"0C841108";
    when 16#005B9# => romdata <= X"81808007";
    when 16#005BA# => romdata <= X"84120C84";
    when 16#005BB# => romdata <= X"1108FEFF";
    when 16#005BC# => romdata <= X"FF068412";
    when 16#005BD# => romdata <= X"0C53900B";
    when 16#005BE# => romdata <= X"893D3494";
    when 16#005BF# => romdata <= X"0284059D";
    when 16#005C0# => romdata <= X"05348002";
    when 16#005C1# => romdata <= X"84059E05";
    when 16#005C2# => romdata <= X"3480E102";
    when 16#005C3# => romdata <= X"84059F05";
    when 16#005C4# => romdata <= X"34883D80";
    when 16#005C5# => romdata <= X"FCC00854";
    when 16#005C6# => romdata <= X"57A41308";
    when 16#005C7# => romdata <= X"70882A81";
    when 16#005C8# => romdata <= X"06515271";
    when 16#005C9# => romdata <= X"802EF238";
    when 16#005CA# => romdata <= X"8751FED6";
    when 16#005CB# => romdata <= X"3F800B80";
    when 16#005CC# => romdata <= X"F7AB3353";
    when 16#005CD# => romdata <= X"53727227";
    when 16#005CE# => romdata <= X"99387154";
    when 16#005CF# => romdata <= X"76137033";
    when 16#005D0# => romdata <= X"5252FEBE";
    when 16#005D1# => romdata <= X"3F811370";
    when 16#005D2# => romdata <= X"81FF0654";
    when 16#005D3# => romdata <= X"52737326";
    when 16#005D4# => romdata <= X"EB38FEC5";
    when 16#005D5# => romdata <= X"3F800B80";
    when 16#005D6# => romdata <= X"F7AB3353";
    when 16#005D7# => romdata <= X"53727227";
    when 16#005D8# => romdata <= X"93387154";
    when 16#005D9# => romdata <= X"FEB33F81";
    when 16#005DA# => romdata <= X"137081FF";
    when 16#005DB# => romdata <= X"06545273";
    when 16#005DC# => romdata <= X"7326F138";
    when 16#005DD# => romdata <= X"74882A54";
    when 16#005DE# => romdata <= X"73893D34";
    when 16#005DF# => romdata <= X"74028405";
    when 16#005E0# => romdata <= X"9D053474";
    when 16#005E1# => romdata <= X"882B7698";
    when 16#005E2# => romdata <= X"2A075271";
    when 16#005E3# => romdata <= X"0284059E";
    when 16#005E4# => romdata <= X"05347490";
    when 16#005E5# => romdata <= X"2B76902A";
    when 16#005E6# => romdata <= X"07547302";
    when 16#005E7# => romdata <= X"84059F05";
    when 16#005E8# => romdata <= X"3474982B";
    when 16#005E9# => romdata <= X"76882A07";
    when 16#005EA# => romdata <= X"53728A3D";
    when 16#005EB# => romdata <= X"34750284";
    when 16#005EC# => romdata <= X"05A10534";
    when 16#005ED# => romdata <= X"80FCC008";
    when 16#005EE# => romdata <= X"53A41308";
    when 16#005EF# => romdata <= X"70882A81";
    when 16#005F0# => romdata <= X"06565274";
    when 16#005F1# => romdata <= X"802EF238";
    when 16#005F2# => romdata <= X"8251FDB6";
    when 16#005F3# => romdata <= X"3F800B80";
    when 16#005F4# => romdata <= X"F7A63353";
    when 16#005F5# => romdata <= X"53727227";
    when 16#005F6# => romdata <= X"99387154";
    when 16#005F7# => romdata <= X"76137033";
    when 16#005F8# => romdata <= X"5256FD9E";
    when 16#005F9# => romdata <= X"3F811370";
    when 16#005FA# => romdata <= X"81FF0654";
    when 16#005FB# => romdata <= X"55737326";
    when 16#005FC# => romdata <= X"EB38FDA5";
    when 16#005FD# => romdata <= X"3F800B80";
    when 16#005FE# => romdata <= X"F7A63353";
    when 16#005FF# => romdata <= X"53727227";
    when 16#00600# => romdata <= X"93387154";
    when 16#00601# => romdata <= X"FD933F81";
    when 16#00602# => romdata <= X"137081FF";
    when 16#00603# => romdata <= X"06545273";
    when 16#00604# => romdata <= X"7326F138";
    when 16#00605# => romdata <= X"8A0B893D";
    when 16#00606# => romdata <= X"34FF8C02";
    when 16#00607# => romdata <= X"84059D05";
    when 16#00608# => romdata <= X"3480FCC0";
    when 16#00609# => romdata <= X"0853A413";
    when 16#0060A# => romdata <= X"0870882A";
    when 16#0060B# => romdata <= X"81065556";
    when 16#0060C# => romdata <= X"73802EF2";
    when 16#0060D# => romdata <= X"388851FC";
    when 16#0060E# => romdata <= X"C93F800B";
    when 16#0060F# => romdata <= X"80F7AC33";
    when 16#00610# => romdata <= X"53537272";
    when 16#00611# => romdata <= X"27993871";
    when 16#00612# => romdata <= X"54761370";
    when 16#00613# => romdata <= X"335255FC";
    when 16#00614# => romdata <= X"B13F8113";
    when 16#00615# => romdata <= X"7081FF06";
    when 16#00616# => romdata <= X"54527373";
    when 16#00617# => romdata <= X"26EB38FC";
    when 16#00618# => romdata <= X"B83F800B";
    when 16#00619# => romdata <= X"80F7AC33";
    when 16#0061A# => romdata <= X"53537272";
    when 16#0061B# => romdata <= X"27933871";
    when 16#0061C# => romdata <= X"54FCA63F";
    when 16#0061D# => romdata <= X"81137081";
    when 16#0061E# => romdata <= X"FF065456";
    when 16#0061F# => romdata <= X"737326F1";
    when 16#00620# => romdata <= X"388A0B89";
    when 16#00621# => romdata <= X"3D34FF8C";
    when 16#00622# => romdata <= X"0284059D";
    when 16#00623# => romdata <= X"053480FC";
    when 16#00624# => romdata <= X"C00853A4";
    when 16#00625# => romdata <= X"13087088";
    when 16#00626# => romdata <= X"2A810655";
    when 16#00627# => romdata <= X"5573802E";
    when 16#00628# => romdata <= X"F2388951";
    when 16#00629# => romdata <= X"FBDC3F80";
    when 16#0062A# => romdata <= X"0B80F7AD";
    when 16#0062B# => romdata <= X"33535372";
    when 16#0062C# => romdata <= X"72279938";
    when 16#0062D# => romdata <= X"71547613";
    when 16#0062E# => romdata <= X"70335252";
    when 16#0062F# => romdata <= X"FBC43F81";
    when 16#00630# => romdata <= X"137081FF";
    when 16#00631# => romdata <= X"06545673";
    when 16#00632# => romdata <= X"7326EB38";
    when 16#00633# => romdata <= X"FBCB3F80";
    when 16#00634# => romdata <= X"0B80F7AD";
    when 16#00635# => romdata <= X"33535372";
    when 16#00636# => romdata <= X"72279338";
    when 16#00637# => romdata <= X"7154FBB9";
    when 16#00638# => romdata <= X"3F811370";
    when 16#00639# => romdata <= X"81FF0654";
    when 16#0063A# => romdata <= X"57737326";
    when 16#0063B# => romdata <= X"F13880FC";
    when 16#0063C# => romdata <= X"E8088411";
    when 16#0063D# => romdata <= X"0880C080";
    when 16#0063E# => romdata <= X"0784120C";
    when 16#0063F# => romdata <= X"841108FF";
    when 16#00640# => romdata <= X"BFFF0684";
    when 16#00641# => romdata <= X"120C5480";
    when 16#00642# => romdata <= X"0BB00C8A";
    when 16#00643# => romdata <= X"3D0D04F8";
    when 16#00644# => romdata <= X"3D0D02AB";
    when 16#00645# => romdata <= X"0533893D";
    when 16#00646# => romdata <= X"80FCC008";
    when 16#00647# => romdata <= X"565856A4";
    when 16#00648# => romdata <= X"14087088";
    when 16#00649# => romdata <= X"2A810651";
    when 16#0064A# => romdata <= X"5372802E";
    when 16#0064B# => romdata <= X"F2387581";
    when 16#0064C# => romdata <= X"800751FA";
    when 16#0064D# => romdata <= X"CD3F800B";
    when 16#0064E# => romdata <= X"80F7A417";
    when 16#0064F# => romdata <= X"33545473";
    when 16#00650# => romdata <= X"73279538";
    when 16#00651# => romdata <= X"72558051";
    when 16#00652# => romdata <= X"FAB83F81";
    when 16#00653# => romdata <= X"147081FF";
    when 16#00654# => romdata <= X"06555374";
    when 16#00655# => romdata <= X"7426EF38";
    when 16#00656# => romdata <= X"FABF3F80";
    when 16#00657# => romdata <= X"0B80F7A4";
    when 16#00658# => romdata <= X"17337081";
    when 16#00659# => romdata <= X"FF065557";
    when 16#0065A# => romdata <= X"54737327";
    when 16#0065B# => romdata <= X"9A387255";
    when 16#0065C# => romdata <= X"761453FA";
    when 16#0065D# => romdata <= X"A43FB008";
    when 16#0065E# => romdata <= X"73348114";
    when 16#0065F# => romdata <= X"7081FF06";
    when 16#00660# => romdata <= X"55537474";
    when 16#00661# => romdata <= X"26EA3875";
    when 16#00662# => romdata <= X"81FF0680";
    when 16#00663# => romdata <= X"F9A85255";
    when 16#00664# => romdata <= X"8B833F80";
    when 16#00665# => romdata <= X"54737527";
    when 16#00666# => romdata <= X"99387317";
    when 16#00667# => romdata <= X"70335353";
    when 16#00668# => romdata <= X"88518B94";
    when 16#00669# => romdata <= X"3F811470";
    when 16#0066A# => romdata <= X"81FF0655";
    when 16#0066B# => romdata <= X"56747426";
    when 16#0066C# => romdata <= X"E9388A51";
    when 16#0066D# => romdata <= X"8AC53F8A";
    when 16#0066E# => romdata <= X"3D0D04FE";
    when 16#0066F# => romdata <= X"3D0D80FC";
    when 16#00670# => romdata <= X"E8088411";
    when 16#00671# => romdata <= X"08708180";
    when 16#00672# => romdata <= X"80078413";
    when 16#00673# => romdata <= X"0C548411";
    when 16#00674# => romdata <= X"0870FEFF";
    when 16#00675# => romdata <= X"FF068413";
    when 16#00676# => romdata <= X"0C5452F9";
    when 16#00677# => romdata <= X"853F80F7";
    when 16#00678# => romdata <= X"B0518AB1";
    when 16#00679# => romdata <= X"3F8751FE";
    when 16#0067A# => romdata <= X"A63F80F7";
    when 16#0067B# => romdata <= X"C0518AA5";
    when 16#0067C# => romdata <= X"3F8251FE";
    when 16#0067D# => romdata <= X"9A3F80F7";
    when 16#0067E# => romdata <= X"D0518A99";
    when 16#0067F# => romdata <= X"3F8551FE";
    when 16#00680# => romdata <= X"8E3F80F7";
    when 16#00681# => romdata <= X"E0518A8D";
    when 16#00682# => romdata <= X"3F8651FE";
    when 16#00683# => romdata <= X"823F80F7";
    when 16#00684# => romdata <= X"F0518A81";
    when 16#00685# => romdata <= X"3F8851FD";
    when 16#00686# => romdata <= X"F63F80F8";
    when 16#00687# => romdata <= X"805189F5";
    when 16#00688# => romdata <= X"3F8951FD";
    when 16#00689# => romdata <= X"EA3F800B";
    when 16#0068A# => romdata <= X"B00C843D";
    when 16#0068B# => romdata <= X"0D04FE3D";
    when 16#0068C# => romdata <= X"0D80FCE8";
    when 16#0068D# => romdata <= X"08841108";
    when 16#0068E# => romdata <= X"820A0784";
    when 16#0068F# => romdata <= X"120C7008";
    when 16#00690# => romdata <= X"70902A84";
    when 16#00691# => romdata <= X"130870FD";
    when 16#00692# => romdata <= X"0A068415";
    when 16#00693# => romdata <= X"0C5481FF";
    when 16#00694# => romdata <= X"FF06B00C";
    when 16#00695# => romdata <= X"5353843D";
    when 16#00696# => romdata <= X"0D04FF3D";
    when 16#00697# => romdata <= X"0D80FCC8";
    when 16#00698# => romdata <= X"08700870";
    when 16#00699# => romdata <= X"81FF0651";
    when 16#0069A# => romdata <= X"51527189";
    when 16#0069B# => romdata <= X"268C3871";
    when 16#0069C# => romdata <= X"101080F9";
    when 16#0069D# => romdata <= X"D0055271";
    when 16#0069E# => romdata <= X"080480F8";
    when 16#0069F# => romdata <= X"90518995";
    when 16#006A0# => romdata <= X"3F8A5188";
    when 16#006A1# => romdata <= X"F63F800B";
    when 16#006A2# => romdata <= X"B00C833D";
    when 16#006A3# => romdata <= X"0D0480E8";
    when 16#006A4# => romdata <= X"AC518981";
    when 16#006A5# => romdata <= X"3F8A5188";
    when 16#006A6# => romdata <= X"E23F800B";
    when 16#006A7# => romdata <= X"B00C833D";
    when 16#006A8# => romdata <= X"0D0480F8";
    when 16#006A9# => romdata <= X"985188ED";
    when 16#006AA# => romdata <= X"3F8A5188";
    when 16#006AB# => romdata <= X"CE3F800B";
    when 16#006AC# => romdata <= X"B00C833D";
    when 16#006AD# => romdata <= X"0D0480F8";
    when 16#006AE# => romdata <= X"A05188D9";
    when 16#006AF# => romdata <= X"3F8A5188";
    when 16#006B0# => romdata <= X"BA3F800B";
    when 16#006B1# => romdata <= X"B00C833D";
    when 16#006B2# => romdata <= X"0D0480F8";
    when 16#006B3# => romdata <= X"AC5188C5";
    when 16#006B4# => romdata <= X"3F8A5188";
    when 16#006B5# => romdata <= X"A63F800B";
    when 16#006B6# => romdata <= X"B00C833D";
    when 16#006B7# => romdata <= X"0D0480F8";
    when 16#006B8# => romdata <= X"B45188B1";
    when 16#006B9# => romdata <= X"3F8A5188";
    when 16#006BA# => romdata <= X"923F800B";
    when 16#006BB# => romdata <= X"B00C833D";
    when 16#006BC# => romdata <= X"0D0480F8";
    when 16#006BD# => romdata <= X"BC51889D";
    when 16#006BE# => romdata <= X"3F8A5187";
    when 16#006BF# => romdata <= X"FE3F800B";
    when 16#006C0# => romdata <= X"B00C833D";
    when 16#006C1# => romdata <= X"0D0480F8";
    when 16#006C2# => romdata <= X"C4518889";
    when 16#006C3# => romdata <= X"3F8A5187";
    when 16#006C4# => romdata <= X"EA3F800B";
    when 16#006C5# => romdata <= X"B00C833D";
    when 16#006C6# => romdata <= X"0D0480F8";
    when 16#006C7# => romdata <= X"CC5187F5";
    when 16#006C8# => romdata <= X"3F8A5187";
    when 16#006C9# => romdata <= X"D63F800B";
    when 16#006CA# => romdata <= X"B00C833D";
    when 16#006CB# => romdata <= X"0D0480F8";
    when 16#006CC# => romdata <= X"D45187E1";
    when 16#006CD# => romdata <= X"3F8A5187";
    when 16#006CE# => romdata <= X"C23F800B";
    when 16#006CF# => romdata <= X"B00C833D";
    when 16#006D0# => romdata <= X"0D04FE3D";
    when 16#006D1# => romdata <= X"0D80FCC8";
    when 16#006D2# => romdata <= X"08841108";
    when 16#006D3# => romdata <= X"80F8DC53";
    when 16#006D4# => romdata <= X"545287C1";
    when 16#006D5# => romdata <= X"3F72822A";
    when 16#006D6# => romdata <= X"81065189";
    when 16#006D7# => romdata <= X"823F80F8";
    when 16#006D8# => romdata <= X"EC5187B1";
    when 16#006D9# => romdata <= X"3F72812A";
    when 16#006DA# => romdata <= X"81065188";
    when 16#006DB# => romdata <= X"F23F80F9";
    when 16#006DC# => romdata <= X"805187A1";
    when 16#006DD# => romdata <= X"3F728106";
    when 16#006DE# => romdata <= X"5188E43F";
    when 16#006DF# => romdata <= X"8A5186FB";
    when 16#006E0# => romdata <= X"3F72B00C";
    when 16#006E1# => romdata <= X"843D0D04";
    when 16#006E2# => romdata <= X"FE3D0D02";
    when 16#006E3# => romdata <= X"93053302";
    when 16#006E4# => romdata <= X"84059705";
    when 16#006E5# => romdata <= X"3380FCC8";
    when 16#006E6# => romdata <= X"08555351";
    when 16#006E7# => romdata <= X"80730C76";
    when 16#006E8# => romdata <= X"88140C70";
    when 16#006E9# => romdata <= X"832B7207";
    when 16#006EA# => romdata <= X"8C140C72";
    when 16#006EB# => romdata <= X"085170FB";
    when 16#006EC# => romdata <= X"3870B00C";
    when 16#006ED# => romdata <= X"843D0D04";
    when 16#006EE# => romdata <= X"FE3D0D80";
    when 16#006EF# => romdata <= X"F9945186";
    when 16#006F0# => romdata <= X"D43F80FC";
    when 16#006F1# => romdata <= X"C808A011";
    when 16#006F2# => romdata <= X"085353A0";
    when 16#006F3# => romdata <= X"5186E93F";
    when 16#006F4# => romdata <= X"80FCC808";
    when 16#006F5# => romdata <= X"A4110853";
    when 16#006F6# => romdata <= X"53A05186";
    when 16#006F7# => romdata <= X"DB3F80F9";
    when 16#006F8# => romdata <= X"AC5186B1";
    when 16#006F9# => romdata <= X"3F80FCC8";
    when 16#006FA# => romdata <= X"08A81108";
    when 16#006FB# => romdata <= X"5353A051";
    when 16#006FC# => romdata <= X"86C63F80";
    when 16#006FD# => romdata <= X"FCC808AC";
    when 16#006FE# => romdata <= X"11085353";
    when 16#006FF# => romdata <= X"A05186B8";
    when 16#00700# => romdata <= X"3F8A5185";
    when 16#00701# => romdata <= X"F63F800B";
    when 16#00702# => romdata <= X"B00C843D";
    when 16#00703# => romdata <= X"0D04FC3D";
    when 16#00704# => romdata <= X"0D80FCC8";
    when 16#00705# => romdata <= X"089C1108";
    when 16#00706# => romdata <= X"7081FF06";
    when 16#00707# => romdata <= X"80F9C454";
    when 16#00708# => romdata <= X"57535385";
    when 16#00709# => romdata <= X"F03F7451";
    when 16#0070A# => romdata <= X"87B53F8A";
    when 16#0070B# => romdata <= X"5185CC3F";
    when 16#0070C# => romdata <= X"800BFF16";
    when 16#0070D# => romdata <= X"55537274";
    when 16#0070E# => romdata <= X"25A23872";
    when 16#0070F# => romdata <= X"101080FC";
    when 16#00710# => romdata <= X"C4080570";
    when 16#00711# => romdata <= X"08525287";
    when 16#00712# => romdata <= X"963F8A51";
    when 16#00713# => romdata <= X"85AD3F81";
    when 16#00714# => romdata <= X"137081FF";
    when 16#00715# => romdata <= X"06545273";
    when 16#00716# => romdata <= X"7324E038";
    when 16#00717# => romdata <= X"74B00C86";
    when 16#00718# => romdata <= X"3D0D04FD";
    when 16#00719# => romdata <= X"3D0D8151";
    when 16#0071A# => romdata <= X"E08C3FB0";
    when 16#0071B# => romdata <= X"0881FF06";
    when 16#0071C# => romdata <= X"528251E1";
    when 16#0071D# => romdata <= X"B33FB008";
    when 16#0071E# => romdata <= X"81FF0653";
    when 16#0071F# => romdata <= X"8351E1A8";
    when 16#00720# => romdata <= X"3F80FCC8";
    when 16#00721# => romdata <= X"08548074";
    when 16#00722# => romdata <= X"0CB00888";
    when 16#00723# => romdata <= X"150C7183";
    when 16#00724# => romdata <= X"2B73078C";
    when 16#00725# => romdata <= X"150C7308";
    when 16#00726# => romdata <= X"5271FB38";
    when 16#00727# => romdata <= X"71B00C85";
    when 16#00728# => romdata <= X"3D0D04FF";
    when 16#00729# => romdata <= X"3D0D8151";
    when 16#0072A# => romdata <= X"DFCC3F80";
    when 16#0072B# => romdata <= X"FCC808B0";
    when 16#0072C# => romdata <= X"0890120C";
    when 16#0072D# => romdata <= X"5282720C";
    when 16#0072E# => romdata <= X"833D0D04";
    when 16#0072F# => romdata <= X"803D0D80";
    when 16#00730# => romdata <= X"FCC80851";
    when 16#00731# => romdata <= X"80710C70";
    when 16#00732# => romdata <= X"B00C823D";
    when 16#00733# => romdata <= X"0D04FD3D";
    when 16#00734# => romdata <= X"0D800B80";
    when 16#00735# => romdata <= X"FCC80854";
    when 16#00736# => romdata <= X"5480730C";
    when 16#00737# => romdata <= X"FECAC090";
    when 16#00738# => romdata <= X"860B8814";
    when 16#00739# => romdata <= X"0C73832B";
    when 16#0073A# => romdata <= X"82078C14";
    when 16#0073B# => romdata <= X"0C720852";
    when 16#0073C# => romdata <= X"71FB3881";
    when 16#0073D# => romdata <= X"147081FF";
    when 16#0073E# => romdata <= X"065551A2";
    when 16#0073F# => romdata <= X"7427DA38";
    when 16#00740# => romdata <= X"71B00C85";
    when 16#00741# => romdata <= X"3D0D04FD";
    when 16#00742# => romdata <= X"3D0D800B";
    when 16#00743# => romdata <= X"80FCC808";
    when 16#00744# => romdata <= X"54548073";
    when 16#00745# => romdata <= X"0C880A0B";
    when 16#00746# => romdata <= X"88140C73";
    when 16#00747# => romdata <= X"832B8107";
    when 16#00748# => romdata <= X"8C140C72";
    when 16#00749# => romdata <= X"085271FB";
    when 16#0074A# => romdata <= X"38811470";
    when 16#0074B# => romdata <= X"81FF0655";
    when 16#0074C# => romdata <= X"51A27427";
    when 16#0074D# => romdata <= X"DD3871B0";
    when 16#0074E# => romdata <= X"0C853D0D";
    when 16#0074F# => romdata <= X"04FE3D0D";
    when 16#00750# => romdata <= X"8151DEB2";
    when 16#00751# => romdata <= X"3F80FCC8";
    when 16#00752# => romdata <= X"08538073";
    when 16#00753# => romdata <= X"0C810B88";
    when 16#00754# => romdata <= X"140CB008";
    when 16#00755# => romdata <= X"832B8FF8";
    when 16#00756# => romdata <= X"06708207";
    when 16#00757# => romdata <= X"8C150C52";
    when 16#00758# => romdata <= X"72085271";
    when 16#00759# => romdata <= X"FB388973";
    when 16#0075A# => romdata <= X"0C71B00C";
    when 16#0075B# => romdata <= X"843D0D04";
    when 16#0075C# => romdata <= X"D88A3F04";
    when 16#0075D# => romdata <= X"FB3D0D77";
    when 16#0075E# => romdata <= X"79555580";
    when 16#0075F# => romdata <= X"56757524";
    when 16#00760# => romdata <= X"AB388074";
    when 16#00761# => romdata <= X"249D3880";
    when 16#00762# => romdata <= X"53735274";
    when 16#00763# => romdata <= X"5180E13F";
    when 16#00764# => romdata <= X"B0085475";
    when 16#00765# => romdata <= X"802E8538";
    when 16#00766# => romdata <= X"B0083054";
    when 16#00767# => romdata <= X"73B00C87";
    when 16#00768# => romdata <= X"3D0D0473";
    when 16#00769# => romdata <= X"30768132";
    when 16#0076A# => romdata <= X"5754DC39";
    when 16#0076B# => romdata <= X"74305581";
    when 16#0076C# => romdata <= X"56738025";
    when 16#0076D# => romdata <= X"D238EC39";
    when 16#0076E# => romdata <= X"FA3D0D78";
    when 16#0076F# => romdata <= X"7A575580";
    when 16#00770# => romdata <= X"57767524";
    when 16#00771# => romdata <= X"A438759F";
    when 16#00772# => romdata <= X"2C548153";
    when 16#00773# => romdata <= X"75743274";
    when 16#00774# => romdata <= X"31527451";
    when 16#00775# => romdata <= X"9B3FB008";
    when 16#00776# => romdata <= X"5476802E";
    when 16#00777# => romdata <= X"8538B008";
    when 16#00778# => romdata <= X"305473B0";
    when 16#00779# => romdata <= X"0C883D0D";
    when 16#0077A# => romdata <= X"04743055";
    when 16#0077B# => romdata <= X"8157D739";
    when 16#0077C# => romdata <= X"FC3D0D76";
    when 16#0077D# => romdata <= X"78535481";
    when 16#0077E# => romdata <= X"53807473";
    when 16#0077F# => romdata <= X"26525572";
    when 16#00780# => romdata <= X"802E9838";
    when 16#00781# => romdata <= X"70802EA9";
    when 16#00782# => romdata <= X"38807224";
    when 16#00783# => romdata <= X"A4387110";
    when 16#00784# => romdata <= X"73107572";
    when 16#00785# => romdata <= X"26535452";
    when 16#00786# => romdata <= X"72EA3873";
    when 16#00787# => romdata <= X"51788338";
    when 16#00788# => romdata <= X"745170B0";
    when 16#00789# => romdata <= X"0C863D0D";
    when 16#0078A# => romdata <= X"0472812A";
    when 16#0078B# => romdata <= X"72812A53";
    when 16#0078C# => romdata <= X"5372802E";
    when 16#0078D# => romdata <= X"E6387174";
    when 16#0078E# => romdata <= X"26EF3873";
    when 16#0078F# => romdata <= X"72317574";
    when 16#00790# => romdata <= X"0774812A";
    when 16#00791# => romdata <= X"74812A55";
    when 16#00792# => romdata <= X"555654E5";
    when 16#00793# => romdata <= X"39101010";
    when 16#00794# => romdata <= X"10101010";
    when 16#00795# => romdata <= X"10101010";
    when 16#00796# => romdata <= X"10101010";
    when 16#00797# => romdata <= X"10101010";
    when 16#00798# => romdata <= X"10101010";
    when 16#00799# => romdata <= X"10101010";
    when 16#0079A# => romdata <= X"10101010";
    when 16#0079B# => romdata <= X"53510473";
    when 16#0079C# => romdata <= X"81FF0673";
    when 16#0079D# => romdata <= X"83060981";
    when 16#0079E# => romdata <= X"05830510";
    when 16#0079F# => romdata <= X"10102B07";
    when 16#007A0# => romdata <= X"72FC060C";
    when 16#007A1# => romdata <= X"5151043C";
    when 16#007A2# => romdata <= X"04727280";
    when 16#007A3# => romdata <= X"728106FF";
    when 16#007A4# => romdata <= X"05097206";
    when 16#007A5# => romdata <= X"05711052";
    when 16#007A6# => romdata <= X"720A100A";
    when 16#007A7# => romdata <= X"5372ED38";
    when 16#007A8# => romdata <= X"51515351";
    when 16#007A9# => romdata <= X"04B008B4";
    when 16#007AA# => romdata <= X"08B80875";
    when 16#007AB# => romdata <= X"75BBB82D";
    when 16#007AC# => romdata <= X"5050B008";
    when 16#007AD# => romdata <= X"56B80CB4";
    when 16#007AE# => romdata <= X"0CB00C51";
    when 16#007AF# => romdata <= X"04B008B4";
    when 16#007B0# => romdata <= X"08B80875";
    when 16#007B1# => romdata <= X"75BAF42D";
    when 16#007B2# => romdata <= X"5050B008";
    when 16#007B3# => romdata <= X"56B80CB4";
    when 16#007B4# => romdata <= X"0CB00C51";
    when 16#007B5# => romdata <= X"04B008B4";
    when 16#007B6# => romdata <= X"08B80890";
    when 16#007B7# => romdata <= X"CB2DB80C";
    when 16#007B8# => romdata <= X"B40CB00C";
    when 16#007B9# => romdata <= X"04FF3D0D";
    when 16#007BA# => romdata <= X"028F0533";
    when 16#007BB# => romdata <= X"80FCF808";
    when 16#007BC# => romdata <= X"52710C80";
    when 16#007BD# => romdata <= X"0BB00C83";
    when 16#007BE# => romdata <= X"3D0D04FF";
    when 16#007BF# => romdata <= X"3D0D028F";
    when 16#007C0# => romdata <= X"05335181";
    when 16#007C1# => romdata <= X"A5900852";
    when 16#007C2# => romdata <= X"712DB008";
    when 16#007C3# => romdata <= X"81FF06B0";
    when 16#007C4# => romdata <= X"0C833D0D";
    when 16#007C5# => romdata <= X"04FE3D0D";
    when 16#007C6# => romdata <= X"74703353";
    when 16#007C7# => romdata <= X"5371802E";
    when 16#007C8# => romdata <= X"93388113";
    when 16#007C9# => romdata <= X"725281A5";
    when 16#007CA# => romdata <= X"90085353";
    when 16#007CB# => romdata <= X"712D7233";
    when 16#007CC# => romdata <= X"5271EF38";
    when 16#007CD# => romdata <= X"843D0D04";
    when 16#007CE# => romdata <= X"F43D0D7F";
    when 16#007CF# => romdata <= X"028405BB";
    when 16#007D0# => romdata <= X"05335557";
    when 16#007D1# => romdata <= X"880B8C3D";
    when 16#007D2# => romdata <= X"5B598953";
    when 16#007D3# => romdata <= X"80FA9C52";
    when 16#007D4# => romdata <= X"795185E6";
    when 16#007D5# => romdata <= X"3F73792E";
    when 16#007D6# => romdata <= X"80FF3878";
    when 16#007D7# => romdata <= X"5673902E";
    when 16#007D8# => romdata <= X"80EC3802";
    when 16#007D9# => romdata <= X"A7055876";
    when 16#007DA# => romdata <= X"8F065473";
    when 16#007DB# => romdata <= X"892680C2";
    when 16#007DC# => romdata <= X"387518B0";
    when 16#007DD# => romdata <= X"15555573";
    when 16#007DE# => romdata <= X"75347684";
    when 16#007DF# => romdata <= X"2AFF1770";
    when 16#007E0# => romdata <= X"81FF0658";
    when 16#007E1# => romdata <= X"555775DF";
    when 16#007E2# => romdata <= X"38781A55";
    when 16#007E3# => romdata <= X"75753479";
    when 16#007E4# => romdata <= X"70335555";
    when 16#007E5# => romdata <= X"73802E93";
    when 16#007E6# => romdata <= X"38811574";
    when 16#007E7# => romdata <= X"5281A590";
    when 16#007E8# => romdata <= X"08575575";
    when 16#007E9# => romdata <= X"2D743354";
    when 16#007EA# => romdata <= X"73EF3878";
    when 16#007EB# => romdata <= X"B00C8E3D";
    when 16#007EC# => romdata <= X"0D047518";
    when 16#007ED# => romdata <= X"B7155555";
    when 16#007EE# => romdata <= X"73753476";
    when 16#007EF# => romdata <= X"842AFF17";
    when 16#007F0# => romdata <= X"7081FF06";
    when 16#007F1# => romdata <= X"58555775";
    when 16#007F2# => romdata <= X"FF9D38FF";
    when 16#007F3# => romdata <= X"BC398470";
    when 16#007F4# => romdata <= X"575902A7";
    when 16#007F5# => romdata <= X"0558FF8F";
    when 16#007F6# => romdata <= X"39827057";
    when 16#007F7# => romdata <= X"59F439F1";
    when 16#007F8# => romdata <= X"3D0D618D";
    when 16#007F9# => romdata <= X"3D705B5C";
    when 16#007FA# => romdata <= X"5A807A56";
    when 16#007FB# => romdata <= X"57767A24";
    when 16#007FC# => romdata <= X"81853878";
    when 16#007FD# => romdata <= X"17548A52";
    when 16#007FE# => romdata <= X"7451848C";
    when 16#007FF# => romdata <= X"3FB008B0";
    when 16#00800# => romdata <= X"05537274";
    when 16#00801# => romdata <= X"34811757";
    when 16#00802# => romdata <= X"8A527451";
    when 16#00803# => romdata <= X"83D53FB0";
    when 16#00804# => romdata <= X"0855B008";
    when 16#00805# => romdata <= X"DE38B008";
    when 16#00806# => romdata <= X"779F2A18";
    when 16#00807# => romdata <= X"70812C5A";
    when 16#00808# => romdata <= X"56568078";
    when 16#00809# => romdata <= X"259E3878";
    when 16#0080A# => romdata <= X"17FF0555";
    when 16#0080B# => romdata <= X"75197033";
    when 16#0080C# => romdata <= X"55537433";
    when 16#0080D# => romdata <= X"73347375";
    when 16#0080E# => romdata <= X"348116FF";
    when 16#0080F# => romdata <= X"16565677";
    when 16#00810# => romdata <= X"7624E938";
    when 16#00811# => romdata <= X"76195880";
    when 16#00812# => romdata <= X"7834807A";
    when 16#00813# => romdata <= X"24177081";
    when 16#00814# => romdata <= X"FF067C70";
    when 16#00815# => romdata <= X"33565755";
    when 16#00816# => romdata <= X"5672802E";
    when 16#00817# => romdata <= X"93388115";
    when 16#00818# => romdata <= X"735281A5";
    when 16#00819# => romdata <= X"90085855";
    when 16#0081A# => romdata <= X"762D7433";
    when 16#0081B# => romdata <= X"5372EF38";
    when 16#0081C# => romdata <= X"73B00C91";
    when 16#0081D# => romdata <= X"3D0D04AD";
    when 16#0081E# => romdata <= X"7B3402AD";
    when 16#0081F# => romdata <= X"057A3071";
    when 16#00820# => romdata <= X"19565659";
    when 16#00821# => romdata <= X"8A527451";
    when 16#00822# => romdata <= X"82FE3FB0";
    when 16#00823# => romdata <= X"08B00553";
    when 16#00824# => romdata <= X"72743481";
    when 16#00825# => romdata <= X"17578A52";
    when 16#00826# => romdata <= X"745182C7";
    when 16#00827# => romdata <= X"3FB00855";
    when 16#00828# => romdata <= X"B008FECF";
    when 16#00829# => romdata <= X"38FEEF39";
    when 16#0082A# => romdata <= X"FD3D0D02";
    when 16#0082B# => romdata <= X"97053302";
    when 16#0082C# => romdata <= X"84059B05";
    when 16#0082D# => romdata <= X"33555372";
    when 16#0082E# => romdata <= X"74279738";
    when 16#0082F# => romdata <= X"A05181A5";
    when 16#00830# => romdata <= X"90085271";
    when 16#00831# => romdata <= X"2D811370";
    when 16#00832# => romdata <= X"81FF0654";
    when 16#00833# => romdata <= X"52737326";
    when 16#00834# => romdata <= X"EB38853D";
    when 16#00835# => romdata <= X"0D04FF3D";
    when 16#00836# => romdata <= X"0D80FCEC";
    when 16#00837# => romdata <= X"08741015";
    when 16#00838# => romdata <= X"70822B94";
    when 16#00839# => romdata <= X"130C5252";
    when 16#0083A# => romdata <= X"850B9813";
    when 16#0083B# => romdata <= X"0C981208";
    when 16#0083C# => romdata <= X"70810651";
    when 16#0083D# => romdata <= X"5170F638";
    when 16#0083E# => romdata <= X"833D0D04";
    when 16#0083F# => romdata <= X"FD3D0D80";
    when 16#00840# => romdata <= X"FCEC0876";
    when 16#00841# => romdata <= X"80E1D429";
    when 16#00842# => romdata <= X"94120C54";
    when 16#00843# => romdata <= X"850B9815";
    when 16#00844# => romdata <= X"0C981408";
    when 16#00845# => romdata <= X"70810651";
    when 16#00846# => romdata <= X"5372F638";
    when 16#00847# => romdata <= X"853D0D04";
    when 16#00848# => romdata <= X"803D0D80";
    when 16#00849# => romdata <= X"FCEC0851";
    when 16#0084A# => romdata <= X"870B8412";
    when 16#0084B# => romdata <= X"0CFF0BA4";
    when 16#0084C# => romdata <= X"120CA70B";
    when 16#0084D# => romdata <= X"A8120C80";
    when 16#0084E# => romdata <= X"E1D40B94";
    when 16#0084F# => romdata <= X"120C870B";
    when 16#00850# => romdata <= X"98120C82";
    when 16#00851# => romdata <= X"3D0D0480";
    when 16#00852# => romdata <= X"3D0D80FC";
    when 16#00853# => romdata <= X"F0085180";
    when 16#00854# => romdata <= X"EC0B8C12";
    when 16#00855# => romdata <= X"0C830B88";
    when 16#00856# => romdata <= X"120C823D";
    when 16#00857# => romdata <= X"0D04803D";
    when 16#00858# => romdata <= X"0D80FCF0";
    when 16#00859# => romdata <= X"08841108";
    when 16#0085A# => romdata <= X"8106B00C";
    when 16#0085B# => romdata <= X"51823D0D";
    when 16#0085C# => romdata <= X"04FF3D0D";
    when 16#0085D# => romdata <= X"80FCF008";
    when 16#0085E# => romdata <= X"52841208";
    when 16#0085F# => romdata <= X"70810651";
    when 16#00860# => romdata <= X"5170802E";
    when 16#00861# => romdata <= X"F4387108";
    when 16#00862# => romdata <= X"7081FF06";
    when 16#00863# => romdata <= X"B00C5183";
    when 16#00864# => romdata <= X"3D0D04FE";
    when 16#00865# => romdata <= X"3D0D0293";
    when 16#00866# => romdata <= X"05335372";
    when 16#00867# => romdata <= X"8A2E9C38";
    when 16#00868# => romdata <= X"80FCF008";
    when 16#00869# => romdata <= X"52841208";
    when 16#0086A# => romdata <= X"70892A70";
    when 16#0086B# => romdata <= X"81065151";
    when 16#0086C# => romdata <= X"5170F238";
    when 16#0086D# => romdata <= X"72720C84";
    when 16#0086E# => romdata <= X"3D0D0480";
    when 16#0086F# => romdata <= X"FCF00852";
    when 16#00870# => romdata <= X"84120870";
    when 16#00871# => romdata <= X"892A7081";
    when 16#00872# => romdata <= X"06515151";
    when 16#00873# => romdata <= X"70F2388D";
    when 16#00874# => romdata <= X"720C8412";
    when 16#00875# => romdata <= X"0870892A";
    when 16#00876# => romdata <= X"70810651";
    when 16#00877# => romdata <= X"515170C5";
    when 16#00878# => romdata <= X"38D239BC";
    when 16#00879# => romdata <= X"0802BC0C";
    when 16#0087A# => romdata <= X"FD3D0D80";
    when 16#0087B# => romdata <= X"53BC088C";
    when 16#0087C# => romdata <= X"050852BC";
    when 16#0087D# => romdata <= X"08880508";
    when 16#0087E# => romdata <= X"51F7F53F";
    when 16#0087F# => romdata <= X"B00870B0";
    when 16#00880# => romdata <= X"0C54853D";
    when 16#00881# => romdata <= X"0DBC0C04";
    when 16#00882# => romdata <= X"BC0802BC";
    when 16#00883# => romdata <= X"0CFD3D0D";
    when 16#00884# => romdata <= X"8153BC08";
    when 16#00885# => romdata <= X"8C050852";
    when 16#00886# => romdata <= X"BC088805";
    when 16#00887# => romdata <= X"0851F7D0";
    when 16#00888# => romdata <= X"3FB00870";
    when 16#00889# => romdata <= X"B00C5485";
    when 16#0088A# => romdata <= X"3D0DBC0C";
    when 16#0088B# => romdata <= X"04803D0D";
    when 16#0088C# => romdata <= X"86518496";
    when 16#0088D# => romdata <= X"3F8151A1";
    when 16#0088E# => romdata <= X"D33FFC3D";
    when 16#0088F# => romdata <= X"0D767079";
    when 16#00890# => romdata <= X"7B555555";
    when 16#00891# => romdata <= X"558F7227";
    when 16#00892# => romdata <= X"8C387275";
    when 16#00893# => romdata <= X"07830651";
    when 16#00894# => romdata <= X"70802EA7";
    when 16#00895# => romdata <= X"38FF1252";
    when 16#00896# => romdata <= X"71FF2E98";
    when 16#00897# => romdata <= X"38727081";
    when 16#00898# => romdata <= X"05543374";
    when 16#00899# => romdata <= X"70810556";
    when 16#0089A# => romdata <= X"34FF1252";
    when 16#0089B# => romdata <= X"71FF2E09";
    when 16#0089C# => romdata <= X"8106EA38";
    when 16#0089D# => romdata <= X"74B00C86";
    when 16#0089E# => romdata <= X"3D0D0474";
    when 16#0089F# => romdata <= X"51727084";
    when 16#008A0# => romdata <= X"05540871";
    when 16#008A1# => romdata <= X"70840553";
    when 16#008A2# => romdata <= X"0C727084";
    when 16#008A3# => romdata <= X"05540871";
    when 16#008A4# => romdata <= X"70840553";
    when 16#008A5# => romdata <= X"0C727084";
    when 16#008A6# => romdata <= X"05540871";
    when 16#008A7# => romdata <= X"70840553";
    when 16#008A8# => romdata <= X"0C727084";
    when 16#008A9# => romdata <= X"05540871";
    when 16#008AA# => romdata <= X"70840553";
    when 16#008AB# => romdata <= X"0CF01252";
    when 16#008AC# => romdata <= X"718F26C9";
    when 16#008AD# => romdata <= X"38837227";
    when 16#008AE# => romdata <= X"95387270";
    when 16#008AF# => romdata <= X"84055408";
    when 16#008B0# => romdata <= X"71708405";
    when 16#008B1# => romdata <= X"530CFC12";
    when 16#008B2# => romdata <= X"52718326";
    when 16#008B3# => romdata <= X"ED387054";
    when 16#008B4# => romdata <= X"FF8339FD";
    when 16#008B5# => romdata <= X"3D0D7553";
    when 16#008B6# => romdata <= X"84D81308";
    when 16#008B7# => romdata <= X"802E8A38";
    when 16#008B8# => romdata <= X"805372B0";
    when 16#008B9# => romdata <= X"0C853D0D";
    when 16#008BA# => romdata <= X"04818052";
    when 16#008BB# => romdata <= X"72518D9B";
    when 16#008BC# => romdata <= X"3FB00884";
    when 16#008BD# => romdata <= X"D8140CFF";
    when 16#008BE# => romdata <= X"53B00880";
    when 16#008BF# => romdata <= X"2EE438B0";
    when 16#008C0# => romdata <= X"08549F53";
    when 16#008C1# => romdata <= X"80747084";
    when 16#008C2# => romdata <= X"05560CFF";
    when 16#008C3# => romdata <= X"13538073";
    when 16#008C4# => romdata <= X"24CE3880";
    when 16#008C5# => romdata <= X"74708405";
    when 16#008C6# => romdata <= X"560CFF13";
    when 16#008C7# => romdata <= X"53728025";
    when 16#008C8# => romdata <= X"E338FFBC";
    when 16#008C9# => romdata <= X"39FD3D0D";
    when 16#008CA# => romdata <= X"75775553";
    when 16#008CB# => romdata <= X"9F74278D";
    when 16#008CC# => romdata <= X"3896730C";
    when 16#008CD# => romdata <= X"FF5271B0";
    when 16#008CE# => romdata <= X"0C853D0D";
    when 16#008CF# => romdata <= X"0484D813";
    when 16#008D0# => romdata <= X"08527180";
    when 16#008D1# => romdata <= X"2E933873";
    when 16#008D2# => romdata <= X"10101270";
    when 16#008D3# => romdata <= X"0879720C";
    when 16#008D4# => romdata <= X"515271B0";
    when 16#008D5# => romdata <= X"0C853D0D";
    when 16#008D6# => romdata <= X"047251FE";
    when 16#008D7# => romdata <= X"F63FFF52";
    when 16#008D8# => romdata <= X"B008D338";
    when 16#008D9# => romdata <= X"84D81308";
    when 16#008DA# => romdata <= X"74101011";
    when 16#008DB# => romdata <= X"70087A72";
    when 16#008DC# => romdata <= X"0C515152";
    when 16#008DD# => romdata <= X"DD39F93D";
    when 16#008DE# => romdata <= X"0D797B58";
    when 16#008DF# => romdata <= X"56769F26";
    when 16#008E0# => romdata <= X"80E83884";
    when 16#008E1# => romdata <= X"D8160854";
    when 16#008E2# => romdata <= X"73802EAA";
    when 16#008E3# => romdata <= X"38761010";
    when 16#008E4# => romdata <= X"14700855";
    when 16#008E5# => romdata <= X"5573802E";
    when 16#008E6# => romdata <= X"BA388058";
    when 16#008E7# => romdata <= X"73812E8F";
    when 16#008E8# => romdata <= X"3873FF2E";
    when 16#008E9# => romdata <= X"A3388075";
    when 16#008EA# => romdata <= X"0C765173";
    when 16#008EB# => romdata <= X"2D805877";
    when 16#008EC# => romdata <= X"B00C893D";
    when 16#008ED# => romdata <= X"0D047551";
    when 16#008EE# => romdata <= X"FE993FFF";
    when 16#008EF# => romdata <= X"58B008EF";
    when 16#008F0# => romdata <= X"3884D816";
    when 16#008F1# => romdata <= X"0854C639";
    when 16#008F2# => romdata <= X"96760C81";
    when 16#008F3# => romdata <= X"0BB00C89";
    when 16#008F4# => romdata <= X"3D0D0475";
    when 16#008F5# => romdata <= X"5181ED3F";
    when 16#008F6# => romdata <= X"7653B008";
    when 16#008F7# => romdata <= X"52755181";
    when 16#008F8# => romdata <= X"AD3FB008";
    when 16#008F9# => romdata <= X"B00C893D";
    when 16#008FA# => romdata <= X"0D049676";
    when 16#008FB# => romdata <= X"0CFF0BB0";
    when 16#008FC# => romdata <= X"0C893D0D";
    when 16#008FD# => romdata <= X"04FC3D0D";
    when 16#008FE# => romdata <= X"76785653";
    when 16#008FF# => romdata <= X"FF54749F";
    when 16#00900# => romdata <= X"26B13884";
    when 16#00901# => romdata <= X"D8130852";
    when 16#00902# => romdata <= X"71802EAE";
    when 16#00903# => romdata <= X"38741010";
    when 16#00904# => romdata <= X"12700853";
    when 16#00905# => romdata <= X"53815471";
    when 16#00906# => romdata <= X"802E9838";
    when 16#00907# => romdata <= X"825471FF";
    when 16#00908# => romdata <= X"2E913883";
    when 16#00909# => romdata <= X"5471812E";
    when 16#0090A# => romdata <= X"8A388073";
    when 16#0090B# => romdata <= X"0C745171";
    when 16#0090C# => romdata <= X"2D805473";
    when 16#0090D# => romdata <= X"B00C863D";
    when 16#0090E# => romdata <= X"0D047251";
    when 16#0090F# => romdata <= X"FD953FB0";
    when 16#00910# => romdata <= X"08F13884";
    when 16#00911# => romdata <= X"D8130852";
    when 16#00912# => romdata <= X"C439FF3D";
    when 16#00913# => romdata <= X"0D735280";
    when 16#00914# => romdata <= X"FCFC0851";
    when 16#00915# => romdata <= X"FEA03F83";
    when 16#00916# => romdata <= X"3D0D04FE";
    when 16#00917# => romdata <= X"3D0D7553";
    when 16#00918# => romdata <= X"745280FC";
    when 16#00919# => romdata <= X"FC0851FD";
    when 16#0091A# => romdata <= X"BC3F843D";
    when 16#0091B# => romdata <= X"0D04803D";
    when 16#0091C# => romdata <= X"0D80FCFC";
    when 16#0091D# => romdata <= X"0851FCDB";
    when 16#0091E# => romdata <= X"3F823D0D";
    when 16#0091F# => romdata <= X"04FF3D0D";
    when 16#00920# => romdata <= X"735280FC";
    when 16#00921# => romdata <= X"FC0851FE";
    when 16#00922# => romdata <= X"EC3F833D";
    when 16#00923# => romdata <= X"0D04FC3D";
    when 16#00924# => romdata <= X"0D800B81";
    when 16#00925# => romdata <= X"A5980C78";
    when 16#00926# => romdata <= X"5277519C";
    when 16#00927# => romdata <= X"AA3FB008";
    when 16#00928# => romdata <= X"54B008FF";
    when 16#00929# => romdata <= X"2E883873";
    when 16#0092A# => romdata <= X"B00C863D";
    when 16#0092B# => romdata <= X"0D0481A5";
    when 16#0092C# => romdata <= X"98085574";
    when 16#0092D# => romdata <= X"802EF038";
    when 16#0092E# => romdata <= X"7675710C";
    when 16#0092F# => romdata <= X"5373B00C";
    when 16#00930# => romdata <= X"863D0D04";
    when 16#00931# => romdata <= X"9BFC3F04";
    when 16#00932# => romdata <= X"FC3D0D76";
    when 16#00933# => romdata <= X"70797073";
    when 16#00934# => romdata <= X"07830654";
    when 16#00935# => romdata <= X"54545570";
    when 16#00936# => romdata <= X"80C33871";
    when 16#00937# => romdata <= X"70087009";
    when 16#00938# => romdata <= X"70F7FBFD";
    when 16#00939# => romdata <= X"FF130670";
    when 16#0093A# => romdata <= X"F8848281";
    when 16#0093B# => romdata <= X"80065151";
    when 16#0093C# => romdata <= X"53535470";
    when 16#0093D# => romdata <= X"A6388414";
    when 16#0093E# => romdata <= X"72747084";
    when 16#0093F# => romdata <= X"05560C70";
    when 16#00940# => romdata <= X"08700970";
    when 16#00941# => romdata <= X"F7FBFDFF";
    when 16#00942# => romdata <= X"130670F8";
    when 16#00943# => romdata <= X"84828180";
    when 16#00944# => romdata <= X"06515153";
    when 16#00945# => romdata <= X"53547080";
    when 16#00946# => romdata <= X"2EDC3873";
    when 16#00947# => romdata <= X"52717081";
    when 16#00948# => romdata <= X"05533351";
    when 16#00949# => romdata <= X"70737081";
    when 16#0094A# => romdata <= X"05553470";
    when 16#0094B# => romdata <= X"F03874B0";
    when 16#0094C# => romdata <= X"0C863D0D";
    when 16#0094D# => romdata <= X"04FD3D0D";
    when 16#0094E# => romdata <= X"75707183";
    when 16#0094F# => romdata <= X"06535552";
    when 16#00950# => romdata <= X"70B83871";
    when 16#00951# => romdata <= X"70087009";
    when 16#00952# => romdata <= X"F7FBFDFF";
    when 16#00953# => romdata <= X"120670F8";
    when 16#00954# => romdata <= X"84828180";
    when 16#00955# => romdata <= X"06515152";
    when 16#00956# => romdata <= X"53709D38";
    when 16#00957# => romdata <= X"84137008";
    when 16#00958# => romdata <= X"7009F7FB";
    when 16#00959# => romdata <= X"FDFF1206";
    when 16#0095A# => romdata <= X"70F88482";
    when 16#0095B# => romdata <= X"81800651";
    when 16#0095C# => romdata <= X"51525370";
    when 16#0095D# => romdata <= X"802EE538";
    when 16#0095E# => romdata <= X"72527133";
    when 16#0095F# => romdata <= X"5170802E";
    when 16#00960# => romdata <= X"8A388112";
    when 16#00961# => romdata <= X"70335252";
    when 16#00962# => romdata <= X"70F83871";
    when 16#00963# => romdata <= X"7431B00C";
    when 16#00964# => romdata <= X"853D0D04";
    when 16#00965# => romdata <= X"FA3D0D78";
    when 16#00966# => romdata <= X"7A7C7054";
    when 16#00967# => romdata <= X"55555272";
    when 16#00968# => romdata <= X"802E80D9";
    when 16#00969# => romdata <= X"38717407";
    when 16#0096A# => romdata <= X"83065170";
    when 16#0096B# => romdata <= X"802E80D4";
    when 16#0096C# => romdata <= X"38FF1353";
    when 16#0096D# => romdata <= X"72FF2EB1";
    when 16#0096E# => romdata <= X"38713374";
    when 16#0096F# => romdata <= X"33565174";
    when 16#00970# => romdata <= X"712E0981";
    when 16#00971# => romdata <= X"06A93872";
    when 16#00972# => romdata <= X"802E8187";
    when 16#00973# => romdata <= X"387081FF";
    when 16#00974# => romdata <= X"06517080";
    when 16#00975# => romdata <= X"2E80FC38";
    when 16#00976# => romdata <= X"81128115";
    when 16#00977# => romdata <= X"FF155555";
    when 16#00978# => romdata <= X"5272FF2E";
    when 16#00979# => romdata <= X"098106D1";
    when 16#0097A# => romdata <= X"38713374";
    when 16#0097B# => romdata <= X"33565170";
    when 16#0097C# => romdata <= X"81FF0675";
    when 16#0097D# => romdata <= X"81FF0671";
    when 16#0097E# => romdata <= X"71315152";
    when 16#0097F# => romdata <= X"5270B00C";
    when 16#00980# => romdata <= X"883D0D04";
    when 16#00981# => romdata <= X"71745755";
    when 16#00982# => romdata <= X"83732788";
    when 16#00983# => romdata <= X"38710874";
    when 16#00984# => romdata <= X"082E8838";
    when 16#00985# => romdata <= X"74765552";
    when 16#00986# => romdata <= X"FF9739FC";
    when 16#00987# => romdata <= X"13537280";
    when 16#00988# => romdata <= X"2EB13874";
    when 16#00989# => romdata <= X"087009F7";
    when 16#0098A# => romdata <= X"FBFDFF12";
    when 16#0098B# => romdata <= X"0670F884";
    when 16#0098C# => romdata <= X"82818006";
    when 16#0098D# => romdata <= X"51515170";
    when 16#0098E# => romdata <= X"9A388415";
    when 16#0098F# => romdata <= X"84175755";
    when 16#00990# => romdata <= X"837327D0";
    when 16#00991# => romdata <= X"38740876";
    when 16#00992# => romdata <= X"082ED038";
    when 16#00993# => romdata <= X"74765552";
    when 16#00994# => romdata <= X"FEDF3980";
    when 16#00995# => romdata <= X"0BB00C88";
    when 16#00996# => romdata <= X"3D0D04F3";
    when 16#00997# => romdata <= X"3D0D6062";
    when 16#00998# => romdata <= X"64725A5A";
    when 16#00999# => romdata <= X"5E5E805C";
    when 16#0099A# => romdata <= X"76708105";
    when 16#0099B# => romdata <= X"583380FA";
    when 16#0099C# => romdata <= X"B1113370";
    when 16#0099D# => romdata <= X"832A7081";
    when 16#0099E# => romdata <= X"06515555";
    when 16#0099F# => romdata <= X"5672E938";
    when 16#009A0# => romdata <= X"75AD2E82";
    when 16#009A1# => romdata <= X"883875AB";
    when 16#009A2# => romdata <= X"2E828438";
    when 16#009A3# => romdata <= X"77307079";
    when 16#009A4# => romdata <= X"07802579";
    when 16#009A5# => romdata <= X"90327030";
    when 16#009A6# => romdata <= X"70720780";
    when 16#009A7# => romdata <= X"25730753";
    when 16#009A8# => romdata <= X"57575153";
    when 16#009A9# => romdata <= X"72802E87";
    when 16#009AA# => romdata <= X"3875B02E";
    when 16#009AB# => romdata <= X"81EB3877";
    when 16#009AC# => romdata <= X"8A388858";
    when 16#009AD# => romdata <= X"75B02E83";
    when 16#009AE# => romdata <= X"388A5881";
    when 16#009AF# => romdata <= X"0A5A7B84";
    when 16#009B0# => romdata <= X"38FE0A5A";
    when 16#009B1# => romdata <= X"77527951";
    when 16#009B2# => romdata <= X"F6BE3FB0";
    when 16#009B3# => romdata <= X"0878537A";
    when 16#009B4# => romdata <= X"525BF68F";
    when 16#009B5# => romdata <= X"3FB0085A";
    when 16#009B6# => romdata <= X"807080FA";
    when 16#009B7# => romdata <= X"B1183370";
    when 16#009B8# => romdata <= X"822A7081";
    when 16#009B9# => romdata <= X"06515656";
    when 16#009BA# => romdata <= X"5A557280";
    when 16#009BB# => romdata <= X"2E80C138";
    when 16#009BC# => romdata <= X"D0165675";
    when 16#009BD# => romdata <= X"782580D7";
    when 16#009BE# => romdata <= X"38807924";
    when 16#009BF# => romdata <= X"757B2607";
    when 16#009C0# => romdata <= X"53729338";
    when 16#009C1# => romdata <= X"747A2E80";
    when 16#009C2# => romdata <= X"EB387A76";
    when 16#009C3# => romdata <= X"2580ED38";
    when 16#009C4# => romdata <= X"72802E80";
    when 16#009C5# => romdata <= X"E738FF77";
    when 16#009C6# => romdata <= X"70810559";
    when 16#009C7# => romdata <= X"33575980";
    when 16#009C8# => romdata <= X"FAB11633";
    when 16#009C9# => romdata <= X"70822A70";
    when 16#009CA# => romdata <= X"81065154";
    when 16#009CB# => romdata <= X"5472C138";
    when 16#009CC# => romdata <= X"73830653";
    when 16#009CD# => romdata <= X"72802E97";
    when 16#009CE# => romdata <= X"38738106";
    when 16#009CF# => romdata <= X"C9175553";
    when 16#009D0# => romdata <= X"728538FF";
    when 16#009D1# => romdata <= X"A9165473";
    when 16#009D2# => romdata <= X"56777624";
    when 16#009D3# => romdata <= X"FFAB3880";
    when 16#009D4# => romdata <= X"792480F0";
    when 16#009D5# => romdata <= X"387B802E";
    when 16#009D6# => romdata <= X"84387430";
    when 16#009D7# => romdata <= X"557C802E";
    when 16#009D8# => romdata <= X"8C38FF17";
    when 16#009D9# => romdata <= X"53788338";
    when 16#009DA# => romdata <= X"7D53727D";
    when 16#009DB# => romdata <= X"0C74B00C";
    when 16#009DC# => romdata <= X"8F3D0D04";
    when 16#009DD# => romdata <= X"8153757B";
    when 16#009DE# => romdata <= X"24FF9538";
    when 16#009DF# => romdata <= X"81757929";
    when 16#009E0# => romdata <= X"17787081";
    when 16#009E1# => romdata <= X"055A3358";
    when 16#009E2# => romdata <= X"5659FF93";
    when 16#009E3# => romdata <= X"39815C76";
    when 16#009E4# => romdata <= X"70810558";
    when 16#009E5# => romdata <= X"3356FDF4";
    when 16#009E6# => romdata <= X"39807733";
    when 16#009E7# => romdata <= X"54547280";
    when 16#009E8# => romdata <= X"F82EB238";
    when 16#009E9# => romdata <= X"7280D832";
    when 16#009EA# => romdata <= X"70307080";
    when 16#009EB# => romdata <= X"25760751";
    when 16#009EC# => romdata <= X"51537280";
    when 16#009ED# => romdata <= X"2EFDF838";
    when 16#009EE# => romdata <= X"81173382";
    when 16#009EF# => romdata <= X"18585690";
    when 16#009F0# => romdata <= X"58FDF839";
    when 16#009F1# => romdata <= X"810A557B";
    when 16#009F2# => romdata <= X"8438FE0A";
    when 16#009F3# => romdata <= X"557F53A2";
    when 16#009F4# => romdata <= X"730CFF89";
    when 16#009F5# => romdata <= X"398154CC";
    when 16#009F6# => romdata <= X"39FD3D0D";
    when 16#009F7# => romdata <= X"77547653";
    when 16#009F8# => romdata <= X"755280FC";
    when 16#009F9# => romdata <= X"FC0851FC";
    when 16#009FA# => romdata <= X"F23F853D";
    when 16#009FB# => romdata <= X"0D04F33D";
    when 16#009FC# => romdata <= X"0D606264";
    when 16#009FD# => romdata <= X"725A5A5D";
    when 16#009FE# => romdata <= X"5D805E76";
    when 16#009FF# => romdata <= X"70810558";
    when 16#00A00# => romdata <= X"3380FAB1";
    when 16#00A01# => romdata <= X"11337083";
    when 16#00A02# => romdata <= X"2A708106";
    when 16#00A03# => romdata <= X"51555556";
    when 16#00A04# => romdata <= X"72E93875";
    when 16#00A05# => romdata <= X"AD2E81FF";
    when 16#00A06# => romdata <= X"3875AB2E";
    when 16#00A07# => romdata <= X"81FB3877";
    when 16#00A08# => romdata <= X"30707907";
    when 16#00A09# => romdata <= X"80257990";
    when 16#00A0A# => romdata <= X"32703070";
    when 16#00A0B# => romdata <= X"72078025";
    when 16#00A0C# => romdata <= X"73075357";
    when 16#00A0D# => romdata <= X"57515372";
    when 16#00A0E# => romdata <= X"802E8738";
    when 16#00A0F# => romdata <= X"75B02E81";
    when 16#00A10# => romdata <= X"E238778A";
    when 16#00A11# => romdata <= X"38885875";
    when 16#00A12# => romdata <= X"B02E8338";
    when 16#00A13# => romdata <= X"8A587752";
    when 16#00A14# => romdata <= X"FF51F38F";
    when 16#00A15# => romdata <= X"3FB00878";
    when 16#00A16# => romdata <= X"535AFF51";
    when 16#00A17# => romdata <= X"F3AA3FB0";
    when 16#00A18# => romdata <= X"085B8070";
    when 16#00A19# => romdata <= X"5A5580FA";
    when 16#00A1A# => romdata <= X"B1163370";
    when 16#00A1B# => romdata <= X"822A7081";
    when 16#00A1C# => romdata <= X"06515454";
    when 16#00A1D# => romdata <= X"72802E80";
    when 16#00A1E# => romdata <= X"C138D016";
    when 16#00A1F# => romdata <= X"56757825";
    when 16#00A20# => romdata <= X"80D73880";
    when 16#00A21# => romdata <= X"7924757B";
    when 16#00A22# => romdata <= X"26075372";
    when 16#00A23# => romdata <= X"9338747A";
    when 16#00A24# => romdata <= X"2E80EB38";
    when 16#00A25# => romdata <= X"7A762580";
    when 16#00A26# => romdata <= X"ED387280";
    when 16#00A27# => romdata <= X"2E80E738";
    when 16#00A28# => romdata <= X"FF777081";
    when 16#00A29# => romdata <= X"05593357";
    when 16#00A2A# => romdata <= X"5980FAB1";
    when 16#00A2B# => romdata <= X"16337082";
    when 16#00A2C# => romdata <= X"2A708106";
    when 16#00A2D# => romdata <= X"51545472";
    when 16#00A2E# => romdata <= X"C1387383";
    when 16#00A2F# => romdata <= X"06537280";
    when 16#00A30# => romdata <= X"2E973873";
    when 16#00A31# => romdata <= X"8106C917";
    when 16#00A32# => romdata <= X"55537285";
    when 16#00A33# => romdata <= X"38FFA916";
    when 16#00A34# => romdata <= X"54735677";
    when 16#00A35# => romdata <= X"7624FFAB";
    when 16#00A36# => romdata <= X"38807924";
    when 16#00A37# => romdata <= X"8189387D";
    when 16#00A38# => romdata <= X"802E8438";
    when 16#00A39# => romdata <= X"7430557B";
    when 16#00A3A# => romdata <= X"802E8C38";
    when 16#00A3B# => romdata <= X"FF175378";
    when 16#00A3C# => romdata <= X"83387C53";
    when 16#00A3D# => romdata <= X"727C0C74";
    when 16#00A3E# => romdata <= X"B00C8F3D";
    when 16#00A3F# => romdata <= X"0D048153";
    when 16#00A40# => romdata <= X"757B24FF";
    when 16#00A41# => romdata <= X"95388175";
    when 16#00A42# => romdata <= X"79291778";
    when 16#00A43# => romdata <= X"7081055A";
    when 16#00A44# => romdata <= X"33585659";
    when 16#00A45# => romdata <= X"FF933981";
    when 16#00A46# => romdata <= X"5E767081";
    when 16#00A47# => romdata <= X"05583356";
    when 16#00A48# => romdata <= X"FDFD3980";
    when 16#00A49# => romdata <= X"77335454";
    when 16#00A4A# => romdata <= X"7280F82E";
    when 16#00A4B# => romdata <= X"80C33872";
    when 16#00A4C# => romdata <= X"80D83270";
    when 16#00A4D# => romdata <= X"30708025";
    when 16#00A4E# => romdata <= X"76075151";
    when 16#00A4F# => romdata <= X"5372802E";
    when 16#00A50# => romdata <= X"FE803881";
    when 16#00A51# => romdata <= X"17338218";
    when 16#00A52# => romdata <= X"58569070";
    when 16#00A53# => romdata <= X"5358FF51";
    when 16#00A54# => romdata <= X"F1913FB0";
    when 16#00A55# => romdata <= X"0878535A";
    when 16#00A56# => romdata <= X"FF51F1AC";
    when 16#00A57# => romdata <= X"3FB0085B";
    when 16#00A58# => romdata <= X"80705A55";
    when 16#00A59# => romdata <= X"FE8039FF";
    when 16#00A5A# => romdata <= X"605455A2";
    when 16#00A5B# => romdata <= X"730CFEF7";
    when 16#00A5C# => romdata <= X"398154FF";
    when 16#00A5D# => romdata <= X"BA39FD3D";
    when 16#00A5E# => romdata <= X"0D775476";
    when 16#00A5F# => romdata <= X"53755280";
    when 16#00A60# => romdata <= X"FCFC0851";
    when 16#00A61# => romdata <= X"FCE83F85";
    when 16#00A62# => romdata <= X"3D0D04F3";
    when 16#00A63# => romdata <= X"3D0D7F61";
    when 16#00A64# => romdata <= X"8B1170F8";
    when 16#00A65# => romdata <= X"065C5555";
    when 16#00A66# => romdata <= X"5E729626";
    when 16#00A67# => romdata <= X"83389059";
    when 16#00A68# => romdata <= X"80792474";
    when 16#00A69# => romdata <= X"7A260753";
    when 16#00A6A# => romdata <= X"80547274";
    when 16#00A6B# => romdata <= X"2E098106";
    when 16#00A6C# => romdata <= X"80CB387D";
    when 16#00A6D# => romdata <= X"518BCA3F";
    when 16#00A6E# => romdata <= X"7883F726";
    when 16#00A6F# => romdata <= X"80C63878";
    when 16#00A70# => romdata <= X"832A7010";
    when 16#00A71# => romdata <= X"10108184";
    when 16#00A72# => romdata <= X"B8058C11";
    when 16#00A73# => romdata <= X"0859595A";
    when 16#00A74# => romdata <= X"76782E83";
    when 16#00A75# => romdata <= X"B0388417";
    when 16#00A76# => romdata <= X"08FC0656";
    when 16#00A77# => romdata <= X"8C170888";
    when 16#00A78# => romdata <= X"1808718C";
    when 16#00A79# => romdata <= X"120C8812";
    when 16#00A7A# => romdata <= X"0C587517";
    when 16#00A7B# => romdata <= X"84110881";
    when 16#00A7C# => romdata <= X"0784120C";
    when 16#00A7D# => romdata <= X"537D518B";
    when 16#00A7E# => romdata <= X"893F8817";
    when 16#00A7F# => romdata <= X"5473B00C";
    when 16#00A80# => romdata <= X"8F3D0D04";
    when 16#00A81# => romdata <= X"78892A79";
    when 16#00A82# => romdata <= X"832A5B53";
    when 16#00A83# => romdata <= X"72802EBF";
    when 16#00A84# => romdata <= X"3878862A";
    when 16#00A85# => romdata <= X"B8055A84";
    when 16#00A86# => romdata <= X"7327B438";
    when 16#00A87# => romdata <= X"80DB135A";
    when 16#00A88# => romdata <= X"947327AB";
    when 16#00A89# => romdata <= X"38788C2A";
    when 16#00A8A# => romdata <= X"80EE055A";
    when 16#00A8B# => romdata <= X"80D47327";
    when 16#00A8C# => romdata <= X"9E38788F";
    when 16#00A8D# => romdata <= X"2A80F705";
    when 16#00A8E# => romdata <= X"5A82D473";
    when 16#00A8F# => romdata <= X"27913878";
    when 16#00A90# => romdata <= X"922A80FC";
    when 16#00A91# => romdata <= X"055A8AD4";
    when 16#00A92# => romdata <= X"73278438";
    when 16#00A93# => romdata <= X"80FE5A79";
    when 16#00A94# => romdata <= X"10101081";
    when 16#00A95# => romdata <= X"84B8058C";
    when 16#00A96# => romdata <= X"11085855";
    when 16#00A97# => romdata <= X"76752EA3";
    when 16#00A98# => romdata <= X"38841708";
    when 16#00A99# => romdata <= X"FC06707A";
    when 16#00A9A# => romdata <= X"31555673";
    when 16#00A9B# => romdata <= X"8F2488D5";
    when 16#00A9C# => romdata <= X"38738025";
    when 16#00A9D# => romdata <= X"FEE6388C";
    when 16#00A9E# => romdata <= X"17085776";
    when 16#00A9F# => romdata <= X"752E0981";
    when 16#00AA0# => romdata <= X"06DF3881";
    when 16#00AA1# => romdata <= X"1A5A8184";
    when 16#00AA2# => romdata <= X"C8085776";
    when 16#00AA3# => romdata <= X"8184C02E";
    when 16#00AA4# => romdata <= X"82C03884";
    when 16#00AA5# => romdata <= X"1708FC06";
    when 16#00AA6# => romdata <= X"707A3155";
    when 16#00AA7# => romdata <= X"56738F24";
    when 16#00AA8# => romdata <= X"81F93881";
    when 16#00AA9# => romdata <= X"84C00B81";
    when 16#00AAA# => romdata <= X"84CC0C81";
    when 16#00AAB# => romdata <= X"84C00B81";
    when 16#00AAC# => romdata <= X"84C80C73";
    when 16#00AAD# => romdata <= X"8025FEB2";
    when 16#00AAE# => romdata <= X"3883FF76";
    when 16#00AAF# => romdata <= X"2783DF38";
    when 16#00AB0# => romdata <= X"75892A76";
    when 16#00AB1# => romdata <= X"832A5553";
    when 16#00AB2# => romdata <= X"72802EBF";
    when 16#00AB3# => romdata <= X"3875862A";
    when 16#00AB4# => romdata <= X"B8055484";
    when 16#00AB5# => romdata <= X"7327B438";
    when 16#00AB6# => romdata <= X"80DB1354";
    when 16#00AB7# => romdata <= X"947327AB";
    when 16#00AB8# => romdata <= X"38758C2A";
    when 16#00AB9# => romdata <= X"80EE0554";
    when 16#00ABA# => romdata <= X"80D47327";
    when 16#00ABB# => romdata <= X"9E38758F";
    when 16#00ABC# => romdata <= X"2A80F705";
    when 16#00ABD# => romdata <= X"5482D473";
    when 16#00ABE# => romdata <= X"27913875";
    when 16#00ABF# => romdata <= X"922A80FC";
    when 16#00AC0# => romdata <= X"05548AD4";
    when 16#00AC1# => romdata <= X"73278438";
    when 16#00AC2# => romdata <= X"80FE5473";
    when 16#00AC3# => romdata <= X"10101081";
    when 16#00AC4# => romdata <= X"84B80588";
    when 16#00AC5# => romdata <= X"11085658";
    when 16#00AC6# => romdata <= X"74782E86";
    when 16#00AC7# => romdata <= X"CF388415";
    when 16#00AC8# => romdata <= X"08FC0653";
    when 16#00AC9# => romdata <= X"7573278D";
    when 16#00ACA# => romdata <= X"38881508";
    when 16#00ACB# => romdata <= X"5574782E";
    when 16#00ACC# => romdata <= X"098106EA";
    when 16#00ACD# => romdata <= X"388C1508";
    when 16#00ACE# => romdata <= X"8184B80B";
    when 16#00ACF# => romdata <= X"84050871";
    when 16#00AD0# => romdata <= X"8C1A0C76";
    when 16#00AD1# => romdata <= X"881A0C78";
    when 16#00AD2# => romdata <= X"88130C78";
    when 16#00AD3# => romdata <= X"8C180C5D";
    when 16#00AD4# => romdata <= X"58795380";
    when 16#00AD5# => romdata <= X"7A2483E6";
    when 16#00AD6# => romdata <= X"3872822C";
    when 16#00AD7# => romdata <= X"81712B5C";
    when 16#00AD8# => romdata <= X"537A7C26";
    when 16#00AD9# => romdata <= X"8198387B";
    when 16#00ADA# => romdata <= X"7B065372";
    when 16#00ADB# => romdata <= X"82F13879";
    when 16#00ADC# => romdata <= X"FC068405";
    when 16#00ADD# => romdata <= X"5A7A1070";
    when 16#00ADE# => romdata <= X"7D06545B";
    when 16#00ADF# => romdata <= X"7282E038";
    when 16#00AE0# => romdata <= X"841A5AF1";
    when 16#00AE1# => romdata <= X"3988178C";
    when 16#00AE2# => romdata <= X"11085858";
    when 16#00AE3# => romdata <= X"76782E09";
    when 16#00AE4# => romdata <= X"8106FCC2";
    when 16#00AE5# => romdata <= X"38821A5A";
    when 16#00AE6# => romdata <= X"FDEC3978";
    when 16#00AE7# => romdata <= X"17798107";
    when 16#00AE8# => romdata <= X"84190C70";
    when 16#00AE9# => romdata <= X"8184CC0C";
    when 16#00AEA# => romdata <= X"708184C8";
    when 16#00AEB# => romdata <= X"0C8184C0";
    when 16#00AEC# => romdata <= X"0B8C120C";
    when 16#00AED# => romdata <= X"8C110888";
    when 16#00AEE# => romdata <= X"120C7481";
    when 16#00AEF# => romdata <= X"0784120C";
    when 16#00AF0# => romdata <= X"74117571";
    when 16#00AF1# => romdata <= X"0C51537D";
    when 16#00AF2# => romdata <= X"5187B73F";
    when 16#00AF3# => romdata <= X"881754FC";
    when 16#00AF4# => romdata <= X"AC398184";
    when 16#00AF5# => romdata <= X"B80B8405";
    when 16#00AF6# => romdata <= X"087A545C";
    when 16#00AF7# => romdata <= X"798025FE";
    when 16#00AF8# => romdata <= X"F83882DA";
    when 16#00AF9# => romdata <= X"397A097C";
    when 16#00AFA# => romdata <= X"06708184";
    when 16#00AFB# => romdata <= X"B80B8405";
    when 16#00AFC# => romdata <= X"0C5C7A10";
    when 16#00AFD# => romdata <= X"5B7A7C26";
    when 16#00AFE# => romdata <= X"85387A85";
    when 16#00AFF# => romdata <= X"B8388184";
    when 16#00B00# => romdata <= X"B80B8805";
    when 16#00B01# => romdata <= X"08708412";
    when 16#00B02# => romdata <= X"08FC0670";
    when 16#00B03# => romdata <= X"7C317C72";
    when 16#00B04# => romdata <= X"268F7225";
    when 16#00B05# => romdata <= X"0757575C";
    when 16#00B06# => romdata <= X"5D557280";
    when 16#00B07# => romdata <= X"2E80DB38";
    when 16#00B08# => romdata <= X"797A1681";
    when 16#00B09# => romdata <= X"84B0081B";
    when 16#00B0A# => romdata <= X"90115A55";
    when 16#00B0B# => romdata <= X"575B8184";
    when 16#00B0C# => romdata <= X"AC08FF2E";
    when 16#00B0D# => romdata <= X"8838A08F";
    when 16#00B0E# => romdata <= X"13E08006";
    when 16#00B0F# => romdata <= X"5776527D";
    when 16#00B10# => romdata <= X"5186C03F";
    when 16#00B11# => romdata <= X"B00854B0";
    when 16#00B12# => romdata <= X"08FF2E90";
    when 16#00B13# => romdata <= X"38B00876";
    when 16#00B14# => romdata <= X"27829938";
    when 16#00B15# => romdata <= X"748184B8";
    when 16#00B16# => romdata <= X"2E829138";
    when 16#00B17# => romdata <= X"8184B80B";
    when 16#00B18# => romdata <= X"88050855";
    when 16#00B19# => romdata <= X"841508FC";
    when 16#00B1A# => romdata <= X"06707A31";
    when 16#00B1B# => romdata <= X"7A72268F";
    when 16#00B1C# => romdata <= X"72250752";
    when 16#00B1D# => romdata <= X"55537283";
    when 16#00B1E# => romdata <= X"E6387479";
    when 16#00B1F# => romdata <= X"81078417";
    when 16#00B20# => romdata <= X"0C791670";
    when 16#00B21# => romdata <= X"8184B80B";
    when 16#00B22# => romdata <= X"88050C75";
    when 16#00B23# => romdata <= X"81078412";
    when 16#00B24# => romdata <= X"0C547E52";
    when 16#00B25# => romdata <= X"5785EB3F";
    when 16#00B26# => romdata <= X"881754FA";
    when 16#00B27# => romdata <= X"E0397583";
    when 16#00B28# => romdata <= X"2A705454";
    when 16#00B29# => romdata <= X"80742481";
    when 16#00B2A# => romdata <= X"9B387282";
    when 16#00B2B# => romdata <= X"2C81712B";
    when 16#00B2C# => romdata <= X"8184BC08";
    when 16#00B2D# => romdata <= X"07708184";
    when 16#00B2E# => romdata <= X"B80B8405";
    when 16#00B2F# => romdata <= X"0C751010";
    when 16#00B30# => romdata <= X"108184B8";
    when 16#00B31# => romdata <= X"05881108";
    when 16#00B32# => romdata <= X"585A5D53";
    when 16#00B33# => romdata <= X"778C180C";
    when 16#00B34# => romdata <= X"7488180C";
    when 16#00B35# => romdata <= X"7688190C";
    when 16#00B36# => romdata <= X"768C160C";
    when 16#00B37# => romdata <= X"FCF33979";
    when 16#00B38# => romdata <= X"7A101010";
    when 16#00B39# => romdata <= X"8184B805";
    when 16#00B3A# => romdata <= X"7057595D";
    when 16#00B3B# => romdata <= X"8C150857";
    when 16#00B3C# => romdata <= X"76752EA3";
    when 16#00B3D# => romdata <= X"38841708";
    when 16#00B3E# => romdata <= X"FC06707A";
    when 16#00B3F# => romdata <= X"31555673";
    when 16#00B40# => romdata <= X"8F2483CA";
    when 16#00B41# => romdata <= X"38738025";
    when 16#00B42# => romdata <= X"8481388C";
    when 16#00B43# => romdata <= X"17085776";
    when 16#00B44# => romdata <= X"752E0981";
    when 16#00B45# => romdata <= X"06DF3888";
    when 16#00B46# => romdata <= X"15811B70";
    when 16#00B47# => romdata <= X"8306555B";
    when 16#00B48# => romdata <= X"5572C938";
    when 16#00B49# => romdata <= X"7C830653";
    when 16#00B4A# => romdata <= X"72802EFD";
    when 16#00B4B# => romdata <= X"B838FF1D";
    when 16#00B4C# => romdata <= X"F819595D";
    when 16#00B4D# => romdata <= X"88180878";
    when 16#00B4E# => romdata <= X"2EEA38FD";
    when 16#00B4F# => romdata <= X"B539831A";
    when 16#00B50# => romdata <= X"53FC9639";
    when 16#00B51# => romdata <= X"83147082";
    when 16#00B52# => romdata <= X"2C81712B";
    when 16#00B53# => romdata <= X"8184BC08";
    when 16#00B54# => romdata <= X"07708184";
    when 16#00B55# => romdata <= X"B80B8405";
    when 16#00B56# => romdata <= X"0C761010";
    when 16#00B57# => romdata <= X"108184B8";
    when 16#00B58# => romdata <= X"05881108";
    when 16#00B59# => romdata <= X"595B5E51";
    when 16#00B5A# => romdata <= X"53FEE139";
    when 16#00B5B# => romdata <= X"8183FC08";
    when 16#00B5C# => romdata <= X"1758B008";
    when 16#00B5D# => romdata <= X"762E818D";
    when 16#00B5E# => romdata <= X"388184AC";
    when 16#00B5F# => romdata <= X"08FF2E83";
    when 16#00B60# => romdata <= X"EC387376";
    when 16#00B61# => romdata <= X"31188183";
    when 16#00B62# => romdata <= X"FC0C7387";
    when 16#00B63# => romdata <= X"06705753";
    when 16#00B64# => romdata <= X"72802E88";
    when 16#00B65# => romdata <= X"38887331";
    when 16#00B66# => romdata <= X"70155556";
    when 16#00B67# => romdata <= X"76149FFF";
    when 16#00B68# => romdata <= X"06A08071";
    when 16#00B69# => romdata <= X"31177054";
    when 16#00B6A# => romdata <= X"7F535753";
    when 16#00B6B# => romdata <= X"83D53FB0";
    when 16#00B6C# => romdata <= X"0853B008";
    when 16#00B6D# => romdata <= X"FF2E81A0";
    when 16#00B6E# => romdata <= X"388183FC";
    when 16#00B6F# => romdata <= X"08167081";
    when 16#00B70# => romdata <= X"83FC0C74";
    when 16#00B71# => romdata <= X"758184B8";
    when 16#00B72# => romdata <= X"0B88050C";
    when 16#00B73# => romdata <= X"74763118";
    when 16#00B74# => romdata <= X"70810751";
    when 16#00B75# => romdata <= X"5556587B";
    when 16#00B76# => romdata <= X"8184B82E";
    when 16#00B77# => romdata <= X"839C3879";
    when 16#00B78# => romdata <= X"8F2682CB";
    when 16#00B79# => romdata <= X"38810B84";
    when 16#00B7A# => romdata <= X"150C8415";
    when 16#00B7B# => romdata <= X"08FC0670";
    when 16#00B7C# => romdata <= X"7A317A72";
    when 16#00B7D# => romdata <= X"268F7225";
    when 16#00B7E# => romdata <= X"07525553";
    when 16#00B7F# => romdata <= X"72802EFC";
    when 16#00B80# => romdata <= X"F93880DB";
    when 16#00B81# => romdata <= X"39B0089F";
    when 16#00B82# => romdata <= X"FF065372";
    when 16#00B83# => romdata <= X"FEEB3877";
    when 16#00B84# => romdata <= X"8183FC0C";
    when 16#00B85# => romdata <= X"8184B80B";
    when 16#00B86# => romdata <= X"8805087B";
    when 16#00B87# => romdata <= X"18810784";
    when 16#00B88# => romdata <= X"120C5581";
    when 16#00B89# => romdata <= X"84A80878";
    when 16#00B8A# => romdata <= X"27863877";
    when 16#00B8B# => romdata <= X"8184A80C";
    when 16#00B8C# => romdata <= X"8184A408";
    when 16#00B8D# => romdata <= X"7827FCAC";
    when 16#00B8E# => romdata <= X"38778184";
    when 16#00B8F# => romdata <= X"A40C8415";
    when 16#00B90# => romdata <= X"08FC0670";
    when 16#00B91# => romdata <= X"7A317A72";
    when 16#00B92# => romdata <= X"268F7225";
    when 16#00B93# => romdata <= X"07525553";
    when 16#00B94# => romdata <= X"72802EFC";
    when 16#00B95# => romdata <= X"A5388839";
    when 16#00B96# => romdata <= X"80745456";
    when 16#00B97# => romdata <= X"FEDB397D";
    when 16#00B98# => romdata <= X"51829F3F";
    when 16#00B99# => romdata <= X"800BB00C";
    when 16#00B9A# => romdata <= X"8F3D0D04";
    when 16#00B9B# => romdata <= X"73538074";
    when 16#00B9C# => romdata <= X"24A93872";
    when 16#00B9D# => romdata <= X"822C8171";
    when 16#00B9E# => romdata <= X"2B8184BC";
    when 16#00B9F# => romdata <= X"08077081";
    when 16#00BA0# => romdata <= X"84B80B84";
    when 16#00BA1# => romdata <= X"050C5D53";
    when 16#00BA2# => romdata <= X"778C180C";
    when 16#00BA3# => romdata <= X"7488180C";
    when 16#00BA4# => romdata <= X"7688190C";
    when 16#00BA5# => romdata <= X"768C160C";
    when 16#00BA6# => romdata <= X"F9B73983";
    when 16#00BA7# => romdata <= X"1470822C";
    when 16#00BA8# => romdata <= X"81712B81";
    when 16#00BA9# => romdata <= X"84BC0807";
    when 16#00BAA# => romdata <= X"708184B8";
    when 16#00BAB# => romdata <= X"0B84050C";
    when 16#00BAC# => romdata <= X"5E5153D4";
    when 16#00BAD# => romdata <= X"397B7B06";
    when 16#00BAE# => romdata <= X"5372FCA3";
    when 16#00BAF# => romdata <= X"38841A7B";
    when 16#00BB0# => romdata <= X"105C5AF1";
    when 16#00BB1# => romdata <= X"39FF1A81";
    when 16#00BB2# => romdata <= X"11515AF7";
    when 16#00BB3# => romdata <= X"B9397817";
    when 16#00BB4# => romdata <= X"79810784";
    when 16#00BB5# => romdata <= X"190C8C18";
    when 16#00BB6# => romdata <= X"08881908";
    when 16#00BB7# => romdata <= X"718C120C";
    when 16#00BB8# => romdata <= X"88120C59";
    when 16#00BB9# => romdata <= X"708184CC";
    when 16#00BBA# => romdata <= X"0C708184";
    when 16#00BBB# => romdata <= X"C80C8184";
    when 16#00BBC# => romdata <= X"C00B8C12";
    when 16#00BBD# => romdata <= X"0C8C1108";
    when 16#00BBE# => romdata <= X"88120C74";
    when 16#00BBF# => romdata <= X"81078412";
    when 16#00BC0# => romdata <= X"0C741175";
    when 16#00BC1# => romdata <= X"710C5153";
    when 16#00BC2# => romdata <= X"F9BD3975";
    when 16#00BC3# => romdata <= X"17841108";
    when 16#00BC4# => romdata <= X"81078412";
    when 16#00BC5# => romdata <= X"0C538C17";
    when 16#00BC6# => romdata <= X"08881808";
    when 16#00BC7# => romdata <= X"718C120C";
    when 16#00BC8# => romdata <= X"88120C58";
    when 16#00BC9# => romdata <= X"7D5180DA";
    when 16#00BCA# => romdata <= X"3F881754";
    when 16#00BCB# => romdata <= X"F5CF3972";
    when 16#00BCC# => romdata <= X"84150CF4";
    when 16#00BCD# => romdata <= X"1AF80670";
    when 16#00BCE# => romdata <= X"841E0881";
    when 16#00BCF# => romdata <= X"0607841E";
    when 16#00BD0# => romdata <= X"0C701D54";
    when 16#00BD1# => romdata <= X"5B850B84";
    when 16#00BD2# => romdata <= X"140C850B";
    when 16#00BD3# => romdata <= X"88140C8F";
    when 16#00BD4# => romdata <= X"7B27FDCF";
    when 16#00BD5# => romdata <= X"38881C52";
    when 16#00BD6# => romdata <= X"7D518290";
    when 16#00BD7# => romdata <= X"3F8184B8";
    when 16#00BD8# => romdata <= X"0B880508";
    when 16#00BD9# => romdata <= X"8183FC08";
    when 16#00BDA# => romdata <= X"5955FDB7";
    when 16#00BDB# => romdata <= X"39778183";
    when 16#00BDC# => romdata <= X"FC0C7381";
    when 16#00BDD# => romdata <= X"84AC0CFC";
    when 16#00BDE# => romdata <= X"91397284";
    when 16#00BDF# => romdata <= X"150CFDA3";
    when 16#00BE0# => romdata <= X"390404FD";
    when 16#00BE1# => romdata <= X"3D0D800B";
    when 16#00BE2# => romdata <= X"81A5980C";
    when 16#00BE3# => romdata <= X"765186CB";
    when 16#00BE4# => romdata <= X"3FB00853";
    when 16#00BE5# => romdata <= X"B008FF2E";
    when 16#00BE6# => romdata <= X"883872B0";
    when 16#00BE7# => romdata <= X"0C853D0D";
    when 16#00BE8# => romdata <= X"0481A598";
    when 16#00BE9# => romdata <= X"08547380";
    when 16#00BEA# => romdata <= X"2EF03875";
    when 16#00BEB# => romdata <= X"74710C52";
    when 16#00BEC# => romdata <= X"72B00C85";
    when 16#00BED# => romdata <= X"3D0D04FB";
    when 16#00BEE# => romdata <= X"3D0D7770";
    when 16#00BEF# => romdata <= X"5256C23F";
    when 16#00BF0# => romdata <= X"8184B80B";
    when 16#00BF1# => romdata <= X"88050884";
    when 16#00BF2# => romdata <= X"1108FC06";
    when 16#00BF3# => romdata <= X"707B319F";
    when 16#00BF4# => romdata <= X"EF05E080";
    when 16#00BF5# => romdata <= X"06E08005";
    when 16#00BF6# => romdata <= X"565653A0";
    when 16#00BF7# => romdata <= X"80742494";
    when 16#00BF8# => romdata <= X"38805275";
    when 16#00BF9# => romdata <= X"51FF9C3F";
    when 16#00BFA# => romdata <= X"8184C008";
    when 16#00BFB# => romdata <= X"155372B0";
    when 16#00BFC# => romdata <= X"082E8F38";
    when 16#00BFD# => romdata <= X"7551FF8A";
    when 16#00BFE# => romdata <= X"3F805372";
    when 16#00BFF# => romdata <= X"B00C873D";
    when 16#00C00# => romdata <= X"0D047330";
    when 16#00C01# => romdata <= X"527551FE";
    when 16#00C02# => romdata <= X"FA3FB008";
    when 16#00C03# => romdata <= X"FF2EA838";
    when 16#00C04# => romdata <= X"8184B80B";
    when 16#00C05# => romdata <= X"88050875";
    when 16#00C06# => romdata <= X"75318107";
    when 16#00C07# => romdata <= X"84120C53";
    when 16#00C08# => romdata <= X"8183FC08";
    when 16#00C09# => romdata <= X"74318183";
    when 16#00C0A# => romdata <= X"FC0C7551";
    when 16#00C0B# => romdata <= X"FED43F81";
    when 16#00C0C# => romdata <= X"0BB00C87";
    when 16#00C0D# => romdata <= X"3D0D0480";
    when 16#00C0E# => romdata <= X"527551FE";
    when 16#00C0F# => romdata <= X"C63F8184";
    when 16#00C10# => romdata <= X"B80B8805";
    when 16#00C11# => romdata <= X"08B00871";
    when 16#00C12# => romdata <= X"3156538F";
    when 16#00C13# => romdata <= X"7525FFA4";
    when 16#00C14# => romdata <= X"38B00881";
    when 16#00C15# => romdata <= X"84AC0831";
    when 16#00C16# => romdata <= X"8183FC0C";
    when 16#00C17# => romdata <= X"74810784";
    when 16#00C18# => romdata <= X"140C7551";
    when 16#00C19# => romdata <= X"FE9C3F80";
    when 16#00C1A# => romdata <= X"53FF9039";
    when 16#00C1B# => romdata <= X"F63D0D7C";
    when 16#00C1C# => romdata <= X"7E545B72";
    when 16#00C1D# => romdata <= X"802E8283";
    when 16#00C1E# => romdata <= X"387A51FE";
    when 16#00C1F# => romdata <= X"843FF813";
    when 16#00C20# => romdata <= X"84110870";
    when 16#00C21# => romdata <= X"FE067013";
    when 16#00C22# => romdata <= X"841108FC";
    when 16#00C23# => romdata <= X"065D5859";
    when 16#00C24# => romdata <= X"54588184";
    when 16#00C25# => romdata <= X"C008752E";
    when 16#00C26# => romdata <= X"82DE3878";
    when 16#00C27# => romdata <= X"84160C80";
    when 16#00C28# => romdata <= X"73810654";
    when 16#00C29# => romdata <= X"5A727A2E";
    when 16#00C2A# => romdata <= X"81D53878";
    when 16#00C2B# => romdata <= X"15841108";
    when 16#00C2C# => romdata <= X"81065153";
    when 16#00C2D# => romdata <= X"72A03878";
    when 16#00C2E# => romdata <= X"17577981";
    when 16#00C2F# => romdata <= X"E6388815";
    when 16#00C30# => romdata <= X"08537281";
    when 16#00C31# => romdata <= X"84C02E82";
    when 16#00C32# => romdata <= X"F9388C15";
    when 16#00C33# => romdata <= X"08708C15";
    when 16#00C34# => romdata <= X"0C738812";
    when 16#00C35# => romdata <= X"0C567681";
    when 16#00C36# => romdata <= X"0784190C";
    when 16#00C37# => romdata <= X"76187771";
    when 16#00C38# => romdata <= X"0C537981";
    when 16#00C39# => romdata <= X"913883FF";
    when 16#00C3A# => romdata <= X"772781C8";
    when 16#00C3B# => romdata <= X"3876892A";
    when 16#00C3C# => romdata <= X"77832A56";
    when 16#00C3D# => romdata <= X"5372802E";
    when 16#00C3E# => romdata <= X"BF387686";
    when 16#00C3F# => romdata <= X"2AB80555";
    when 16#00C40# => romdata <= X"847327B4";
    when 16#00C41# => romdata <= X"3880DB13";
    when 16#00C42# => romdata <= X"55947327";
    when 16#00C43# => romdata <= X"AB38768C";
    when 16#00C44# => romdata <= X"2A80EE05";
    when 16#00C45# => romdata <= X"5580D473";
    when 16#00C46# => romdata <= X"279E3876";
    when 16#00C47# => romdata <= X"8F2A80F7";
    when 16#00C48# => romdata <= X"055582D4";
    when 16#00C49# => romdata <= X"73279138";
    when 16#00C4A# => romdata <= X"76922A80";
    when 16#00C4B# => romdata <= X"FC05558A";
    when 16#00C4C# => romdata <= X"D4732784";
    when 16#00C4D# => romdata <= X"3880FE55";
    when 16#00C4E# => romdata <= X"74101010";
    when 16#00C4F# => romdata <= X"8184B805";
    when 16#00C50# => romdata <= X"88110855";
    when 16#00C51# => romdata <= X"5673762E";
    when 16#00C52# => romdata <= X"82B33884";
    when 16#00C53# => romdata <= X"1408FC06";
    when 16#00C54# => romdata <= X"53767327";
    when 16#00C55# => romdata <= X"8D388814";
    when 16#00C56# => romdata <= X"08547376";
    when 16#00C57# => romdata <= X"2E098106";
    when 16#00C58# => romdata <= X"EA388C14";
    when 16#00C59# => romdata <= X"08708C1A";
    when 16#00C5A# => romdata <= X"0C74881A";
    when 16#00C5B# => romdata <= X"0C788812";
    when 16#00C5C# => romdata <= X"0C56778C";
    when 16#00C5D# => romdata <= X"150C7A51";
    when 16#00C5E# => romdata <= X"FC883F8C";
    when 16#00C5F# => romdata <= X"3D0D0477";
    when 16#00C60# => romdata <= X"08787131";
    when 16#00C61# => romdata <= X"59770588";
    when 16#00C62# => romdata <= X"19085457";
    when 16#00C63# => romdata <= X"728184C0";
    when 16#00C64# => romdata <= X"2E80E038";
    when 16#00C65# => romdata <= X"8C180870";
    when 16#00C66# => romdata <= X"8C150C73";
    when 16#00C67# => romdata <= X"88120C56";
    when 16#00C68# => romdata <= X"FE893988";
    when 16#00C69# => romdata <= X"15088C16";
    when 16#00C6A# => romdata <= X"08708C13";
    when 16#00C6B# => romdata <= X"0C578817";
    when 16#00C6C# => romdata <= X"0CFEA339";
    when 16#00C6D# => romdata <= X"76832A70";
    when 16#00C6E# => romdata <= X"54558075";
    when 16#00C6F# => romdata <= X"24819838";
    when 16#00C70# => romdata <= X"72822C81";
    when 16#00C71# => romdata <= X"712B8184";
    when 16#00C72# => romdata <= X"BC080781";
    when 16#00C73# => romdata <= X"84B80B84";
    when 16#00C74# => romdata <= X"050C5374";
    when 16#00C75# => romdata <= X"10101081";
    when 16#00C76# => romdata <= X"84B80588";
    when 16#00C77# => romdata <= X"11085556";
    when 16#00C78# => romdata <= X"758C190C";
    when 16#00C79# => romdata <= X"7388190C";
    when 16#00C7A# => romdata <= X"7788170C";
    when 16#00C7B# => romdata <= X"778C150C";
    when 16#00C7C# => romdata <= X"FF843981";
    when 16#00C7D# => romdata <= X"5AFDB439";
    when 16#00C7E# => romdata <= X"78177381";
    when 16#00C7F# => romdata <= X"06545772";
    when 16#00C80# => romdata <= X"98387708";
    when 16#00C81# => romdata <= X"78713159";
    when 16#00C82# => romdata <= X"77058C19";
    when 16#00C83# => romdata <= X"08881A08";
    when 16#00C84# => romdata <= X"718C120C";
    when 16#00C85# => romdata <= X"88120C57";
    when 16#00C86# => romdata <= X"57768107";
    when 16#00C87# => romdata <= X"84190C77";
    when 16#00C88# => romdata <= X"8184B80B";
    when 16#00C89# => romdata <= X"88050C81";
    when 16#00C8A# => romdata <= X"84B40877";
    when 16#00C8B# => romdata <= X"26FEC738";
    when 16#00C8C# => romdata <= X"8184B008";
    when 16#00C8D# => romdata <= X"527A51FA";
    when 16#00C8E# => romdata <= X"FE3F7A51";
    when 16#00C8F# => romdata <= X"FAC43FFE";
    when 16#00C90# => romdata <= X"BA398178";
    when 16#00C91# => romdata <= X"8C150C78";
    when 16#00C92# => romdata <= X"88150C73";
    when 16#00C93# => romdata <= X"8C1A0C73";
    when 16#00C94# => romdata <= X"881A0C5A";
    when 16#00C95# => romdata <= X"FD803983";
    when 16#00C96# => romdata <= X"1570822C";
    when 16#00C97# => romdata <= X"81712B81";
    when 16#00C98# => romdata <= X"84BC0807";
    when 16#00C99# => romdata <= X"8184B80B";
    when 16#00C9A# => romdata <= X"84050C51";
    when 16#00C9B# => romdata <= X"53741010";
    when 16#00C9C# => romdata <= X"108184B8";
    when 16#00C9D# => romdata <= X"05881108";
    when 16#00C9E# => romdata <= X"5556FEE4";
    when 16#00C9F# => romdata <= X"39745380";
    when 16#00CA0# => romdata <= X"7524A738";
    when 16#00CA1# => romdata <= X"72822C81";
    when 16#00CA2# => romdata <= X"712B8184";
    when 16#00CA3# => romdata <= X"BC080781";
    when 16#00CA4# => romdata <= X"84B80B84";
    when 16#00CA5# => romdata <= X"050C5375";
    when 16#00CA6# => romdata <= X"8C190C73";
    when 16#00CA7# => romdata <= X"88190C77";
    when 16#00CA8# => romdata <= X"88170C77";
    when 16#00CA9# => romdata <= X"8C150CFD";
    when 16#00CAA# => romdata <= X"CD398315";
    when 16#00CAB# => romdata <= X"70822C81";
    when 16#00CAC# => romdata <= X"712B8184";
    when 16#00CAD# => romdata <= X"BC080781";
    when 16#00CAE# => romdata <= X"84B80B84";
    when 16#00CAF# => romdata <= X"050C5153";
    when 16#00CB0# => romdata <= X"D639810B";
    when 16#00CB1# => romdata <= X"B00C0480";
    when 16#00CB2# => romdata <= X"3D0D7281";
    when 16#00CB3# => romdata <= X"2E893880";
    when 16#00CB4# => romdata <= X"0BB00C82";
    when 16#00CB5# => romdata <= X"3D0D0473";
    when 16#00CB6# => romdata <= X"51B23FFE";
    when 16#00CB7# => romdata <= X"3D0D81A5";
    when 16#00CB8# => romdata <= X"94085170";
    when 16#00CB9# => romdata <= X"8A3881A5";
    when 16#00CBA# => romdata <= X"9C7081A5";
    when 16#00CBB# => romdata <= X"940C5170";
    when 16#00CBC# => romdata <= X"75125252";
    when 16#00CBD# => romdata <= X"FF537087";
    when 16#00CBE# => romdata <= X"FB808026";
    when 16#00CBF# => romdata <= X"88387081";
    when 16#00CC0# => romdata <= X"A5940C71";
    when 16#00CC1# => romdata <= X"5372B00C";
    when 16#00CC2# => romdata <= X"843D0D04";
    when 16#00CC3# => romdata <= X"00FF3900";
    when 16#00CC4# => romdata <= X"68656C70";
    when 16#00CC5# => romdata <= X"00000000";
    when 16#00CC6# => romdata <= X"73797374";
    when 16#00CC7# => romdata <= X"656D2072";
    when 16#00CC8# => romdata <= X"65736574";
    when 16#00CC9# => romdata <= X"00000000";
    when 16#00CCA# => romdata <= X"72657365";
    when 16#00CCB# => romdata <= X"74000000";
    when 16#00CCC# => romdata <= X"73686F77";
    when 16#00CCD# => romdata <= X"20737973";
    when 16#00CCE# => romdata <= X"74656D20";
    when 16#00CCF# => romdata <= X"696E666F";
    when 16#00CD0# => romdata <= X"203C7665";
    when 16#00CD1# => romdata <= X"72626F73";
    when 16#00CD2# => romdata <= X"653E0000";
    when 16#00CD3# => romdata <= X"73797369";
    when 16#00CD4# => romdata <= X"6E666F00";
    when 16#00CD5# => romdata <= X"7265706F";
    when 16#00CD6# => romdata <= X"72742076";
    when 16#00CD7# => romdata <= X"65727369";
    when 16#00CD8# => romdata <= X"6F6E0000";
    when 16#00CD9# => romdata <= X"76657273";
    when 16#00CDA# => romdata <= X"696F6E00";
    when 16#00CDB# => romdata <= X"72656E61";
    when 16#00CDC# => romdata <= X"20636F6E";
    when 16#00CDD# => romdata <= X"74726F6C";
    when 16#00CDE# => romdata <= X"6C657220";
    when 16#00CDF# => romdata <= X"73746174";
    when 16#00CE0# => romdata <= X"75730000";
    when 16#00CE1# => romdata <= X"72656E61";
    when 16#00CE2# => romdata <= X"20737461";
    when 16#00CE3# => romdata <= X"74757300";
    when 16#00CE4# => romdata <= X"3C636861";
    when 16#00CE5# => romdata <= X"6E6E656C";
    when 16#00CE6# => romdata <= X"3E203C68";
    when 16#00CE7# => romdata <= X"6967683E";
    when 16#00CE8# => romdata <= X"203C6C6F";
    when 16#00CE9# => romdata <= X"775F636F";
    when 16#00CEA# => romdata <= X"6E666967";
    when 16#00CEB# => romdata <= X"3E000000";
    when 16#00CEC# => romdata <= X"636F6E66";
    when 16#00CED# => romdata <= X"69670000";
    when 16#00CEE# => romdata <= X"646F2063";
    when 16#00CEF# => romdata <= X"6F6D706C";
    when 16#00CF0# => romdata <= X"65746520";
    when 16#00CF1# => romdata <= X"64656D6F";
    when 16#00CF2# => romdata <= X"20636F6E";
    when 16#00CF3# => romdata <= X"66696720";
    when 16#00CF4# => romdata <= X"666F7220";
    when 16#00CF5# => romdata <= X"52454E41";
    when 16#00CF6# => romdata <= X"00000000";
    when 16#00CF7# => romdata <= X"64656D6F";
    when 16#00CF8# => romdata <= X"00000000";
    when 16#00CF9# => romdata <= X"73657420";
    when 16#00CFA# => romdata <= X"52454E41";
    when 16#00CFB# => romdata <= X"20746F20";
    when 16#00CFC# => romdata <= X"706F7765";
    when 16#00CFD# => romdata <= X"7220646F";
    when 16#00CFE# => romdata <= X"776E206D";
    when 16#00CFF# => romdata <= X"6F646500";
    when 16#00D00# => romdata <= X"706F6666";
    when 16#00D01# => romdata <= X"00000000";
    when 16#00D02# => romdata <= X"73657420";
    when 16#00D03# => romdata <= X"72656E61";
    when 16#00D04# => romdata <= X"20636861";
    when 16#00D05# => romdata <= X"6E6E656C";
    when 16#00D06# => romdata <= X"20302074";
    when 16#00D07# => romdata <= X"6F20666F";
    when 16#00D08# => romdata <= X"6C6C6F77";
    when 16#00D09# => romdata <= X"6572206D";
    when 16#00D0A# => romdata <= X"6F646500";
    when 16#00D0B# => romdata <= X"666F6C6C";
    when 16#00D0C# => romdata <= X"6F770000";
    when 16#00D0D# => romdata <= X"3C74696D";
    when 16#00D0E# => romdata <= X"653E2061";
    when 16#00D0F# => romdata <= X"63746976";
    when 16#00D10# => romdata <= X"61746520";
    when 16#00D11# => romdata <= X"52454E41";
    when 16#00D12# => romdata <= X"00000000";
    when 16#00D13# => romdata <= X"61637175";
    when 16#00D14# => romdata <= X"69726500";
    when 16#00D15# => romdata <= X"73657420";
    when 16#00D16# => romdata <= X"52454E41";
    when 16#00D17# => romdata <= X"20636F6E";
    when 16#00D18# => romdata <= X"74726F6C";
    when 16#00D19# => romdata <= X"6C657220";
    when 16#00D1A# => romdata <= X"746F2049";
    when 16#00D1B# => romdata <= X"444C4500";
    when 16#00D1C# => romdata <= X"73746F70";
    when 16#00D1D# => romdata <= X"00000000";
    when 16#00D1E# => romdata <= X"7072696E";
    when 16#00D1F# => romdata <= X"74207472";
    when 16#00D20# => romdata <= X"69676765";
    when 16#00D21# => romdata <= X"72206368";
    when 16#00D22# => romdata <= X"61696E73";
    when 16#00D23# => romdata <= X"00000000";
    when 16#00D24# => romdata <= X"63686169";
    when 16#00D25# => romdata <= X"6E730000";
    when 16#00D26# => romdata <= X"7072696E";
    when 16#00D27# => romdata <= X"74207361";
    when 16#00D28# => romdata <= X"6D706C65";
    when 16#00D29# => romdata <= X"64205245";
    when 16#00D2A# => romdata <= X"4E412074";
    when 16#00D2B# => romdata <= X"6F6B656E";
    when 16#00D2C# => romdata <= X"73000000";
    when 16#00D2D# => romdata <= X"746F6B65";
    when 16#00D2E# => romdata <= X"6E000000";
    when 16#00D2F# => romdata <= X"74726F75";
    when 16#00D30# => romdata <= X"626C6573";
    when 16#00D31# => romdata <= X"65617263";
    when 16#00D32# => romdata <= X"68205245";
    when 16#00D33# => romdata <= X"4E410000";
    when 16#00D34# => romdata <= X"74726F75";
    when 16#00D35# => romdata <= X"626C6500";
    when 16#00D36# => romdata <= X"696E6974";
    when 16#00D37# => romdata <= X"616C697A";
    when 16#00D38# => romdata <= X"65204444";
    when 16#00D39# => romdata <= X"53206368";
    when 16#00D3A# => romdata <= X"6970203C";
    when 16#00D3B# => romdata <= X"66726571";
    when 16#00D3C# => romdata <= X"2074756E";
    when 16#00D3D# => romdata <= X"696E6720";
    when 16#00D3E# => romdata <= X"776F7264";
    when 16#00D3F# => romdata <= X"3E000000";
    when 16#00D40# => romdata <= X"64647369";
    when 16#00D41# => romdata <= X"6E697400";
    when 16#00D42# => romdata <= X"72656164";
    when 16#00D43# => romdata <= X"20646473";
    when 16#00D44# => romdata <= X"20726567";
    when 16#00D45# => romdata <= X"69737465";
    when 16#00D46# => romdata <= X"72730000";
    when 16#00D47# => romdata <= X"64647369";
    when 16#00D48# => romdata <= X"6E666F00";
    when 16#00D49# => romdata <= X"72756E6E";
    when 16#00D4A# => romdata <= X"696E6720";
    when 16#00D4B# => romdata <= X"6C696768";
    when 16#00D4C# => romdata <= X"74000000";
    when 16#00D4D# => romdata <= X"72756E00";
    when 16#00D4E# => romdata <= X"63686563";
    when 16#00D4F# => romdata <= X"6B204932";
    when 16#00D50# => romdata <= X"43206164";
    when 16#00D51# => romdata <= X"64726573";
    when 16#00D52# => romdata <= X"73000000";
    when 16#00D53# => romdata <= X"69326300";
    when 16#00D54# => romdata <= X"72656164";
    when 16#00D55# => romdata <= X"20454550";
    when 16#00D56# => romdata <= X"524F4D20";
    when 16#00D57# => romdata <= X"3C627573";
    when 16#00D58# => romdata <= X"3E203C69";
    when 16#00D59# => romdata <= X"32635F61";
    when 16#00D5A# => romdata <= X"6464723E";
    when 16#00D5B# => romdata <= X"203C6C65";
    when 16#00D5C# => romdata <= X"6E677468";
    when 16#00D5D# => romdata <= X"3E000000";
    when 16#00D5E# => romdata <= X"65657072";
    when 16#00D5F# => romdata <= X"6F6D0000";
    when 16#00D60# => romdata <= X"72656164";
    when 16#00D61# => romdata <= X"20616463";
    when 16#00D62# => romdata <= X"2076616C";
    when 16#00D63# => romdata <= X"75650000";
    when 16#00D64# => romdata <= X"61646300";
    when 16#00D65# => romdata <= X"67656E65";
    when 16#00D66# => romdata <= X"72617465";
    when 16#00D67# => romdata <= X"20746573";
    when 16#00D68# => romdata <= X"7420696D";
    when 16#00D69# => romdata <= X"70756C73";
    when 16#00D6A# => romdata <= X"65000000";
    when 16#00D6B# => romdata <= X"74657374";
    when 16#00D6C# => romdata <= X"67656E00";
    when 16#00D6D# => romdata <= X"616C6961";
    when 16#00D6E# => romdata <= X"7320666F";
    when 16#00D6F# => romdata <= X"72207800";
    when 16#00D70# => romdata <= X"6D656D00";
    when 16#00D71# => romdata <= X"77726974";
    when 16#00D72# => romdata <= X"6520776F";
    when 16#00D73# => romdata <= X"7264203C";
    when 16#00D74# => romdata <= X"61646472";
    when 16#00D75# => romdata <= X"3E203C6C";
    when 16#00D76# => romdata <= X"656E6774";
    when 16#00D77# => romdata <= X"683E203C";
    when 16#00D78# => romdata <= X"76616C75";
    when 16#00D79# => romdata <= X"65287329";
    when 16#00D7A# => romdata <= X"3E000000";
    when 16#00D7B# => romdata <= X"776D656D";
    when 16#00D7C# => romdata <= X"00000000";
    when 16#00D7D# => romdata <= X"6558616D";
    when 16#00D7E# => romdata <= X"696E6520";
    when 16#00D7F# => romdata <= X"6D656D6F";
    when 16#00D80# => romdata <= X"7279203C";
    when 16#00D81# => romdata <= X"61646472";
    when 16#00D82# => romdata <= X"3E203C6C";
    when 16#00D83# => romdata <= X"656E6774";
    when 16#00D84# => romdata <= X"683E0000";
    when 16#00D85# => romdata <= X"78000000";
    when 16#00D86# => romdata <= X"636C6561";
    when 16#00D87# => romdata <= X"72207363";
    when 16#00D88# => romdata <= X"7265656E";
    when 16#00D89# => romdata <= X"00000000";
    when 16#00D8A# => romdata <= X"636C6561";
    when 16#00D8B# => romdata <= X"72000000";
    when 16#00D8C# => romdata <= X"0A0A0000";
    when 16#00D8D# => romdata <= X"72656E61";
    when 16#00D8E# => romdata <= X"3320636F";
    when 16#00D8F# => romdata <= X"6E74726F";
    when 16#00D90# => romdata <= X"6C6C6572";
    when 16#00D91# => romdata <= X"20626F61";
    when 16#00D92# => romdata <= X"72640000";
    when 16#00D93# => romdata <= X"20286F6E";
    when 16#00D94# => romdata <= X"2073696D";
    when 16#00D95# => romdata <= X"290A0000";
    when 16#00D96# => romdata <= X"0A485720";
    when 16#00D97# => romdata <= X"73796E74";
    when 16#00D98# => romdata <= X"68657369";
    when 16#00D99# => romdata <= X"7A65643A";
    when 16#00D9A# => romdata <= X"20000000";
    when 16#00D9B# => romdata <= X"0A535720";
    when 16#00D9C# => romdata <= X"636F6D70";
    when 16#00D9D# => romdata <= X"696C6564";
    when 16#00D9E# => romdata <= X"2020203A";
    when 16#00D9F# => romdata <= X"204A616E";
    when 16#00DA0# => romdata <= X"20203220";
    when 16#00DA1# => romdata <= X"32303132";
    when 16#00DA2# => romdata <= X"20203134";
    when 16#00DA3# => romdata <= X"3A32313A";
    when 16#00DA4# => romdata <= X"30320000";
    when 16#00DA5# => romdata <= X"0A737973";
    when 16#00DA6# => romdata <= X"74656D20";
    when 16#00DA7# => romdata <= X"636C6F63";
    when 16#00DA8# => romdata <= X"6B20203A";
    when 16#00DA9# => romdata <= X"20000000";
    when 16#00DAA# => romdata <= X"204D487A";
    when 16#00DAB# => romdata <= X"0A000000";
    when 16#00DAC# => romdata <= X"44454255";
    when 16#00DAD# => romdata <= X"47204D4F";
    when 16#00DAE# => romdata <= X"44450000";
    when 16#00DAF# => romdata <= X"204F4E0A";
    when 16#00DB0# => romdata <= X"00000000";
    when 16#00DB1# => romdata <= X"56312E30";
    when 16#00DB2# => romdata <= X"2D31322E";
    when 16#00DB3# => romdata <= X"32303131";
    when 16#00DB4# => romdata <= X"5F524F45";
    when 16#00DB5# => romdata <= X"5F5A5055";
    when 16#00DB6# => romdata <= X"00000000";
    when 16#00DB7# => romdata <= X"4552524F";
    when 16#00DB8# => romdata <= X"523A2074";
    when 16#00DB9# => romdata <= X"6F6F206D";
    when 16#00DBA# => romdata <= X"75636820";
    when 16#00DBB# => romdata <= X"636F6D6D";
    when 16#00DBC# => romdata <= X"616E6473";
    when 16#00DBD# => romdata <= X"2E0A0000";
    when 16#00DBE# => romdata <= X"3E200000";
    when 16#00DBF# => romdata <= X"636F6D6D";
    when 16#00DC0# => romdata <= X"616E6420";
    when 16#00DC1# => romdata <= X"6E6F7420";
    when 16#00DC2# => romdata <= X"666F756E";
    when 16#00DC3# => romdata <= X"642E0A00";
    when 16#00DC4# => romdata <= X"73757070";
    when 16#00DC5# => romdata <= X"6F727465";
    when 16#00DC6# => romdata <= X"6420636F";
    when 16#00DC7# => romdata <= X"6D6D616E";
    when 16#00DC8# => romdata <= X"64733A0A";
    when 16#00DC9# => romdata <= X"0A000000";
    when 16#00DCA# => romdata <= X"202D2000";
    when 16#00DCB# => romdata <= X"76656E64";
    when 16#00DCC# => romdata <= X"6F723F20";
    when 16#00DCD# => romdata <= X"20000000";
    when 16#00DCE# => romdata <= X"485A4452";
    when 16#00DCF# => romdata <= X"20202020";
    when 16#00DD0# => romdata <= X"20000000";
    when 16#00DD1# => romdata <= X"67616973";
    when 16#00DD2# => romdata <= X"6C657220";
    when 16#00DD3# => romdata <= X"20000000";
    when 16#00DD4# => romdata <= X"45534120";
    when 16#00DD5# => romdata <= X"20202020";
    when 16#00DD6# => romdata <= X"20000000";
    when 16#00DD7# => romdata <= X"756E6B6E";
    when 16#00DD8# => romdata <= X"6F776E20";
    when 16#00DD9# => romdata <= X"64657669";
    when 16#00DDA# => romdata <= X"63650000";
    when 16#00DDB# => romdata <= X"4C656F6E";
    when 16#00DDC# => romdata <= X"32204D65";
    when 16#00DDD# => romdata <= X"6D6F7279";
    when 16#00DDE# => romdata <= X"20436F6E";
    when 16#00DDF# => romdata <= X"74726F6C";
    when 16#00DE0# => romdata <= X"6C657200";
    when 16#00DE1# => romdata <= X"56474120";
    when 16#00DE2# => romdata <= X"636F6E74";
    when 16#00DE3# => romdata <= X"726F6C6C";
    when 16#00DE4# => romdata <= X"65720000";
    when 16#00DE5# => romdata <= X"53504920";
    when 16#00DE6# => romdata <= X"4D656D6F";
    when 16#00DE7# => romdata <= X"72792043";
    when 16#00DE8# => romdata <= X"6F6E7472";
    when 16#00DE9# => romdata <= X"6F6C6C65";
    when 16#00DEA# => romdata <= X"72000000";
    when 16#00DEB# => romdata <= X"53504920";
    when 16#00DEC# => romdata <= X"436F6E74";
    when 16#00DED# => romdata <= X"726F6C6C";
    when 16#00DEE# => romdata <= X"65720000";
    when 16#00DEF# => romdata <= X"414D4241";
    when 16#00DF0# => romdata <= X"20577261";
    when 16#00DF1# => romdata <= X"70706572";
    when 16#00DF2# => romdata <= X"20666F72";
    when 16#00DF3# => romdata <= X"204F4320";
    when 16#00DF4# => romdata <= X"4932432D";
    when 16#00DF5# => romdata <= X"6D617374";
    when 16#00DF6# => romdata <= X"65720000";
    when 16#00DF7# => romdata <= X"47522031";
    when 16#00DF8# => romdata <= X"302F3130";
    when 16#00DF9# => romdata <= X"30204D62";
    when 16#00DFA# => romdata <= X"69742045";
    when 16#00DFB# => romdata <= X"74686572";
    when 16#00DFC# => romdata <= X"6E657420";
    when 16#00DFD# => romdata <= X"4D414300";
    when 16#00DFE# => romdata <= X"47656E65";
    when 16#00DFF# => romdata <= X"72616C20";
    when 16#00E00# => romdata <= X"50757270";
    when 16#00E01# => romdata <= X"6F736520";
    when 16#00E02# => romdata <= X"492F4F20";
    when 16#00E03# => romdata <= X"706F7274";
    when 16#00E04# => romdata <= X"00000000";
    when 16#00E05# => romdata <= X"4D6F6475";
    when 16#00E06# => romdata <= X"6C617220";
    when 16#00E07# => romdata <= X"54696D65";
    when 16#00E08# => romdata <= X"7220556E";
    when 16#00E09# => romdata <= X"69740000";
    when 16#00E0A# => romdata <= X"4475616C";
    when 16#00E0B# => romdata <= X"2D706F72";
    when 16#00E0C# => romdata <= X"74204148";
    when 16#00E0D# => romdata <= X"42205352";
    when 16#00E0E# => romdata <= X"414D206D";
    when 16#00E0F# => romdata <= X"6F64756C";
    when 16#00E10# => romdata <= X"65000000";
    when 16#00E11# => romdata <= X"47656E65";
    when 16#00E12# => romdata <= X"72696320";
    when 16#00E13# => romdata <= X"55415254";
    when 16#00E14# => romdata <= X"00000000";
    when 16#00E15# => romdata <= X"4148422F";
    when 16#00E16# => romdata <= X"41504220";
    when 16#00E17# => romdata <= X"42726964";
    when 16#00E18# => romdata <= X"67650000";
    when 16#00E19# => romdata <= X"64696666";
    when 16#00E1A# => romdata <= X"6572656E";
    when 16#00E1B# => romdata <= X"7469616C";
    when 16#00E1C# => romdata <= X"20637572";
    when 16#00E1D# => romdata <= X"72656E74";
    when 16#00E1E# => romdata <= X"206D6F6E";
    when 16#00E1F# => romdata <= X"69746F72";
    when 16#00E20# => romdata <= X"00000000";
    when 16#00E21# => romdata <= X"64656275";
    when 16#00E22# => romdata <= X"67207472";
    when 16#00E23# => romdata <= X"61636572";
    when 16#00E24# => romdata <= X"206D656D";
    when 16#00E25# => romdata <= X"6F727900";
    when 16#00E26# => romdata <= X"4541444F";
    when 16#00E27# => romdata <= X"47533130";
    when 16#00E28# => romdata <= X"32206469";
    when 16#00E29# => romdata <= X"73706C61";
    when 16#00E2A# => romdata <= X"79206472";
    when 16#00E2B# => romdata <= X"69766572";
    when 16#00E2C# => romdata <= X"00000000";
    when 16#00E2D# => romdata <= X"64656275";
    when 16#00E2E# => romdata <= X"67206275";
    when 16#00E2F# => romdata <= X"66666572";
    when 16#00E30# => romdata <= X"20636F6E";
    when 16#00E31# => romdata <= X"74726F6C";
    when 16#00E32# => romdata <= X"00000000";
    when 16#00E33# => romdata <= X"52454E41";
    when 16#00E34# => romdata <= X"3320636F";
    when 16#00E35# => romdata <= X"6E74726F";
    when 16#00E36# => romdata <= X"6C6C6572";
    when 16#00E37# => romdata <= X"00000000";
    when 16#00E38# => romdata <= X"53465020";
    when 16#00E39# => romdata <= X"636F6E74";
    when 16#00E3A# => romdata <= X"726F6C6C";
    when 16#00E3B# => romdata <= X"65720000";
    when 16#00E3C# => romdata <= X"5A505520";
    when 16#00E3D# => romdata <= X"4D656D6F";
    when 16#00E3E# => romdata <= X"72792077";
    when 16#00E3F# => romdata <= X"72617070";
    when 16#00E40# => romdata <= X"65720000";
    when 16#00E41# => romdata <= X"5A505520";
    when 16#00E42# => romdata <= X"41484220";
    when 16#00E43# => romdata <= X"57726170";
    when 16#00E44# => romdata <= X"70657200";
    when 16#00E45# => romdata <= X"6265616D";
    when 16#00E46# => romdata <= X"20706F73";
    when 16#00E47# => romdata <= X"6974696F";
    when 16#00E48# => romdata <= X"6E206D6F";
    when 16#00E49# => romdata <= X"6E69746F";
    when 16#00E4A# => romdata <= X"72000000";
    when 16#00E4B# => romdata <= X"74726967";
    when 16#00E4C# => romdata <= X"67657220";
    when 16#00E4D# => romdata <= X"67656E65";
    when 16#00E4E# => romdata <= X"7261746F";
    when 16#00E4F# => romdata <= X"72000000";
    when 16#00E50# => romdata <= X"64656275";
    when 16#00E51# => romdata <= X"6720636F";
    when 16#00E52# => romdata <= X"6E736F6C";
    when 16#00E53# => romdata <= X"65000000";
    when 16#00E54# => romdata <= X"44434D20";
    when 16#00E55# => romdata <= X"70686173";
    when 16#00E56# => romdata <= X"65207368";
    when 16#00E57# => romdata <= X"69667420";
    when 16#00E58# => romdata <= X"636F6E74";
    when 16#00E59# => romdata <= X"726F6C00";
    when 16#00E5A# => romdata <= X"20206170";
    when 16#00E5B# => romdata <= X"62736C76";
    when 16#00E5C# => romdata <= X"00000000";
    when 16#00E5D# => romdata <= X"76656E64";
    when 16#00E5E# => romdata <= X"20307800";
    when 16#00E5F# => romdata <= X"64657620";
    when 16#00E60# => romdata <= X"30780000";
    when 16#00E61# => romdata <= X"76657220";
    when 16#00E62# => romdata <= X"00000000";
    when 16#00E63# => romdata <= X"69727120";
    when 16#00E64# => romdata <= X"00000000";
    when 16#00E65# => romdata <= X"61646472";
    when 16#00E66# => romdata <= X"20307800";
    when 16#00E67# => romdata <= X"6168626D";
    when 16#00E68# => romdata <= X"73740000";
    when 16#00E69# => romdata <= X"61686273";
    when 16#00E6A# => romdata <= X"6C760000";
    when 16#00E6B# => romdata <= X"00000F71";
    when 16#00E6C# => romdata <= X"00001042";
    when 16#00E6D# => romdata <= X"00001037";
    when 16#00E6E# => romdata <= X"0000106E";
    when 16#00E6F# => romdata <= X"00001063";
    when 16#00E70# => romdata <= X"00001058";
    when 16#00E71# => romdata <= X"0000104D";
    when 16#00E72# => romdata <= X"00001016";
    when 16#00E73# => romdata <= X"0000100B";
    when 16#00E74# => romdata <= X"00001000";
    when 16#00E75# => romdata <= X"00000FF5";
    when 16#00E76# => romdata <= X"0000102C";
    when 16#00E77# => romdata <= X"00001021";
    when 16#00E78# => romdata <= X"00000FEA";
    when 16#00E79# => romdata <= X"00000F71";
    when 16#00E7A# => romdata <= X"00000F71";
    when 16#00E7B# => romdata <= X"00000F71";
    when 16#00E7C# => romdata <= X"00000F71";
    when 16#00E7D# => romdata <= X"00000F71";
    when 16#00E7E# => romdata <= X"00000FDF";
    when 16#00E7F# => romdata <= X"00000F71";
    when 16#00E80# => romdata <= X"00000F71";
    when 16#00E81# => romdata <= X"00000FD4";
    when 16#00E82# => romdata <= X"00000F71";
    when 16#00E83# => romdata <= X"00000FC9";
    when 16#00E84# => romdata <= X"00000F71";
    when 16#00E85# => romdata <= X"00000F71";
    when 16#00E86# => romdata <= X"00000F71";
    when 16#00E87# => romdata <= X"00000F71";
    when 16#00E88# => romdata <= X"00000F71";
    when 16#00E89# => romdata <= X"00000F71";
    when 16#00E8A# => romdata <= X"00000F71";
    when 16#00E8B# => romdata <= X"00000F71";
    when 16#00E8C# => romdata <= X"00000FBE";
    when 16#00E8D# => romdata <= X"00000F71";
    when 16#00E8E# => romdata <= X"00000F71";
    when 16#00E8F# => romdata <= X"00000FB3";
    when 16#00E90# => romdata <= X"00000F71";
    when 16#00E91# => romdata <= X"00000F71";
    when 16#00E92# => romdata <= X"00000F71";
    when 16#00E93# => romdata <= X"00000F71";
    when 16#00E94# => romdata <= X"00000F71";
    when 16#00E95# => romdata <= X"00000F71";
    when 16#00E96# => romdata <= X"00000F71";
    when 16#00E97# => romdata <= X"00000F71";
    when 16#00E98# => romdata <= X"00000F71";
    when 16#00E99# => romdata <= X"00000F71";
    when 16#00E9A# => romdata <= X"00000FA8";
    when 16#00E9B# => romdata <= X"00000F71";
    when 16#00E9C# => romdata <= X"00000F71";
    when 16#00E9D# => romdata <= X"00000F71";
    when 16#00E9E# => romdata <= X"00000F71";
    when 16#00E9F# => romdata <= X"00000F9D";
    when 16#00EA0# => romdata <= X"00000F71";
    when 16#00EA1# => romdata <= X"00000F71";
    when 16#00EA2# => romdata <= X"00000F71";
    when 16#00EA3# => romdata <= X"00000F71";
    when 16#00EA4# => romdata <= X"00000F71";
    when 16#00EA5# => romdata <= X"00000F71";
    when 16#00EA6# => romdata <= X"00000F71";
    when 16#00EA7# => romdata <= X"00000F71";
    when 16#00EA8# => romdata <= X"00000F71";
    when 16#00EA9# => romdata <= X"00000F71";
    when 16#00EAA# => romdata <= X"00000F71";
    when 16#00EAB# => romdata <= X"00000F71";
    when 16#00EAC# => romdata <= X"00000F71";
    when 16#00EAD# => romdata <= X"00000F71";
    when 16#00EAE# => romdata <= X"00000F71";
    when 16#00EAF# => romdata <= X"00000F71";
    when 16#00EB0# => romdata <= X"00000F71";
    when 16#00EB1# => romdata <= X"00000F71";
    when 16#00EB2# => romdata <= X"00000F71";
    when 16#00EB3# => romdata <= X"00000F71";
    when 16#00EB4# => romdata <= X"00000F71";
    when 16#00EB5# => romdata <= X"00000F71";
    when 16#00EB6# => romdata <= X"00000F71";
    when 16#00EB7# => romdata <= X"00000F92";
    when 16#00EB8# => romdata <= X"00000F71";
    when 16#00EB9# => romdata <= X"00000F71";
    when 16#00EBA# => romdata <= X"00000F71";
    when 16#00EBB# => romdata <= X"00000F71";
    when 16#00EBC# => romdata <= X"00000F71";
    when 16#00EBD# => romdata <= X"00000F71";
    when 16#00EBE# => romdata <= X"00000F71";
    when 16#00EBF# => romdata <= X"00000F71";
    when 16#00EC0# => romdata <= X"00000F71";
    when 16#00EC1# => romdata <= X"00000F71";
    when 16#00EC2# => romdata <= X"00000F71";
    when 16#00EC3# => romdata <= X"00000F71";
    when 16#00EC4# => romdata <= X"00000F71";
    when 16#00EC5# => romdata <= X"00000F71";
    when 16#00EC6# => romdata <= X"00000F71";
    when 16#00EC7# => romdata <= X"00000F71";
    when 16#00EC8# => romdata <= X"00000F71";
    when 16#00EC9# => romdata <= X"00000F71";
    when 16#00ECA# => romdata <= X"00000F71";
    when 16#00ECB# => romdata <= X"00000F71";
    when 16#00ECC# => romdata <= X"00000F71";
    when 16#00ECD# => romdata <= X"00000F71";
    when 16#00ECE# => romdata <= X"00000F71";
    when 16#00ECF# => romdata <= X"00000F71";
    when 16#00ED0# => romdata <= X"00000F71";
    when 16#00ED1# => romdata <= X"00000F71";
    when 16#00ED2# => romdata <= X"00000F71";
    when 16#00ED3# => romdata <= X"00000F87";
    when 16#00ED4# => romdata <= X"69326320";
    when 16#00ED5# => romdata <= X"464D430A";
    when 16#00ED6# => romdata <= X"00000000";
    when 16#00ED7# => romdata <= X"61646472";
    when 16#00ED8# => romdata <= X"6573733A";
    when 16#00ED9# => romdata <= X"20307800";
    when 16#00EDA# => romdata <= X"2020202D";
    when 16#00EDB# => romdata <= X"2D3E2020";
    when 16#00EDC# => romdata <= X"2041434B";
    when 16#00EDD# => romdata <= X"0A000000";
    when 16#00EDE# => romdata <= X"72656164";
    when 16#00EDF# => romdata <= X"20646174";
    when 16#00EE0# => romdata <= X"61202800";
    when 16#00EE1# => romdata <= X"20627974";
    when 16#00EE2# => romdata <= X"65732920";
    when 16#00EE3# => romdata <= X"66726F6D";
    when 16#00EE4# => romdata <= X"20493243";
    when 16#00EE5# => romdata <= X"2D616464";
    when 16#00EE6# => romdata <= X"72657373";
    when 16#00EE7# => romdata <= X"20307800";
    when 16#00EE8# => romdata <= X"0A307800";
    when 16#00EE9# => romdata <= X"02020606";
    when 16#00EEA# => romdata <= X"06040304";
    when 16#00EEB# => romdata <= X"02020102";
    when 16#00EEC# => romdata <= X"636F6E74";
    when 16#00EED# => romdata <= X"726F6C20";
    when 16#00EEE# => romdata <= X"2020203A";
    when 16#00EEF# => romdata <= X"20000000";
    when 16#00EF0# => romdata <= X"66726571";
    when 16#00EF1# => romdata <= X"75656E63";
    when 16#00EF2# => romdata <= X"7920203A";
    when 16#00EF3# => romdata <= X"20000000";
    when 16#00EF4# => romdata <= X"75706461";
    when 16#00EF5# => romdata <= X"74652063";
    when 16#00EF6# => romdata <= X"6C6B203A";
    when 16#00EF7# => romdata <= X"20000000";
    when 16#00EF8# => romdata <= X"72616D70";
    when 16#00EF9# => romdata <= X"20726174";
    when 16#00EFA# => romdata <= X"6520203A";
    when 16#00EFB# => romdata <= X"20000000";
    when 16#00EFC# => romdata <= X"49206D75";
    when 16#00EFD# => romdata <= X"6C742072";
    when 16#00EFE# => romdata <= X"6567203A";
    when 16#00EFF# => romdata <= X"20000000";
    when 16#00F00# => romdata <= X"51206D75";
    when 16#00F01# => romdata <= X"6C742072";
    when 16#00F02# => romdata <= X"6567203A";
    when 16#00F03# => romdata <= X"20000000";
    when 16#00F04# => romdata <= X"554E4B4E";
    when 16#00F05# => romdata <= X"4F574E00";
    when 16#00F06# => romdata <= X"69646C65";
    when 16#00F07# => romdata <= X"00000000";
    when 16#00F08# => romdata <= X"636F6E66";
    when 16#00F09# => romdata <= X"69677572";
    when 16#00F0A# => romdata <= X"65000000";
    when 16#00F0B# => romdata <= X"64657465";
    when 16#00F0C# => romdata <= X"63740000";
    when 16#00F0D# => romdata <= X"61717569";
    when 16#00F0E# => romdata <= X"72650000";
    when 16#00F0F# => romdata <= X"616E616C";
    when 16#00F10# => romdata <= X"797A6500";
    when 16#00F11# => romdata <= X"64657369";
    when 16#00F12# => romdata <= X"72650000";
    when 16#00F13# => romdata <= X"72656164";
    when 16#00F14# => romdata <= X"6F757400";
    when 16#00F15# => romdata <= X"72656164";
    when 16#00F16# => romdata <= X"6C616700";
    when 16#00F17# => romdata <= X"66617374";
    when 16#00F18# => romdata <= X"20747269";
    when 16#00F19# => romdata <= X"67676572";
    when 16#00F1A# => romdata <= X"203A2000";
    when 16#00F1B# => romdata <= X"0A736C6F";
    when 16#00F1C# => romdata <= X"77207472";
    when 16#00F1D# => romdata <= X"69676765";
    when 16#00F1E# => romdata <= X"72203A20";
    when 16#00F1F# => romdata <= X"00000000";
    when 16#00F20# => romdata <= X"0A6F7665";
    when 16#00F21# => romdata <= X"72666C6F";
    when 16#00F22# => romdata <= X"77202020";
    when 16#00F23# => romdata <= X"20203A20";
    when 16#00F24# => romdata <= X"00000000";
    when 16#00F25# => romdata <= X"66617374";
    when 16#00F26# => romdata <= X"20747269";
    when 16#00F27# => romdata <= X"67676572";
    when 16#00F28# => romdata <= X"20636861";
    when 16#00F29# => romdata <= X"696E3A20";
    when 16#00F2A# => romdata <= X"30780000";
    when 16#00F2B# => romdata <= X"0A736C6F";
    when 16#00F2C# => romdata <= X"77207472";
    when 16#00F2D# => romdata <= X"69676765";
    when 16#00F2E# => romdata <= X"72206368";
    when 16#00F2F# => romdata <= X"61696E3A";
    when 16#00F30# => romdata <= X"20307800";
    when 16#00F31# => romdata <= X"746F6B65";
    when 16#00F32# => romdata <= X"6E733A20";
    when 16#00F33# => romdata <= X"00000000";
    when 16#00F34# => romdata <= X"00001AA2";
    when 16#00F35# => romdata <= X"00001AB6";
    when 16#00F36# => romdata <= X"00001A7A";
    when 16#00F37# => romdata <= X"00001ACA";
    when 16#00F38# => romdata <= X"00001ADE";
    when 16#00F39# => romdata <= X"00001AF2";
    when 16#00F3A# => romdata <= X"00001B06";
    when 16#00F3B# => romdata <= X"00001B1A";
    when 16#00F3C# => romdata <= X"00001B2E";
    when 16#00F3D# => romdata <= X"00001A8E";
    when 16#00F3E# => romdata <= X"30622020";
    when 16#00F3F# => romdata <= X"20202020";
    when 16#00F40# => romdata <= X"20202020";
    when 16#00F41# => romdata <= X"20202020";
    when 16#00F42# => romdata <= X"20202020";
    when 16#00F43# => romdata <= X"20202020";
    when 16#00F44# => romdata <= X"20202020";
    when 16#00F45# => romdata <= X"20202020";
    when 16#00F46# => romdata <= X"20200000";
    when 16#00F47# => romdata <= X"20202020";
    when 16#00F48# => romdata <= X"20202020";
    when 16#00F49# => romdata <= X"00000000";
    when 16#00F4A# => romdata <= X"79657300";
    when 16#00F4B# => romdata <= X"6E6F0000";
    when 16#00F4C# => romdata <= X"00202020";
    when 16#00F4D# => romdata <= X"20202020";
    when 16#00F4E# => romdata <= X"20202828";
    when 16#00F4F# => romdata <= X"28282820";
    when 16#00F50# => romdata <= X"20202020";
    when 16#00F51# => romdata <= X"20202020";
    when 16#00F52# => romdata <= X"20202020";
    when 16#00F53# => romdata <= X"20202020";
    when 16#00F54# => romdata <= X"20881010";
    when 16#00F55# => romdata <= X"10101010";
    when 16#00F56# => romdata <= X"10101010";
    when 16#00F57# => romdata <= X"10101010";
    when 16#00F58# => romdata <= X"10040404";
    when 16#00F59# => romdata <= X"04040404";
    when 16#00F5A# => romdata <= X"04040410";
    when 16#00F5B# => romdata <= X"10101010";
    when 16#00F5C# => romdata <= X"10104141";
    when 16#00F5D# => romdata <= X"41414141";
    when 16#00F5E# => romdata <= X"01010101";
    when 16#00F5F# => romdata <= X"01010101";
    when 16#00F60# => romdata <= X"01010101";
    when 16#00F61# => romdata <= X"01010101";
    when 16#00F62# => romdata <= X"01010101";
    when 16#00F63# => romdata <= X"10101010";
    when 16#00F64# => romdata <= X"10104242";
    when 16#00F65# => romdata <= X"42424242";
    when 16#00F66# => romdata <= X"02020202";
    when 16#00F67# => romdata <= X"02020202";
    when 16#00F68# => romdata <= X"02020202";
    when 16#00F69# => romdata <= X"02020202";
    when 16#00F6A# => romdata <= X"02020202";
    when 16#00F6B# => romdata <= X"10101010";
    when 16#00F6C# => romdata <= X"20000000";
    when 16#00F6D# => romdata <= X"00000000";
    when 16#00F6E# => romdata <= X"00000000";
    when 16#00F6F# => romdata <= X"00000000";
    when 16#00F70# => romdata <= X"00000000";
    when 16#00F71# => romdata <= X"00000000";
    when 16#00F72# => romdata <= X"00000000";
    when 16#00F73# => romdata <= X"00000000";
    when 16#00F74# => romdata <= X"00000000";
    when 16#00F75# => romdata <= X"00000000";
    when 16#00F76# => romdata <= X"00000000";
    when 16#00F77# => romdata <= X"00000000";
    when 16#00F78# => romdata <= X"00000000";
    when 16#00F79# => romdata <= X"00000000";
    when 16#00F7A# => romdata <= X"00000000";
    when 16#00F7B# => romdata <= X"00000000";
    when 16#00F7C# => romdata <= X"00000000";
    when 16#00F7D# => romdata <= X"00000000";
    when 16#00F7E# => romdata <= X"00000000";
    when 16#00F7F# => romdata <= X"00000000";
    when 16#00F80# => romdata <= X"00000000";
    when 16#00F81# => romdata <= X"00000000";
    when 16#00F82# => romdata <= X"00000000";
    when 16#00F83# => romdata <= X"00000000";
    when 16#00F84# => romdata <= X"00000000";
    when 16#00F85# => romdata <= X"00000000";
    when 16#00F86# => romdata <= X"00000000";
    when 16#00F87# => romdata <= X"00000000";
    when 16#00F88# => romdata <= X"00000000";
    when 16#00F89# => romdata <= X"00000000";
    when 16#00F8A# => romdata <= X"00000000";
    when 16#00F8B# => romdata <= X"00000000";
    when 16#00F8C# => romdata <= X"00000000";
    when 16#00F8D# => romdata <= X"43000000";
    when 16#00F8E# => romdata <= X"00000000";
    when 16#00F8F# => romdata <= X"00000000";
    when 16#00F90# => romdata <= X"80000B00";
    when 16#00F91# => romdata <= X"10000000";
    when 16#00F92# => romdata <= X"80000D00";
    when 16#00F93# => romdata <= X"00FFFFFF";
    when 16#00F94# => romdata <= X"FF00FFFF";
    when 16#00F95# => romdata <= X"FFFF00FF";
    when 16#00F96# => romdata <= X"FFFFFF00";
    when 16#00F97# => romdata <= X"00000000";
    when 16#00F98# => romdata <= X"00000000";
    when 16#00F99# => romdata <= X"80000A00";
    when 16#00F9A# => romdata <= X"80000400";
    when 16#00F9B# => romdata <= X"80000200";
    when 16#00F9C# => romdata <= X"80000100";
    when 16#00F9D# => romdata <= X"80000004";
    when 16#00F9E# => romdata <= X"80000000";
    when 16#00F9F# => romdata <= X"00003E80";
    when 16#00FA0# => romdata <= X"00000000";
    when 16#00FA1# => romdata <= X"000040E8";
    when 16#00FA2# => romdata <= X"00004144";
    when 16#00FA3# => romdata <= X"000041A0";
    when 16#00FA4# => romdata <= X"00000000";
    when 16#00FA5# => romdata <= X"00000000";
    when 16#00FA6# => romdata <= X"00000000";
    when 16#00FA7# => romdata <= X"00000000";
    when 16#00FA8# => romdata <= X"00000000";
    when 16#00FA9# => romdata <= X"00000000";
    when 16#00FAA# => romdata <= X"00000000";
    when 16#00FAB# => romdata <= X"00000000";
    when 16#00FAC# => romdata <= X"00000000";
    when 16#00FAD# => romdata <= X"00003E34";
    when 16#00FAE# => romdata <= X"00000000";
    when 16#00FAF# => romdata <= X"00000000";
    when 16#00FB0# => romdata <= X"00000000";
    when 16#00FB1# => romdata <= X"00000000";
    when 16#00FB2# => romdata <= X"00000000";
    when 16#00FB3# => romdata <= X"00000000";
    when 16#00FB4# => romdata <= X"00000000";
    when 16#00FB5# => romdata <= X"00000000";
    when 16#00FB6# => romdata <= X"00000000";
    when 16#00FB7# => romdata <= X"00000000";
    when 16#00FB8# => romdata <= X"00000000";
    when 16#00FB9# => romdata <= X"00000000";
    when 16#00FBA# => romdata <= X"00000000";
    when 16#00FBB# => romdata <= X"00000000";
    when 16#00FBC# => romdata <= X"00000000";
    when 16#00FBD# => romdata <= X"00000000";
    when 16#00FBE# => romdata <= X"00000000";
    when 16#00FBF# => romdata <= X"00000000";
    when 16#00FC0# => romdata <= X"00000000";
    when 16#00FC1# => romdata <= X"00000000";
    when 16#00FC2# => romdata <= X"00000000";
    when 16#00FC3# => romdata <= X"00000000";
    when 16#00FC4# => romdata <= X"00000000";
    when 16#00FC5# => romdata <= X"00000000";
    when 16#00FC6# => romdata <= X"00000000";
    when 16#00FC7# => romdata <= X"00000000";
    when 16#00FC8# => romdata <= X"00000000";
    when 16#00FC9# => romdata <= X"00000000";
    when 16#00FCA# => romdata <= X"00000001";
    when 16#00FCB# => romdata <= X"330EABCD";
    when 16#00FCC# => romdata <= X"1234E66D";
    when 16#00FCD# => romdata <= X"DEEC0005";
    when 16#00FCE# => romdata <= X"000B0000";
    when 16#00FCF# => romdata <= X"00000000";
    when 16#00FD0# => romdata <= X"00000000";
    when 16#00FD1# => romdata <= X"00000000";
    when 16#00FD2# => romdata <= X"00000000";
    when 16#00FD3# => romdata <= X"00000000";
    when 16#00FD4# => romdata <= X"00000000";
    when 16#00FD5# => romdata <= X"00000000";
    when 16#00FD6# => romdata <= X"00000000";
    when 16#00FD7# => romdata <= X"00000000";
    when 16#00FD8# => romdata <= X"00000000";
    when 16#00FD9# => romdata <= X"00000000";
    when 16#00FDA# => romdata <= X"00000000";
    when 16#00FDB# => romdata <= X"00000000";
    when 16#00FDC# => romdata <= X"00000000";
    when 16#00FDD# => romdata <= X"00000000";
    when 16#00FDE# => romdata <= X"00000000";
    when 16#00FDF# => romdata <= X"00000000";
    when 16#00FE0# => romdata <= X"00000000";
    when 16#00FE1# => romdata <= X"00000000";
    when 16#00FE2# => romdata <= X"00000000";
    when 16#00FE3# => romdata <= X"00000000";
    when 16#00FE4# => romdata <= X"00000000";
    when 16#00FE5# => romdata <= X"00000000";
    when 16#00FE6# => romdata <= X"00000000";
    when 16#00FE7# => romdata <= X"00000000";
    when 16#00FE8# => romdata <= X"00000000";
    when 16#00FE9# => romdata <= X"00000000";
    when 16#00FEA# => romdata <= X"00000000";
    when 16#00FEB# => romdata <= X"00000000";
    when 16#00FEC# => romdata <= X"00000000";
    when 16#00FED# => romdata <= X"00000000";
    when 16#00FEE# => romdata <= X"00000000";
    when 16#00FEF# => romdata <= X"00000000";
    when 16#00FF0# => romdata <= X"00000000";
    when 16#00FF1# => romdata <= X"00000000";
    when 16#00FF2# => romdata <= X"00000000";
    when 16#00FF3# => romdata <= X"00000000";
    when 16#00FF4# => romdata <= X"00000000";
    when 16#00FF5# => romdata <= X"00000000";
    when 16#00FF6# => romdata <= X"00000000";
    when 16#00FF7# => romdata <= X"00000000";
    when 16#00FF8# => romdata <= X"00000000";
    when 16#00FF9# => romdata <= X"00000000";
    when 16#00FFA# => romdata <= X"00000000";
    when 16#00FFB# => romdata <= X"00000000";
    when 16#00FFC# => romdata <= X"00000000";
    when 16#00FFD# => romdata <= X"00000000";
    when 16#00FFE# => romdata <= X"00000000";
    when 16#00FFF# => romdata <= X"00000000";
    when 16#01000# => romdata <= X"00000000";
    when 16#01001# => romdata <= X"00000000";
    when 16#01002# => romdata <= X"00000000";
    when 16#01003# => romdata <= X"00000000";
    when 16#01004# => romdata <= X"00000000";
    when 16#01005# => romdata <= X"00000000";
    when 16#01006# => romdata <= X"00000000";
    when 16#01007# => romdata <= X"00000000";
    when 16#01008# => romdata <= X"00000000";
    when 16#01009# => romdata <= X"00000000";
    when 16#0100A# => romdata <= X"00000000";
    when 16#0100B# => romdata <= X"00000000";
    when 16#0100C# => romdata <= X"00000000";
    when 16#0100D# => romdata <= X"00000000";
    when 16#0100E# => romdata <= X"00000000";
    when 16#0100F# => romdata <= X"00000000";
    when 16#01010# => romdata <= X"00000000";
    when 16#01011# => romdata <= X"00000000";
    when 16#01012# => romdata <= X"00000000";
    when 16#01013# => romdata <= X"00000000";
    when 16#01014# => romdata <= X"00000000";
    when 16#01015# => romdata <= X"00000000";
    when 16#01016# => romdata <= X"00000000";
    when 16#01017# => romdata <= X"00000000";
    when 16#01018# => romdata <= X"00000000";
    when 16#01019# => romdata <= X"00000000";
    when 16#0101A# => romdata <= X"00000000";
    when 16#0101B# => romdata <= X"00000000";
    when 16#0101C# => romdata <= X"00000000";
    when 16#0101D# => romdata <= X"00000000";
    when 16#0101E# => romdata <= X"00000000";
    when 16#0101F# => romdata <= X"00000000";
    when 16#01020# => romdata <= X"00000000";
    when 16#01021# => romdata <= X"00000000";
    when 16#01022# => romdata <= X"00000000";
    when 16#01023# => romdata <= X"00000000";
    when 16#01024# => romdata <= X"00000000";
    when 16#01025# => romdata <= X"00000000";
    when 16#01026# => romdata <= X"00000000";
    when 16#01027# => romdata <= X"00000000";
    when 16#01028# => romdata <= X"00000000";
    when 16#01029# => romdata <= X"00000000";
    when 16#0102A# => romdata <= X"00000000";
    when 16#0102B# => romdata <= X"00000000";
    when 16#0102C# => romdata <= X"00000000";
    when 16#0102D# => romdata <= X"00000000";
    when 16#0102E# => romdata <= X"00000000";
    when 16#0102F# => romdata <= X"00000000";
    when 16#01030# => romdata <= X"00000000";
    when 16#01031# => romdata <= X"00000000";
    when 16#01032# => romdata <= X"00000000";
    when 16#01033# => romdata <= X"00000000";
    when 16#01034# => romdata <= X"00000000";
    when 16#01035# => romdata <= X"00000000";
    when 16#01036# => romdata <= X"00000000";
    when 16#01037# => romdata <= X"00000000";
    when 16#01038# => romdata <= X"00000000";
    when 16#01039# => romdata <= X"00000000";
    when 16#0103A# => romdata <= X"00000000";
    when 16#0103B# => romdata <= X"00000000";
    when 16#0103C# => romdata <= X"00000000";
    when 16#0103D# => romdata <= X"00000000";
    when 16#0103E# => romdata <= X"00000000";
    when 16#0103F# => romdata <= X"00000000";
    when 16#01040# => romdata <= X"00000000";
    when 16#01041# => romdata <= X"00000000";
    when 16#01042# => romdata <= X"00000000";
    when 16#01043# => romdata <= X"00000000";
    when 16#01044# => romdata <= X"00000000";
    when 16#01045# => romdata <= X"00000000";
    when 16#01046# => romdata <= X"00000000";
    when 16#01047# => romdata <= X"00000000";
    when 16#01048# => romdata <= X"00000000";
    when 16#01049# => romdata <= X"00000000";
    when 16#0104A# => romdata <= X"00000000";
    when 16#0104B# => romdata <= X"00000000";
    when 16#0104C# => romdata <= X"00000000";
    when 16#0104D# => romdata <= X"00000000";
    when 16#0104E# => romdata <= X"00000000";
    when 16#0104F# => romdata <= X"00000000";
    when 16#01050# => romdata <= X"00000000";
    when 16#01051# => romdata <= X"00000000";
    when 16#01052# => romdata <= X"00000000";
    when 16#01053# => romdata <= X"00000000";
    when 16#01054# => romdata <= X"00000000";
    when 16#01055# => romdata <= X"00000000";
    when 16#01056# => romdata <= X"00000000";
    when 16#01057# => romdata <= X"00000000";
    when 16#01058# => romdata <= X"00000000";
    when 16#01059# => romdata <= X"00000000";
    when 16#0105A# => romdata <= X"00000000";
    when 16#0105B# => romdata <= X"00000000";
    when 16#0105C# => romdata <= X"00000000";
    when 16#0105D# => romdata <= X"00000000";
    when 16#0105E# => romdata <= X"00000000";
    when 16#0105F# => romdata <= X"00000000";
    when 16#01060# => romdata <= X"00000000";
    when 16#01061# => romdata <= X"00000000";
    when 16#01062# => romdata <= X"00000000";
    when 16#01063# => romdata <= X"00000000";
    when 16#01064# => romdata <= X"00000000";
    when 16#01065# => romdata <= X"00000000";
    when 16#01066# => romdata <= X"00000000";
    when 16#01067# => romdata <= X"00000000";
    when 16#01068# => romdata <= X"00000000";
    when 16#01069# => romdata <= X"00000000";
    when 16#0106A# => romdata <= X"00000000";
    when 16#0106B# => romdata <= X"00000000";
    when 16#0106C# => romdata <= X"00000000";
    when 16#0106D# => romdata <= X"00000000";
    when 16#0106E# => romdata <= X"00000000";
    when 16#0106F# => romdata <= X"00000000";
    when 16#01070# => romdata <= X"00000000";
    when 16#01071# => romdata <= X"00000000";
    when 16#01072# => romdata <= X"00000000";
    when 16#01073# => romdata <= X"00000000";
    when 16#01074# => romdata <= X"00000000";
    when 16#01075# => romdata <= X"00000000";
    when 16#01076# => romdata <= X"00000000";
    when 16#01077# => romdata <= X"00000000";
    when 16#01078# => romdata <= X"00000000";
    when 16#01079# => romdata <= X"00000000";
    when 16#0107A# => romdata <= X"00000000";
    when 16#0107B# => romdata <= X"00000000";
    when 16#0107C# => romdata <= X"00000000";
    when 16#0107D# => romdata <= X"00000000";
    when 16#0107E# => romdata <= X"00000000";
    when 16#0107F# => romdata <= X"00000000";
    when 16#01080# => romdata <= X"00000000";
    when 16#01081# => romdata <= X"00000000";
    when 16#01082# => romdata <= X"00000000";
    when 16#01083# => romdata <= X"00000000";
    when 16#01084# => romdata <= X"00000000";
    when 16#01085# => romdata <= X"00000000";
    when 16#01086# => romdata <= X"00000000";
    when 16#01087# => romdata <= X"00000000";
    when 16#01088# => romdata <= X"00000000";
    when 16#01089# => romdata <= X"00000000";
    when 16#0108A# => romdata <= X"00000000";
    when 16#0108B# => romdata <= X"FFFFFFFF";
    when 16#0108C# => romdata <= X"00000000";
    when 16#0108D# => romdata <= X"00020000";
    when 16#0108E# => romdata <= X"00000000";
    when 16#0108F# => romdata <= X"00000000";
    when 16#01090# => romdata <= X"00004238";
    when 16#01091# => romdata <= X"00004238";
    when 16#01092# => romdata <= X"00004240";
    when 16#01093# => romdata <= X"00004240";
    when 16#01094# => romdata <= X"00004248";
    when 16#01095# => romdata <= X"00004248";
    when 16#01096# => romdata <= X"00004250";
    when 16#01097# => romdata <= X"00004250";
    when 16#01098# => romdata <= X"00004258";
    when 16#01099# => romdata <= X"00004258";
    when 16#0109A# => romdata <= X"00004260";
    when 16#0109B# => romdata <= X"00004260";
    when 16#0109C# => romdata <= X"00004268";
    when 16#0109D# => romdata <= X"00004268";
    when 16#0109E# => romdata <= X"00004270";
    when 16#0109F# => romdata <= X"00004270";
    when 16#010A0# => romdata <= X"00004278";
    when 16#010A1# => romdata <= X"00004278";
    when 16#010A2# => romdata <= X"00004280";
    when 16#010A3# => romdata <= X"00004280";
    when 16#010A4# => romdata <= X"00004288";
    when 16#010A5# => romdata <= X"00004288";
    when 16#010A6# => romdata <= X"00004290";
    when 16#010A7# => romdata <= X"00004290";
    when 16#010A8# => romdata <= X"00004298";
    when 16#010A9# => romdata <= X"00004298";
    when 16#010AA# => romdata <= X"000042A0";
    when 16#010AB# => romdata <= X"000042A0";
    when 16#010AC# => romdata <= X"000042A8";
    when 16#010AD# => romdata <= X"000042A8";
    when 16#010AE# => romdata <= X"000042B0";
    when 16#010AF# => romdata <= X"000042B0";
    when 16#010B0# => romdata <= X"000042B8";
    when 16#010B1# => romdata <= X"000042B8";
    when 16#010B2# => romdata <= X"000042C0";
    when 16#010B3# => romdata <= X"000042C0";
    when 16#010B4# => romdata <= X"000042C8";
    when 16#010B5# => romdata <= X"000042C8";
    when 16#010B6# => romdata <= X"000042D0";
    when 16#010B7# => romdata <= X"000042D0";
    when 16#010B8# => romdata <= X"000042D8";
    when 16#010B9# => romdata <= X"000042D8";
    when 16#010BA# => romdata <= X"000042E0";
    when 16#010BB# => romdata <= X"000042E0";
    when 16#010BC# => romdata <= X"000042E8";
    when 16#010BD# => romdata <= X"000042E8";
    when 16#010BE# => romdata <= X"000042F0";
    when 16#010BF# => romdata <= X"000042F0";
    when 16#010C0# => romdata <= X"000042F8";
    when 16#010C1# => romdata <= X"000042F8";
    when 16#010C2# => romdata <= X"00004300";
    when 16#010C3# => romdata <= X"00004300";
    when 16#010C4# => romdata <= X"00004308";
    when 16#010C5# => romdata <= X"00004308";
    when 16#010C6# => romdata <= X"00004310";
    when 16#010C7# => romdata <= X"00004310";
    when 16#010C8# => romdata <= X"00004318";
    when 16#010C9# => romdata <= X"00004318";
    when 16#010CA# => romdata <= X"00004320";
    when 16#010CB# => romdata <= X"00004320";
    when 16#010CC# => romdata <= X"00004328";
    when 16#010CD# => romdata <= X"00004328";
    when 16#010CE# => romdata <= X"00004330";
    when 16#010CF# => romdata <= X"00004330";
    when 16#010D0# => romdata <= X"00004338";
    when 16#010D1# => romdata <= X"00004338";
    when 16#010D2# => romdata <= X"00004340";
    when 16#010D3# => romdata <= X"00004340";
    when 16#010D4# => romdata <= X"00004348";
    when 16#010D5# => romdata <= X"00004348";
    when 16#010D6# => romdata <= X"00004350";
    when 16#010D7# => romdata <= X"00004350";
    when 16#010D8# => romdata <= X"00004358";
    when 16#010D9# => romdata <= X"00004358";
    when 16#010DA# => romdata <= X"00004360";
    when 16#010DB# => romdata <= X"00004360";
    when 16#010DC# => romdata <= X"00004368";
    when 16#010DD# => romdata <= X"00004368";
    when 16#010DE# => romdata <= X"00004370";
    when 16#010DF# => romdata <= X"00004370";
    when 16#010E0# => romdata <= X"00004378";
    when 16#010E1# => romdata <= X"00004378";
    when 16#010E2# => romdata <= X"00004380";
    when 16#010E3# => romdata <= X"00004380";
    when 16#010E4# => romdata <= X"00004388";
    when 16#010E5# => romdata <= X"00004388";
    when 16#010E6# => romdata <= X"00004390";
    when 16#010E7# => romdata <= X"00004390";
    when 16#010E8# => romdata <= X"00004398";
    when 16#010E9# => romdata <= X"00004398";
    when 16#010EA# => romdata <= X"000043A0";
    when 16#010EB# => romdata <= X"000043A0";
    when 16#010EC# => romdata <= X"000043A8";
    when 16#010ED# => romdata <= X"000043A8";
    when 16#010EE# => romdata <= X"000043B0";
    when 16#010EF# => romdata <= X"000043B0";
    when 16#010F0# => romdata <= X"000043B8";
    when 16#010F1# => romdata <= X"000043B8";
    when 16#010F2# => romdata <= X"000043C0";
    when 16#010F3# => romdata <= X"000043C0";
    when 16#010F4# => romdata <= X"000043C8";
    when 16#010F5# => romdata <= X"000043C8";
    when 16#010F6# => romdata <= X"000043D0";
    when 16#010F7# => romdata <= X"000043D0";
    when 16#010F8# => romdata <= X"000043D8";
    when 16#010F9# => romdata <= X"000043D8";
    when 16#010FA# => romdata <= X"000043E0";
    when 16#010FB# => romdata <= X"000043E0";
    when 16#010FC# => romdata <= X"000043E8";
    when 16#010FD# => romdata <= X"000043E8";
    when 16#010FE# => romdata <= X"000043F0";
    when 16#010FF# => romdata <= X"000043F0";
    when 16#01100# => romdata <= X"000043F8";
    when 16#01101# => romdata <= X"000043F8";
    when 16#01102# => romdata <= X"00004400";
    when 16#01103# => romdata <= X"00004400";
    when 16#01104# => romdata <= X"00004408";
    when 16#01105# => romdata <= X"00004408";
    when 16#01106# => romdata <= X"00004410";
    when 16#01107# => romdata <= X"00004410";
    when 16#01108# => romdata <= X"00004418";
    when 16#01109# => romdata <= X"00004418";
    when 16#0110A# => romdata <= X"00004420";
    when 16#0110B# => romdata <= X"00004420";
    when 16#0110C# => romdata <= X"00004428";
    when 16#0110D# => romdata <= X"00004428";
    when 16#0110E# => romdata <= X"00004430";
    when 16#0110F# => romdata <= X"00004430";
    when 16#01110# => romdata <= X"00004438";
    when 16#01111# => romdata <= X"00004438";
    when 16#01112# => romdata <= X"00004440";
    when 16#01113# => romdata <= X"00004440";
    when 16#01114# => romdata <= X"00004448";
    when 16#01115# => romdata <= X"00004448";
    when 16#01116# => romdata <= X"00004450";
    when 16#01117# => romdata <= X"00004450";
    when 16#01118# => romdata <= X"00004458";
    when 16#01119# => romdata <= X"00004458";
    when 16#0111A# => romdata <= X"00004460";
    when 16#0111B# => romdata <= X"00004460";
    when 16#0111C# => romdata <= X"00004468";
    when 16#0111D# => romdata <= X"00004468";
    when 16#0111E# => romdata <= X"00004470";
    when 16#0111F# => romdata <= X"00004470";
    when 16#01120# => romdata <= X"00004478";
    when 16#01121# => romdata <= X"00004478";
    when 16#01122# => romdata <= X"00004480";
    when 16#01123# => romdata <= X"00004480";
    when 16#01124# => romdata <= X"00004488";
    when 16#01125# => romdata <= X"00004488";
    when 16#01126# => romdata <= X"00004490";
    when 16#01127# => romdata <= X"00004490";
    when 16#01128# => romdata <= X"00004498";
    when 16#01129# => romdata <= X"00004498";
    when 16#0112A# => romdata <= X"000044A0";
    when 16#0112B# => romdata <= X"000044A0";
    when 16#0112C# => romdata <= X"000044A8";
    when 16#0112D# => romdata <= X"000044A8";
    when 16#0112E# => romdata <= X"000044B0";
    when 16#0112F# => romdata <= X"000044B0";
    when 16#01130# => romdata <= X"000044B8";
    when 16#01131# => romdata <= X"000044B8";
    when 16#01132# => romdata <= X"000044C0";
    when 16#01133# => romdata <= X"000044C0";
    when 16#01134# => romdata <= X"000044C8";
    when 16#01135# => romdata <= X"000044C8";
    when 16#01136# => romdata <= X"000044D0";
    when 16#01137# => romdata <= X"000044D0";
    when 16#01138# => romdata <= X"000044D8";
    when 16#01139# => romdata <= X"000044D8";
    when 16#0113A# => romdata <= X"000044E0";
    when 16#0113B# => romdata <= X"000044E0";
    when 16#0113C# => romdata <= X"000044E8";
    when 16#0113D# => romdata <= X"000044E8";
    when 16#0113E# => romdata <= X"000044F0";
    when 16#0113F# => romdata <= X"000044F0";
    when 16#01140# => romdata <= X"000044F8";
    when 16#01141# => romdata <= X"000044F8";
    when 16#01142# => romdata <= X"00004500";
    when 16#01143# => romdata <= X"00004500";
    when 16#01144# => romdata <= X"00004508";
    when 16#01145# => romdata <= X"00004508";
    when 16#01146# => romdata <= X"00004510";
    when 16#01147# => romdata <= X"00004510";
    when 16#01148# => romdata <= X"00004518";
    when 16#01149# => romdata <= X"00004518";
    when 16#0114A# => romdata <= X"00004520";
    when 16#0114B# => romdata <= X"00004520";
    when 16#0114C# => romdata <= X"00004528";
    when 16#0114D# => romdata <= X"00004528";
    when 16#0114E# => romdata <= X"00004530";
    when 16#0114F# => romdata <= X"00004530";
    when 16#01150# => romdata <= X"00004538";
    when 16#01151# => romdata <= X"00004538";
    when 16#01152# => romdata <= X"00004540";
    when 16#01153# => romdata <= X"00004540";
    when 16#01154# => romdata <= X"00004548";
    when 16#01155# => romdata <= X"00004548";
    when 16#01156# => romdata <= X"00004550";
    when 16#01157# => romdata <= X"00004550";
    when 16#01158# => romdata <= X"00004558";
    when 16#01159# => romdata <= X"00004558";
    when 16#0115A# => romdata <= X"00004560";
    when 16#0115B# => romdata <= X"00004560";
    when 16#0115C# => romdata <= X"00004568";
    when 16#0115D# => romdata <= X"00004568";
    when 16#0115E# => romdata <= X"00004570";
    when 16#0115F# => romdata <= X"00004570";
    when 16#01160# => romdata <= X"00004578";
    when 16#01161# => romdata <= X"00004578";
    when 16#01162# => romdata <= X"00004580";
    when 16#01163# => romdata <= X"00004580";
    when 16#01164# => romdata <= X"00004588";
    when 16#01165# => romdata <= X"00004588";
    when 16#01166# => romdata <= X"00004590";
    when 16#01167# => romdata <= X"00004590";
    when 16#01168# => romdata <= X"00004598";
    when 16#01169# => romdata <= X"00004598";
    when 16#0116A# => romdata <= X"000045A0";
    when 16#0116B# => romdata <= X"000045A0";
    when 16#0116C# => romdata <= X"000045A8";
    when 16#0116D# => romdata <= X"000045A8";
    when 16#0116E# => romdata <= X"000045B0";
    when 16#0116F# => romdata <= X"000045B0";
    when 16#01170# => romdata <= X"000045B8";
    when 16#01171# => romdata <= X"000045B8";
    when 16#01172# => romdata <= X"000045C0";
    when 16#01173# => romdata <= X"000045C0";
    when 16#01174# => romdata <= X"000045C8";
    when 16#01175# => romdata <= X"000045C8";
    when 16#01176# => romdata <= X"000045D0";
    when 16#01177# => romdata <= X"000045D0";
    when 16#01178# => romdata <= X"000045D8";
    when 16#01179# => romdata <= X"000045D8";
    when 16#0117A# => romdata <= X"000045E0";
    when 16#0117B# => romdata <= X"000045E0";
    when 16#0117C# => romdata <= X"000045E8";
    when 16#0117D# => romdata <= X"000045E8";
    when 16#0117E# => romdata <= X"000045F0";
    when 16#0117F# => romdata <= X"000045F0";
    when 16#01180# => romdata <= X"000045F8";
    when 16#01181# => romdata <= X"000045F8";
    when 16#01182# => romdata <= X"00004600";
    when 16#01183# => romdata <= X"00004600";
    when 16#01184# => romdata <= X"00004608";
    when 16#01185# => romdata <= X"00004608";
    when 16#01186# => romdata <= X"00004610";
    when 16#01187# => romdata <= X"00004610";
    when 16#01188# => romdata <= X"00004618";
    when 16#01189# => romdata <= X"00004618";
    when 16#0118A# => romdata <= X"00004620";
    when 16#0118B# => romdata <= X"00004620";
    when 16#0118C# => romdata <= X"00004628";
    when 16#0118D# => romdata <= X"00004628";
    when 16#0118E# => romdata <= X"00004630";
    when 16#0118F# => romdata <= X"00004630";
    when 16#01190# => romdata <= X"00004630";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
