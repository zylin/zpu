-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0bbbd80c",
     3 => x"3a0b0b0b",
     4 => x"aefc0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0bafbe2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bbb",
   162 => x"c4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0ba9",
   171 => x"e72d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bab",
   179 => x"992d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bbbd40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81fb3fa8",
   257 => x"de3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104bb",
   280 => x"d408802e",
   281 => x"a338bbd8",
   282 => x"08822ebd",
   283 => x"38838080",
   284 => x"0b0b0b80",
   285 => x"c3940c82",
   286 => x"a0800b80",
   287 => x"c3980c82",
   288 => x"90800b80",
   289 => x"c39c0c04",
   290 => x"f8808080",
   291 => x"a40b0b0b",
   292 => x"80c3940c",
   293 => x"f8808082",
   294 => x"800b80c3",
   295 => x"980cf880",
   296 => x"8084800b",
   297 => x"80c39c0c",
   298 => x"0480c0a8",
   299 => x"808c0b0b",
   300 => x"0b80c394",
   301 => x"0c80c0a8",
   302 => x"80940b80",
   303 => x"c3980c0b",
   304 => x"0b0bb190",
   305 => x"0b80c39c",
   306 => x"0c04ff3d",
   307 => x"0d80c3a0",
   308 => x"335170a4",
   309 => x"38bbe008",
   310 => x"70085252",
   311 => x"70802e92",
   312 => x"388412bb",
   313 => x"e00c702d",
   314 => x"bbe00870",
   315 => x"08525270",
   316 => x"f038810b",
   317 => x"80c3a034",
   318 => x"833d0d04",
   319 => x"04803d0d",
   320 => x"0b0b80c3",
   321 => x"9008802e",
   322 => x"8e380b0b",
   323 => x"0b0b800b",
   324 => x"802e0981",
   325 => x"06853882",
   326 => x"3d0d040b",
   327 => x"0b80c390",
   328 => x"510b0b0b",
   329 => x"f5da3f82",
   330 => x"3d0d0404",
   331 => x"f83d0d7a",
   332 => x"7c595380",
   333 => x"73565776",
   334 => x"732480dc",
   335 => x"38771754",
   336 => x"8a527451",
   337 => x"9efc3f80",
   338 => x"08b00553",
   339 => x"72743481",
   340 => x"17578a52",
   341 => x"74519ec5",
   342 => x"3f800855",
   343 => x"8008de38",
   344 => x"8008779f",
   345 => x"2a187081",
   346 => x"2c5b5656",
   347 => x"8079259e",
   348 => x"387717ff",
   349 => x"05557518",
   350 => x"70335553",
   351 => x"74337334",
   352 => x"73753481",
   353 => x"16ff1656",
   354 => x"56787624",
   355 => x"e9387618",
   356 => x"56807634",
   357 => x"8a3d0d04",
   358 => x"ad787081",
   359 => x"055a3472",
   360 => x"30781855",
   361 => x"558a5274",
   362 => x"519e973f",
   363 => x"8008b005",
   364 => x"53727434",
   365 => x"8117578a",
   366 => x"5274519d",
   367 => x"e03f8008",
   368 => x"558008fe",
   369 => x"f838ff98",
   370 => x"39f93d0d",
   371 => x"79707133",
   372 => x"7081ff06",
   373 => x"54555555",
   374 => x"70802eb0",
   375 => x"38bbf808",
   376 => x"527281ff",
   377 => x"06811555",
   378 => x"53728a2e",
   379 => x"80f43884",
   380 => x"12087082",
   381 => x"2a810652",
   382 => x"5770802e",
   383 => x"f2387272",
   384 => x"0c733370",
   385 => x"81ff0659",
   386 => x"5377d638",
   387 => x"74753352",
   388 => x"5670802e",
   389 => x"80c83870",
   390 => x"bbf00859",
   391 => x"53811680",
   392 => x"c3a83370",
   393 => x"81ff0670",
   394 => x"10101180",
   395 => x"c3ac3370",
   396 => x"81ff0672",
   397 => x"90291170",
   398 => x"882b7a07",
   399 => x"7f0c5359",
   400 => x"59545458",
   401 => x"56728a2e",
   402 => x"be387380",
   403 => x"cf2eb838",
   404 => x"81155372",
   405 => x"80c3ac34",
   406 => x"75335372",
   407 => x"c038893d",
   408 => x"0d048412",
   409 => x"0870822a",
   410 => x"81065758",
   411 => x"75802ef2",
   412 => x"388d720c",
   413 => x"84120870",
   414 => x"822a8106",
   415 => x"52577080",
   416 => x"2efeec38",
   417 => x"fef83971",
   418 => x"a3269938",
   419 => x"81175271",
   420 => x"80c3a834",
   421 => x"800b80c3",
   422 => x"ac347533",
   423 => x"5372fefd",
   424 => x"38ffbb39",
   425 => x"800b80c3",
   426 => x"a834800b",
   427 => x"80c3ac34",
   428 => x"e939e93d",
   429 => x"0dbbf008",
   430 => x"55800b84",
   431 => x"160cfe80",
   432 => x"0a0b8816",
   433 => x"0c800b80",
   434 => x"c3a83480",
   435 => x"0b80c3ac",
   436 => x"34943d70",
   437 => x"53bbe408",
   438 => x"84110853",
   439 => x"555cfccc",
   440 => x"3fb4980b",
   441 => x"b4983355",
   442 => x"5a73802e",
   443 => x"80cb38bb",
   444 => x"f0087457",
   445 => x"5b811a80",
   446 => x"c3a83370",
   447 => x"81ff0670",
   448 => x"10101180",
   449 => x"c3ac3370",
   450 => x"81ff0672",
   451 => x"90291170",
   452 => x"882b7d07",
   453 => x"620c445c",
   454 => x"5c42575a",
   455 => x"5a758a2e",
   456 => x"87d03876",
   457 => x"80cf2e87",
   458 => x"c9388118",
   459 => x"577680c3",
   460 => x"ac347933",
   461 => x"5675ffbd",
   462 => x"387b7c33",
   463 => x"555a7380",
   464 => x"2e80cb38",
   465 => x"bbf00874",
   466 => x"575b811a",
   467 => x"80c3a833",
   468 => x"7081ff06",
   469 => x"70101011",
   470 => x"80c3ac33",
   471 => x"7081ff06",
   472 => x"72902911",
   473 => x"70882b7d",
   474 => x"07620c46",
   475 => x"5c5c5757",
   476 => x"5a5a758a",
   477 => x"2e879938",
   478 => x"7680cf2e",
   479 => x"87923881",
   480 => x"18597880",
   481 => x"c3ac3479",
   482 => x"335675ff",
   483 => x"bd38b4a8",
   484 => x"0bb4a833",
   485 => x"555a7380",
   486 => x"2e80cb38",
   487 => x"bbf00874",
   488 => x"575b811a",
   489 => x"80c3a833",
   490 => x"7081ff06",
   491 => x"70101011",
   492 => x"80c3ac33",
   493 => x"7081ff06",
   494 => x"72902911",
   495 => x"70882b7d",
   496 => x"07620c44",
   497 => x"5c5c4257",
   498 => x"5a5a758a",
   499 => x"2e868538",
   500 => x"7680cf2e",
   501 => x"85fe3881",
   502 => x"18567580",
   503 => x"c3ac3479",
   504 => x"335675ff",
   505 => x"bd38890a",
   506 => x"5c807093",
   507 => x"3d028c05",
   508 => x"80c10541",
   509 => x"425e5f7c",
   510 => x"bf065a79",
   511 => x"82b638b4",
   512 => x"900bb490",
   513 => x"33555a73",
   514 => x"802e80cb",
   515 => x"38bbf008",
   516 => x"74575b81",
   517 => x"1a80c3a8",
   518 => x"337081ff",
   519 => x"06701010",
   520 => x"1180c3ac",
   521 => x"337081ff",
   522 => x"06729029",
   523 => x"1170882b",
   524 => x"7d07620c",
   525 => x"535c5c57",
   526 => x"575a5a75",
   527 => x"8a2e8386",
   528 => x"387680cf",
   529 => x"2e82ff38",
   530 => x"81185978",
   531 => x"80c3ac34",
   532 => x"79335675",
   533 => x"ffbd387b",
   534 => x"568b53b1",
   535 => x"94527f51",
   536 => x"9d813f88",
   537 => x"57758f06",
   538 => x"54738926",
   539 => x"82bc3876",
   540 => x"1eb01555",
   541 => x"55737534",
   542 => x"75842aff",
   543 => x"187081ff",
   544 => x"06595c56",
   545 => x"76df387f",
   546 => x"6033555a",
   547 => x"73802e80",
   548 => x"cb38bbf0",
   549 => x"0874575b",
   550 => x"811a80c3",
   551 => x"a8337081",
   552 => x"ff067010",
   553 => x"101180c3",
   554 => x"ac337081",
   555 => x"ff067290",
   556 => x"29117088",
   557 => x"2b7d0762",
   558 => x"0c535c5c",
   559 => x"57575a5a",
   560 => x"758a2e85",
   561 => x"94387680",
   562 => x"cf2e858d",
   563 => x"38811855",
   564 => x"7480c3ac",
   565 => x"34793356",
   566 => x"75ffbd38",
   567 => x"b4ac0bb4",
   568 => x"ac33555a",
   569 => x"73802e80",
   570 => x"cb38bbf0",
   571 => x"0874575b",
   572 => x"811a80c3",
   573 => x"a8337081",
   574 => x"ff067010",
   575 => x"101180c3",
   576 => x"ac337081",
   577 => x"ff067290",
   578 => x"29117088",
   579 => x"2b7d0762",
   580 => x"0c535c5c",
   581 => x"57575a5a",
   582 => x"758a2e84",
   583 => x"da387680",
   584 => x"cf2e84d3",
   585 => x"38811857",
   586 => x"7680c3ac",
   587 => x"34793356",
   588 => x"75ffbd38",
   589 => x"7b7c082e",
   590 => x"81aa38b4",
   591 => x"b00bb4b0",
   592 => x"33555a73",
   593 => x"802e80cb",
   594 => x"38bbf008",
   595 => x"74575b81",
   596 => x"1a80c3a8",
   597 => x"337081ff",
   598 => x"06701010",
   599 => x"1180c3ac",
   600 => x"337081ff",
   601 => x"06729029",
   602 => x"1170882b",
   603 => x"7d07620c",
   604 => x"535c5c57",
   605 => x"575a5a75",
   606 => x"8a2e829e",
   607 => x"387680cf",
   608 => x"2e829738",
   609 => x"81185675",
   610 => x"80c3ac34",
   611 => x"79335675",
   612 => x"ffbd3881",
   613 => x"1f5f821c",
   614 => x"811e5e5c",
   615 => x"8fff7d27",
   616 => x"fcd5387e",
   617 => x"800c993d",
   618 => x"0d04761e",
   619 => x"b7155555",
   620 => x"73753475",
   621 => x"842aff18",
   622 => x"7081ff06",
   623 => x"595c5676",
   624 => x"fda338fd",
   625 => x"c23974a3",
   626 => x"2681fa38",
   627 => x"81195776",
   628 => x"80c3a834",
   629 => x"800b80c3",
   630 => x"ac347933",
   631 => x"5675fcb3",
   632 => x"38fcf439",
   633 => x"841c5a79",
   634 => x"7a082e09",
   635 => x"8106fecb",
   636 => x"38b4b40b",
   637 => x"b4b43355",
   638 => x"5a73802e",
   639 => x"ff9838bb",
   640 => x"f0087481",
   641 => x"1c80c3a8",
   642 => x"337081ff",
   643 => x"06701010",
   644 => x"1180c3ac",
   645 => x"337081ff",
   646 => x"06729029",
   647 => x"1170882b",
   648 => x"7807790c",
   649 => x"535e5e59",
   650 => x"595c5c57",
   651 => x"5b758a2e",
   652 => x"80ca3876",
   653 => x"80cf2e80",
   654 => x"c3388118",
   655 => x"597880c3",
   656 => x"ac347933",
   657 => x"5675802e",
   658 => x"fecc3881",
   659 => x"1a80c3a8",
   660 => x"337081ff",
   661 => x"06701010",
   662 => x"1180c3ac",
   663 => x"337081ff",
   664 => x"06729029",
   665 => x"1170882b",
   666 => x"7d07620c",
   667 => x"535c5c57",
   668 => x"575a5a75",
   669 => x"8a2e0981",
   670 => x"06ffb838",
   671 => x"74a32682",
   672 => x"b0388119",
   673 => x"587780c3",
   674 => x"a834800b",
   675 => x"80c3ac34",
   676 => x"79335675",
   677 => x"ffb538fd",
   678 => x"fd3974a3",
   679 => x"26993881",
   680 => x"19557480",
   681 => x"c3a83480",
   682 => x"0b80c3ac",
   683 => x"34793356",
   684 => x"75fd9c38",
   685 => x"fddd3980",
   686 => x"0b80c3a8",
   687 => x"34800b80",
   688 => x"c3ac34e9",
   689 => x"39800b80",
   690 => x"c3a83480",
   691 => x"0b80c3ac",
   692 => x"34fe8739",
   693 => x"74a32680",
   694 => x"f1388119",
   695 => x"557480c3",
   696 => x"a834800b",
   697 => x"80c3ac34",
   698 => x"79335675",
   699 => x"f9b438f9",
   700 => x"f53974a3",
   701 => x"2680c438",
   702 => x"81195675",
   703 => x"80c3a834",
   704 => x"800b80c3",
   705 => x"ac347933",
   706 => x"5675f7e9",
   707 => x"38f8aa39",
   708 => x"74a32699",
   709 => x"38811958",
   710 => x"7780c3a8",
   711 => x"34800b80",
   712 => x"c3ac3479",
   713 => x"335675f8",
   714 => x"a138f8e2",
   715 => x"39800b80",
   716 => x"c3a83480",
   717 => x"0b80c3ac",
   718 => x"34e93980",
   719 => x"0b80c3a8",
   720 => x"34800b80",
   721 => x"c3ac34ff",
   722 => x"bd39800b",
   723 => x"80c3a834",
   724 => x"800b80c3",
   725 => x"ac34ff90",
   726 => x"3974a326",
   727 => x"80c43881",
   728 => x"19587780",
   729 => x"c3a83480",
   730 => x"0b80c3ac",
   731 => x"34793356",
   732 => x"75faa538",
   733 => x"fae63974",
   734 => x"a3269938",
   735 => x"81195675",
   736 => x"80c3a834",
   737 => x"800b80c3",
   738 => x"ac347933",
   739 => x"5675fae0",
   740 => x"38fba139",
   741 => x"800b80c3",
   742 => x"a834800b",
   743 => x"80c3ac34",
   744 => x"e939800b",
   745 => x"80c3a834",
   746 => x"800b80c3",
   747 => x"ac34ffbd",
   748 => x"39800b80",
   749 => x"c3a83480",
   750 => x"0b80c3ac",
   751 => x"34fdd139",
   752 => x"ed3d0db9",
   753 => x"c451f481",
   754 => x"3fb9e051",
   755 => x"f3fb3f90",
   756 => x"3d7053bb",
   757 => x"e4088411",
   758 => x"0853555c",
   759 => x"f2ce3f7b",
   760 => x"51f3e63f",
   761 => x"b4ac51f3",
   762 => x"e03ff5c6",
   763 => x"3f80088e",
   764 => x"3d5a568b",
   765 => x"53b19452",
   766 => x"785195e7",
   767 => x"3f880284",
   768 => x"05b10559",
   769 => x"57758f06",
   770 => x"54738926",
   771 => x"84c53876",
   772 => x"18b01555",
   773 => x"55737534",
   774 => x"75842aff",
   775 => x"187081ff",
   776 => x"06595656",
   777 => x"76df3878",
   778 => x"79335557",
   779 => x"73802ea8",
   780 => x"3873bbf8",
   781 => x"08565681",
   782 => x"1757758a",
   783 => x"2e84b038",
   784 => x"84150870",
   785 => x"822a8106",
   786 => x"555a7380",
   787 => x"2ef23875",
   788 => x"750c7633",
   789 => x"5675e038",
   790 => x"78793355",
   791 => x"5a73802e",
   792 => x"80cb3873",
   793 => x"bbf0085c",
   794 => x"56811a80",
   795 => x"c3a83370",
   796 => x"81ff0670",
   797 => x"10101180",
   798 => x"c3ac3370",
   799 => x"81ff0672",
   800 => x"90291170",
   801 => x"882b7d07",
   802 => x"620c535c",
   803 => x"5c57575a",
   804 => x"5a758a2e",
   805 => x"83fe3876",
   806 => x"80cf2e83",
   807 => x"f7388118",
   808 => x"577680c3",
   809 => x"ac347933",
   810 => x"5675ffbd",
   811 => x"38bbe408",
   812 => x"8411085a",
   813 => x"55fe8179",
   814 => x"25993880",
   815 => x"0b84160c",
   816 => x"815186ff",
   817 => x"3fbbe408",
   818 => x"8411085a",
   819 => x"5578fe81",
   820 => x"24e93883",
   821 => x"ffff58fe",
   822 => x"810b8416",
   823 => x"085c597a",
   824 => x"81fe2480",
   825 => x"c638800b",
   826 => x"88160cf3",
   827 => x"c53f8008",
   828 => x"83ffff06",
   829 => x"55747827",
   830 => x"8b3874bb",
   831 => x"e4088411",
   832 => x"085b5b58",
   833 => x"b49051f1",
   834 => x"c03f7b52",
   835 => x"7451f09c",
   836 => x"3f7b51f1",
   837 => x"b43f7480",
   838 => x"2e83a438",
   839 => x"bbe40884",
   840 => x"11085c55",
   841 => x"81fe7b25",
   842 => x"ffbc3884",
   843 => x"15085a84",
   844 => x"15085473",
   845 => x"81fe2480",
   846 => x"c438800b",
   847 => x"88160cf2",
   848 => x"f13f8008",
   849 => x"83ffff06",
   850 => x"55747827",
   851 => x"8b3874bb",
   852 => x"e4088411",
   853 => x"085b5758",
   854 => x"b49051f0",
   855 => x"ec3f7b52",
   856 => x"7451efc8",
   857 => x"3f7b51f0",
   858 => x"e03f7482",
   859 => x"dd38bbe4",
   860 => x"08841108",
   861 => x"555581fe",
   862 => x"7425ffbe",
   863 => x"38841508",
   864 => x"5780777a",
   865 => x"31575473",
   866 => x"7625b538",
   867 => x"800b8416",
   868 => x"0c815185",
   869 => x"ae3f8114",
   870 => x"7083ffff",
   871 => x"06555573",
   872 => x"76259d38",
   873 => x"bbe40855",
   874 => x"800b8416",
   875 => x"0c815185",
   876 => x"923f8114",
   877 => x"7083ffff",
   878 => x"06555575",
   879 => x"7424e538",
   880 => x"b9ec51f0",
   881 => x"843f7b52",
   882 => x"7951eee0",
   883 => x"3f7b51ef",
   884 => x"f83fb9fc",
   885 => x"51eff23f",
   886 => x"7b527651",
   887 => x"eece3f7b",
   888 => x"51efe63f",
   889 => x"ba8c51ef",
   890 => x"e03f7b52",
   891 => x"767a3170",
   892 => x"525beeb8",
   893 => x"3f7b51ef",
   894 => x"d03fba9c",
   895 => x"51efca3f",
   896 => x"7b527a9f",
   897 => x"2a1b7081",
   898 => x"2c5257ee",
   899 => x"9f3f7b51",
   900 => x"efb73fba",
   901 => x"ac51efb1",
   902 => x"3f7b5277",
   903 => x"51ee8d3f",
   904 => x"7b51efa5",
   905 => x"3fbabc51",
   906 => x"ef9f3f7b",
   907 => x"527851ed",
   908 => x"fb3f7b51",
   909 => x"ef933fba",
   910 => x"cc51ef8d",
   911 => x"3f7b52bb",
   912 => x"e4088411",
   913 => x"085258ed",
   914 => x"e33f7b51",
   915 => x"eefb3f95",
   916 => x"3d0d0476",
   917 => x"18b71555",
   918 => x"55737534",
   919 => x"75842aff",
   920 => x"187081ff",
   921 => x"06595656",
   922 => x"76fb9a38",
   923 => x"fbb93984",
   924 => x"15087082",
   925 => x"2a810659",
   926 => x"5b77802e",
   927 => x"f2388d75",
   928 => x"0c841508",
   929 => x"70822a81",
   930 => x"06555a73",
   931 => x"802efbb0",
   932 => x"38fbbc39",
   933 => x"74a32699",
   934 => x"38811956",
   935 => x"7580c3a8",
   936 => x"34800b80",
   937 => x"c3ac3479",
   938 => x"335675fb",
   939 => x"bc38fbfd",
   940 => x"39800b80",
   941 => x"c3a83480",
   942 => x"0b80c3ac",
   943 => x"34e939bb",
   944 => x"e4088411",
   945 => x"085b55fc",
   946 => x"e639bbe4",
   947 => x"08841108",
   948 => x"58558077",
   949 => x"7a315754",
   950 => x"757424fd",
   951 => x"af38fde0",
   952 => x"39f83d0d",
   953 => x"bbec0870",
   954 => x"08810a06",
   955 => x"80c3a40c",
   956 => x"53890a52",
   957 => x"83ffff53",
   958 => x"71720c84",
   959 => x"12ff1454",
   960 => x"52728025",
   961 => x"f33884a9",
   962 => x"3f84b63f",
   963 => x"bbf00852",
   964 => x"800b8413",
   965 => x"0cfe800a",
   966 => x"0b88130c",
   967 => x"800b80c3",
   968 => x"a834800b",
   969 => x"80c3ac34",
   970 => x"bbf80854",
   971 => x"b60b8c15",
   972 => x"0c830b88",
   973 => x"150cbbec",
   974 => x"08881108",
   975 => x"81ff0788",
   976 => x"120c54bb",
   977 => x"e80853ff",
   978 => x"0b84140c",
   979 => x"fc94800b",
   980 => x"88140c82",
   981 => x"d0affdfb",
   982 => x"0b8c140c",
   983 => x"80c0730c",
   984 => x"72087086",
   985 => x"2a810651",
   986 => x"5473f538",
   987 => x"90130870",
   988 => x"832a8106",
   989 => x"515271f4",
   990 => x"3881fc80",
   991 => x"810b9014",
   992 => x"0c901308",
   993 => x"70832a81",
   994 => x"06515271",
   995 => x"f43880fd",
   996 => x"c0810b90",
   997 => x"140cbadc",
   998 => x"5188e53f",
   999 => x"b3e051ec",
  1000 => x"a83f71bb",
  1001 => x"f0085553",
  1002 => x"72882b74",
  1003 => x"0c811353",
  1004 => x"97907326",
  1005 => x"f338800b",
  1006 => x"80c3a834",
  1007 => x"800b80c3",
  1008 => x"ac34bae8",
  1009 => x"51ec823f",
  1010 => x"80c3a408",
  1011 => x"802e80ed",
  1012 => x"38baf051",
  1013 => x"ebf33fbb",
  1014 => x"8051ebed",
  1015 => x"3ff7e13f",
  1016 => x"8a518181",
  1017 => x"3f800bbb",
  1018 => x"f0085553",
  1019 => x"72882b74",
  1020 => x"0c811353",
  1021 => x"97907326",
  1022 => x"f338800b",
  1023 => x"80c3a834",
  1024 => x"800b80c3",
  1025 => x"ac34edaa",
  1026 => x"3fbbec08",
  1027 => x"70087087",
  1028 => x"2a810651",
  1029 => x"55537380",
  1030 => x"2e8a38bb",
  1031 => x"e4085280",
  1032 => x"0b84130c",
  1033 => x"72087084",
  1034 => x"2a810654",
  1035 => x"5272802e",
  1036 => x"d538bbe4",
  1037 => x"0853800b",
  1038 => x"88140cca",
  1039 => x"39bba451",
  1040 => x"ff9239fd",
  1041 => x"3d0dbbf4",
  1042 => x"0876b0ea",
  1043 => x"2994120c",
  1044 => x"54850b98",
  1045 => x"150c9814",
  1046 => x"08708106",
  1047 => x"515372f6",
  1048 => x"38853d0d",
  1049 => x"04fb3d0d",
  1050 => x"77568055",
  1051 => x"74762781",
  1052 => x"9838bbf4",
  1053 => x"0854bfa9",
  1054 => x"bc0b9415",
  1055 => x"0c850b98",
  1056 => x"150c9814",
  1057 => x"08708106",
  1058 => x"515372f6",
  1059 => x"38bfa9bc",
  1060 => x"0b94150c",
  1061 => x"850b9815",
  1062 => x"0c981408",
  1063 => x"70810651",
  1064 => x"5372f638",
  1065 => x"bfa9bc0b",
  1066 => x"94150c85",
  1067 => x"0b98150c",
  1068 => x"98140870",
  1069 => x"81065153",
  1070 => x"72f638bf",
  1071 => x"a9bc0b94",
  1072 => x"150c850b",
  1073 => x"98150c98",
  1074 => x"14087081",
  1075 => x"06515372",
  1076 => x"f638bfa9",
  1077 => x"bc0b9415",
  1078 => x"0c850b98",
  1079 => x"150c9814",
  1080 => x"08708106",
  1081 => x"515372f6",
  1082 => x"38bfa9bc",
  1083 => x"0b94150c",
  1084 => x"850b9815",
  1085 => x"0c981408",
  1086 => x"70810651",
  1087 => x"5372f638",
  1088 => x"81155575",
  1089 => x"7526feee",
  1090 => x"38873d0d",
  1091 => x"04ff3d0d",
  1092 => x"bbf40874",
  1093 => x"10107510",
  1094 => x"0594120c",
  1095 => x"52850b98",
  1096 => x"130c9812",
  1097 => x"08708106",
  1098 => x"515170f6",
  1099 => x"38833d0d",
  1100 => x"04803d0d",
  1101 => x"bbf40851",
  1102 => x"870b8412",
  1103 => x"0c823d0d",
  1104 => x"04fd3d0d",
  1105 => x"bbec0888",
  1106 => x"110883de",
  1107 => x"80078812",
  1108 => x"0c841108",
  1109 => x"fca1ff06",
  1110 => x"84120c53",
  1111 => x"8f51fde3",
  1112 => x"3fbbec08",
  1113 => x"841108e1",
  1114 => x"ff068412",
  1115 => x"0c841108",
  1116 => x"86800784",
  1117 => x"120c8411",
  1118 => x"0880c080",
  1119 => x"0784120c",
  1120 => x"538151ff",
  1121 => x"883fbbec",
  1122 => x"08841108",
  1123 => x"ffbfff06",
  1124 => x"84120c53",
  1125 => x"8551fdab",
  1126 => x"3fbbec08",
  1127 => x"84110880",
  1128 => x"c0800784",
  1129 => x"120c5381",
  1130 => x"51fee23f",
  1131 => x"bbec0884",
  1132 => x"1108ffbf",
  1133 => x"ff068412",
  1134 => x"0c538151",
  1135 => x"fd853fbb",
  1136 => x"ec088411",
  1137 => x"0880c080",
  1138 => x"0784120c",
  1139 => x"538151fe",
  1140 => x"bc3fbbec",
  1141 => x"08841108",
  1142 => x"ffbfff06",
  1143 => x"84120c53",
  1144 => x"8151fcdf",
  1145 => x"3fbbec08",
  1146 => x"841108e1",
  1147 => x"ff068412",
  1148 => x"0c538480",
  1149 => x"0b841408",
  1150 => x"70720784",
  1151 => x"160c5384",
  1152 => x"14087080",
  1153 => x"c0800784",
  1154 => x"160c5354",
  1155 => x"8151fdfd",
  1156 => x"3fbbec08",
  1157 => x"84110870",
  1158 => x"ffbfff06",
  1159 => x"84130c53",
  1160 => x"538551fc",
  1161 => x"9e3fbbec",
  1162 => x"08841108",
  1163 => x"70feffff",
  1164 => x"0684130c",
  1165 => x"53841108",
  1166 => x"70e1ff06",
  1167 => x"84130c53",
  1168 => x"84110870",
  1169 => x"76078413",
  1170 => x"0c538411",
  1171 => x"0880c080",
  1172 => x"0784120c",
  1173 => x"538151fd",
  1174 => x"b43fbbec",
  1175 => x"08841108",
  1176 => x"ffbfff06",
  1177 => x"84120c84",
  1178 => x"1108e1ff",
  1179 => x"0684120c",
  1180 => x"84110890",
  1181 => x"80078412",
  1182 => x"0c841108",
  1183 => x"80c08007",
  1184 => x"84120c54",
  1185 => x"8151fd85",
  1186 => x"3fbbec08",
  1187 => x"841108ff",
  1188 => x"bfff0684",
  1189 => x"120c54aa",
  1190 => x"51fcf23f",
  1191 => x"bbec0884",
  1192 => x"1108feff",
  1193 => x"ff068412",
  1194 => x"0c841108",
  1195 => x"e1ff0684",
  1196 => x"120c8411",
  1197 => x"0884120c",
  1198 => x"84110880",
  1199 => x"c0800784",
  1200 => x"120c5481",
  1201 => x"51fcc63f",
  1202 => x"bbec0884",
  1203 => x"1108ffbf",
  1204 => x"ff068412",
  1205 => x"0c841108",
  1206 => x"e1ff0684",
  1207 => x"120c8411",
  1208 => x"08988007",
  1209 => x"84120c84",
  1210 => x"110880c0",
  1211 => x"80078412",
  1212 => x"0c548151",
  1213 => x"fc973fbb",
  1214 => x"ec088411",
  1215 => x"08ffbfff",
  1216 => x"0684120c",
  1217 => x"54aa51fc",
  1218 => x"843fbbec",
  1219 => x"08841108",
  1220 => x"feffff06",
  1221 => x"84120c84",
  1222 => x"1108e1ff",
  1223 => x"0684120c",
  1224 => x"84110884",
  1225 => x"120c8411",
  1226 => x"0880c080",
  1227 => x"0784120c",
  1228 => x"548151fb",
  1229 => x"d83fbbec",
  1230 => x"08841108",
  1231 => x"ffbfff06",
  1232 => x"84120c84",
  1233 => x"1108e1ff",
  1234 => x"0684120c",
  1235 => x"8411088c",
  1236 => x"80078412",
  1237 => x"0c841108",
  1238 => x"80c08007",
  1239 => x"84120c54",
  1240 => x"8151fba9",
  1241 => x"3fbbec08",
  1242 => x"841108ff",
  1243 => x"bfff0684",
  1244 => x"120c54aa",
  1245 => x"51fb963f",
  1246 => x"810bbbec",
  1247 => x"08841108",
  1248 => x"70feffff",
  1249 => x"0684130c",
  1250 => x"54841108",
  1251 => x"70e1ff06",
  1252 => x"84130c54",
  1253 => x"84110884",
  1254 => x"120c8411",
  1255 => x"087080c0",
  1256 => x"80078413",
  1257 => x"0c545470",
  1258 => x"5254fae1",
  1259 => x"3fbbec08",
  1260 => x"84110870",
  1261 => x"ffbfff06",
  1262 => x"84130c53",
  1263 => x"84110870",
  1264 => x"e1ff0684",
  1265 => x"130c5384",
  1266 => x"11087082",
  1267 => x"80078413",
  1268 => x"0c538411",
  1269 => x"087080c0",
  1270 => x"80078413",
  1271 => x"0c535373",
  1272 => x"51faaa3f",
  1273 => x"bbec0884",
  1274 => x"1108ffbf",
  1275 => x"ff068412",
  1276 => x"0c53aa51",
  1277 => x"fa973f82",
  1278 => x"51f8c83f",
  1279 => x"853d0d04",
  1280 => x"fb3d0d77",
  1281 => x"70335356",
  1282 => x"71802e81",
  1283 => x"8c387155",
  1284 => x"8116bbec",
  1285 => x"08841108",
  1286 => x"81808007",
  1287 => x"84120c84",
  1288 => x"1108e1ff",
  1289 => x"0684120c",
  1290 => x"76842b9e",
  1291 => x"80068412",
  1292 => x"08707207",
  1293 => x"84140c55",
  1294 => x"84120880",
  1295 => x"c0800784",
  1296 => x"130c5654",
  1297 => x"568151f9",
  1298 => x"c43fbbec",
  1299 => x"08841108",
  1300 => x"ffbfff06",
  1301 => x"84120c84",
  1302 => x"1108e1ff",
  1303 => x"0684120c",
  1304 => x"75882b9e",
  1305 => x"80068412",
  1306 => x"08710784",
  1307 => x"130c8412",
  1308 => x"0880c080",
  1309 => x"0784130c",
  1310 => x"55538151",
  1311 => x"f98f3fbb",
  1312 => x"ec088411",
  1313 => x"08ffbfff",
  1314 => x"0684120c",
  1315 => x"53ae51f8",
  1316 => x"fc3f7533",
  1317 => x"5574fef8",
  1318 => x"38873d0d",
  1319 => x"048c0802",
  1320 => x"8c0cfd3d",
  1321 => x"0d80538c",
  1322 => x"088c0508",
  1323 => x"528c0888",
  1324 => x"05085182",
  1325 => x"de3f8008",
  1326 => x"70800c54",
  1327 => x"853d0d8c",
  1328 => x"0c048c08",
  1329 => x"028c0cfd",
  1330 => x"3d0d8153",
  1331 => x"8c088c05",
  1332 => x"08528c08",
  1333 => x"88050851",
  1334 => x"82b93f80",
  1335 => x"0870800c",
  1336 => x"54853d0d",
  1337 => x"8c0c048c",
  1338 => x"08028c0c",
  1339 => x"f93d0d80",
  1340 => x"0b8c08fc",
  1341 => x"050c8c08",
  1342 => x"88050880",
  1343 => x"25ab388c",
  1344 => x"08880508",
  1345 => x"308c0888",
  1346 => x"050c800b",
  1347 => x"8c08f405",
  1348 => x"0c8c08fc",
  1349 => x"05088838",
  1350 => x"810b8c08",
  1351 => x"f4050c8c",
  1352 => x"08f40508",
  1353 => x"8c08fc05",
  1354 => x"0c8c088c",
  1355 => x"05088025",
  1356 => x"ab388c08",
  1357 => x"8c050830",
  1358 => x"8c088c05",
  1359 => x"0c800b8c",
  1360 => x"08f0050c",
  1361 => x"8c08fc05",
  1362 => x"08883881",
  1363 => x"0b8c08f0",
  1364 => x"050c8c08",
  1365 => x"f005088c",
  1366 => x"08fc050c",
  1367 => x"80538c08",
  1368 => x"8c050852",
  1369 => x"8c088805",
  1370 => x"085181a7",
  1371 => x"3f800870",
  1372 => x"8c08f805",
  1373 => x"0c548c08",
  1374 => x"fc050880",
  1375 => x"2e8c388c",
  1376 => x"08f80508",
  1377 => x"308c08f8",
  1378 => x"050c8c08",
  1379 => x"f8050870",
  1380 => x"800c5489",
  1381 => x"3d0d8c0c",
  1382 => x"048c0802",
  1383 => x"8c0cfb3d",
  1384 => x"0d800b8c",
  1385 => x"08fc050c",
  1386 => x"8c088805",
  1387 => x"08802593",
  1388 => x"388c0888",
  1389 => x"0508308c",
  1390 => x"0888050c",
  1391 => x"810b8c08",
  1392 => x"fc050c8c",
  1393 => x"088c0508",
  1394 => x"80258c38",
  1395 => x"8c088c05",
  1396 => x"08308c08",
  1397 => x"8c050c81",
  1398 => x"538c088c",
  1399 => x"0508528c",
  1400 => x"08880508",
  1401 => x"51ad3f80",
  1402 => x"08708c08",
  1403 => x"f8050c54",
  1404 => x"8c08fc05",
  1405 => x"08802e8c",
  1406 => x"388c08f8",
  1407 => x"0508308c",
  1408 => x"08f8050c",
  1409 => x"8c08f805",
  1410 => x"0870800c",
  1411 => x"54873d0d",
  1412 => x"8c0c048c",
  1413 => x"08028c0c",
  1414 => x"fd3d0d81",
  1415 => x"0b8c08fc",
  1416 => x"050c800b",
  1417 => x"8c08f805",
  1418 => x"0c8c088c",
  1419 => x"05088c08",
  1420 => x"88050827",
  1421 => x"ac388c08",
  1422 => x"fc050880",
  1423 => x"2ea33880",
  1424 => x"0b8c088c",
  1425 => x"05082499",
  1426 => x"388c088c",
  1427 => x"0508108c",
  1428 => x"088c050c",
  1429 => x"8c08fc05",
  1430 => x"08108c08",
  1431 => x"fc050cc9",
  1432 => x"398c08fc",
  1433 => x"0508802e",
  1434 => x"80c9388c",
  1435 => x"088c0508",
  1436 => x"8c088805",
  1437 => x"0826a138",
  1438 => x"8c088805",
  1439 => x"088c088c",
  1440 => x"0508318c",
  1441 => x"0888050c",
  1442 => x"8c08f805",
  1443 => x"088c08fc",
  1444 => x"0508078c",
  1445 => x"08f8050c",
  1446 => x"8c08fc05",
  1447 => x"08812a8c",
  1448 => x"08fc050c",
  1449 => x"8c088c05",
  1450 => x"08812a8c",
  1451 => x"088c050c",
  1452 => x"ffaf398c",
  1453 => x"08900508",
  1454 => x"802e8f38",
  1455 => x"8c088805",
  1456 => x"08708c08",
  1457 => x"f4050c51",
  1458 => x"8d398c08",
  1459 => x"f8050870",
  1460 => x"8c08f405",
  1461 => x"0c518c08",
  1462 => x"f4050880",
  1463 => x"0c853d0d",
  1464 => x"8c0c04fc",
  1465 => x"3d0d7670",
  1466 => x"797b5555",
  1467 => x"55558f72",
  1468 => x"278c3872",
  1469 => x"75078306",
  1470 => x"5170802e",
  1471 => x"a738ff12",
  1472 => x"5271ff2e",
  1473 => x"98387270",
  1474 => x"81055433",
  1475 => x"74708105",
  1476 => x"5634ff12",
  1477 => x"5271ff2e",
  1478 => x"098106ea",
  1479 => x"3874800c",
  1480 => x"863d0d04",
  1481 => x"74517270",
  1482 => x"84055408",
  1483 => x"71708405",
  1484 => x"530c7270",
  1485 => x"84055408",
  1486 => x"71708405",
  1487 => x"530c7270",
  1488 => x"84055408",
  1489 => x"71708405",
  1490 => x"530c7270",
  1491 => x"84055408",
  1492 => x"71708405",
  1493 => x"530cf012",
  1494 => x"52718f26",
  1495 => x"c9388372",
  1496 => x"27953872",
  1497 => x"70840554",
  1498 => x"08717084",
  1499 => x"05530cfc",
  1500 => x"12527183",
  1501 => x"26ed3870",
  1502 => x"54ff8339",
  1503 => x"fd3d0d80",
  1504 => x"0bbbd808",
  1505 => x"54547281",
  1506 => x"2e993873",
  1507 => x"80c3b00c",
  1508 => x"d9cd3fd8",
  1509 => x"eb3fbbfc",
  1510 => x"528151ee",
  1511 => x"c43f8008",
  1512 => x"519f3f72",
  1513 => x"80c3b00c",
  1514 => x"d9b53fd8",
  1515 => x"d33fbbfc",
  1516 => x"528151ee",
  1517 => x"ac3f8008",
  1518 => x"51873f00",
  1519 => x"ff3900ff",
  1520 => x"39f73d0d",
  1521 => x"7bbc8008",
  1522 => x"82c81108",
  1523 => x"5a545a77",
  1524 => x"802e80d9",
  1525 => x"38818818",
  1526 => x"841908ff",
  1527 => x"0581712b",
  1528 => x"59555980",
  1529 => x"742480e9",
  1530 => x"38807424",
  1531 => x"b5387382",
  1532 => x"2b781188",
  1533 => x"05565681",
  1534 => x"80190877",
  1535 => x"06537280",
  1536 => x"2eb53878",
  1537 => x"16700853",
  1538 => x"53795174",
  1539 => x"0853722d",
  1540 => x"ff14fc17",
  1541 => x"fc177981",
  1542 => x"2c5a5757",
  1543 => x"54738025",
  1544 => x"d6387708",
  1545 => x"5877ffad",
  1546 => x"38bc8008",
  1547 => x"53bc1308",
  1548 => x"a5387951",
  1549 => x"ff853f74",
  1550 => x"0853722d",
  1551 => x"ff14fc17",
  1552 => x"fc177981",
  1553 => x"2c5a5757",
  1554 => x"54738025",
  1555 => x"ffa938d2",
  1556 => x"398057ff",
  1557 => x"94397251",
  1558 => x"bc130853",
  1559 => x"722d7951",
  1560 => x"fed93fff",
  1561 => x"3d0d80c3",
  1562 => x"840bfc05",
  1563 => x"70085252",
  1564 => x"70ff2e91",
  1565 => x"38702dfc",
  1566 => x"12700852",
  1567 => x"5270ff2e",
  1568 => x"098106f1",
  1569 => x"38833d0d",
  1570 => x"0404d8be",
  1571 => x"3f040000",
  1572 => x"00000040",
  1573 => x"30782020",
  1574 => x"20202020",
  1575 => x"20200000",
  1576 => x"0a677265",
  1577 => x"74682072",
  1578 => x"65676973",
  1579 => x"74657273",
  1580 => x"3a000000",
  1581 => x"0a636f6e",
  1582 => x"74726f6c",
  1583 => x"3a202020",
  1584 => x"20202000",
  1585 => x"0a737461",
  1586 => x"7475733a",
  1587 => x"20202020",
  1588 => x"20202000",
  1589 => x"0a6d6163",
  1590 => x"5f6d7362",
  1591 => x"3a202020",
  1592 => x"20202000",
  1593 => x"0a6d6163",
  1594 => x"5f6c7362",
  1595 => x"3a202020",
  1596 => x"20202000",
  1597 => x"0a6d6469",
  1598 => x"6f5f636f",
  1599 => x"6e74726f",
  1600 => x"6c3a2000",
  1601 => x"0a74785f",
  1602 => x"706f696e",
  1603 => x"7465723a",
  1604 => x"20202000",
  1605 => x"0a72785f",
  1606 => x"706f696e",
  1607 => x"7465723a",
  1608 => x"20202000",
  1609 => x"0a656463",
  1610 => x"6c5f6970",
  1611 => x"3a202020",
  1612 => x"20202000",
  1613 => x"0a686173",
  1614 => x"685f6d73",
  1615 => x"623a2020",
  1616 => x"20202000",
  1617 => x"0a686173",
  1618 => x"685f6c73",
  1619 => x"623a2020",
  1620 => x"20202000",
  1621 => x"0a6d6469",
  1622 => x"6f207068",
  1623 => x"79207265",
  1624 => x"67697374",
  1625 => x"65727300",
  1626 => x"0a206d64",
  1627 => x"696f2070",
  1628 => x"68793a20",
  1629 => x"00000000",
  1630 => x"0a202072",
  1631 => x"65673a20",
  1632 => x"00000000",
  1633 => x"2d3e2000",
  1634 => x"0a677265",
  1635 => x"74682d3e",
  1636 => x"636f6e74",
  1637 => x"726f6c20",
  1638 => x"3a000000",
  1639 => x"0a677265",
  1640 => x"74682d3e",
  1641 => x"73746174",
  1642 => x"75732020",
  1643 => x"3a000000",
  1644 => x"0a646573",
  1645 => x"63722d3e",
  1646 => x"636f6e74",
  1647 => x"726f6c20",
  1648 => x"3a000000",
  1649 => x"77726974",
  1650 => x"65206164",
  1651 => x"64726573",
  1652 => x"733a2000",
  1653 => x"20206c65",
  1654 => x"6e677468",
  1655 => x"3a200000",
  1656 => x"0a0a0000",
  1657 => x"72656164",
  1658 => x"20206164",
  1659 => x"64726573",
  1660 => x"733a2000",
  1661 => x"20206578",
  1662 => x"70656374",
  1663 => x"3a200000",
  1664 => x"2020676f",
  1665 => x"743a2000",
  1666 => x"20657272",
  1667 => x"6f720000",
  1668 => x"0a000000",
  1669 => x"206f6b00",
  1670 => x"70686173",
  1671 => x"65207368",
  1672 => x"69667420",
  1673 => x"3a200000",
  1674 => x"20202020",
  1675 => x"20000000",
  1676 => x"21000000",
  1677 => x"2e000000",
  1678 => x"44445220",
  1679 => x"6d656d6f",
  1680 => x"72792069",
  1681 => x"6e666f00",
  1682 => x"0a617574",
  1683 => x"6f20745f",
  1684 => x"52455245",
  1685 => x"5348203a",
  1686 => x"00000000",
  1687 => x"0a636c6f",
  1688 => x"636b2065",
  1689 => x"6e61626c",
  1690 => x"6520203a",
  1691 => x"00000000",
  1692 => x"0a696e69",
  1693 => x"74616c69",
  1694 => x"7a652020",
  1695 => x"2020203a",
  1696 => x"00000000",
  1697 => x"0a636f6c",
  1698 => x"756d6e20",
  1699 => x"73697a65",
  1700 => x"2020203a",
  1701 => x"00000000",
  1702 => x"0a62616e",
  1703 => x"6b73697a",
  1704 => x"65202020",
  1705 => x"2020203a",
  1706 => x"00000000",
  1707 => x"4d627974",
  1708 => x"65000000",
  1709 => x"0a745f52",
  1710 => x"43442020",
  1711 => x"20202020",
  1712 => x"2020203a",
  1713 => x"00000000",
  1714 => x"0a745f52",
  1715 => x"46432020",
  1716 => x"20202020",
  1717 => x"2020203a",
  1718 => x"00000000",
  1719 => x"0a745f52",
  1720 => x"50202020",
  1721 => x"20202020",
  1722 => x"2020203a",
  1723 => x"00000000",
  1724 => x"0a726566",
  1725 => x"72657368",
  1726 => x"20656e2e",
  1727 => x"2020203a",
  1728 => x"00000000",
  1729 => x"0a444452",
  1730 => x"20667265",
  1731 => x"7175656e",
  1732 => x"6379203a",
  1733 => x"00000000",
  1734 => x"0a444452",
  1735 => x"20646174",
  1736 => x"61207769",
  1737 => x"6474683a",
  1738 => x"00000000",
  1739 => x"0a6d6f62",
  1740 => x"696c6520",
  1741 => x"73757070",
  1742 => x"6f72743a",
  1743 => x"00000000",
  1744 => x"0a73656c",
  1745 => x"66207265",
  1746 => x"66726573",
  1747 => x"6820203a",
  1748 => x"00000000",
  1749 => x"756e6b6e",
  1750 => x"6f776e00",
  1751 => x"20617272",
  1752 => x"61790000",
  1753 => x"0a74656d",
  1754 => x"702d636f",
  1755 => x"6d702072",
  1756 => x"6566723a",
  1757 => x"00000000",
  1758 => x"c2b04300",
  1759 => x"0a647269",
  1760 => x"76652073",
  1761 => x"7472656e",
  1762 => x"6774683a",
  1763 => x"00000000",
  1764 => x"0a706f77",
  1765 => x"65722073",
  1766 => x"6176696e",
  1767 => x"6720203a",
  1768 => x"00000000",
  1769 => x"0a745f58",
  1770 => x"50202020",
  1771 => x"20202020",
  1772 => x"2020203a",
  1773 => x"00000000",
  1774 => x"0a745f58",
  1775 => x"53522020",
  1776 => x"20202020",
  1777 => x"2020203a",
  1778 => x"00000000",
  1779 => x"0a745f43",
  1780 => x"4b452020",
  1781 => x"20202020",
  1782 => x"2020203a",
  1783 => x"00000000",
  1784 => x"0a434153",
  1785 => x"206c6174",
  1786 => x"656e6379",
  1787 => x"2020203a",
  1788 => x"00000000",
  1789 => x"0a6d6f62",
  1790 => x"696c6520",
  1791 => x"656e6162",
  1792 => x"6c65643a",
  1793 => x"00000000",
  1794 => x"0a737461",
  1795 => x"74757320",
  1796 => x"72656164",
  1797 => x"2020203a",
  1798 => x"00000000",
  1799 => x"332f3400",
  1800 => x"38350000",
  1801 => x"68616c66",
  1802 => x"00000000",
  1803 => x"34303639",
  1804 => x"00000000",
  1805 => x"20353132",
  1806 => x"00000000",
  1807 => x"66756c6c",
  1808 => x"00000000",
  1809 => x"37300000",
  1810 => x"34350000",
  1811 => x"31303234",
  1812 => x"00000000",
  1813 => x"31350000",
  1814 => x"312f3400",
  1815 => x"32303438",
  1816 => x"00000000",
  1817 => x"312f3800",
  1818 => x"312f3200",
  1819 => x"312f3100",
  1820 => x"64656570",
  1821 => x"20706f77",
  1822 => x"65722064",
  1823 => x"6f776e00",
  1824 => x"636c6f63",
  1825 => x"6b207374",
  1826 => x"6f700000",
  1827 => x"73656c66",
  1828 => x"20726566",
  1829 => x"72657368",
  1830 => x"00000000",
  1831 => x"706f7765",
  1832 => x"7220646f",
  1833 => x"776e0000",
  1834 => x"6e6f6e65",
  1835 => x"00000000",
  1836 => x"61646472",
  1837 => x"6573733a",
  1838 => x"20000000",
  1839 => x"20646174",
  1840 => x"613a2000",
  1841 => x"0a0a4443",
  1842 => x"4d207068",
  1843 => x"61736520",
  1844 => x"73686966",
  1845 => x"74207465",
  1846 => x"7374696e",
  1847 => x"67000000",
  1848 => x"0a696e69",
  1849 => x"7469616c",
  1850 => x"3a200000",
  1851 => x"0a6c6f77",
  1852 => x"3a202020",
  1853 => x"20202020",
  1854 => x"20200000",
  1855 => x"0a686967",
  1856 => x"683a2020",
  1857 => x"20202020",
  1858 => x"20200000",
  1859 => x"0a646966",
  1860 => x"663a2020",
  1861 => x"20202020",
  1862 => x"20200000",
  1863 => x"0a646966",
  1864 => x"662f323a",
  1865 => x"20202020",
  1866 => x"20200000",
  1867 => x"0a6d696e",
  1868 => x"5f657272",
  1869 => x"3a202020",
  1870 => x"20200000",
  1871 => x"0a6d696e",
  1872 => x"5f657272",
  1873 => x"5f706f73",
  1874 => x"3a200000",
  1875 => x"0a66696e",
  1876 => x"616c3a20",
  1877 => x"20202020",
  1878 => x"20200000",
  1879 => x"696e6974",
  1880 => x"20646f6e",
  1881 => x"652e0000",
  1882 => x"74657374",
  1883 => x"2e632000",
  1884 => x"286f6e20",
  1885 => x"73696d75",
  1886 => x"6c61746f",
  1887 => x"72290a00",
  1888 => x"636f6d70",
  1889 => x"696c6564",
  1890 => x"3a205365",
  1891 => x"70203133",
  1892 => x"20323031",
  1893 => x"30202031",
  1894 => x"373a3233",
  1895 => x"3a33370a",
  1896 => x"00000000",
  1897 => x"286f6e20",
  1898 => x"68617264",
  1899 => x"77617265",
  1900 => x"290a0000",
  1901 => x"64756d6d",
  1902 => x"792e6578",
  1903 => x"65000000",
  1904 => x"43000000",
  1905 => x"00ffffff",
  1906 => x"ff00ffff",
  1907 => x"ffff00ff",
  1908 => x"ffffff00",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"0000218c",
  1913 => x"80000e00",
  1914 => x"80000c00",
  1915 => x"80000800",
  1916 => x"80000600",
  1917 => x"80000200",
  1918 => x"80000100",
  1919 => x"00001db4",
  1920 => x"00001e04",
  1921 => x"00000000",
  1922 => x"0000206c",
  1923 => x"000020c8",
  1924 => x"00002124",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"00000000",
  1931 => x"00000000",
  1932 => x"00000000",
  1933 => x"00000000",
  1934 => x"00001dc0",
  1935 => x"00000000",
  1936 => x"00000000",
  1937 => x"00000000",
  1938 => x"00000000",
  1939 => x"00000000",
  1940 => x"00000000",
  1941 => x"00000000",
  1942 => x"00000000",
  1943 => x"00000000",
  1944 => x"00000000",
  1945 => x"00000000",
  1946 => x"00000000",
  1947 => x"00000000",
  1948 => x"00000000",
  1949 => x"00000000",
  1950 => x"00000000",
  1951 => x"00000000",
  1952 => x"00000000",
  1953 => x"00000000",
  1954 => x"00000000",
  1955 => x"00000000",
  1956 => x"00000000",
  1957 => x"00000000",
  1958 => x"00000000",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00000000",
  1962 => x"00000000",
  1963 => x"00000001",
  1964 => x"330eabcd",
  1965 => x"1234e66d",
  1966 => x"deec0005",
  1967 => x"000b0000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00000000",
  1984 => x"00000000",
  1985 => x"00000000",
  1986 => x"00000000",
  1987 => x"00000000",
  1988 => x"00000000",
  1989 => x"00000000",
  1990 => x"00000000",
  1991 => x"00000000",
  1992 => x"00000000",
  1993 => x"00000000",
  1994 => x"00000000",
  1995 => x"00000000",
  1996 => x"00000000",
  1997 => x"00000000",
  1998 => x"00000000",
  1999 => x"00000000",
  2000 => x"00000000",
  2001 => x"00000000",
  2002 => x"00000000",
  2003 => x"00000000",
  2004 => x"00000000",
  2005 => x"00000000",
  2006 => x"00000000",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00000000",
  2010 => x"00000000",
  2011 => x"00000000",
  2012 => x"00000000",
  2013 => x"00000000",
  2014 => x"00000000",
  2015 => x"00000000",
  2016 => x"00000000",
  2017 => x"00000000",
  2018 => x"00000000",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00000000",
  2026 => x"00000000",
  2027 => x"00000000",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000000",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"00000000",
  2049 => x"00000000",
  2050 => x"00000000",
  2051 => x"00000000",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"ffffffff",
  2145 => x"00000000",
  2146 => x"ffffffff",
  2147 => x"00000000",
  2148 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
