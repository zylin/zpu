-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0bbccc0c",
     3 => x"3a0b0b0b",
     4 => x"b5860400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0bb5c82d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bbc",
   162 => x"b8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0bb1",
   171 => x"8a2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bb2",
   179 => x"bc2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bbcc80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81fb3fae",
   257 => x"e83f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104bc",
   280 => x"c808802e",
   281 => x"a338bccc",
   282 => x"08822ebd",
   283 => x"38838080",
   284 => x"0b0b0b80",
   285 => x"c4800c82",
   286 => x"a0800b80",
   287 => x"c4840c82",
   288 => x"90800b80",
   289 => x"c4880c04",
   290 => x"f8808080",
   291 => x"a40b0b0b",
   292 => x"80c4800c",
   293 => x"f8808082",
   294 => x"800b80c4",
   295 => x"840cf880",
   296 => x"8084800b",
   297 => x"80c4880c",
   298 => x"0480c0a8",
   299 => x"808c0b0b",
   300 => x"0b80c480",
   301 => x"0c80c0a8",
   302 => x"80940b80",
   303 => x"c4840c0b",
   304 => x"0b0bb798",
   305 => x"0b80c488",
   306 => x"0c04ff3d",
   307 => x"0d80c48c",
   308 => x"335170a4",
   309 => x"38bcd408",
   310 => x"70085252",
   311 => x"70802e92",
   312 => x"388412bc",
   313 => x"d40c702d",
   314 => x"bcd40870",
   315 => x"08525270",
   316 => x"f038810b",
   317 => x"80c48c34",
   318 => x"833d0d04",
   319 => x"04803d0d",
   320 => x"0b0b80c3",
   321 => x"fc08802e",
   322 => x"8e380b0b",
   323 => x"0b0b800b",
   324 => x"802e0981",
   325 => x"06853882",
   326 => x"3d0d040b",
   327 => x"0b80c3fc",
   328 => x"510b0b0b",
   329 => x"f5da3f82",
   330 => x"3d0d0404",
   331 => x"fd3d0dbc",
   332 => x"e00876b0",
   333 => x"ea299412",
   334 => x"0c54850b",
   335 => x"98150c98",
   336 => x"14087081",
   337 => x"06515372",
   338 => x"f638853d",
   339 => x"0d04ff3d",
   340 => x"0dbce008",
   341 => x"74101075",
   342 => x"10059412",
   343 => x"0c52850b",
   344 => x"98130c98",
   345 => x"12087081",
   346 => x"06515170",
   347 => x"f638833d",
   348 => x"0d04803d",
   349 => x"0d725180",
   350 => x"71278738",
   351 => x"ff115170",
   352 => x"fb38823d",
   353 => x"0d04803d",
   354 => x"0dbce008",
   355 => x"51870b84",
   356 => x"120c823d",
   357 => x"0d04803d",
   358 => x"0dbce408",
   359 => x"51b60b8c",
   360 => x"120c830b",
   361 => x"88120c82",
   362 => x"3d0d04ff",
   363 => x"3d0dbce4",
   364 => x"08528412",
   365 => x"08708106",
   366 => x"51517080",
   367 => x"2ef43871",
   368 => x"087081ff",
   369 => x"06800c51",
   370 => x"833d0d04",
   371 => x"fe3d0d02",
   372 => x"930533bc",
   373 => x"e4085353",
   374 => x"84120870",
   375 => x"892a7081",
   376 => x"06515151",
   377 => x"70f23872",
   378 => x"720c843d",
   379 => x"0d04fe3d",
   380 => x"0d029305",
   381 => x"3353728a",
   382 => x"2e9b38bc",
   383 => x"e4085284",
   384 => x"12087089",
   385 => x"2a708106",
   386 => x"51515170",
   387 => x"f2387272",
   388 => x"0c843d0d",
   389 => x"04bce408",
   390 => x"52841208",
   391 => x"70892a70",
   392 => x"81065151",
   393 => x"5170f238",
   394 => x"8d720c84",
   395 => x"12087089",
   396 => x"2a708106",
   397 => x"51515170",
   398 => x"c638d339",
   399 => x"fd3d0d75",
   400 => x"70335254",
   401 => x"70802ea7",
   402 => x"3870bce4",
   403 => x"08535381",
   404 => x"1454728a",
   405 => x"2e9d3884",
   406 => x"12087089",
   407 => x"2a708106",
   408 => x"51515170",
   409 => x"f2387272",
   410 => x"0c733353",
   411 => x"72e13885",
   412 => x"3d0d0484",
   413 => x"12087089",
   414 => x"2a708106",
   415 => x"51515170",
   416 => x"f2388d72",
   417 => x"0c841208",
   418 => x"70892a70",
   419 => x"81065151",
   420 => x"5170c438",
   421 => x"d139f83d",
   422 => x"0d7a7c59",
   423 => x"53807356",
   424 => x"57767324",
   425 => x"80dc3877",
   426 => x"17548a52",
   427 => x"7451a3b5",
   428 => x"3f8008b0",
   429 => x"05537274",
   430 => x"34811757",
   431 => x"8a527451",
   432 => x"a2fe3f80",
   433 => x"08558008",
   434 => x"de388008",
   435 => x"779f2a18",
   436 => x"70812c5b",
   437 => x"56568079",
   438 => x"259e3877",
   439 => x"17ff0555",
   440 => x"75187033",
   441 => x"55537433",
   442 => x"73347375",
   443 => x"348116ff",
   444 => x"16565678",
   445 => x"7624e938",
   446 => x"76185680",
   447 => x"76348a3d",
   448 => x"0d04ad78",
   449 => x"7081055a",
   450 => x"34723078",
   451 => x"1855558a",
   452 => x"527451a2",
   453 => x"d03f8008",
   454 => x"b0055372",
   455 => x"74348117",
   456 => x"578a5274",
   457 => x"51a2993f",
   458 => x"80085580",
   459 => x"08fef838",
   460 => x"ff983980",
   461 => x"3d0dbcdc",
   462 => x"085181ff",
   463 => x"0b88120c",
   464 => x"823d0d04",
   465 => x"fb3d0d88",
   466 => x"80e0870b",
   467 => x"bcdc08bc",
   468 => x"e0087284",
   469 => x"130c5657",
   470 => x"55afd7c2",
   471 => x"0b94150c",
   472 => x"850b9815",
   473 => x"0c981408",
   474 => x"70810651",
   475 => x"5372f638",
   476 => x"749f2a75",
   477 => x"10077084",
   478 => x"180c55af",
   479 => x"d7c20b94",
   480 => x"150c850b",
   481 => x"98150cdd",
   482 => x"39fd3d0d",
   483 => x"bcdc0854",
   484 => x"80d50b84",
   485 => x"150cbce4",
   486 => x"08528412",
   487 => x"08810651",
   488 => x"70802ef6",
   489 => x"38710870",
   490 => x"81ff06f6",
   491 => x"11525451",
   492 => x"70ae268b",
   493 => x"38701010",
   494 => x"b79c0551",
   495 => x"70080484",
   496 => x"12087089",
   497 => x"2a708106",
   498 => x"51515170",
   499 => x"f238ab72",
   500 => x"0c728a2e",
   501 => x"a6388412",
   502 => x"0870892a",
   503 => x"70810651",
   504 => x"515170f2",
   505 => x"3872720c",
   506 => x"84120870",
   507 => x"892a8106",
   508 => x"515372f4",
   509 => x"38ad720c",
   510 => x"ffa03984",
   511 => x"12087089",
   512 => x"2a708106",
   513 => x"51515170",
   514 => x"f2388d72",
   515 => x"0c841208",
   516 => x"70892a70",
   517 => x"81065151",
   518 => x"5170ffba",
   519 => x"38c73981",
   520 => x"ff0b8415",
   521 => x"0cfef339",
   522 => x"80ff0b84",
   523 => x"150cfeea",
   524 => x"39bf0b84",
   525 => x"150cfee2",
   526 => x"399f0b84",
   527 => x"150cfeda",
   528 => x"398f0b84",
   529 => x"150cfed2",
   530 => x"39870b84",
   531 => x"150cfeca",
   532 => x"39830b84",
   533 => x"150cfec2",
   534 => x"39810b84",
   535 => x"150cfeba",
   536 => x"39800b84",
   537 => x"150cfeb2",
   538 => x"39ff3d0d",
   539 => x"bcdc0852",
   540 => x"7108708f",
   541 => x"06707184",
   542 => x"2b078415",
   543 => x"0c515171",
   544 => x"08708f06",
   545 => x"7071842b",
   546 => x"0784150c",
   547 => x"5151e139",
   548 => x"f23d0dba",
   549 => x"940bba94",
   550 => x"33545672",
   551 => x"802ea638",
   552 => x"72bce408",
   553 => x"55558116",
   554 => x"56748a2e",
   555 => x"90b63884",
   556 => x"14087089",
   557 => x"2a81065a",
   558 => x"5378f438",
   559 => x"74740c75",
   560 => x"335574e2",
   561 => x"38baa80b",
   562 => x"baa83354",
   563 => x"5672802e",
   564 => x"a638bce4",
   565 => x"08735654",
   566 => x"81165674",
   567 => x"8a2e90a5",
   568 => x"38841408",
   569 => x"70892a81",
   570 => x"065b5779",
   571 => x"f4387474",
   572 => x"0c753355",
   573 => x"74e238bc",
   574 => x"d8087008",
   575 => x"8d3d705c",
   576 => x"5c545480",
   577 => x"73565776",
   578 => x"7324909a",
   579 => x"38781756",
   580 => x"8a527451",
   581 => x"9ecf3f80",
   582 => x"08b00558",
   583 => x"77763481",
   584 => x"17578a52",
   585 => x"74519e98",
   586 => x"3f800855",
   587 => x"8008de38",
   588 => x"8008779f",
   589 => x"2a187081",
   590 => x"2c5a5656",
   591 => x"8078259e",
   592 => x"387817ff",
   593 => x"05557519",
   594 => x"70335553",
   595 => x"74337334",
   596 => x"73753481",
   597 => x"16ff1656",
   598 => x"56777624",
   599 => x"e9387619",
   600 => x"56807634",
   601 => x"797a3354",
   602 => x"5672802e",
   603 => x"a638bce4",
   604 => x"08735654",
   605 => x"81165674",
   606 => x"8a2e8fdb",
   607 => x"38841408",
   608 => x"70892a81",
   609 => x"06545772",
   610 => x"f4387474",
   611 => x"0c753355",
   612 => x"74e238ba",
   613 => x"b80bbab8",
   614 => x"33545672",
   615 => x"802ea638",
   616 => x"bce40873",
   617 => x"56548116",
   618 => x"56748a2e",
   619 => x"8fca3884",
   620 => x"14087089",
   621 => x"2a810658",
   622 => x"5376f438",
   623 => x"74740c75",
   624 => x"335574e2",
   625 => x"38bcd808",
   626 => x"8411087b",
   627 => x"5b545580",
   628 => x"73565776",
   629 => x"732496fa",
   630 => x"38781754",
   631 => x"8a527451",
   632 => x"9d833f80",
   633 => x"08b00556",
   634 => x"75743481",
   635 => x"17578a52",
   636 => x"74519ccc",
   637 => x"3f800855",
   638 => x"8008de38",
   639 => x"8008779f",
   640 => x"2a187081",
   641 => x"2c5a5456",
   642 => x"8078259e",
   643 => x"387817ff",
   644 => x"05557519",
   645 => x"70335553",
   646 => x"74337334",
   647 => x"73753481",
   648 => x"16ff1656",
   649 => x"56777624",
   650 => x"e9387619",
   651 => x"58807834",
   652 => x"797a3354",
   653 => x"5672802e",
   654 => x"a638bce4",
   655 => x"08735654",
   656 => x"81165674",
   657 => x"8a2e8ed1",
   658 => x"38841408",
   659 => x"70892a81",
   660 => x"06595777",
   661 => x"f4387474",
   662 => x"0c753355",
   663 => x"74e238ba",
   664 => x"c80bbac8",
   665 => x"33545672",
   666 => x"802ea638",
   667 => x"bce40873",
   668 => x"56548116",
   669 => x"56748a2e",
   670 => x"8ec03884",
   671 => x"14087089",
   672 => x"2a810658",
   673 => x"5876f438",
   674 => x"74740c75",
   675 => x"335574e2",
   676 => x"38bcd808",
   677 => x"8811087b",
   678 => x"5b545580",
   679 => x"73565776",
   680 => x"732494fd",
   681 => x"38781756",
   682 => x"8a527451",
   683 => x"9bb73f80",
   684 => x"08b00554",
   685 => x"73763481",
   686 => x"17578a52",
   687 => x"74519b80",
   688 => x"3f800855",
   689 => x"8008de38",
   690 => x"8008779f",
   691 => x"2a187081",
   692 => x"2c5a5456",
   693 => x"8078259e",
   694 => x"387817ff",
   695 => x"05557519",
   696 => x"70335553",
   697 => x"74337334",
   698 => x"73753481",
   699 => x"16ff1656",
   700 => x"56777624",
   701 => x"e9387619",
   702 => x"58807834",
   703 => x"797a3354",
   704 => x"5672802e",
   705 => x"a638bce4",
   706 => x"08735654",
   707 => x"81165674",
   708 => x"8a2e8dc7",
   709 => x"38841408",
   710 => x"70892a81",
   711 => x"06595777",
   712 => x"f4387474",
   713 => x"0c753355",
   714 => x"74e238ba",
   715 => x"d80bbad8",
   716 => x"33545672",
   717 => x"802ea638",
   718 => x"bce40873",
   719 => x"56548116",
   720 => x"56748a2e",
   721 => x"8db63884",
   722 => x"14087089",
   723 => x"2a810658",
   724 => x"5876f438",
   725 => x"74740c75",
   726 => x"335574e2",
   727 => x"38bcd808",
   728 => x"8c11087b",
   729 => x"5b545580",
   730 => x"73565776",
   731 => x"73249380",
   732 => x"38781756",
   733 => x"8a527451",
   734 => x"99eb3f80",
   735 => x"08b00554",
   736 => x"73763481",
   737 => x"17578a52",
   738 => x"745199b4",
   739 => x"3f800855",
   740 => x"8008de38",
   741 => x"8008779f",
   742 => x"2a187081",
   743 => x"2c5a5456",
   744 => x"8078259e",
   745 => x"387817ff",
   746 => x"05557519",
   747 => x"70335553",
   748 => x"74337334",
   749 => x"73753481",
   750 => x"16ff1656",
   751 => x"56777624",
   752 => x"e9387619",
   753 => x"58807834",
   754 => x"797a3354",
   755 => x"5672802e",
   756 => x"a638bce4",
   757 => x"08735654",
   758 => x"81165674",
   759 => x"8a2e8cbd",
   760 => x"38841408",
   761 => x"70892a81",
   762 => x"06595777",
   763 => x"f4387474",
   764 => x"0c753355",
   765 => x"74e238ba",
   766 => x"e80bbae8",
   767 => x"33545672",
   768 => x"802ea638",
   769 => x"bce40873",
   770 => x"56548116",
   771 => x"56748a2e",
   772 => x"8cac3884",
   773 => x"14087089",
   774 => x"2a810658",
   775 => x"5876f438",
   776 => x"74740c75",
   777 => x"335574e2",
   778 => x"38bcd808",
   779 => x"9011087b",
   780 => x"5b545580",
   781 => x"73565776",
   782 => x"73249183",
   783 => x"38781756",
   784 => x"8a527451",
   785 => x"989f3f80",
   786 => x"08b00554",
   787 => x"73763481",
   788 => x"17578a52",
   789 => x"745197e8",
   790 => x"3f800855",
   791 => x"8008de38",
   792 => x"8008779f",
   793 => x"2a187081",
   794 => x"2c5a5456",
   795 => x"8078259e",
   796 => x"387817ff",
   797 => x"05557519",
   798 => x"70335553",
   799 => x"74337334",
   800 => x"73753481",
   801 => x"16ff1656",
   802 => x"56777624",
   803 => x"e9387619",
   804 => x"58807834",
   805 => x"797a3354",
   806 => x"5672802e",
   807 => x"a638bce4",
   808 => x"08735654",
   809 => x"81165674",
   810 => x"8a2e8bb3",
   811 => x"38841408",
   812 => x"70892a81",
   813 => x"06595777",
   814 => x"f4387474",
   815 => x"0c753355",
   816 => x"74e238ba",
   817 => x"f80bbaf8",
   818 => x"33545672",
   819 => x"802ea638",
   820 => x"bce40873",
   821 => x"56548116",
   822 => x"56748a2e",
   823 => x"8ba23884",
   824 => x"14087089",
   825 => x"2a810658",
   826 => x"5876f438",
   827 => x"74740c75",
   828 => x"335574e2",
   829 => x"38bcd808",
   830 => x"9411087b",
   831 => x"5b545580",
   832 => x"73565776",
   833 => x"73248f86",
   834 => x"38781756",
   835 => x"8a527451",
   836 => x"96d33f80",
   837 => x"08b00554",
   838 => x"73763481",
   839 => x"17578a52",
   840 => x"7451969c",
   841 => x"3f800855",
   842 => x"8008de38",
   843 => x"8008779f",
   844 => x"2a187081",
   845 => x"2c5a5456",
   846 => x"8078259e",
   847 => x"387817ff",
   848 => x"05557519",
   849 => x"70335553",
   850 => x"74337334",
   851 => x"73753481",
   852 => x"16ff1656",
   853 => x"56777624",
   854 => x"e9387619",
   855 => x"58807834",
   856 => x"797a3354",
   857 => x"5672802e",
   858 => x"a638bce4",
   859 => x"08735654",
   860 => x"81165674",
   861 => x"8a2e8aa9",
   862 => x"38841408",
   863 => x"70892a81",
   864 => x"06595777",
   865 => x"f4387474",
   866 => x"0c753355",
   867 => x"74e238bb",
   868 => x"880bbb88",
   869 => x"33545672",
   870 => x"802ea638",
   871 => x"bce40873",
   872 => x"56548116",
   873 => x"56748a2e",
   874 => x"8a983884",
   875 => x"14087089",
   876 => x"2a810658",
   877 => x"5876f438",
   878 => x"74740c75",
   879 => x"335574e2",
   880 => x"38bcd808",
   881 => x"9811087b",
   882 => x"5b545580",
   883 => x"73565776",
   884 => x"73248d89",
   885 => x"38781756",
   886 => x"8a527451",
   887 => x"95873f80",
   888 => x"08b00554",
   889 => x"73763481",
   890 => x"17578a52",
   891 => x"745194d0",
   892 => x"3f800855",
   893 => x"8008de38",
   894 => x"8008779f",
   895 => x"2a187081",
   896 => x"2c5a5456",
   897 => x"8078259e",
   898 => x"387817ff",
   899 => x"05557519",
   900 => x"70335553",
   901 => x"74337334",
   902 => x"73753481",
   903 => x"16ff1656",
   904 => x"56777624",
   905 => x"e9387619",
   906 => x"58807834",
   907 => x"797a3354",
   908 => x"5672802e",
   909 => x"a638bce4",
   910 => x"08735654",
   911 => x"81165674",
   912 => x"8a2e899f",
   913 => x"38841408",
   914 => x"70892a81",
   915 => x"06595777",
   916 => x"f4387474",
   917 => x"0c753355",
   918 => x"74e238bb",
   919 => x"980bbb98",
   920 => x"33545672",
   921 => x"802ea638",
   922 => x"bce40873",
   923 => x"56548116",
   924 => x"56748a2e",
   925 => x"898e3884",
   926 => x"14087089",
   927 => x"2a810658",
   928 => x"5876f438",
   929 => x"74740c75",
   930 => x"335574e2",
   931 => x"38bcd808",
   932 => x"9c11087b",
   933 => x"5b545580",
   934 => x"73565776",
   935 => x"73248b8c",
   936 => x"38781756",
   937 => x"8a527451",
   938 => x"93bb3f80",
   939 => x"08b00554",
   940 => x"73763481",
   941 => x"17578a52",
   942 => x"74519384",
   943 => x"3f800855",
   944 => x"8008de38",
   945 => x"8008779f",
   946 => x"2a187081",
   947 => x"2c5a5456",
   948 => x"8078259e",
   949 => x"387817ff",
   950 => x"05557519",
   951 => x"70335553",
   952 => x"74337334",
   953 => x"73753481",
   954 => x"16ff1656",
   955 => x"56777624",
   956 => x"e9387619",
   957 => x"58807834",
   958 => x"797a3354",
   959 => x"5672802e",
   960 => x"a638bce4",
   961 => x"08735654",
   962 => x"81165674",
   963 => x"8a2e8895",
   964 => x"38841408",
   965 => x"70892a81",
   966 => x"06595777",
   967 => x"f4387474",
   968 => x"0c753355",
   969 => x"74e238bb",
   970 => x"a80bbba8",
   971 => x"33545672",
   972 => x"802ea638",
   973 => x"bce40873",
   974 => x"56548116",
   975 => x"56748a2e",
   976 => x"88843884",
   977 => x"14087089",
   978 => x"2a810658",
   979 => x"5876f438",
   980 => x"74740c75",
   981 => x"335574e2",
   982 => x"38bcd808",
   983 => x"a011087b",
   984 => x"5b545580",
   985 => x"73565776",
   986 => x"7324898f",
   987 => x"38781756",
   988 => x"8a527451",
   989 => x"91ef3f80",
   990 => x"08b00554",
   991 => x"73763481",
   992 => x"17578a52",
   993 => x"745191b8",
   994 => x"3f800855",
   995 => x"8008de38",
   996 => x"8008779f",
   997 => x"2a187081",
   998 => x"2c5a5456",
   999 => x"8078259e",
  1000 => x"387817ff",
  1001 => x"05557519",
  1002 => x"70335553",
  1003 => x"74337334",
  1004 => x"73753481",
  1005 => x"16ff1656",
  1006 => x"56777624",
  1007 => x"e9387619",
  1008 => x"58807834",
  1009 => x"797a3354",
  1010 => x"5672802e",
  1011 => x"a638bce4",
  1012 => x"08735654",
  1013 => x"81165674",
  1014 => x"8a2e878b",
  1015 => x"38841408",
  1016 => x"70892a81",
  1017 => x"06595777",
  1018 => x"f4387474",
  1019 => x"0c753355",
  1020 => x"74e238bb",
  1021 => x"b80bbbb8",
  1022 => x"33545672",
  1023 => x"802ea638",
  1024 => x"bce40873",
  1025 => x"56548116",
  1026 => x"56748a2e",
  1027 => x"86fa3884",
  1028 => x"14087089",
  1029 => x"2a810658",
  1030 => x"5876f438",
  1031 => x"74740c75",
  1032 => x"335574e2",
  1033 => x"38bcd808",
  1034 => x"a411087b",
  1035 => x"5b545580",
  1036 => x"73565776",
  1037 => x"73248792",
  1038 => x"38781756",
  1039 => x"8a527451",
  1040 => x"90a33f80",
  1041 => x"08b00554",
  1042 => x"73763481",
  1043 => x"17578a52",
  1044 => x"74518fec",
  1045 => x"3f800855",
  1046 => x"8008de38",
  1047 => x"8008779f",
  1048 => x"2a187081",
  1049 => x"2c5a5456",
  1050 => x"8078259e",
  1051 => x"387817ff",
  1052 => x"05557519",
  1053 => x"70335553",
  1054 => x"74337334",
  1055 => x"73753481",
  1056 => x"16ff1656",
  1057 => x"56777624",
  1058 => x"e9387619",
  1059 => x"58807834",
  1060 => x"797a3354",
  1061 => x"5672802e",
  1062 => x"89e938bc",
  1063 => x"e4087356",
  1064 => x"54811656",
  1065 => x"748a2e86",
  1066 => x"80388414",
  1067 => x"0870892a",
  1068 => x"8106545a",
  1069 => x"72f43874",
  1070 => x"740c7533",
  1071 => x"5574e238",
  1072 => x"84140870",
  1073 => x"892a8106",
  1074 => x"565974f4",
  1075 => x"388d740c",
  1076 => x"84140870",
  1077 => x"892a8106",
  1078 => x"585876f4",
  1079 => x"388a740c",
  1080 => x"903d0d04",
  1081 => x"84140870",
  1082 => x"892a8106",
  1083 => x"545872f4",
  1084 => x"388d740c",
  1085 => x"84140870",
  1086 => x"892a8106",
  1087 => x"5a5378ef",
  1088 => x"ae38efb8",
  1089 => x"39841408",
  1090 => x"70892a81",
  1091 => x"06585976",
  1092 => x"f4388d74",
  1093 => x"0c841408",
  1094 => x"70892a81",
  1095 => x"065b5779",
  1096 => x"efbf38ef",
  1097 => x"c939ad7a",
  1098 => x"3402a905",
  1099 => x"73307119",
  1100 => x"5856598a",
  1101 => x"5274518e",
  1102 => x"ac3f8008",
  1103 => x"b0055877",
  1104 => x"76348117",
  1105 => x"578a5274",
  1106 => x"518df53f",
  1107 => x"80085580",
  1108 => x"08efba38",
  1109 => x"efda3984",
  1110 => x"14087089",
  1111 => x"2a81065a",
  1112 => x"5878f438",
  1113 => x"8d740c84",
  1114 => x"14087089",
  1115 => x"2a810654",
  1116 => x"5772f089",
  1117 => x"38f09339",
  1118 => x"84140870",
  1119 => x"892a8106",
  1120 => x"595977f4",
  1121 => x"388d740c",
  1122 => x"84140870",
  1123 => x"892a8106",
  1124 => x"585376f0",
  1125 => x"9a38f0a4",
  1126 => x"39841408",
  1127 => x"70892a81",
  1128 => x"065a5378",
  1129 => x"f4388d74",
  1130 => x"0c841408",
  1131 => x"70892a81",
  1132 => x"06595777",
  1133 => x"f19338f1",
  1134 => x"9d398414",
  1135 => x"0870892a",
  1136 => x"81065459",
  1137 => x"72f4388d",
  1138 => x"740c8414",
  1139 => x"0870892a",
  1140 => x"81065858",
  1141 => x"76f1a438",
  1142 => x"f1ae3984",
  1143 => x"14087089",
  1144 => x"2a81065a",
  1145 => x"5378f438",
  1146 => x"8d740c84",
  1147 => x"14087089",
  1148 => x"2a810659",
  1149 => x"5777f29d",
  1150 => x"38f2a739",
  1151 => x"84140870",
  1152 => x"892a8106",
  1153 => x"545972f4",
  1154 => x"388d740c",
  1155 => x"84140870",
  1156 => x"892a8106",
  1157 => x"585876f2",
  1158 => x"ae38f2b8",
  1159 => x"39841408",
  1160 => x"70892a81",
  1161 => x"065a5378",
  1162 => x"f4388d74",
  1163 => x"0c841408",
  1164 => x"70892a81",
  1165 => x"06595777",
  1166 => x"f3a738f3",
  1167 => x"b1398414",
  1168 => x"0870892a",
  1169 => x"81065459",
  1170 => x"72f4388d",
  1171 => x"740c8414",
  1172 => x"0870892a",
  1173 => x"81065858",
  1174 => x"76f3b838",
  1175 => x"f3c23984",
  1176 => x"14087089",
  1177 => x"2a81065a",
  1178 => x"5378f438",
  1179 => x"8d740c84",
  1180 => x"14087089",
  1181 => x"2a810659",
  1182 => x"5777f4b1",
  1183 => x"38f4bb39",
  1184 => x"84140870",
  1185 => x"892a8106",
  1186 => x"545972f4",
  1187 => x"388d740c",
  1188 => x"84140870",
  1189 => x"892a8106",
  1190 => x"585876f4",
  1191 => x"c238f4cc",
  1192 => x"39841408",
  1193 => x"70892a81",
  1194 => x"065a5378",
  1195 => x"f4388d74",
  1196 => x"0c841408",
  1197 => x"70892a81",
  1198 => x"06595777",
  1199 => x"f5bb38f5",
  1200 => x"c5398414",
  1201 => x"0870892a",
  1202 => x"81065459",
  1203 => x"72f4388d",
  1204 => x"740c8414",
  1205 => x"0870892a",
  1206 => x"81065858",
  1207 => x"76f5cc38",
  1208 => x"f5d63984",
  1209 => x"14087089",
  1210 => x"2a81065a",
  1211 => x"5378f438",
  1212 => x"8d740c84",
  1213 => x"14087089",
  1214 => x"2a810659",
  1215 => x"5777f6c5",
  1216 => x"38f6cf39",
  1217 => x"84140870",
  1218 => x"892a8106",
  1219 => x"545972f4",
  1220 => x"388d740c",
  1221 => x"84140870",
  1222 => x"892a8106",
  1223 => x"585876f6",
  1224 => x"d638f6e0",
  1225 => x"39841408",
  1226 => x"70892a81",
  1227 => x"065a5378",
  1228 => x"f4388d74",
  1229 => x"0c841408",
  1230 => x"70892a81",
  1231 => x"06595777",
  1232 => x"f7cf38f7",
  1233 => x"d9398414",
  1234 => x"0870892a",
  1235 => x"81065459",
  1236 => x"72f4388d",
  1237 => x"740c8414",
  1238 => x"0870892a",
  1239 => x"81065858",
  1240 => x"76f7e038",
  1241 => x"f7ea3984",
  1242 => x"14087089",
  1243 => x"2a81065a",
  1244 => x"5378f438",
  1245 => x"8d740c84",
  1246 => x"14087089",
  1247 => x"2a810659",
  1248 => x"5777f8d9",
  1249 => x"38f8e339",
  1250 => x"84140870",
  1251 => x"892a8106",
  1252 => x"545972f4",
  1253 => x"388d740c",
  1254 => x"84140870",
  1255 => x"892a8106",
  1256 => x"585876f8",
  1257 => x"ea38f8f4",
  1258 => x"39841408",
  1259 => x"70892a81",
  1260 => x"065b5779",
  1261 => x"f4388d74",
  1262 => x"0c841408",
  1263 => x"70892a81",
  1264 => x"06545a72",
  1265 => x"f9e438f9",
  1266 => x"ee39ad7a",
  1267 => x"3402a905",
  1268 => x"73307119",
  1269 => x"5856598a",
  1270 => x"52745189",
  1271 => x"883f8008",
  1272 => x"b0055473",
  1273 => x"76348117",
  1274 => x"578a5274",
  1275 => x"5188d13f",
  1276 => x"80085580",
  1277 => x"08f8c238",
  1278 => x"f8e239ad",
  1279 => x"7a3402a9",
  1280 => x"05733071",
  1281 => x"19585659",
  1282 => x"8a527451",
  1283 => x"88d73f80",
  1284 => x"08b00554",
  1285 => x"73763481",
  1286 => x"17578a52",
  1287 => x"745188a0",
  1288 => x"3f800855",
  1289 => x"8008f6c5",
  1290 => x"38f6e539",
  1291 => x"ad7a3402",
  1292 => x"a9057330",
  1293 => x"71195856",
  1294 => x"598a5274",
  1295 => x"5188a63f",
  1296 => x"8008b005",
  1297 => x"54737634",
  1298 => x"8117578a",
  1299 => x"52745187",
  1300 => x"ef3f8008",
  1301 => x"558008f4",
  1302 => x"c838f4e8",
  1303 => x"39ad7a34",
  1304 => x"02a90573",
  1305 => x"30711958",
  1306 => x"56598a52",
  1307 => x"745187f5",
  1308 => x"3f8008b0",
  1309 => x"05547376",
  1310 => x"34811757",
  1311 => x"8a527451",
  1312 => x"87be3f80",
  1313 => x"08558008",
  1314 => x"f2cb38f2",
  1315 => x"eb39ad7a",
  1316 => x"3402a905",
  1317 => x"73307119",
  1318 => x"5856598a",
  1319 => x"52745187",
  1320 => x"c43f8008",
  1321 => x"b0055473",
  1322 => x"76348117",
  1323 => x"578a5274",
  1324 => x"51878d3f",
  1325 => x"80085580",
  1326 => x"08f0ce38",
  1327 => x"f0ee39ad",
  1328 => x"7a3402a9",
  1329 => x"05733071",
  1330 => x"19585659",
  1331 => x"8a527451",
  1332 => x"87933f80",
  1333 => x"08b00554",
  1334 => x"73763481",
  1335 => x"17578a52",
  1336 => x"745186dc",
  1337 => x"3f800855",
  1338 => x"8008eed1",
  1339 => x"38eef139",
  1340 => x"ad7a3402",
  1341 => x"a9057330",
  1342 => x"71195856",
  1343 => x"598a5274",
  1344 => x"5186e23f",
  1345 => x"8008b005",
  1346 => x"54737634",
  1347 => x"8117578a",
  1348 => x"52745186",
  1349 => x"ab3f8008",
  1350 => x"558008ec",
  1351 => x"d438ecf4",
  1352 => x"39ad7a34",
  1353 => x"02a90573",
  1354 => x"30711958",
  1355 => x"56598a52",
  1356 => x"745186b1",
  1357 => x"3f8008b0",
  1358 => x"05547376",
  1359 => x"34811757",
  1360 => x"8a527451",
  1361 => x"85fa3f80",
  1362 => x"08558008",
  1363 => x"ead738ea",
  1364 => x"f739ad7a",
  1365 => x"3402a905",
  1366 => x"73307119",
  1367 => x"5656598a",
  1368 => x"52745186",
  1369 => x"803f8008",
  1370 => x"b0055675",
  1371 => x"74348117",
  1372 => x"578a5274",
  1373 => x"5185c93f",
  1374 => x"80085580",
  1375 => x"08e8da38",
  1376 => x"e8fa39bc",
  1377 => x"e4088411",
  1378 => x"0870892a",
  1379 => x"8106575a",
  1380 => x"5474f6ac",
  1381 => x"38f6b639",
  1382 => x"fa3d0dbc",
  1383 => x"dc087008",
  1384 => x"810a06bc",
  1385 => x"e0085558",
  1386 => x"55870b84",
  1387 => x"140cbce4",
  1388 => x"0854b60b",
  1389 => x"8c150c83",
  1390 => x"0b88150c",
  1391 => x"bbc80bbb",
  1392 => x"c8335456",
  1393 => x"72802ea4",
  1394 => x"38725581",
  1395 => x"1656748a",
  1396 => x"2e81e238",
  1397 => x"84140870",
  1398 => x"892a7081",
  1399 => x"06515153",
  1400 => x"72f23874",
  1401 => x"740c7533",
  1402 => x"5574e038",
  1403 => x"bbcc0bbb",
  1404 => x"cc335456",
  1405 => x"72802ea4",
  1406 => x"38725581",
  1407 => x"1656748a",
  1408 => x"2e81d738",
  1409 => x"84140870",
  1410 => x"892a7081",
  1411 => x"06515153",
  1412 => x"72f23874",
  1413 => x"740c7533",
  1414 => x"5574e038",
  1415 => x"76802e82",
  1416 => x"d938bbe4",
  1417 => x"0bbbe433",
  1418 => x"54567280",
  1419 => x"2ea23872",
  1420 => x"55811656",
  1421 => x"748a2e81",
  1422 => x"c6388414",
  1423 => x"0870892a",
  1424 => x"81065153",
  1425 => x"72f43874",
  1426 => x"740c7533",
  1427 => x"5574e238",
  1428 => x"bbf40bbb",
  1429 => x"f4335456",
  1430 => x"72802ea2",
  1431 => x"38725581",
  1432 => x"1656748a",
  1433 => x"2e81b938",
  1434 => x"84140870",
  1435 => x"892a8106",
  1436 => x"515372f4",
  1437 => x"3874740c",
  1438 => x"75335574",
  1439 => x"e238e490",
  1440 => x"3fbcdc08",
  1441 => x"5680d50b",
  1442 => x"84170cbc",
  1443 => x"e4085484",
  1444 => x"14088106",
  1445 => x"5574802e",
  1446 => x"f6387308",
  1447 => x"7081ff06",
  1448 => x"f6115256",
  1449 => x"5372ae26",
  1450 => x"81973872",
  1451 => x"1010b8d8",
  1452 => x"05577608",
  1453 => x"04841408",
  1454 => x"70892a70",
  1455 => x"81065151",
  1456 => x"5372f238",
  1457 => x"8d740c84",
  1458 => x"14087089",
  1459 => x"2a708106",
  1460 => x"51515372",
  1461 => x"fdfe38fe",
  1462 => x"8a398414",
  1463 => x"0870892a",
  1464 => x"70810651",
  1465 => x"515372f2",
  1466 => x"388d740c",
  1467 => x"84140870",
  1468 => x"892a7081",
  1469 => x"06515153",
  1470 => x"72fe8938",
  1471 => x"fe953984",
  1472 => x"14087089",
  1473 => x"2a810651",
  1474 => x"5776f438",
  1475 => x"8d740c84",
  1476 => x"14087089",
  1477 => x"2a810651",
  1478 => x"5372fe9e",
  1479 => x"38fea839",
  1480 => x"84140870",
  1481 => x"892a8106",
  1482 => x"515776f4",
  1483 => x"388d740c",
  1484 => x"84140870",
  1485 => x"892a8106",
  1486 => x"515372fe",
  1487 => x"ab38feb5",
  1488 => x"39841408",
  1489 => x"70892a81",
  1490 => x"06515372",
  1491 => x"f438ab74",
  1492 => x"0c748a2e",
  1493 => x"80ff3884",
  1494 => x"14087089",
  1495 => x"2a810651",
  1496 => x"5372f438",
  1497 => x"74740c84",
  1498 => x"14087089",
  1499 => x"2a810656",
  1500 => x"5374f438",
  1501 => x"ad740cfe",
  1502 => x"9639bc98",
  1503 => x"0bbc9833",
  1504 => x"54567280",
  1505 => x"2efdc938",
  1506 => x"72811757",
  1507 => x"55748a2e",
  1508 => x"a5388414",
  1509 => x"0870892a",
  1510 => x"81065153",
  1511 => x"72f43874",
  1512 => x"740c7533",
  1513 => x"5574802e",
  1514 => x"fda63881",
  1515 => x"1656748a",
  1516 => x"2e098106",
  1517 => x"dd388414",
  1518 => x"0870892a",
  1519 => x"81065157",
  1520 => x"76f4388d",
  1521 => x"740c8414",
  1522 => x"0870892a",
  1523 => x"81065153",
  1524 => x"72c038cb",
  1525 => x"39841408",
  1526 => x"70892a81",
  1527 => x"06515776",
  1528 => x"f4388d74",
  1529 => x"0c841408",
  1530 => x"70892a81",
  1531 => x"06515372",
  1532 => x"fee538fe",
  1533 => x"ef3981ff",
  1534 => x"0b84170c",
  1535 => x"fd913980",
  1536 => x"ff0b8417",
  1537 => x"0cfd8839",
  1538 => x"bf0b8417",
  1539 => x"0cfd8039",
  1540 => x"9f0b8417",
  1541 => x"0cfcf839",
  1542 => x"8f0b8417",
  1543 => x"0cfcf039",
  1544 => x"870b8417",
  1545 => x"0cfce839",
  1546 => x"830b8417",
  1547 => x"0cfce039",
  1548 => x"810b8417",
  1549 => x"0cfcd839",
  1550 => x"800b8417",
  1551 => x"0cfcd039",
  1552 => x"8c08028c",
  1553 => x"0cfd3d0d",
  1554 => x"80538c08",
  1555 => x"8c050852",
  1556 => x"8c088805",
  1557 => x"085182de",
  1558 => x"3f800870",
  1559 => x"800c5485",
  1560 => x"3d0d8c0c",
  1561 => x"048c0802",
  1562 => x"8c0cfd3d",
  1563 => x"0d81538c",
  1564 => x"088c0508",
  1565 => x"528c0888",
  1566 => x"05085182",
  1567 => x"b93f8008",
  1568 => x"70800c54",
  1569 => x"853d0d8c",
  1570 => x"0c048c08",
  1571 => x"028c0cf9",
  1572 => x"3d0d800b",
  1573 => x"8c08fc05",
  1574 => x"0c8c0888",
  1575 => x"05088025",
  1576 => x"ab388c08",
  1577 => x"88050830",
  1578 => x"8c088805",
  1579 => x"0c800b8c",
  1580 => x"08f4050c",
  1581 => x"8c08fc05",
  1582 => x"08883881",
  1583 => x"0b8c08f4",
  1584 => x"050c8c08",
  1585 => x"f405088c",
  1586 => x"08fc050c",
  1587 => x"8c088c05",
  1588 => x"088025ab",
  1589 => x"388c088c",
  1590 => x"0508308c",
  1591 => x"088c050c",
  1592 => x"800b8c08",
  1593 => x"f0050c8c",
  1594 => x"08fc0508",
  1595 => x"8838810b",
  1596 => x"8c08f005",
  1597 => x"0c8c08f0",
  1598 => x"05088c08",
  1599 => x"fc050c80",
  1600 => x"538c088c",
  1601 => x"0508528c",
  1602 => x"08880508",
  1603 => x"5181a73f",
  1604 => x"8008708c",
  1605 => x"08f8050c",
  1606 => x"548c08fc",
  1607 => x"0508802e",
  1608 => x"8c388c08",
  1609 => x"f8050830",
  1610 => x"8c08f805",
  1611 => x"0c8c08f8",
  1612 => x"05087080",
  1613 => x"0c54893d",
  1614 => x"0d8c0c04",
  1615 => x"8c08028c",
  1616 => x"0cfb3d0d",
  1617 => x"800b8c08",
  1618 => x"fc050c8c",
  1619 => x"08880508",
  1620 => x"80259338",
  1621 => x"8c088805",
  1622 => x"08308c08",
  1623 => x"88050c81",
  1624 => x"0b8c08fc",
  1625 => x"050c8c08",
  1626 => x"8c050880",
  1627 => x"258c388c",
  1628 => x"088c0508",
  1629 => x"308c088c",
  1630 => x"050c8153",
  1631 => x"8c088c05",
  1632 => x"08528c08",
  1633 => x"88050851",
  1634 => x"ad3f8008",
  1635 => x"708c08f8",
  1636 => x"050c548c",
  1637 => x"08fc0508",
  1638 => x"802e8c38",
  1639 => x"8c08f805",
  1640 => x"08308c08",
  1641 => x"f8050c8c",
  1642 => x"08f80508",
  1643 => x"70800c54",
  1644 => x"873d0d8c",
  1645 => x"0c048c08",
  1646 => x"028c0cfd",
  1647 => x"3d0d810b",
  1648 => x"8c08fc05",
  1649 => x"0c800b8c",
  1650 => x"08f8050c",
  1651 => x"8c088c05",
  1652 => x"088c0888",
  1653 => x"050827ac",
  1654 => x"388c08fc",
  1655 => x"0508802e",
  1656 => x"a338800b",
  1657 => x"8c088c05",
  1658 => x"08249938",
  1659 => x"8c088c05",
  1660 => x"08108c08",
  1661 => x"8c050c8c",
  1662 => x"08fc0508",
  1663 => x"108c08fc",
  1664 => x"050cc939",
  1665 => x"8c08fc05",
  1666 => x"08802e80",
  1667 => x"c9388c08",
  1668 => x"8c05088c",
  1669 => x"08880508",
  1670 => x"26a1388c",
  1671 => x"08880508",
  1672 => x"8c088c05",
  1673 => x"08318c08",
  1674 => x"88050c8c",
  1675 => x"08f80508",
  1676 => x"8c08fc05",
  1677 => x"08078c08",
  1678 => x"f8050c8c",
  1679 => x"08fc0508",
  1680 => x"812a8c08",
  1681 => x"fc050c8c",
  1682 => x"088c0508",
  1683 => x"812a8c08",
  1684 => x"8c050cff",
  1685 => x"af398c08",
  1686 => x"90050880",
  1687 => x"2e8f388c",
  1688 => x"08880508",
  1689 => x"708c08f4",
  1690 => x"050c518d",
  1691 => x"398c08f8",
  1692 => x"0508708c",
  1693 => x"08f4050c",
  1694 => x"518c08f4",
  1695 => x"0508800c",
  1696 => x"853d0d8c",
  1697 => x"0c04fd3d",
  1698 => x"0d800bbc",
  1699 => x"cc085454",
  1700 => x"72812e99",
  1701 => x"387380c4",
  1702 => x"900cd3c3",
  1703 => x"3fd2e13f",
  1704 => x"bce85281",
  1705 => x"51f5f13f",
  1706 => x"8008519f",
  1707 => x"3f7280c4",
  1708 => x"900cd3ab",
  1709 => x"3fd2c93f",
  1710 => x"bce85281",
  1711 => x"51f5d93f",
  1712 => x"80085187",
  1713 => x"3f00ff39",
  1714 => x"00ff39f7",
  1715 => x"3d0d7bbc",
  1716 => x"ec0882c8",
  1717 => x"11085a54",
  1718 => x"5a77802e",
  1719 => x"80d93881",
  1720 => x"88188419",
  1721 => x"08ff0581",
  1722 => x"712b5955",
  1723 => x"59807424",
  1724 => x"80e93880",
  1725 => x"7424b538",
  1726 => x"73822b78",
  1727 => x"11880556",
  1728 => x"56818019",
  1729 => x"08770653",
  1730 => x"72802eb5",
  1731 => x"38781670",
  1732 => x"08535379",
  1733 => x"51740853",
  1734 => x"722dff14",
  1735 => x"fc17fc17",
  1736 => x"79812c5a",
  1737 => x"57575473",
  1738 => x"8025d638",
  1739 => x"77085877",
  1740 => x"ffad38bc",
  1741 => x"ec0853bc",
  1742 => x"1308a538",
  1743 => x"7951ff85",
  1744 => x"3f740853",
  1745 => x"722dff14",
  1746 => x"fc17fc17",
  1747 => x"79812c5a",
  1748 => x"57575473",
  1749 => x"8025ffa9",
  1750 => x"38d23980",
  1751 => x"57ff9439",
  1752 => x"7251bc13",
  1753 => x"0853722d",
  1754 => x"7951fed9",
  1755 => x"3fff3d0d",
  1756 => x"80c3f00b",
  1757 => x"fc057008",
  1758 => x"525270ff",
  1759 => x"2e913870",
  1760 => x"2dfc1270",
  1761 => x"08525270",
  1762 => x"ff2e0981",
  1763 => x"06f13883",
  1764 => x"3d0d0404",
  1765 => x"d2b43f04",
  1766 => x"00000040",
  1767 => x"0000079a",
  1768 => x"000007bf",
  1769 => x"000007bf",
  1770 => x"0000079a",
  1771 => x"000007bf",
  1772 => x"000007bf",
  1773 => x"000007bf",
  1774 => x"000007bf",
  1775 => x"000007bf",
  1776 => x"000007bf",
  1777 => x"000007bf",
  1778 => x"000007bf",
  1779 => x"000007bf",
  1780 => x"000007bf",
  1781 => x"000007bf",
  1782 => x"000007bf",
  1783 => x"000007bf",
  1784 => x"000007bf",
  1785 => x"000007bf",
  1786 => x"000007bf",
  1787 => x"000007bf",
  1788 => x"000007bf",
  1789 => x"000007bf",
  1790 => x"000007bf",
  1791 => x"000007bf",
  1792 => x"000007bf",
  1793 => x"000007bf",
  1794 => x"000007bf",
  1795 => x"000007bf",
  1796 => x"000007bf",
  1797 => x"000007bf",
  1798 => x"000007bf",
  1799 => x"000007bf",
  1800 => x"000007bf",
  1801 => x"000007bf",
  1802 => x"000007bf",
  1803 => x"000007bf",
  1804 => x"000007bf",
  1805 => x"00000861",
  1806 => x"00000859",
  1807 => x"00000851",
  1808 => x"00000849",
  1809 => x"00000841",
  1810 => x"00000839",
  1811 => x"00000831",
  1812 => x"00000828",
  1813 => x"0000081f",
  1814 => x"0000168f",
  1815 => x"00001741",
  1816 => x"00001741",
  1817 => x"0000168f",
  1818 => x"00001741",
  1819 => x"00001741",
  1820 => x"00001741",
  1821 => x"00001741",
  1822 => x"00001741",
  1823 => x"00001741",
  1824 => x"00001741",
  1825 => x"00001741",
  1826 => x"00001741",
  1827 => x"00001741",
  1828 => x"00001741",
  1829 => x"00001741",
  1830 => x"00001741",
  1831 => x"00001741",
  1832 => x"00001741",
  1833 => x"00001741",
  1834 => x"00001741",
  1835 => x"00001741",
  1836 => x"00001741",
  1837 => x"00001741",
  1838 => x"00001741",
  1839 => x"00001741",
  1840 => x"00001741",
  1841 => x"00001741",
  1842 => x"00001741",
  1843 => x"00001741",
  1844 => x"00001741",
  1845 => x"00001741",
  1846 => x"00001741",
  1847 => x"00001741",
  1848 => x"00001741",
  1849 => x"00001741",
  1850 => x"00001741",
  1851 => x"00001741",
  1852 => x"00001838",
  1853 => x"00001830",
  1854 => x"00001828",
  1855 => x"00001820",
  1856 => x"00001818",
  1857 => x"00001810",
  1858 => x"00001808",
  1859 => x"000017ff",
  1860 => x"000017f6",
  1861 => x"0a677265",
  1862 => x"74682072",
  1863 => x"65676973",
  1864 => x"74657273",
  1865 => x"3a000000",
  1866 => x"0a636f6e",
  1867 => x"74726f6c",
  1868 => x"3a202020",
  1869 => x"20202000",
  1870 => x"0a737461",
  1871 => x"7475733a",
  1872 => x"20202020",
  1873 => x"20202000",
  1874 => x"0a6d6163",
  1875 => x"5f6d7362",
  1876 => x"3a202020",
  1877 => x"20202000",
  1878 => x"0a6d6163",
  1879 => x"5f6c7362",
  1880 => x"3a202020",
  1881 => x"20202000",
  1882 => x"0a6d6469",
  1883 => x"6f5f636f",
  1884 => x"6e74726f",
  1885 => x"6c3a2000",
  1886 => x"0a74785f",
  1887 => x"706f696e",
  1888 => x"7465723a",
  1889 => x"20202000",
  1890 => x"0a72785f",
  1891 => x"706f696e",
  1892 => x"7465723a",
  1893 => x"20202000",
  1894 => x"0a656463",
  1895 => x"6c5f6970",
  1896 => x"3a202020",
  1897 => x"20202000",
  1898 => x"0a686173",
  1899 => x"685f6d73",
  1900 => x"623a2020",
  1901 => x"20202000",
  1902 => x"0a686173",
  1903 => x"685f6c73",
  1904 => x"623a2020",
  1905 => x"20202000",
  1906 => x"0a0a0000",
  1907 => x"536f432c",
  1908 => x"205a5055",
  1909 => x"20746573",
  1910 => x"74207072",
  1911 => x"6f677261",
  1912 => x"6d200000",
  1913 => x"286f6e20",
  1914 => x"73696d75",
  1915 => x"6c61746f",
  1916 => x"72290a00",
  1917 => x"636f6d70",
  1918 => x"696c6564",
  1919 => x"3a204175",
  1920 => x"67202035",
  1921 => x"20323031",
  1922 => x"30202020",
  1923 => x"31383a30",
  1924 => x"323a3437",
  1925 => x"0a000000",
  1926 => x"286f6e20",
  1927 => x"68617264",
  1928 => x"77617265",
  1929 => x"290a0000",
  1930 => x"64756d6d",
  1931 => x"792e6578",
  1932 => x"65000000",
  1933 => x"43000000",
  1934 => x"00ffffff",
  1935 => x"ff00ffff",
  1936 => x"ffff00ff",
  1937 => x"ffffff00",
  1938 => x"00000000",
  1939 => x"00000000",
  1940 => x"00000000",
  1941 => x"000021f8",
  1942 => x"80000c00",
  1943 => x"80000800",
  1944 => x"80000200",
  1945 => x"80000100",
  1946 => x"00001e28",
  1947 => x"00001e70",
  1948 => x"00000000",
  1949 => x"000020d8",
  1950 => x"00002134",
  1951 => x"00002190",
  1952 => x"00000000",
  1953 => x"00000000",
  1954 => x"00000000",
  1955 => x"00000000",
  1956 => x"00000000",
  1957 => x"00000000",
  1958 => x"00000000",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00001e34",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00000000",
  1984 => x"00000000",
  1985 => x"00000000",
  1986 => x"00000000",
  1987 => x"00000000",
  1988 => x"00000000",
  1989 => x"00000000",
  1990 => x"00000001",
  1991 => x"330eabcd",
  1992 => x"1234e66d",
  1993 => x"deec0005",
  1994 => x"000b0000",
  1995 => x"00000000",
  1996 => x"00000000",
  1997 => x"00000000",
  1998 => x"00000000",
  1999 => x"00000000",
  2000 => x"00000000",
  2001 => x"00000000",
  2002 => x"00000000",
  2003 => x"00000000",
  2004 => x"00000000",
  2005 => x"00000000",
  2006 => x"00000000",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00000000",
  2010 => x"00000000",
  2011 => x"00000000",
  2012 => x"00000000",
  2013 => x"00000000",
  2014 => x"00000000",
  2015 => x"00000000",
  2016 => x"00000000",
  2017 => x"00000000",
  2018 => x"00000000",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00000000",
  2026 => x"00000000",
  2027 => x"00000000",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000000",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"00000000",
  2049 => x"00000000",
  2050 => x"00000000",
  2051 => x"00000000",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"ffffffff",
  2172 => x"00000000",
  2173 => x"ffffffff",
  2174 => x"00000000",
  2175 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
