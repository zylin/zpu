-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


--type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);
type ram_type is array(natural range 0 to bram_words-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80db8c0c",
     3 => x"3a0b0b80",
     4 => x"d2d00400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"90040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80da",
   162 => x"f8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f8040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"e0040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80db880c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82d33f80",
   257 => x"ccbe3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80088408",
   281 => x"88087575",
   282 => x"b2cb2d50",
   283 => x"50800856",
   284 => x"880c840c",
   285 => x"800c5104",
   286 => x"80088408",
   287 => x"88087575",
   288 => x"b1992d50",
   289 => x"50800856",
   290 => x"880c840c",
   291 => x"800c5104",
   292 => x"80088408",
   293 => x"880880d3",
   294 => x"9d2d880c",
   295 => x"840c800c",
   296 => x"0480db88",
   297 => x"08802ea9",
   298 => x"3880db8c",
   299 => x"08822e80",
   300 => x"c5388380",
   301 => x"800b8180",
   302 => x"8080800c",
   303 => x"82a0800b",
   304 => x"81808080",
   305 => x"840c8290",
   306 => x"800b8180",
   307 => x"8080880c",
   308 => x"04f88080",
   309 => x"80a40b81",
   310 => x"80808080",
   311 => x"0cf88080",
   312 => x"82800b81",
   313 => x"80808084",
   314 => x"0cf88080",
   315 => x"84800b81",
   316 => x"80808088",
   317 => x"0c0480c0",
   318 => x"a8808c0b",
   319 => x"81808080",
   320 => x"800c80c0",
   321 => x"a880940b",
   322 => x"81808080",
   323 => x"840c0b0b",
   324 => x"80d4f00b",
   325 => x"81808080",
   326 => x"880c04ff",
   327 => x"3d0d8180",
   328 => x"80808c33",
   329 => x"5170a938",
   330 => x"80db9408",
   331 => x"70085252",
   332 => x"70802e94",
   333 => x"38841280",
   334 => x"db940c70",
   335 => x"2d80db94",
   336 => x"08700852",
   337 => x"5270ee38",
   338 => x"810b8180",
   339 => x"80808c34",
   340 => x"833d0d04",
   341 => x"04803d0d",
   342 => x"0b0b80eb",
   343 => x"8808802e",
   344 => x"8e380b0b",
   345 => x"0b0b800b",
   346 => x"802e0981",
   347 => x"06853882",
   348 => x"3d0d040b",
   349 => x"0b80eb88",
   350 => x"510b0b0b",
   351 => x"f5823f82",
   352 => x"3d0d0404",
   353 => x"fd3d0d80",
   354 => x"dba00888",
   355 => x"110883de",
   356 => x"80078812",
   357 => x"0c841108",
   358 => x"fca1ff06",
   359 => x"84120c53",
   360 => x"8f51a2b4",
   361 => x"3f80dba0",
   362 => x"08841108",
   363 => x"e1ff0684",
   364 => x"120c8411",
   365 => x"08868007",
   366 => x"84120c84",
   367 => x"110880c0",
   368 => x"80078412",
   369 => x"0c538151",
   370 => x"a1e93f80",
   371 => x"dba00884",
   372 => x"1108ffbf",
   373 => x"ff068412",
   374 => x"0c538551",
   375 => x"a1fa3f80",
   376 => x"dba00884",
   377 => x"110880c0",
   378 => x"80078412",
   379 => x"0c538151",
   380 => x"a1c13f80",
   381 => x"dba00884",
   382 => x"1108ffbf",
   383 => x"ff068412",
   384 => x"0c538151",
   385 => x"a1d23f80",
   386 => x"dba00884",
   387 => x"110880c0",
   388 => x"80078412",
   389 => x"0c538151",
   390 => x"a1993f80",
   391 => x"dba00884",
   392 => x"1108ffbf",
   393 => x"ff068412",
   394 => x"0c538151",
   395 => x"a1aa3f80",
   396 => x"dba00884",
   397 => x"1108e1ff",
   398 => x"0684120c",
   399 => x"5384800b",
   400 => x"84140870",
   401 => x"72078416",
   402 => x"0c538414",
   403 => x"087080c0",
   404 => x"80078416",
   405 => x"0c535481",
   406 => x"51a0d83f",
   407 => x"80dba008",
   408 => x"84110870",
   409 => x"ffbfff06",
   410 => x"84130c53",
   411 => x"538551a0",
   412 => x"e73f80db",
   413 => x"a0088411",
   414 => x"0870feff",
   415 => x"ff068413",
   416 => x"0c538411",
   417 => x"0870e1ff",
   418 => x"0684130c",
   419 => x"53841108",
   420 => x"70760784",
   421 => x"130c5384",
   422 => x"110880c0",
   423 => x"80078412",
   424 => x"0c538151",
   425 => x"a08d3f80",
   426 => x"dba00884",
   427 => x"1108ffbf",
   428 => x"ff068412",
   429 => x"0c841108",
   430 => x"e1ff0684",
   431 => x"120c8411",
   432 => x"08908007",
   433 => x"84120c84",
   434 => x"110880c0",
   435 => x"80078412",
   436 => x"0c548151",
   437 => x"9fdd3f80",
   438 => x"dba00884",
   439 => x"1108ffbf",
   440 => x"ff068412",
   441 => x"0c54aa51",
   442 => x"9fc93f80",
   443 => x"dba00884",
   444 => x"1108feff",
   445 => x"ff068412",
   446 => x"0c841108",
   447 => x"e1ff0684",
   448 => x"120c8411",
   449 => x"0884120c",
   450 => x"84110880",
   451 => x"c0800784",
   452 => x"120c5481",
   453 => x"519f9c3f",
   454 => x"80dba008",
   455 => x"841108ff",
   456 => x"bfff0684",
   457 => x"120c8411",
   458 => x"08e1ff06",
   459 => x"84120c84",
   460 => x"11089880",
   461 => x"0784120c",
   462 => x"84110880",
   463 => x"c0800784",
   464 => x"120c5481",
   465 => x"519eec3f",
   466 => x"80dba008",
   467 => x"841108ff",
   468 => x"bfff0684",
   469 => x"120c54aa",
   470 => x"519ed83f",
   471 => x"80dba008",
   472 => x"841108fe",
   473 => x"ffff0684",
   474 => x"120c8411",
   475 => x"08e1ff06",
   476 => x"84120c84",
   477 => x"11088412",
   478 => x"0c841108",
   479 => x"80c08007",
   480 => x"84120c54",
   481 => x"81519eab",
   482 => x"3f80dba0",
   483 => x"08841108",
   484 => x"ffbfff06",
   485 => x"84120c84",
   486 => x"1108e1ff",
   487 => x"0684120c",
   488 => x"8411088c",
   489 => x"80078412",
   490 => x"0c841108",
   491 => x"80c08007",
   492 => x"84120c54",
   493 => x"81519dfb",
   494 => x"3f80dba0",
   495 => x"08841108",
   496 => x"ffbfff06",
   497 => x"84120c54",
   498 => x"aa519de7",
   499 => x"3f810b80",
   500 => x"dba00884",
   501 => x"110870fe",
   502 => x"ffff0684",
   503 => x"130c5484",
   504 => x"110870e1",
   505 => x"ff068413",
   506 => x"0c548411",
   507 => x"0884120c",
   508 => x"84110870",
   509 => x"80c08007",
   510 => x"84130c54",
   511 => x"54705254",
   512 => x"9db13f80",
   513 => x"dba00884",
   514 => x"110870ff",
   515 => x"bfff0684",
   516 => x"130c5384",
   517 => x"110870e1",
   518 => x"ff068413",
   519 => x"0c538411",
   520 => x"08708280",
   521 => x"0784130c",
   522 => x"53841108",
   523 => x"7080c080",
   524 => x"0784130c",
   525 => x"53537351",
   526 => x"9cf93f80",
   527 => x"dba00884",
   528 => x"1108ffbf",
   529 => x"ff068412",
   530 => x"0c53aa51",
   531 => x"9ce53f82",
   532 => x"519d853f",
   533 => x"853d0d04",
   534 => x"fc3d0d02",
   535 => x"9b053302",
   536 => x"84059f05",
   537 => x"33545272",
   538 => x"822e81ad",
   539 => x"38827325",
   540 => x"91387283",
   541 => x"2e83bc38",
   542 => x"72842e82",
   543 => x"a938863d",
   544 => x"0d047281",
   545 => x"2e098106",
   546 => x"f538ff80",
   547 => x"127081ff",
   548 => x"0680dba0",
   549 => x"08841108",
   550 => x"feffff06",
   551 => x"84120c84",
   552 => x"1108e1ff",
   553 => x"0684120c",
   554 => x"71842b9e",
   555 => x"80068412",
   556 => x"08707207",
   557 => x"84140c54",
   558 => x"84120880",
   559 => x"c0800784",
   560 => x"130c5755",
   561 => x"56528151",
   562 => x"9be93f80",
   563 => x"dba00884",
   564 => x"1108ffbf",
   565 => x"ff068412",
   566 => x"0c841108",
   567 => x"e1ff0684",
   568 => x"120c7588",
   569 => x"2b9e8006",
   570 => x"84120871",
   571 => x"0784130c",
   572 => x"84120880",
   573 => x"c0800784",
   574 => x"130c5553",
   575 => x"81519bb3",
   576 => x"3f80dba0",
   577 => x"08841108",
   578 => x"ffbfff06",
   579 => x"84120c53",
   580 => x"aa519b9f",
   581 => x"3f863d0d",
   582 => x"04c01270",
   583 => x"81ff0680",
   584 => x"dba00884",
   585 => x"1108feff",
   586 => x"ff068412",
   587 => x"0c841108",
   588 => x"e1ff0684",
   589 => x"120c7184",
   590 => x"2b9e8006",
   591 => x"84120870",
   592 => x"72078414",
   593 => x"0c548412",
   594 => x"0880c080",
   595 => x"0784130c",
   596 => x"57555652",
   597 => x"81519adb",
   598 => x"3f80dba0",
   599 => x"08841108",
   600 => x"ffbfff06",
   601 => x"84120c84",
   602 => x"1108e1ff",
   603 => x"0684120c",
   604 => x"75882b9e",
   605 => x"80068412",
   606 => x"08710784",
   607 => x"130c8412",
   608 => x"0880c080",
   609 => x"0784130c",
   610 => x"55538151",
   611 => x"9aa53f80",
   612 => x"dba00884",
   613 => x"1108ffbf",
   614 => x"ff068412",
   615 => x"0c53aa51",
   616 => x"9a913ffe",
   617 => x"f039d012",
   618 => x"7081ff06",
   619 => x"80dba008",
   620 => x"841108fe",
   621 => x"ffff0684",
   622 => x"120c8411",
   623 => x"08e1ff06",
   624 => x"84120c71",
   625 => x"842b9e80",
   626 => x"06841208",
   627 => x"70720784",
   628 => x"140c5484",
   629 => x"120880c0",
   630 => x"80078413",
   631 => x"0c575556",
   632 => x"52815199",
   633 => x"ce3f80db",
   634 => x"a0088411",
   635 => x"08ffbfff",
   636 => x"0684120c",
   637 => x"841108e1",
   638 => x"ff068412",
   639 => x"0c75882b",
   640 => x"9e800684",
   641 => x"12087107",
   642 => x"84130c84",
   643 => x"120880c0",
   644 => x"80078413",
   645 => x"0c555381",
   646 => x"5199983f",
   647 => x"80dba008",
   648 => x"841108ff",
   649 => x"bfff0684",
   650 => x"120c53aa",
   651 => x"5199843f",
   652 => x"fde339ff",
   653 => x"90127081",
   654 => x"ff0680db",
   655 => x"a0088411",
   656 => x"08feffff",
   657 => x"0684120c",
   658 => x"841108e1",
   659 => x"ff068412",
   660 => x"0c71842b",
   661 => x"9e800684",
   662 => x"12087072",
   663 => x"0784140c",
   664 => x"54841208",
   665 => x"80c08007",
   666 => x"84130c57",
   667 => x"55565281",
   668 => x"5198c03f",
   669 => x"80dba008",
   670 => x"841108ff",
   671 => x"bfff0684",
   672 => x"120c8411",
   673 => x"08e1ff06",
   674 => x"84120c75",
   675 => x"882b9e80",
   676 => x"06841208",
   677 => x"71078413",
   678 => x"0c841208",
   679 => x"80c08007",
   680 => x"84130c55",
   681 => x"53815198",
   682 => x"8a3f80db",
   683 => x"a0088411",
   684 => x"08ffbfff",
   685 => x"0684120c",
   686 => x"53aa5197",
   687 => x"f63ffcd5",
   688 => x"39fb3d0d",
   689 => x"77703353",
   690 => x"5671802e",
   691 => x"818f3871",
   692 => x"55811680",
   693 => x"dba00884",
   694 => x"11088180",
   695 => x"80078412",
   696 => x"0c841108",
   697 => x"e1ff0684",
   698 => x"120c7684",
   699 => x"2b9e8006",
   700 => x"84120870",
   701 => x"72078414",
   702 => x"0c558412",
   703 => x"0880c080",
   704 => x"0784130c",
   705 => x"56545681",
   706 => x"5197a83f",
   707 => x"80dba008",
   708 => x"841108ff",
   709 => x"bfff0684",
   710 => x"120c8411",
   711 => x"08e1ff06",
   712 => x"84120c75",
   713 => x"882b9e80",
   714 => x"06841208",
   715 => x"71078413",
   716 => x"0c841208",
   717 => x"80c08007",
   718 => x"84130c55",
   719 => x"53815196",
   720 => x"f23f80db",
   721 => x"a0088411",
   722 => x"08ffbfff",
   723 => x"0684120c",
   724 => x"53ae5196",
   725 => x"de3f7533",
   726 => x"5574fef5",
   727 => x"38873d0d",
   728 => x"04ff3d0d",
   729 => x"028f0533",
   730 => x"70525297",
   731 => x"d93f7151",
   732 => x"98cc3f71",
   733 => x"800c833d",
   734 => x"0d04fa3d",
   735 => x"0d02a305",
   736 => x"3356758d",
   737 => x"2e818238",
   738 => x"75883270",
   739 => x"307780ff",
   740 => x"32703072",
   741 => x"80257180",
   742 => x"25075451",
   743 => x"56585574",
   744 => x"97389f76",
   745 => x"278e3881",
   746 => x"808087c8",
   747 => x"335580ce",
   748 => x"7527b438",
   749 => x"883d0d04",
   750 => x"81808087",
   751 => x"c8335675",
   752 => x"802ef138",
   753 => x"885193ec",
   754 => x"3fa05193",
   755 => x"e73f8851",
   756 => x"93e23f81",
   757 => x"808087c8",
   758 => x"33ff0557",
   759 => x"76818080",
   760 => x"87c83488",
   761 => x"3d0d0475",
   762 => x"5193c93f",
   763 => x"81808087",
   764 => x"c8338111",
   765 => x"55577381",
   766 => x"808087c8",
   767 => x"34758180",
   768 => x"8086f418",
   769 => x"34883d0d",
   770 => x"048a5193",
   771 => x"a73f8180",
   772 => x"8087c833",
   773 => x"81115654",
   774 => x"74818080",
   775 => x"87c83480",
   776 => x"0b818080",
   777 => x"86f41534",
   778 => x"8056800b",
   779 => x"81808086",
   780 => x"f4173356",
   781 => x"5474a02e",
   782 => x"83388154",
   783 => x"74802e90",
   784 => x"3873802e",
   785 => x"8b388116",
   786 => x"7081ff06",
   787 => x"5757db39",
   788 => x"75802e80",
   789 => x"c538800b",
   790 => x"81808087",
   791 => x"c4335555",
   792 => x"747427af",
   793 => x"38735774",
   794 => x"10101075",
   795 => x"10057654",
   796 => x"81808086",
   797 => x"f4538180",
   798 => x"80809405",
   799 => x"51a1e83f",
   800 => x"8008802e",
   801 => x"a8388115",
   802 => x"7081ff06",
   803 => x"56547675",
   804 => x"26d53880",
   805 => x"d4f85192",
   806 => x"b73f80d4",
   807 => x"f45192b0",
   808 => x"3f800b81",
   809 => x"808087c8",
   810 => x"34883d0d",
   811 => x"04741010",
   812 => x"81808086",
   813 => x"b4057008",
   814 => x"81808087",
   815 => x"cc0c5680",
   816 => x"0b818080",
   817 => x"87c834e1",
   818 => x"39fc3d0d",
   819 => x"8a5191e4",
   820 => x"3f800b81",
   821 => x"808087c8",
   822 => x"34800b81",
   823 => x"808087c4",
   824 => x"34800b81",
   825 => x"808087cc",
   826 => x"0c80d58c",
   827 => x"52818080",
   828 => x"8094519f",
   829 => x"a63f80d5",
   830 => x"90528180",
   831 => x"8087c433",
   832 => x"70101011",
   833 => x"70101010",
   834 => x"81808081",
   835 => x"b4055356",
   836 => x"549f883f",
   837 => x"81808087",
   838 => x"c4337010",
   839 => x"10818080",
   840 => x"86b405a0",
   841 => x"f8710c54",
   842 => x"81115155",
   843 => x"74818080",
   844 => x"87c43480",
   845 => x"d5b85274",
   846 => x"81ff0670",
   847 => x"8a298180",
   848 => x"80809405",
   849 => x"52539ed3",
   850 => x"3f80d5c0",
   851 => x"52818080",
   852 => x"87c43370",
   853 => x"10101170",
   854 => x"10101081",
   855 => x"808081b4",
   856 => x"05535555",
   857 => x"9eb53f81",
   858 => x"808087c4",
   859 => x"33701010",
   860 => x"81808086",
   861 => x"b405a0dd",
   862 => x"710c5481",
   863 => x"11515473",
   864 => x"81808087",
   865 => x"c43480d5",
   866 => x"dc527381",
   867 => x"ff06708a",
   868 => x"29818080",
   869 => x"80940552",
   870 => x"539e803f",
   871 => x"80d5e052",
   872 => x"81808087",
   873 => x"c4337010",
   874 => x"10117010",
   875 => x"10108180",
   876 => x"8081b405",
   877 => x"5356549d",
   878 => x"e23f8180",
   879 => x"8087c433",
   880 => x"70101081",
   881 => x"808086b4",
   882 => x"05a8ac71",
   883 => x"0c548111",
   884 => x"51557481",
   885 => x"808087c4",
   886 => x"3480d680",
   887 => x"527481ff",
   888 => x"06708a29",
   889 => x"81808080",
   890 => x"94055253",
   891 => x"9dad3f80",
   892 => x"d6885281",
   893 => x"808087c4",
   894 => x"33701010",
   895 => x"11701010",
   896 => x"10818080",
   897 => x"81b40553",
   898 => x"55559d8f",
   899 => x"3f818080",
   900 => x"87c43370",
   901 => x"10108180",
   902 => x"8086b405",
   903 => x"a8df710c",
   904 => x"54811151",
   905 => x"54738180",
   906 => x"8087c434",
   907 => x"80d69c52",
   908 => x"7381ff06",
   909 => x"708a2981",
   910 => x"80808094",
   911 => x"0552539c",
   912 => x"da3f80d6",
   913 => x"a4528180",
   914 => x"8087c433",
   915 => x"70101011",
   916 => x"70101010",
   917 => x"81808081",
   918 => x"b4055356",
   919 => x"549cbc3f",
   920 => x"81808087",
   921 => x"c4337010",
   922 => x"10818080",
   923 => x"86b4059f",
   924 => x"cd710c54",
   925 => x"81115155",
   926 => x"74818080",
   927 => x"87c43480",
   928 => x"d6b45274",
   929 => x"81ff0670",
   930 => x"8a298180",
   931 => x"80809405",
   932 => x"52539c87",
   933 => x"3f80d6ec",
   934 => x"52818080",
   935 => x"87c43370",
   936 => x"10101170",
   937 => x"10101081",
   938 => x"808081b4",
   939 => x"05535555",
   940 => x"9be93f81",
   941 => x"808087c4",
   942 => x"33701010",
   943 => x"81808086",
   944 => x"b4059eab",
   945 => x"710c5481",
   946 => x"05537281",
   947 => x"808087c4",
   948 => x"3480d4f4",
   949 => x"518df93f",
   950 => x"810b8180",
   951 => x"8087d034",
   952 => x"90af3f80",
   953 => x"08b63881",
   954 => x"808087cc",
   955 => x"0853728f",
   956 => x"38818080",
   957 => x"87d03353",
   958 => x"72e63886",
   959 => x"3d0d0472",
   960 => x"2d800b81",
   961 => x"808087cc",
   962 => x"0c80d4f4",
   963 => x"518dc13f",
   964 => x"81808087",
   965 => x"d0335372",
   966 => x"c738e039",
   967 => x"90863f80",
   968 => x"0881ff06",
   969 => x"51f8d33f",
   970 => x"ffb639fc",
   971 => x"3d0d8a51",
   972 => x"8d823f80",
   973 => x"d6bc518d",
   974 => x"973f800b",
   975 => x"81808087",
   976 => x"c4335353",
   977 => x"72722780",
   978 => x"fb387210",
   979 => x"10107310",
   980 => x"05818080",
   981 => x"80940570",
   982 => x"52548cf4",
   983 => x"3f72822b",
   984 => x"7311832b",
   985 => x"81808081",
   986 => x"b4113351",
   987 => x"53557180",
   988 => x"2eb83873",
   989 => x"519b913f",
   990 => x"800881ff",
   991 => x"06527189",
   992 => x"269338a0",
   993 => x"518cad3f",
   994 => x"81127081",
   995 => x"ff065354",
   996 => x"897227ef",
   997 => x"3880d6d4",
   998 => x"518cb53f",
   999 => x"7215832b",
  1000 => x"81808081",
  1001 => x"b405518c",
  1002 => x"a73f8a51",
  1003 => x"8c863f81",
  1004 => x"137081ff",
  1005 => x"06818080",
  1006 => x"87c43354",
  1007 => x"54557173",
  1008 => x"26ff8738",
  1009 => x"8a518bec",
  1010 => x"3f863d0d",
  1011 => x"04803d0d",
  1012 => x"8c518be0",
  1013 => x"3f823d0d",
  1014 => x"04fe3d0d",
  1015 => x"02930533",
  1016 => x"80d6e452",
  1017 => x"538be93f",
  1018 => x"72518c89",
  1019 => x"3f80d6f0",
  1020 => x"518bdd3f",
  1021 => x"72882b80",
  1022 => x"db980811",
  1023 => x"70085353",
  1024 => x"538bf23f",
  1025 => x"80d6fc51",
  1026 => x"8bc63f80",
  1027 => x"db980813",
  1028 => x"84110852",
  1029 => x"528bde3f",
  1030 => x"80d78851",
  1031 => x"8bb23f80",
  1032 => x"db980813",
  1033 => x"88110852",
  1034 => x"528bca3f",
  1035 => x"80d79451",
  1036 => x"8b9e3f80",
  1037 => x"db980813",
  1038 => x"8c110852",
  1039 => x"528bb63f",
  1040 => x"80d7a051",
  1041 => x"8b8a3f80",
  1042 => x"db980813",
  1043 => x"90110852",
  1044 => x"538ba23f",
  1045 => x"8a518adc",
  1046 => x"3f843d0d",
  1047 => x"04ff3d0d",
  1048 => x"80527151",
  1049 => x"fef33f81",
  1050 => x"127081ff",
  1051 => x"06515283",
  1052 => x"7227ef38",
  1053 => x"833d0d04",
  1054 => x"f03d0d80",
  1055 => x"0b818080",
  1056 => x"86f43381",
  1057 => x"808086f4",
  1058 => x"59555673",
  1059 => x"a02e0981",
  1060 => x"06983881",
  1061 => x"167081ff",
  1062 => x"06818080",
  1063 => x"86f41170",
  1064 => x"33535957",
  1065 => x"5473a02e",
  1066 => x"ea388058",
  1067 => x"80773356",
  1068 => x"5474742e",
  1069 => x"83388154",
  1070 => x"74a02e83",
  1071 => x"f5387384",
  1072 => x"a63874a0",
  1073 => x"2e83eb38",
  1074 => x"81187081",
  1075 => x"ff06595a",
  1076 => x"817826d8",
  1077 => x"388a5392",
  1078 => x"3dfc0552",
  1079 => x"76519dcc",
  1080 => x"3f800881",
  1081 => x"ff065980",
  1082 => x"0b818080",
  1083 => x"86f43381",
  1084 => x"808086f4",
  1085 => x"59555673",
  1086 => x"a02e0981",
  1087 => x"06983881",
  1088 => x"167081ff",
  1089 => x"06818080",
  1090 => x"86f41170",
  1091 => x"33575957",
  1092 => x"5873a02e",
  1093 => x"ea388058",
  1094 => x"80773356",
  1095 => x"5474742e",
  1096 => x"83388154",
  1097 => x"74a02e83",
  1098 => x"d0387384",
  1099 => x"813874a0",
  1100 => x"2e83c638",
  1101 => x"81187081",
  1102 => x"ff065955",
  1103 => x"827826d8",
  1104 => x"388a5392",
  1105 => x"3df80552",
  1106 => x"76519ce0",
  1107 => x"3f80085c",
  1108 => x"800b8180",
  1109 => x"8086f433",
  1110 => x"81808086",
  1111 => x"f4595556",
  1112 => x"73a02e09",
  1113 => x"81069838",
  1114 => x"81167081",
  1115 => x"ff068180",
  1116 => x"8086f411",
  1117 => x"70335752",
  1118 => x"575773a0",
  1119 => x"2eea3880",
  1120 => x"58807733",
  1121 => x"56547474",
  1122 => x"2e833881",
  1123 => x"5474a02e",
  1124 => x"83ae3873",
  1125 => x"83df3874",
  1126 => x"a02e83a4",
  1127 => x"38811870",
  1128 => x"81ff0659",
  1129 => x"5a837826",
  1130 => x"d8388a53",
  1131 => x"923df405",
  1132 => x"5276519b",
  1133 => x"f73f8008",
  1134 => x"5b800b81",
  1135 => x"808086f4",
  1136 => x"33818080",
  1137 => x"86f45955",
  1138 => x"5673a02e",
  1139 => x"09810698",
  1140 => x"38811670",
  1141 => x"81ff0681",
  1142 => x"808086f4",
  1143 => x"11703357",
  1144 => x"59575873",
  1145 => x"a02eea38",
  1146 => x"80588077",
  1147 => x"33565474",
  1148 => x"742e8338",
  1149 => x"815474a0",
  1150 => x"2e838c38",
  1151 => x"7383bd38",
  1152 => x"74a02e83",
  1153 => x"82388118",
  1154 => x"7081ff06",
  1155 => x"595a8478",
  1156 => x"26d8388a",
  1157 => x"53923df0",
  1158 => x"05527651",
  1159 => x"9b8e3f80",
  1160 => x"085a800b",
  1161 => x"81808086",
  1162 => x"f4338180",
  1163 => x"8086f459",
  1164 => x"555673a0",
  1165 => x"2e098106",
  1166 => x"98388116",
  1167 => x"7081ff06",
  1168 => x"81808086",
  1169 => x"f4117033",
  1170 => x"57595758",
  1171 => x"73a02eea",
  1172 => x"38805880",
  1173 => x"77335654",
  1174 => x"74742e83",
  1175 => x"38815474",
  1176 => x"a02e82ea",
  1177 => x"3873839b",
  1178 => x"3874a02e",
  1179 => x"82e03881",
  1180 => x"187081ff",
  1181 => x"06595485",
  1182 => x"7826d838",
  1183 => x"8a53923d",
  1184 => x"ec055276",
  1185 => x"519aa53f",
  1186 => x"78832683",
  1187 => x"88387882",
  1188 => x"802980db",
  1189 => x"9808057c",
  1190 => x"84120c7b",
  1191 => x"88120c7a",
  1192 => x"8c120c80",
  1193 => x"0890120c",
  1194 => x"587851fa",
  1195 => x"ac3f923d",
  1196 => x"0d048116",
  1197 => x"7081ff06",
  1198 => x"81808086",
  1199 => x"f4117033",
  1200 => x"5c525757",
  1201 => x"78a02e09",
  1202 => x"8106fbfc",
  1203 => x"38811670",
  1204 => x"81ff0681",
  1205 => x"808086f4",
  1206 => x"1170335c",
  1207 => x"52575778",
  1208 => x"a02ecf38",
  1209 => x"fbe23981",
  1210 => x"167081ff",
  1211 => x"06818080",
  1212 => x"86f41159",
  1213 => x"5755fbb4",
  1214 => x"39811670",
  1215 => x"81ff0681",
  1216 => x"808086f4",
  1217 => x"1170335f",
  1218 => x"5957547b",
  1219 => x"a02e0981",
  1220 => x"06fca138",
  1221 => x"81167081",
  1222 => x"ff068180",
  1223 => x"8086f411",
  1224 => x"70335f59",
  1225 => x"57547ba0",
  1226 => x"2ecf38fc",
  1227 => x"87398116",
  1228 => x"7081ff06",
  1229 => x"81808086",
  1230 => x"f4115957",
  1231 => x"5bfbd939",
  1232 => x"81167081",
  1233 => x"ff068180",
  1234 => x"8086f411",
  1235 => x"70335759",
  1236 => x"575573a0",
  1237 => x"2e098106",
  1238 => x"fcc33881",
  1239 => x"167081ff",
  1240 => x"06818080",
  1241 => x"86f41170",
  1242 => x"33575957",
  1243 => x"5573a02e",
  1244 => x"cf38fca9",
  1245 => x"39811670",
  1246 => x"81ff0681",
  1247 => x"808086f4",
  1248 => x"1159575b",
  1249 => x"fbfb3981",
  1250 => x"167081ff",
  1251 => x"06818080",
  1252 => x"86f41170",
  1253 => x"33575957",
  1254 => x"5573a02e",
  1255 => x"098106fc",
  1256 => x"e5388116",
  1257 => x"7081ff06",
  1258 => x"81808086",
  1259 => x"f4117033",
  1260 => x"57595755",
  1261 => x"73a02ecf",
  1262 => x"38fccb39",
  1263 => x"81167081",
  1264 => x"ff068180",
  1265 => x"8086f411",
  1266 => x"525757fc",
  1267 => x"9d398116",
  1268 => x"7081ff06",
  1269 => x"81808086",
  1270 => x"f4117033",
  1271 => x"57595755",
  1272 => x"73a02e09",
  1273 => x"8106fd87",
  1274 => x"38811670",
  1275 => x"81ff0681",
  1276 => x"808086f4",
  1277 => x"11703357",
  1278 => x"59575573",
  1279 => x"a02ecf38",
  1280 => x"fced3981",
  1281 => x"167081ff",
  1282 => x"06818080",
  1283 => x"86f41152",
  1284 => x"5757fcbf",
  1285 => x"3980d7ac",
  1286 => x"5183b53f",
  1287 => x"785183d5",
  1288 => x"3f80d7cc",
  1289 => x"5183a93f",
  1290 => x"923d0d04",
  1291 => x"fe3d0d80",
  1292 => x"0b80db98",
  1293 => x"08545271",
  1294 => x"82802913",
  1295 => x"5181710c",
  1296 => x"81127081",
  1297 => x"ff065351",
  1298 => x"837227eb",
  1299 => x"3880dba0",
  1300 => x"08841108",
  1301 => x"810a0784",
  1302 => x"120c5284",
  1303 => x"3d0d04ff",
  1304 => x"3d0d80db",
  1305 => x"a0088411",
  1306 => x"0870fe0a",
  1307 => x"0684130c",
  1308 => x"5252833d",
  1309 => x"0d04fd3d",
  1310 => x"0d80dba0",
  1311 => x"08700881",
  1312 => x"0a068180",
  1313 => x"8080900c",
  1314 => x"5484f03f",
  1315 => x"81808080",
  1316 => x"9008ab9e",
  1317 => x"55537284",
  1318 => x"3896e154",
  1319 => x"73818080",
  1320 => x"87d40c72",
  1321 => x"802e81f0",
  1322 => x"3885eb3f",
  1323 => x"80d7f451",
  1324 => x"829e3f8c",
  1325 => x"5181fd3f",
  1326 => x"80d7f851",
  1327 => x"82923f81",
  1328 => x"80808090",
  1329 => x"08802e81",
  1330 => x"a43880d8",
  1331 => x"94518280",
  1332 => x"3f818080",
  1333 => x"80900880",
  1334 => x"2e81a238",
  1335 => x"80db9808",
  1336 => x"54820b84",
  1337 => x"150c800b",
  1338 => x"88150c80",
  1339 => x"0b8c150c",
  1340 => x"840b9015",
  1341 => x"0c800b82",
  1342 => x"84150c81",
  1343 => x"0b828815",
  1344 => x"0c810b82",
  1345 => x"8c150c80",
  1346 => x"0b829015",
  1347 => x"0c810b82",
  1348 => x"80150c81",
  1349 => x"0b848415",
  1350 => x"0c820b84",
  1351 => x"88150c82",
  1352 => x"0b848c15",
  1353 => x"0c800b84",
  1354 => x"90150c81",
  1355 => x"0b848015",
  1356 => x"0c820b86",
  1357 => x"84150c82",
  1358 => x"0b868815",
  1359 => x"0c820b86",
  1360 => x"8c150c83",
  1361 => x"0b869015",
  1362 => x"0c810b86",
  1363 => x"80150c80",
  1364 => x"dba00884",
  1365 => x"11087081",
  1366 => x"0a078413",
  1367 => x"0c548411",
  1368 => x"0870fe0a",
  1369 => x"0684130c",
  1370 => x"54548aa9",
  1371 => x"3f80d8a0",
  1372 => x"5180dd3f",
  1373 => x"81808080",
  1374 => x"9008fee0",
  1375 => x"3880d8c4",
  1376 => x"51eabe3f",
  1377 => x"82528351",
  1378 => x"e5ce3f80",
  1379 => x"d8d851ea",
  1380 => x"b03feeb5",
  1381 => x"3f89fe3f",
  1382 => x"dfea3ffe",
  1383 => x"8c39ff3d",
  1384 => x"0d028f05",
  1385 => x"3380dbac",
  1386 => x"0852710c",
  1387 => x"800b800c",
  1388 => x"833d0d04",
  1389 => x"ff3d0d02",
  1390 => x"8f053351",
  1391 => x"81808087",
  1392 => x"d4085271",
  1393 => x"2d800881",
  1394 => x"ff06800c",
  1395 => x"833d0d04",
  1396 => x"fe3d0d74",
  1397 => x"70335353",
  1398 => x"71802e95",
  1399 => x"38811372",
  1400 => x"52818080",
  1401 => x"87d40853",
  1402 => x"53712d72",
  1403 => x"335271ed",
  1404 => x"38843d0d",
  1405 => x"04f23d0d",
  1406 => x"608c3d70",
  1407 => x"5b5b5380",
  1408 => x"73565776",
  1409 => x"732480fa",
  1410 => x"38781754",
  1411 => x"8a527451",
  1412 => x"84e23f80",
  1413 => x"08b00553",
  1414 => x"72743481",
  1415 => x"17578a52",
  1416 => x"745184ab",
  1417 => x"3f800855",
  1418 => x"8008de38",
  1419 => x"8008779f",
  1420 => x"2a187081",
  1421 => x"2c5a5656",
  1422 => x"8078259e",
  1423 => x"387817ff",
  1424 => x"05557519",
  1425 => x"70335553",
  1426 => x"74337334",
  1427 => x"73753481",
  1428 => x"16ff1656",
  1429 => x"56777624",
  1430 => x"e9387619",
  1431 => x"56807634",
  1432 => x"79703354",
  1433 => x"5472802e",
  1434 => x"95388114",
  1435 => x"73528180",
  1436 => x"8087d408",
  1437 => x"5854762d",
  1438 => x"73335372",
  1439 => x"ed38903d",
  1440 => x"0d04ad7a",
  1441 => x"3402a905",
  1442 => x"73307119",
  1443 => x"5656598a",
  1444 => x"52745183",
  1445 => x"df3f8008",
  1446 => x"b0055372",
  1447 => x"74348117",
  1448 => x"578a5274",
  1449 => x"5183a83f",
  1450 => x"80085580",
  1451 => x"08feda38",
  1452 => x"fefa39ff",
  1453 => x"3d0d80db",
  1454 => x"a4087410",
  1455 => x"10751005",
  1456 => x"94120c52",
  1457 => x"850b9813",
  1458 => x"0c981208",
  1459 => x"70810651",
  1460 => x"5170f638",
  1461 => x"833d0d04",
  1462 => x"fd3d0d80",
  1463 => x"dba40876",
  1464 => x"b0ea2994",
  1465 => x"120c5485",
  1466 => x"0b98150c",
  1467 => x"98140870",
  1468 => x"81065153",
  1469 => x"72f63885",
  1470 => x"3d0d0480",
  1471 => x"3d0d80db",
  1472 => x"a80851b6",
  1473 => x"0b8c120c",
  1474 => x"830b8812",
  1475 => x"0c823d0d",
  1476 => x"04803d0d",
  1477 => x"80dba808",
  1478 => x"84110881",
  1479 => x"06800c51",
  1480 => x"823d0d04",
  1481 => x"ff3d0d80",
  1482 => x"dba80852",
  1483 => x"84120870",
  1484 => x"81065151",
  1485 => x"70802ef4",
  1486 => x"38710870",
  1487 => x"81ff0680",
  1488 => x"0c51833d",
  1489 => x"0d04fe3d",
  1490 => x"0d029305",
  1491 => x"3353728a",
  1492 => x"2e9c3880",
  1493 => x"dba80852",
  1494 => x"84120870",
  1495 => x"892a7081",
  1496 => x"06515151",
  1497 => x"70f23872",
  1498 => x"720c843d",
  1499 => x"0d0480db",
  1500 => x"a8085284",
  1501 => x"12087089",
  1502 => x"2a708106",
  1503 => x"51515170",
  1504 => x"f2388d72",
  1505 => x"0c841208",
  1506 => x"70892a70",
  1507 => x"81065151",
  1508 => x"5170c538",
  1509 => x"d239803d",
  1510 => x"0d80db9c",
  1511 => x"0851800b",
  1512 => x"84120c83",
  1513 => x"fe800b88",
  1514 => x"120c800b",
  1515 => x"81808087",
  1516 => x"d834800b",
  1517 => x"81808087",
  1518 => x"dc34823d",
  1519 => x"0d04fa3d",
  1520 => x"0d02a305",
  1521 => x"3380db9c",
  1522 => x"08818080",
  1523 => x"87d83370",
  1524 => x"81ff0670",
  1525 => x"10101181",
  1526 => x"808087dc",
  1527 => x"337081ff",
  1528 => x"06729029",
  1529 => x"1170882b",
  1530 => x"7807770c",
  1531 => x"535b5b55",
  1532 => x"55595454",
  1533 => x"738a2e9a",
  1534 => x"387480cf",
  1535 => x"2e943873",
  1536 => x"8c2eaa38",
  1537 => x"81165372",
  1538 => x"81808087",
  1539 => x"dc34883d",
  1540 => x"0d0471a3",
  1541 => x"26a73881",
  1542 => x"17527181",
  1543 => x"808087d8",
  1544 => x"34800b81",
  1545 => x"808087dc",
  1546 => x"34883d0d",
  1547 => x"04805271",
  1548 => x"882b730c",
  1549 => x"81125297",
  1550 => x"907226f3",
  1551 => x"38800b81",
  1552 => x"808087d8",
  1553 => x"34800b81",
  1554 => x"808087dc",
  1555 => x"34db398c",
  1556 => x"08028c0c",
  1557 => x"fd3d0d80",
  1558 => x"538c088c",
  1559 => x"0508528c",
  1560 => x"08880508",
  1561 => x"5182de3f",
  1562 => x"80087080",
  1563 => x"0c54853d",
  1564 => x"0d8c0c04",
  1565 => x"8c08028c",
  1566 => x"0cfd3d0d",
  1567 => x"81538c08",
  1568 => x"8c050852",
  1569 => x"8c088805",
  1570 => x"085182b9",
  1571 => x"3f800870",
  1572 => x"800c5485",
  1573 => x"3d0d8c0c",
  1574 => x"048c0802",
  1575 => x"8c0cf93d",
  1576 => x"0d800b8c",
  1577 => x"08fc050c",
  1578 => x"8c088805",
  1579 => x"088025ab",
  1580 => x"388c0888",
  1581 => x"0508308c",
  1582 => x"0888050c",
  1583 => x"800b8c08",
  1584 => x"f4050c8c",
  1585 => x"08fc0508",
  1586 => x"8838810b",
  1587 => x"8c08f405",
  1588 => x"0c8c08f4",
  1589 => x"05088c08",
  1590 => x"fc050c8c",
  1591 => x"088c0508",
  1592 => x"8025ab38",
  1593 => x"8c088c05",
  1594 => x"08308c08",
  1595 => x"8c050c80",
  1596 => x"0b8c08f0",
  1597 => x"050c8c08",
  1598 => x"fc050888",
  1599 => x"38810b8c",
  1600 => x"08f0050c",
  1601 => x"8c08f005",
  1602 => x"088c08fc",
  1603 => x"050c8053",
  1604 => x"8c088c05",
  1605 => x"08528c08",
  1606 => x"88050851",
  1607 => x"81a73f80",
  1608 => x"08708c08",
  1609 => x"f8050c54",
  1610 => x"8c08fc05",
  1611 => x"08802e8c",
  1612 => x"388c08f8",
  1613 => x"0508308c",
  1614 => x"08f8050c",
  1615 => x"8c08f805",
  1616 => x"0870800c",
  1617 => x"54893d0d",
  1618 => x"8c0c048c",
  1619 => x"08028c0c",
  1620 => x"fb3d0d80",
  1621 => x"0b8c08fc",
  1622 => x"050c8c08",
  1623 => x"88050880",
  1624 => x"2593388c",
  1625 => x"08880508",
  1626 => x"308c0888",
  1627 => x"050c810b",
  1628 => x"8c08fc05",
  1629 => x"0c8c088c",
  1630 => x"05088025",
  1631 => x"8c388c08",
  1632 => x"8c050830",
  1633 => x"8c088c05",
  1634 => x"0c81538c",
  1635 => x"088c0508",
  1636 => x"528c0888",
  1637 => x"050851ad",
  1638 => x"3f800870",
  1639 => x"8c08f805",
  1640 => x"0c548c08",
  1641 => x"fc050880",
  1642 => x"2e8c388c",
  1643 => x"08f80508",
  1644 => x"308c08f8",
  1645 => x"050c8c08",
  1646 => x"f8050870",
  1647 => x"800c5487",
  1648 => x"3d0d8c0c",
  1649 => x"048c0802",
  1650 => x"8c0cfd3d",
  1651 => x"0d810b8c",
  1652 => x"08fc050c",
  1653 => x"800b8c08",
  1654 => x"f8050c8c",
  1655 => x"088c0508",
  1656 => x"8c088805",
  1657 => x"0827ac38",
  1658 => x"8c08fc05",
  1659 => x"08802ea3",
  1660 => x"38800b8c",
  1661 => x"088c0508",
  1662 => x"2499388c",
  1663 => x"088c0508",
  1664 => x"108c088c",
  1665 => x"050c8c08",
  1666 => x"fc050810",
  1667 => x"8c08fc05",
  1668 => x"0cc9398c",
  1669 => x"08fc0508",
  1670 => x"802e80c9",
  1671 => x"388c088c",
  1672 => x"05088c08",
  1673 => x"88050826",
  1674 => x"a1388c08",
  1675 => x"8805088c",
  1676 => x"088c0508",
  1677 => x"318c0888",
  1678 => x"050c8c08",
  1679 => x"f805088c",
  1680 => x"08fc0508",
  1681 => x"078c08f8",
  1682 => x"050c8c08",
  1683 => x"fc050881",
  1684 => x"2a8c08fc",
  1685 => x"050c8c08",
  1686 => x"8c050881",
  1687 => x"2a8c088c",
  1688 => x"050cffaf",
  1689 => x"398c0890",
  1690 => x"0508802e",
  1691 => x"8f388c08",
  1692 => x"88050870",
  1693 => x"8c08f405",
  1694 => x"0c518d39",
  1695 => x"8c08f805",
  1696 => x"08708c08",
  1697 => x"f4050c51",
  1698 => x"8c08f405",
  1699 => x"08800c85",
  1700 => x"3d0d8c0c",
  1701 => x"04803d0d",
  1702 => x"865182fd",
  1703 => x"3f81519d",
  1704 => x"f93ffd3d",
  1705 => x"0d755384",
  1706 => x"d8130880",
  1707 => x"2e8a3880",
  1708 => x"5372800c",
  1709 => x"853d0d04",
  1710 => x"81805272",
  1711 => x"518a823f",
  1712 => x"800884d8",
  1713 => x"140cff53",
  1714 => x"8008802e",
  1715 => x"e4388008",
  1716 => x"549f5380",
  1717 => x"74708405",
  1718 => x"560cff13",
  1719 => x"53807324",
  1720 => x"ce388074",
  1721 => x"70840556",
  1722 => x"0cff1353",
  1723 => x"728025e3",
  1724 => x"38ffbc39",
  1725 => x"fd3d0d75",
  1726 => x"7755539f",
  1727 => x"74278d38",
  1728 => x"96730cff",
  1729 => x"5271800c",
  1730 => x"853d0d04",
  1731 => x"84d81308",
  1732 => x"5271802e",
  1733 => x"93387310",
  1734 => x"10127008",
  1735 => x"79720c51",
  1736 => x"5271800c",
  1737 => x"853d0d04",
  1738 => x"7251fef6",
  1739 => x"3fff5280",
  1740 => x"08d33884",
  1741 => x"d8130874",
  1742 => x"10101170",
  1743 => x"087a720c",
  1744 => x"515152dd",
  1745 => x"39f93d0d",
  1746 => x"797b5856",
  1747 => x"769f2680",
  1748 => x"e83884d8",
  1749 => x"16085473",
  1750 => x"802eaa38",
  1751 => x"76101014",
  1752 => x"70085555",
  1753 => x"73802eba",
  1754 => x"38805873",
  1755 => x"812e8f38",
  1756 => x"73ff2ea3",
  1757 => x"3880750c",
  1758 => x"7651732d",
  1759 => x"80587780",
  1760 => x"0c893d0d",
  1761 => x"047551fe",
  1762 => x"993fff58",
  1763 => x"8008ef38",
  1764 => x"84d81608",
  1765 => x"54c63996",
  1766 => x"760c810b",
  1767 => x"800c893d",
  1768 => x"0d047551",
  1769 => x"81f13f76",
  1770 => x"53800852",
  1771 => x"755181ad",
  1772 => x"3f800880",
  1773 => x"0c893d0d",
  1774 => x"0496760c",
  1775 => x"ff0b800c",
  1776 => x"893d0d04",
  1777 => x"fc3d0d76",
  1778 => x"785653ff",
  1779 => x"54749f26",
  1780 => x"b13884d8",
  1781 => x"13085271",
  1782 => x"802eae38",
  1783 => x"74101012",
  1784 => x"70085353",
  1785 => x"81547180",
  1786 => x"2e983882",
  1787 => x"5471ff2e",
  1788 => x"91388354",
  1789 => x"71812e8a",
  1790 => x"3880730c",
  1791 => x"7451712d",
  1792 => x"80547380",
  1793 => x"0c863d0d",
  1794 => x"047251fd",
  1795 => x"953f8008",
  1796 => x"f13884d8",
  1797 => x"130852c4",
  1798 => x"39ff3d0d",
  1799 => x"735280db",
  1800 => x"b00851fe",
  1801 => x"a03f833d",
  1802 => x"0d04fe3d",
  1803 => x"0d755374",
  1804 => x"5280dbb0",
  1805 => x"0851fdbc",
  1806 => x"3f843d0d",
  1807 => x"04803d0d",
  1808 => x"80dbb008",
  1809 => x"51fcdb3f",
  1810 => x"823d0d04",
  1811 => x"ff3d0d73",
  1812 => x"5280dbb0",
  1813 => x"0851feec",
  1814 => x"3f833d0d",
  1815 => x"04fc3d0d",
  1816 => x"800b8180",
  1817 => x"8087e80c",
  1818 => x"78527751",
  1819 => x"99943f80",
  1820 => x"08548008",
  1821 => x"ff2e8838",
  1822 => x"73800c86",
  1823 => x"3d0d0481",
  1824 => x"808087e8",
  1825 => x"08557480",
  1826 => x"2eee3876",
  1827 => x"75710c53",
  1828 => x"73800c86",
  1829 => x"3d0d0498",
  1830 => x"e43f04fc",
  1831 => x"3d0d7670",
  1832 => x"79707307",
  1833 => x"83065454",
  1834 => x"54557080",
  1835 => x"c3387170",
  1836 => x"08700970",
  1837 => x"f7fbfdff",
  1838 => x"130670f8",
  1839 => x"84828180",
  1840 => x"06515153",
  1841 => x"535470a6",
  1842 => x"38841472",
  1843 => x"74708405",
  1844 => x"560c7008",
  1845 => x"700970f7",
  1846 => x"fbfdff13",
  1847 => x"0670f884",
  1848 => x"82818006",
  1849 => x"51515353",
  1850 => x"5470802e",
  1851 => x"dc387352",
  1852 => x"71708105",
  1853 => x"53335170",
  1854 => x"73708105",
  1855 => x"553470f0",
  1856 => x"3874800c",
  1857 => x"863d0d04",
  1858 => x"fd3d0d75",
  1859 => x"70718306",
  1860 => x"53555270",
  1861 => x"b8387170",
  1862 => x"087009f7",
  1863 => x"fbfdff12",
  1864 => x"0670f884",
  1865 => x"82818006",
  1866 => x"51515253",
  1867 => x"709d3884",
  1868 => x"13700870",
  1869 => x"09f7fbfd",
  1870 => x"ff120670",
  1871 => x"f8848281",
  1872 => x"80065151",
  1873 => x"52537080",
  1874 => x"2ee53872",
  1875 => x"52713351",
  1876 => x"70802e8a",
  1877 => x"38811270",
  1878 => x"33525270",
  1879 => x"f8387174",
  1880 => x"31800c85",
  1881 => x"3d0d04fa",
  1882 => x"3d0d787a",
  1883 => x"7c705455",
  1884 => x"55527280",
  1885 => x"2e80d938",
  1886 => x"71740783",
  1887 => x"06517080",
  1888 => x"2e80d438",
  1889 => x"ff135372",
  1890 => x"ff2eb138",
  1891 => x"71337433",
  1892 => x"56517471",
  1893 => x"2e098106",
  1894 => x"a9387280",
  1895 => x"2e818738",
  1896 => x"7081ff06",
  1897 => x"5170802e",
  1898 => x"80fc3881",
  1899 => x"128115ff",
  1900 => x"15555552",
  1901 => x"72ff2e09",
  1902 => x"8106d138",
  1903 => x"71337433",
  1904 => x"56517081",
  1905 => x"ff067581",
  1906 => x"ff067171",
  1907 => x"31515252",
  1908 => x"70800c88",
  1909 => x"3d0d0471",
  1910 => x"74575583",
  1911 => x"73278838",
  1912 => x"71087408",
  1913 => x"2e883874",
  1914 => x"765552ff",
  1915 => x"9739fc13",
  1916 => x"5372802e",
  1917 => x"b1387408",
  1918 => x"7009f7fb",
  1919 => x"fdff1206",
  1920 => x"70f88482",
  1921 => x"81800651",
  1922 => x"5151709a",
  1923 => x"38841584",
  1924 => x"17575583",
  1925 => x"7327d038",
  1926 => x"74087608",
  1927 => x"2ed03874",
  1928 => x"765552fe",
  1929 => x"df39800b",
  1930 => x"800c883d",
  1931 => x"0d04f33d",
  1932 => x"0d606264",
  1933 => x"725a5a5e",
  1934 => x"5e805c76",
  1935 => x"70810558",
  1936 => x"3380d8e5",
  1937 => x"11337083",
  1938 => x"2a708106",
  1939 => x"51555556",
  1940 => x"72e93875",
  1941 => x"ad2e8288",
  1942 => x"3875ab2e",
  1943 => x"82843877",
  1944 => x"30707907",
  1945 => x"80257990",
  1946 => x"32703070",
  1947 => x"72078025",
  1948 => x"73075357",
  1949 => x"57515372",
  1950 => x"802e8738",
  1951 => x"75b02e81",
  1952 => x"eb38778a",
  1953 => x"38885875",
  1954 => x"b02e8338",
  1955 => x"8a58810a",
  1956 => x"5a7b8438",
  1957 => x"fe0a5a77",
  1958 => x"527951f3",
  1959 => x"d73f8008",
  1960 => x"78537a52",
  1961 => x"5bf3a83f",
  1962 => x"80085a80",
  1963 => x"7080d8e5",
  1964 => x"18337082",
  1965 => x"2a708106",
  1966 => x"5156565a",
  1967 => x"5572802e",
  1968 => x"80c138d0",
  1969 => x"16567578",
  1970 => x"2580d738",
  1971 => x"80792475",
  1972 => x"7b260753",
  1973 => x"72933874",
  1974 => x"7a2e80eb",
  1975 => x"387a7625",
  1976 => x"80ed3872",
  1977 => x"802e80e7",
  1978 => x"38ff7770",
  1979 => x"81055933",
  1980 => x"575980d8",
  1981 => x"e5163370",
  1982 => x"822a7081",
  1983 => x"06515454",
  1984 => x"72c13873",
  1985 => x"83065372",
  1986 => x"802e9738",
  1987 => x"738106c9",
  1988 => x"17555372",
  1989 => x"8538ffa9",
  1990 => x"16547356",
  1991 => x"777624ff",
  1992 => x"ab388079",
  1993 => x"2480f038",
  1994 => x"7b802e84",
  1995 => x"38743055",
  1996 => x"7c802e8c",
  1997 => x"38ff1753",
  1998 => x"7883387d",
  1999 => x"53727d0c",
  2000 => x"74800c8f",
  2001 => x"3d0d0481",
  2002 => x"53757b24",
  2003 => x"ff953881",
  2004 => x"75792917",
  2005 => x"78708105",
  2006 => x"5a335856",
  2007 => x"59ff9339",
  2008 => x"815c7670",
  2009 => x"81055833",
  2010 => x"56fdf439",
  2011 => x"80773354",
  2012 => x"547280f8",
  2013 => x"2eb23872",
  2014 => x"80d83270",
  2015 => x"30708025",
  2016 => x"76075151",
  2017 => x"5372802e",
  2018 => x"fdf83881",
  2019 => x"17338218",
  2020 => x"58569058",
  2021 => x"fdf83981",
  2022 => x"0a557b84",
  2023 => x"38fe0a55",
  2024 => x"7f53a273",
  2025 => x"0cff8939",
  2026 => x"8154cc39",
  2027 => x"fd3d0d77",
  2028 => x"54765375",
  2029 => x"5280dbb0",
  2030 => x"0851fcf2",
  2031 => x"3f853d0d",
  2032 => x"04f33d0d",
  2033 => x"7f618b11",
  2034 => x"70f8065c",
  2035 => x"55555e72",
  2036 => x"96268338",
  2037 => x"90598079",
  2038 => x"24747a26",
  2039 => x"07538054",
  2040 => x"72742e09",
  2041 => x"810680cb",
  2042 => x"387d518b",
  2043 => x"ca3f7883",
  2044 => x"f72680c6",
  2045 => x"3878832a",
  2046 => x"70101010",
  2047 => x"80e2ec05",
  2048 => x"8c110859",
  2049 => x"595a7678",
  2050 => x"2e83b038",
  2051 => x"841708fc",
  2052 => x"06568c17",
  2053 => x"08881808",
  2054 => x"718c120c",
  2055 => x"88120c58",
  2056 => x"75178411",
  2057 => x"08810784",
  2058 => x"120c537d",
  2059 => x"518b893f",
  2060 => x"88175473",
  2061 => x"800c8f3d",
  2062 => x"0d047889",
  2063 => x"2a79832a",
  2064 => x"5b537280",
  2065 => x"2ebf3878",
  2066 => x"862ab805",
  2067 => x"5a847327",
  2068 => x"b43880db",
  2069 => x"135a9473",
  2070 => x"27ab3878",
  2071 => x"8c2a80ee",
  2072 => x"055a80d4",
  2073 => x"73279e38",
  2074 => x"788f2a80",
  2075 => x"f7055a82",
  2076 => x"d4732791",
  2077 => x"3878922a",
  2078 => x"80fc055a",
  2079 => x"8ad47327",
  2080 => x"843880fe",
  2081 => x"5a791010",
  2082 => x"1080e2ec",
  2083 => x"058c1108",
  2084 => x"58557675",
  2085 => x"2ea33884",
  2086 => x"1708fc06",
  2087 => x"707a3155",
  2088 => x"56738f24",
  2089 => x"88d53873",
  2090 => x"8025fee6",
  2091 => x"388c1708",
  2092 => x"5776752e",
  2093 => x"098106df",
  2094 => x"38811a5a",
  2095 => x"80e2fc08",
  2096 => x"577680e2",
  2097 => x"f42e82c0",
  2098 => x"38841708",
  2099 => x"fc06707a",
  2100 => x"31555673",
  2101 => x"8f2481f9",
  2102 => x"3880e2f4",
  2103 => x"0b80e380",
  2104 => x"0c80e2f4",
  2105 => x"0b80e2fc",
  2106 => x"0c738025",
  2107 => x"feb23883",
  2108 => x"ff762783",
  2109 => x"df387589",
  2110 => x"2a76832a",
  2111 => x"55537280",
  2112 => x"2ebf3875",
  2113 => x"862ab805",
  2114 => x"54847327",
  2115 => x"b43880db",
  2116 => x"13549473",
  2117 => x"27ab3875",
  2118 => x"8c2a80ee",
  2119 => x"055480d4",
  2120 => x"73279e38",
  2121 => x"758f2a80",
  2122 => x"f7055482",
  2123 => x"d4732791",
  2124 => x"3875922a",
  2125 => x"80fc0554",
  2126 => x"8ad47327",
  2127 => x"843880fe",
  2128 => x"54731010",
  2129 => x"1080e2ec",
  2130 => x"05881108",
  2131 => x"56587478",
  2132 => x"2e86cf38",
  2133 => x"841508fc",
  2134 => x"06537573",
  2135 => x"278d3888",
  2136 => x"15085574",
  2137 => x"782e0981",
  2138 => x"06ea388c",
  2139 => x"150880e2",
  2140 => x"ec0b8405",
  2141 => x"08718c1a",
  2142 => x"0c76881a",
  2143 => x"0c788813",
  2144 => x"0c788c18",
  2145 => x"0c5d5879",
  2146 => x"53807a24",
  2147 => x"83e63872",
  2148 => x"822c8171",
  2149 => x"2b5c537a",
  2150 => x"7c268198",
  2151 => x"387b7b06",
  2152 => x"537282f1",
  2153 => x"3879fc06",
  2154 => x"84055a7a",
  2155 => x"10707d06",
  2156 => x"545b7282",
  2157 => x"e038841a",
  2158 => x"5af13988",
  2159 => x"178c1108",
  2160 => x"58587678",
  2161 => x"2e098106",
  2162 => x"fcc23882",
  2163 => x"1a5afdec",
  2164 => x"39781779",
  2165 => x"81078419",
  2166 => x"0c7080e3",
  2167 => x"800c7080",
  2168 => x"e2fc0c80",
  2169 => x"e2f40b8c",
  2170 => x"120c8c11",
  2171 => x"0888120c",
  2172 => x"74810784",
  2173 => x"120c7411",
  2174 => x"75710c51",
  2175 => x"537d5187",
  2176 => x"b73f8817",
  2177 => x"54fcac39",
  2178 => x"80e2ec0b",
  2179 => x"8405087a",
  2180 => x"545c7980",
  2181 => x"25fef838",
  2182 => x"82da397a",
  2183 => x"097c0670",
  2184 => x"80e2ec0b",
  2185 => x"84050c5c",
  2186 => x"7a105b7a",
  2187 => x"7c268538",
  2188 => x"7a85b838",
  2189 => x"80e2ec0b",
  2190 => x"88050870",
  2191 => x"841208fc",
  2192 => x"06707c31",
  2193 => x"7c72268f",
  2194 => x"72250757",
  2195 => x"575c5d55",
  2196 => x"72802e80",
  2197 => x"db38797a",
  2198 => x"1680e2e4",
  2199 => x"081b9011",
  2200 => x"5a55575b",
  2201 => x"80e2e008",
  2202 => x"ff2e8838",
  2203 => x"a08f13e0",
  2204 => x"80065776",
  2205 => x"527d5186",
  2206 => x"c03f8008",
  2207 => x"548008ff",
  2208 => x"2e903880",
  2209 => x"08762782",
  2210 => x"99387480",
  2211 => x"e2ec2e82",
  2212 => x"913880e2",
  2213 => x"ec0b8805",
  2214 => x"08558415",
  2215 => x"08fc0670",
  2216 => x"7a317a72",
  2217 => x"268f7225",
  2218 => x"07525553",
  2219 => x"7283e638",
  2220 => x"74798107",
  2221 => x"84170c79",
  2222 => x"167080e2",
  2223 => x"ec0b8805",
  2224 => x"0c758107",
  2225 => x"84120c54",
  2226 => x"7e525785",
  2227 => x"eb3f8817",
  2228 => x"54fae039",
  2229 => x"75832a70",
  2230 => x"54548074",
  2231 => x"24819b38",
  2232 => x"72822c81",
  2233 => x"712b80e2",
  2234 => x"f0080770",
  2235 => x"80e2ec0b",
  2236 => x"84050c75",
  2237 => x"10101080",
  2238 => x"e2ec0588",
  2239 => x"1108585a",
  2240 => x"5d53778c",
  2241 => x"180c7488",
  2242 => x"180c7688",
  2243 => x"190c768c",
  2244 => x"160cfcf3",
  2245 => x"39797a10",
  2246 => x"101080e2",
  2247 => x"ec057057",
  2248 => x"595d8c15",
  2249 => x"08577675",
  2250 => x"2ea33884",
  2251 => x"1708fc06",
  2252 => x"707a3155",
  2253 => x"56738f24",
  2254 => x"83ca3873",
  2255 => x"80258481",
  2256 => x"388c1708",
  2257 => x"5776752e",
  2258 => x"098106df",
  2259 => x"38881581",
  2260 => x"1b708306",
  2261 => x"555b5572",
  2262 => x"c9387c83",
  2263 => x"06537280",
  2264 => x"2efdb838",
  2265 => x"ff1df819",
  2266 => x"595d8818",
  2267 => x"08782eea",
  2268 => x"38fdb539",
  2269 => x"831a53fc",
  2270 => x"96398314",
  2271 => x"70822c81",
  2272 => x"712b80e2",
  2273 => x"f0080770",
  2274 => x"80e2ec0b",
  2275 => x"84050c76",
  2276 => x"10101080",
  2277 => x"e2ec0588",
  2278 => x"1108595b",
  2279 => x"5e5153fe",
  2280 => x"e13980e2",
  2281 => x"b0081758",
  2282 => x"8008762e",
  2283 => x"818d3880",
  2284 => x"e2e008ff",
  2285 => x"2e83ec38",
  2286 => x"73763118",
  2287 => x"80e2b00c",
  2288 => x"73870670",
  2289 => x"57537280",
  2290 => x"2e883888",
  2291 => x"73317015",
  2292 => x"55567614",
  2293 => x"9fff06a0",
  2294 => x"80713117",
  2295 => x"70547f53",
  2296 => x"575383d5",
  2297 => x"3f800853",
  2298 => x"8008ff2e",
  2299 => x"81a03880",
  2300 => x"e2b00816",
  2301 => x"7080e2b0",
  2302 => x"0c747580",
  2303 => x"e2ec0b88",
  2304 => x"050c7476",
  2305 => x"31187081",
  2306 => x"07515556",
  2307 => x"587b80e2",
  2308 => x"ec2e839c",
  2309 => x"38798f26",
  2310 => x"82cb3881",
  2311 => x"0b84150c",
  2312 => x"841508fc",
  2313 => x"06707a31",
  2314 => x"7a72268f",
  2315 => x"72250752",
  2316 => x"55537280",
  2317 => x"2efcf938",
  2318 => x"80db3980",
  2319 => x"089fff06",
  2320 => x"5372feeb",
  2321 => x"387780e2",
  2322 => x"b00c80e2",
  2323 => x"ec0b8805",
  2324 => x"087b1881",
  2325 => x"0784120c",
  2326 => x"5580e2dc",
  2327 => x"08782786",
  2328 => x"387780e2",
  2329 => x"dc0c80e2",
  2330 => x"d8087827",
  2331 => x"fcac3877",
  2332 => x"80e2d80c",
  2333 => x"841508fc",
  2334 => x"06707a31",
  2335 => x"7a72268f",
  2336 => x"72250752",
  2337 => x"55537280",
  2338 => x"2efca538",
  2339 => x"88398074",
  2340 => x"5456fedb",
  2341 => x"397d5182",
  2342 => x"9f3f800b",
  2343 => x"800c8f3d",
  2344 => x"0d047353",
  2345 => x"807424a9",
  2346 => x"3872822c",
  2347 => x"81712b80",
  2348 => x"e2f00807",
  2349 => x"7080e2ec",
  2350 => x"0b84050c",
  2351 => x"5d53778c",
  2352 => x"180c7488",
  2353 => x"180c7688",
  2354 => x"190c768c",
  2355 => x"160cf9b7",
  2356 => x"39831470",
  2357 => x"822c8171",
  2358 => x"2b80e2f0",
  2359 => x"08077080",
  2360 => x"e2ec0b84",
  2361 => x"050c5e51",
  2362 => x"53d4397b",
  2363 => x"7b065372",
  2364 => x"fca33884",
  2365 => x"1a7b105c",
  2366 => x"5af139ff",
  2367 => x"1a811151",
  2368 => x"5af7b939",
  2369 => x"78177981",
  2370 => x"0784190c",
  2371 => x"8c180888",
  2372 => x"1908718c",
  2373 => x"120c8812",
  2374 => x"0c597080",
  2375 => x"e3800c70",
  2376 => x"80e2fc0c",
  2377 => x"80e2f40b",
  2378 => x"8c120c8c",
  2379 => x"11088812",
  2380 => x"0c748107",
  2381 => x"84120c74",
  2382 => x"1175710c",
  2383 => x"5153f9bd",
  2384 => x"39751784",
  2385 => x"11088107",
  2386 => x"84120c53",
  2387 => x"8c170888",
  2388 => x"1808718c",
  2389 => x"120c8812",
  2390 => x"0c587d51",
  2391 => x"80da3f88",
  2392 => x"1754f5cf",
  2393 => x"39728415",
  2394 => x"0cf41af8",
  2395 => x"0670841e",
  2396 => x"08810607",
  2397 => x"841e0c70",
  2398 => x"1d545b85",
  2399 => x"0b84140c",
  2400 => x"850b8814",
  2401 => x"0c8f7b27",
  2402 => x"fdcf3888",
  2403 => x"1c527d51",
  2404 => x"82953f80",
  2405 => x"e2ec0b88",
  2406 => x"050880e2",
  2407 => x"b0085955",
  2408 => x"fdb73977",
  2409 => x"80e2b00c",
  2410 => x"7380e2e0",
  2411 => x"0cfc9139",
  2412 => x"7284150c",
  2413 => x"fda33904",
  2414 => x"04fd3d0d",
  2415 => x"800b8180",
  2416 => x"8087e80c",
  2417 => x"765186cf",
  2418 => x"3f800853",
  2419 => x"8008ff2e",
  2420 => x"88387280",
  2421 => x"0c853d0d",
  2422 => x"04818080",
  2423 => x"87e80854",
  2424 => x"73802eee",
  2425 => x"38757471",
  2426 => x"0c527280",
  2427 => x"0c853d0d",
  2428 => x"04fb3d0d",
  2429 => x"77705256",
  2430 => x"ffbd3f80",
  2431 => x"e2ec0b88",
  2432 => x"05088411",
  2433 => x"08fc0670",
  2434 => x"7b319fef",
  2435 => x"05e08006",
  2436 => x"e0800556",
  2437 => x"5653a080",
  2438 => x"74249438",
  2439 => x"80527551",
  2440 => x"ff973f80",
  2441 => x"e2f40815",
  2442 => x"53728008",
  2443 => x"2e8f3875",
  2444 => x"51ff853f",
  2445 => x"80537280",
  2446 => x"0c873d0d",
  2447 => x"04733052",
  2448 => x"7551fef5",
  2449 => x"3f8008ff",
  2450 => x"2ea83880",
  2451 => x"e2ec0b88",
  2452 => x"05087575",
  2453 => x"31810784",
  2454 => x"120c5380",
  2455 => x"e2b00874",
  2456 => x"3180e2b0",
  2457 => x"0c7551fe",
  2458 => x"cf3f810b",
  2459 => x"800c873d",
  2460 => x"0d048052",
  2461 => x"7551fec1",
  2462 => x"3f80e2ec",
  2463 => x"0b880508",
  2464 => x"80087131",
  2465 => x"56538f75",
  2466 => x"25ffa438",
  2467 => x"800880e2",
  2468 => x"e0083180",
  2469 => x"e2b00c74",
  2470 => x"81078414",
  2471 => x"0c7551fe",
  2472 => x"973f8053",
  2473 => x"ff9039f6",
  2474 => x"3d0d7c7e",
  2475 => x"545b7280",
  2476 => x"2e828338",
  2477 => x"7a51fdff",
  2478 => x"3ff81384",
  2479 => x"110870fe",
  2480 => x"06701384",
  2481 => x"1108fc06",
  2482 => x"5d585954",
  2483 => x"5880e2f4",
  2484 => x"08752e82",
  2485 => x"de387884",
  2486 => x"160c8073",
  2487 => x"8106545a",
  2488 => x"727a2e81",
  2489 => x"d5387815",
  2490 => x"84110881",
  2491 => x"06515372",
  2492 => x"a0387817",
  2493 => x"577981e6",
  2494 => x"38881508",
  2495 => x"537280e2",
  2496 => x"f42e82f9",
  2497 => x"388c1508",
  2498 => x"708c150c",
  2499 => x"7388120c",
  2500 => x"56768107",
  2501 => x"84190c76",
  2502 => x"1877710c",
  2503 => x"53798191",
  2504 => x"3883ff77",
  2505 => x"2781c838",
  2506 => x"76892a77",
  2507 => x"832a5653",
  2508 => x"72802ebf",
  2509 => x"3876862a",
  2510 => x"b8055584",
  2511 => x"7327b438",
  2512 => x"80db1355",
  2513 => x"947327ab",
  2514 => x"38768c2a",
  2515 => x"80ee0555",
  2516 => x"80d47327",
  2517 => x"9e38768f",
  2518 => x"2a80f705",
  2519 => x"5582d473",
  2520 => x"27913876",
  2521 => x"922a80fc",
  2522 => x"05558ad4",
  2523 => x"73278438",
  2524 => x"80fe5574",
  2525 => x"10101080",
  2526 => x"e2ec0588",
  2527 => x"11085556",
  2528 => x"73762e82",
  2529 => x"b3388414",
  2530 => x"08fc0653",
  2531 => x"7673278d",
  2532 => x"38881408",
  2533 => x"5473762e",
  2534 => x"098106ea",
  2535 => x"388c1408",
  2536 => x"708c1a0c",
  2537 => x"74881a0c",
  2538 => x"7888120c",
  2539 => x"56778c15",
  2540 => x"0c7a51fc",
  2541 => x"833f8c3d",
  2542 => x"0d047708",
  2543 => x"78713159",
  2544 => x"77058819",
  2545 => x"08545772",
  2546 => x"80e2f42e",
  2547 => x"80e0388c",
  2548 => x"1808708c",
  2549 => x"150c7388",
  2550 => x"120c56fe",
  2551 => x"89398815",
  2552 => x"088c1608",
  2553 => x"708c130c",
  2554 => x"5788170c",
  2555 => x"fea33976",
  2556 => x"832a7054",
  2557 => x"55807524",
  2558 => x"81983872",
  2559 => x"822c8171",
  2560 => x"2b80e2f0",
  2561 => x"080780e2",
  2562 => x"ec0b8405",
  2563 => x"0c537410",
  2564 => x"101080e2",
  2565 => x"ec058811",
  2566 => x"08555675",
  2567 => x"8c190c73",
  2568 => x"88190c77",
  2569 => x"88170c77",
  2570 => x"8c150cff",
  2571 => x"8439815a",
  2572 => x"fdb43978",
  2573 => x"17738106",
  2574 => x"54577298",
  2575 => x"38770878",
  2576 => x"71315977",
  2577 => x"058c1908",
  2578 => x"881a0871",
  2579 => x"8c120c88",
  2580 => x"120c5757",
  2581 => x"76810784",
  2582 => x"190c7780",
  2583 => x"e2ec0b88",
  2584 => x"050c80e2",
  2585 => x"e8087726",
  2586 => x"fec73880",
  2587 => x"e2e40852",
  2588 => x"7a51fafd",
  2589 => x"3f7a51fa",
  2590 => x"bf3ffeba",
  2591 => x"3981788c",
  2592 => x"150c7888",
  2593 => x"150c738c",
  2594 => x"1a0c7388",
  2595 => x"1a0c5afd",
  2596 => x"80398315",
  2597 => x"70822c81",
  2598 => x"712b80e2",
  2599 => x"f0080780",
  2600 => x"e2ec0b84",
  2601 => x"050c5153",
  2602 => x"74101010",
  2603 => x"80e2ec05",
  2604 => x"88110855",
  2605 => x"56fee439",
  2606 => x"74538075",
  2607 => x"24a73872",
  2608 => x"822c8171",
  2609 => x"2b80e2f0",
  2610 => x"080780e2",
  2611 => x"ec0b8405",
  2612 => x"0c53758c",
  2613 => x"190c7388",
  2614 => x"190c7788",
  2615 => x"170c778c",
  2616 => x"150cfdcd",
  2617 => x"39831570",
  2618 => x"822c8171",
  2619 => x"2b80e2f0",
  2620 => x"080780e2",
  2621 => x"ec0b8405",
  2622 => x"0c5153d6",
  2623 => x"39810b80",
  2624 => x"0c04803d",
  2625 => x"0d72812e",
  2626 => x"8938800b",
  2627 => x"800c823d",
  2628 => x"0d047351",
  2629 => x"81843ffe",
  2630 => x"3d0d8180",
  2631 => x"8087e008",
  2632 => x"51708e38",
  2633 => x"81808087",
  2634 => x"ec708180",
  2635 => x"8087e00c",
  2636 => x"51707512",
  2637 => x"5252ff53",
  2638 => x"7087fb80",
  2639 => x"80268a38",
  2640 => x"70818080",
  2641 => x"87e00c71",
  2642 => x"5372800c",
  2643 => x"843d0d04",
  2644 => x"fd3d0d80",
  2645 => x"0b80db8c",
  2646 => x"08545472",
  2647 => x"812e9e38",
  2648 => x"73818080",
  2649 => x"87e40cff",
  2650 => x"b6b73fff",
  2651 => x"b5923f80",
  2652 => x"eaf45281",
  2653 => x"51d5ff3f",
  2654 => x"800851a4",
  2655 => x"3f728180",
  2656 => x"8087e40c",
  2657 => x"ffb69a3f",
  2658 => x"ffb4f53f",
  2659 => x"80eaf452",
  2660 => x"8151d5e2",
  2661 => x"3f800851",
  2662 => x"873f00ff",
  2663 => x"3900ff39",
  2664 => x"f73d0d7b",
  2665 => x"80dbb008",
  2666 => x"82c81108",
  2667 => x"5a545a77",
  2668 => x"802e80da",
  2669 => x"38818818",
  2670 => x"841908ff",
  2671 => x"0581712b",
  2672 => x"59555980",
  2673 => x"742480ea",
  2674 => x"38807424",
  2675 => x"b5387382",
  2676 => x"2b781188",
  2677 => x"05565681",
  2678 => x"80190877",
  2679 => x"06537280",
  2680 => x"2eb63878",
  2681 => x"16700853",
  2682 => x"53795174",
  2683 => x"0853722d",
  2684 => x"ff14fc17",
  2685 => x"fc177981",
  2686 => x"2c5a5757",
  2687 => x"54738025",
  2688 => x"d6387708",
  2689 => x"5877ffad",
  2690 => x"3880dbb0",
  2691 => x"0853bc13",
  2692 => x"08a53879",
  2693 => x"51ff833f",
  2694 => x"74085372",
  2695 => x"2dff14fc",
  2696 => x"17fc1779",
  2697 => x"812c5a57",
  2698 => x"57547380",
  2699 => x"25ffa838",
  2700 => x"d1398057",
  2701 => x"ff933972",
  2702 => x"51bc1308",
  2703 => x"53722d79",
  2704 => x"51fed73f",
  2705 => x"ff3d0d80",
  2706 => x"eafc0bfc",
  2707 => x"05700852",
  2708 => x"5270ff2e",
  2709 => x"9138702d",
  2710 => x"fc127008",
  2711 => x"525270ff",
  2712 => x"2e098106",
  2713 => x"f138833d",
  2714 => x"0d0404ff",
  2715 => x"b5ad3f04",
  2716 => x"00000040",
  2717 => x"3e200000",
  2718 => x"636f6d6d",
  2719 => x"616e6420",
  2720 => x"6e6f7420",
  2721 => x"666f756e",
  2722 => x"642e0a00",
  2723 => x"73657400",
  2724 => x"73657420",
  2725 => x"3c636861",
  2726 => x"6e6e656c",
  2727 => x"3e203c77",
  2728 => x"6169743e",
  2729 => x"203c6f6e",
  2730 => x"3e203c6f",
  2731 => x"66663e20",
  2732 => x"3c636f75",
  2733 => x"6e743e00",
  2734 => x"73746174",
  2735 => x"75730000",
  2736 => x"67657420",
  2737 => x"616c6c20",
  2738 => x"6368616e",
  2739 => x"6e656c20",
  2740 => x"73657474",
  2741 => x"696e6773",
  2742 => x"00000000",
  2743 => x"72756e00",
  2744 => x"67656e65",
  2745 => x"72617465",
  2746 => x"20736967",
  2747 => x"6e616c20",
  2748 => x"6f6e2061",
  2749 => x"6c6c2063",
  2750 => x"68616e6e",
  2751 => x"656c7300",
  2752 => x"73746f70",
  2753 => x"00000000",
  2754 => x"73746f70",
  2755 => x"20616c6c",
  2756 => x"20636861",
  2757 => x"6e6e656c",
  2758 => x"73000000",
  2759 => x"636c6561",
  2760 => x"72000000",
  2761 => x"636c6561",
  2762 => x"72207363",
  2763 => x"7265656e",
  2764 => x"00000000",
  2765 => x"68656c70",
  2766 => x"00000000",
  2767 => x"73757070",
  2768 => x"6f727465",
  2769 => x"6420636f",
  2770 => x"6d6d616e",
  2771 => x"64733a0a",
  2772 => x"0a000000",
  2773 => x"202d2000",
  2774 => x"30780000",
  2775 => x"0a307800",
  2776 => x"203a2000",
  2777 => x"6368616e",
  2778 => x"6e656c20",
  2779 => x"00000000",
  2780 => x"09202073",
  2781 => x"74617475",
  2782 => x"733a2000",
  2783 => x"09202020",
  2784 => x"20776169",
  2785 => x"743a2000",
  2786 => x"09202020",
  2787 => x"2020206f",
  2788 => x"6e3a2000",
  2789 => x"09202020",
  2790 => x"20206f66",
  2791 => x"663a2000",
  2792 => x"09202020",
  2793 => x"636f756e",
  2794 => x"743a2000",
  2795 => x"4572726f",
  2796 => x"723a2077",
  2797 => x"726f6e67",
  2798 => x"20636861",
  2799 => x"6e6e656c",
  2800 => x"206e756d",
  2801 => x"62657220",
  2802 => x"28000000",
  2803 => x"290a0000",
  2804 => x"68656170",
  2805 => x"20707472",
  2806 => x"3a200000",
  2807 => x"66726565",
  2808 => x"206d656d",
  2809 => x"3a200000",
  2810 => x"656e643a",
  2811 => x"20202020",
  2812 => x"20200000",
  2813 => x"0a0a0000",
  2814 => x"63656e74",
  2815 => x"72616c20",
  2816 => x"74726967",
  2817 => x"67657220",
  2818 => x"67656e65",
  2819 => x"7261746f",
  2820 => x"72200000",
  2821 => x"286f6e20",
  2822 => x"73696d29",
  2823 => x"0a000000",
  2824 => x"0a636f6d",
  2825 => x"70696c65",
  2826 => x"643a204d",
  2827 => x"61722032",
  2828 => x"35203230",
  2829 => x"31312020",
  2830 => x"31343a34",
  2831 => x"313a3230",
  2832 => x"0a000000",
  2833 => x"63656e74",
  2834 => x"72616c20",
  2835 => x"20747269",
  2836 => x"67676572",
  2837 => x"00000000",
  2838 => x"67656e65",
  2839 => x"7261746f",
  2840 => x"72000000",
  2841 => x"00202020",
  2842 => x"20202020",
  2843 => x"20202828",
  2844 => x"28282820",
  2845 => x"20202020",
  2846 => x"20202020",
  2847 => x"20202020",
  2848 => x"20202020",
  2849 => x"20881010",
  2850 => x"10101010",
  2851 => x"10101010",
  2852 => x"10101010",
  2853 => x"10040404",
  2854 => x"04040404",
  2855 => x"04040410",
  2856 => x"10101010",
  2857 => x"10104141",
  2858 => x"41414141",
  2859 => x"01010101",
  2860 => x"01010101",
  2861 => x"01010101",
  2862 => x"01010101",
  2863 => x"01010101",
  2864 => x"10101010",
  2865 => x"10104242",
  2866 => x"42424242",
  2867 => x"02020202",
  2868 => x"02020202",
  2869 => x"02020202",
  2870 => x"02020202",
  2871 => x"02020202",
  2872 => x"10101010",
  2873 => x"20000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000000",
  2884 => x"00000000",
  2885 => x"00000000",
  2886 => x"00000000",
  2887 => x"00000000",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000000",
  2895 => x"00000000",
  2896 => x"00000000",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000000",
  2900 => x"00000000",
  2901 => x"00000000",
  2902 => x"00000000",
  2903 => x"00000000",
  2904 => x"00000000",
  2905 => x"00000000",
  2906 => x"43000000",
  2907 => x"64756d6d",
  2908 => x"792e6578",
  2909 => x"65000000",
  2910 => x"00ffffff",
  2911 => x"ff00ffff",
  2912 => x"ffff00ff",
  2913 => x"ffffff00",
  2914 => x"00000000",
  2915 => x"00000000",
  2916 => x"00000000",
  2917 => x"00003584",
  2918 => x"80000800",
  2919 => x"80000600",
  2920 => x"80000400",
  2921 => x"80000200",
  2922 => x"80000100",
  2923 => x"80000000",
  2924 => x"00002db4",
  2925 => x"00000000",
  2926 => x"0000301c",
  2927 => x"00003078",
  2928 => x"000030d4",
  2929 => x"00000000",
  2930 => x"00000000",
  2931 => x"00000000",
  2932 => x"00000000",
  2933 => x"00000000",
  2934 => x"00000000",
  2935 => x"00000000",
  2936 => x"00000000",
  2937 => x"00000000",
  2938 => x"00002d68",
  2939 => x"00000000",
  2940 => x"00000000",
  2941 => x"00000000",
  2942 => x"00000000",
  2943 => x"00000000",
  2944 => x"00000000",
  2945 => x"00000000",
  2946 => x"00000000",
  2947 => x"00000000",
  2948 => x"00000000",
  2949 => x"00000000",
  2950 => x"00000000",
  2951 => x"00000000",
  2952 => x"00000000",
  2953 => x"00000000",
  2954 => x"00000000",
  2955 => x"00000000",
  2956 => x"00000000",
  2957 => x"00000000",
  2958 => x"00000000",
  2959 => x"00000000",
  2960 => x"00000000",
  2961 => x"00000000",
  2962 => x"00000000",
  2963 => x"00000000",
  2964 => x"00000000",
  2965 => x"00000000",
  2966 => x"00000000",
  2967 => x"00000001",
  2968 => x"330eabcd",
  2969 => x"1234e66d",
  2970 => x"deec0005",
  2971 => x"000b0000",
  2972 => x"00000000",
  2973 => x"00000000",
  2974 => x"00000000",
  2975 => x"00000000",
  2976 => x"00000000",
  2977 => x"00000000",
  2978 => x"00000000",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00000000",
  2983 => x"00000000",
  2984 => x"00000000",
  2985 => x"00000000",
  2986 => x"00000000",
  2987 => x"00000000",
  2988 => x"00000000",
  2989 => x"00000000",
  2990 => x"00000000",
  2991 => x"00000000",
  2992 => x"00000000",
  2993 => x"00000000",
  2994 => x"00000000",
  2995 => x"00000000",
  2996 => x"00000000",
  2997 => x"00000000",
  2998 => x"00000000",
  2999 => x"00000000",
  3000 => x"00000000",
  3001 => x"00000000",
  3002 => x"00000000",
  3003 => x"00000000",
  3004 => x"00000000",
  3005 => x"00000000",
  3006 => x"00000000",
  3007 => x"00000000",
  3008 => x"00000000",
  3009 => x"00000000",
  3010 => x"00000000",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"00000000",
  3015 => x"00000000",
  3016 => x"00000000",
  3017 => x"00000000",
  3018 => x"00000000",
  3019 => x"00000000",
  3020 => x"00000000",
  3021 => x"00000000",
  3022 => x"00000000",
  3023 => x"00000000",
  3024 => x"00000000",
  3025 => x"00000000",
  3026 => x"00000000",
  3027 => x"00000000",
  3028 => x"00000000",
  3029 => x"00000000",
  3030 => x"00000000",
  3031 => x"00000000",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"00000000",
  3041 => x"00000000",
  3042 => x"00000000",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000000",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00000000",
  3050 => x"00000000",
  3051 => x"00000000",
  3052 => x"00000000",
  3053 => x"00000000",
  3054 => x"00000000",
  3055 => x"00000000",
  3056 => x"00000000",
  3057 => x"00000000",
  3058 => x"00000000",
  3059 => x"00000000",
  3060 => x"00000000",
  3061 => x"00000000",
  3062 => x"00000000",
  3063 => x"00000000",
  3064 => x"00000000",
  3065 => x"00000000",
  3066 => x"00000000",
  3067 => x"00000000",
  3068 => x"00000000",
  3069 => x"00000000",
  3070 => x"00000000",
  3071 => x"00000000",
  3072 => x"00000000",
  3073 => x"00000000",
  3074 => x"00000000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000000",
  3084 => x"00000000",
  3085 => x"00000000",
  3086 => x"00000000",
  3087 => x"00000000",
  3088 => x"00000000",
  3089 => x"00000000",
  3090 => x"00000000",
  3091 => x"00000000",
  3092 => x"00000000",
  3093 => x"00000000",
  3094 => x"00000000",
  3095 => x"00000000",
  3096 => x"00000000",
  3097 => x"00000000",
  3098 => x"00000000",
  3099 => x"00000000",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00000000",
  3103 => x"00000000",
  3104 => x"00000000",
  3105 => x"00000000",
  3106 => x"00000000",
  3107 => x"00000000",
  3108 => x"00000000",
  3109 => x"00000000",
  3110 => x"00000000",
  3111 => x"00000000",
  3112 => x"00000000",
  3113 => x"00000000",
  3114 => x"00000000",
  3115 => x"00000000",
  3116 => x"00000000",
  3117 => x"00000000",
  3118 => x"00000000",
  3119 => x"00000000",
  3120 => x"00000000",
  3121 => x"00000000",
  3122 => x"00000000",
  3123 => x"00000000",
  3124 => x"00000000",
  3125 => x"00000000",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000000",
  3151 => x"00000000",
  3152 => x"00000000",
  3153 => x"00000000",
  3154 => x"00000000",
  3155 => x"00000000",
  3156 => x"00000000",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"ffffffff",
  3161 => x"00000000",
  3162 => x"00020000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"0000316c",
  3166 => x"0000316c",
  3167 => x"00003174",
  3168 => x"00003174",
  3169 => x"0000317c",
  3170 => x"0000317c",
  3171 => x"00003184",
  3172 => x"00003184",
  3173 => x"0000318c",
  3174 => x"0000318c",
  3175 => x"00003194",
  3176 => x"00003194",
  3177 => x"0000319c",
  3178 => x"0000319c",
  3179 => x"000031a4",
  3180 => x"000031a4",
  3181 => x"000031ac",
  3182 => x"000031ac",
  3183 => x"000031b4",
  3184 => x"000031b4",
  3185 => x"000031bc",
  3186 => x"000031bc",
  3187 => x"000031c4",
  3188 => x"000031c4",
  3189 => x"000031cc",
  3190 => x"000031cc",
  3191 => x"000031d4",
  3192 => x"000031d4",
  3193 => x"000031dc",
  3194 => x"000031dc",
  3195 => x"000031e4",
  3196 => x"000031e4",
  3197 => x"000031ec",
  3198 => x"000031ec",
  3199 => x"000031f4",
  3200 => x"000031f4",
  3201 => x"000031fc",
  3202 => x"000031fc",
  3203 => x"00003204",
  3204 => x"00003204",
  3205 => x"0000320c",
  3206 => x"0000320c",
  3207 => x"00003214",
  3208 => x"00003214",
  3209 => x"0000321c",
  3210 => x"0000321c",
  3211 => x"00003224",
  3212 => x"00003224",
  3213 => x"0000322c",
  3214 => x"0000322c",
  3215 => x"00003234",
  3216 => x"00003234",
  3217 => x"0000323c",
  3218 => x"0000323c",
  3219 => x"00003244",
  3220 => x"00003244",
  3221 => x"0000324c",
  3222 => x"0000324c",
  3223 => x"00003254",
  3224 => x"00003254",
  3225 => x"0000325c",
  3226 => x"0000325c",
  3227 => x"00003264",
  3228 => x"00003264",
  3229 => x"0000326c",
  3230 => x"0000326c",
  3231 => x"00003274",
  3232 => x"00003274",
  3233 => x"0000327c",
  3234 => x"0000327c",
  3235 => x"00003284",
  3236 => x"00003284",
  3237 => x"0000328c",
  3238 => x"0000328c",
  3239 => x"00003294",
  3240 => x"00003294",
  3241 => x"0000329c",
  3242 => x"0000329c",
  3243 => x"000032a4",
  3244 => x"000032a4",
  3245 => x"000032ac",
  3246 => x"000032ac",
  3247 => x"000032b4",
  3248 => x"000032b4",
  3249 => x"000032bc",
  3250 => x"000032bc",
  3251 => x"000032c4",
  3252 => x"000032c4",
  3253 => x"000032cc",
  3254 => x"000032cc",
  3255 => x"000032d4",
  3256 => x"000032d4",
  3257 => x"000032dc",
  3258 => x"000032dc",
  3259 => x"000032e4",
  3260 => x"000032e4",
  3261 => x"000032ec",
  3262 => x"000032ec",
  3263 => x"000032f4",
  3264 => x"000032f4",
  3265 => x"000032fc",
  3266 => x"000032fc",
  3267 => x"00003304",
  3268 => x"00003304",
  3269 => x"0000330c",
  3270 => x"0000330c",
  3271 => x"00003314",
  3272 => x"00003314",
  3273 => x"0000331c",
  3274 => x"0000331c",
  3275 => x"00003324",
  3276 => x"00003324",
  3277 => x"0000332c",
  3278 => x"0000332c",
  3279 => x"00003334",
  3280 => x"00003334",
  3281 => x"0000333c",
  3282 => x"0000333c",
  3283 => x"00003344",
  3284 => x"00003344",
  3285 => x"0000334c",
  3286 => x"0000334c",
  3287 => x"00003354",
  3288 => x"00003354",
  3289 => x"0000335c",
  3290 => x"0000335c",
  3291 => x"00003364",
  3292 => x"00003364",
  3293 => x"0000336c",
  3294 => x"0000336c",
  3295 => x"00003374",
  3296 => x"00003374",
  3297 => x"0000337c",
  3298 => x"0000337c",
  3299 => x"00003384",
  3300 => x"00003384",
  3301 => x"0000338c",
  3302 => x"0000338c",
  3303 => x"00003394",
  3304 => x"00003394",
  3305 => x"0000339c",
  3306 => x"0000339c",
  3307 => x"000033a4",
  3308 => x"000033a4",
  3309 => x"000033ac",
  3310 => x"000033ac",
  3311 => x"000033b4",
  3312 => x"000033b4",
  3313 => x"000033bc",
  3314 => x"000033bc",
  3315 => x"000033c4",
  3316 => x"000033c4",
  3317 => x"000033cc",
  3318 => x"000033cc",
  3319 => x"000033d4",
  3320 => x"000033d4",
  3321 => x"000033dc",
  3322 => x"000033dc",
  3323 => x"000033e4",
  3324 => x"000033e4",
  3325 => x"000033ec",
  3326 => x"000033ec",
  3327 => x"000033f4",
  3328 => x"000033f4",
  3329 => x"000033fc",
  3330 => x"000033fc",
  3331 => x"00003404",
  3332 => x"00003404",
  3333 => x"0000340c",
  3334 => x"0000340c",
  3335 => x"00003414",
  3336 => x"00003414",
  3337 => x"0000341c",
  3338 => x"0000341c",
  3339 => x"00003424",
  3340 => x"00003424",
  3341 => x"0000342c",
  3342 => x"0000342c",
  3343 => x"00003434",
  3344 => x"00003434",
  3345 => x"0000343c",
  3346 => x"0000343c",
  3347 => x"00003444",
  3348 => x"00003444",
  3349 => x"0000344c",
  3350 => x"0000344c",
  3351 => x"00003454",
  3352 => x"00003454",
  3353 => x"0000345c",
  3354 => x"0000345c",
  3355 => x"00003464",
  3356 => x"00003464",
  3357 => x"0000346c",
  3358 => x"0000346c",
  3359 => x"00003474",
  3360 => x"00003474",
  3361 => x"0000347c",
  3362 => x"0000347c",
  3363 => x"00003484",
  3364 => x"00003484",
  3365 => x"0000348c",
  3366 => x"0000348c",
  3367 => x"00003494",
  3368 => x"00003494",
  3369 => x"0000349c",
  3370 => x"0000349c",
  3371 => x"000034a4",
  3372 => x"000034a4",
  3373 => x"000034ac",
  3374 => x"000034ac",
  3375 => x"000034b4",
  3376 => x"000034b4",
  3377 => x"000034bc",
  3378 => x"000034bc",
  3379 => x"000034c4",
  3380 => x"000034c4",
  3381 => x"000034cc",
  3382 => x"000034cc",
  3383 => x"000034d4",
  3384 => x"000034d4",
  3385 => x"000034dc",
  3386 => x"000034dc",
  3387 => x"000034e4",
  3388 => x"000034e4",
  3389 => x"000034ec",
  3390 => x"000034ec",
  3391 => x"000034f4",
  3392 => x"000034f4",
  3393 => x"000034fc",
  3394 => x"000034fc",
  3395 => x"00003504",
  3396 => x"00003504",
  3397 => x"0000350c",
  3398 => x"0000350c",
  3399 => x"00003514",
  3400 => x"00003514",
  3401 => x"0000351c",
  3402 => x"0000351c",
  3403 => x"00003524",
  3404 => x"00003524",
  3405 => x"0000352c",
  3406 => x"0000352c",
  3407 => x"00003534",
  3408 => x"00003534",
  3409 => x"0000353c",
  3410 => x"0000353c",
  3411 => x"00003544",
  3412 => x"00003544",
  3413 => x"0000354c",
  3414 => x"0000354c",
  3415 => x"00003554",
  3416 => x"00003554",
  3417 => x"0000355c",
  3418 => x"0000355c",
  3419 => x"00003564",
  3420 => x"00003564",
  3421 => x"00002d6c",
  3422 => x"ffffffff",
  3423 => x"00000000",
  3424 => x"ffffffff",
  3425 => x"00000000",
  3426 => x"00000000",
	others => x"aaaaaaaa" -- mask for mem check
	--others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
