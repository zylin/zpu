-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80dee40c",
     3 => x"3a0b0b80",
     4 => x"cbdb0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b91bf2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80de",
   162 => x"d0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0ba9",
   171 => x"922d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0baa",
   179 => x"c42d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80dee00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"c5c23f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80dee008",
   281 => x"802ea438",
   282 => x"80dee408",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80ee",
   286 => x"e80c82a0",
   287 => x"800b80ee",
   288 => x"ec0c8290",
   289 => x"800b80ee",
   290 => x"f00c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"eee80cf8",
   294 => x"80808280",
   295 => x"0b80eeec",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"eef00c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80eee80c",
   302 => x"80c0a880",
   303 => x"940b80ee",
   304 => x"ec0c0b0b",
   305 => x"80cdf40b",
   306 => x"80eef00c",
   307 => x"04ff3d0d",
   308 => x"80eef433",
   309 => x"5170a738",
   310 => x"80deec08",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"deec0c70",
   315 => x"2d80deec",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80ee",
   319 => x"f434833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80eee408",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"eee4510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404fd3d",
   333 => x"0d80def8",
   334 => x"08881108",
   335 => x"83de8007",
   336 => x"88120c84",
   337 => x"1108fca1",
   338 => x"ff068412",
   339 => x"0c538f51",
   340 => x"9ae03f80",
   341 => x"def80884",
   342 => x"1108e1ff",
   343 => x"0684120c",
   344 => x"84110886",
   345 => x"80078412",
   346 => x"0c841108",
   347 => x"80c08007",
   348 => x"84120c53",
   349 => x"81519a95",
   350 => x"3f80def8",
   351 => x"08841108",
   352 => x"ffbfff06",
   353 => x"84120c53",
   354 => x"85519aa6",
   355 => x"3f80def8",
   356 => x"08841108",
   357 => x"80c08007",
   358 => x"84120c53",
   359 => x"815199ed",
   360 => x"3f80def8",
   361 => x"08841108",
   362 => x"ffbfff06",
   363 => x"84120c53",
   364 => x"815199fe",
   365 => x"3f80def8",
   366 => x"08841108",
   367 => x"80c08007",
   368 => x"84120c53",
   369 => x"815199c5",
   370 => x"3f80def8",
   371 => x"08841108",
   372 => x"ffbfff06",
   373 => x"84120c53",
   374 => x"815199d6",
   375 => x"3f80def8",
   376 => x"08841108",
   377 => x"e1ff0684",
   378 => x"120c5384",
   379 => x"800b8414",
   380 => x"08707207",
   381 => x"84160c53",
   382 => x"84140870",
   383 => x"80c08007",
   384 => x"84160c53",
   385 => x"54815199",
   386 => x"843f80de",
   387 => x"f8088411",
   388 => x"0870ffbf",
   389 => x"ff068413",
   390 => x"0c535385",
   391 => x"5199933f",
   392 => x"80def808",
   393 => x"84110870",
   394 => x"feffff06",
   395 => x"84130c53",
   396 => x"84110870",
   397 => x"e1ff0684",
   398 => x"130c5384",
   399 => x"11087076",
   400 => x"0784130c",
   401 => x"53841108",
   402 => x"80c08007",
   403 => x"84120c53",
   404 => x"815198b9",
   405 => x"3f80def8",
   406 => x"08841108",
   407 => x"ffbfff06",
   408 => x"84120c84",
   409 => x"1108e1ff",
   410 => x"0684120c",
   411 => x"84110890",
   412 => x"80078412",
   413 => x"0c841108",
   414 => x"80c08007",
   415 => x"84120c54",
   416 => x"81519889",
   417 => x"3f80def8",
   418 => x"08841108",
   419 => x"ffbfff06",
   420 => x"84120c54",
   421 => x"aa5197f5",
   422 => x"3f80def8",
   423 => x"08841108",
   424 => x"feffff06",
   425 => x"84120c84",
   426 => x"1108e1ff",
   427 => x"0684120c",
   428 => x"84110884",
   429 => x"120c8411",
   430 => x"0880c080",
   431 => x"0784120c",
   432 => x"54815197",
   433 => x"c83f80de",
   434 => x"f8088411",
   435 => x"08ffbfff",
   436 => x"0684120c",
   437 => x"841108e1",
   438 => x"ff068412",
   439 => x"0c841108",
   440 => x"98800784",
   441 => x"120c8411",
   442 => x"0880c080",
   443 => x"0784120c",
   444 => x"54815197",
   445 => x"983f80de",
   446 => x"f8088411",
   447 => x"08ffbfff",
   448 => x"0684120c",
   449 => x"54aa5197",
   450 => x"843f80de",
   451 => x"f8088411",
   452 => x"08feffff",
   453 => x"0684120c",
   454 => x"841108e1",
   455 => x"ff068412",
   456 => x"0c841108",
   457 => x"84120c84",
   458 => x"110880c0",
   459 => x"80078412",
   460 => x"0c548151",
   461 => x"96d73f80",
   462 => x"def80884",
   463 => x"1108ffbf",
   464 => x"ff068412",
   465 => x"0c841108",
   466 => x"e1ff0684",
   467 => x"120c8411",
   468 => x"088c8007",
   469 => x"84120c84",
   470 => x"110880c0",
   471 => x"80078412",
   472 => x"0c548151",
   473 => x"96a73f80",
   474 => x"def80884",
   475 => x"1108ffbf",
   476 => x"ff068412",
   477 => x"0c54aa51",
   478 => x"96933f81",
   479 => x"0b80def8",
   480 => x"08841108",
   481 => x"70feffff",
   482 => x"0684130c",
   483 => x"54841108",
   484 => x"70e1ff06",
   485 => x"84130c54",
   486 => x"84110884",
   487 => x"120c8411",
   488 => x"087080c0",
   489 => x"80078413",
   490 => x"0c545470",
   491 => x"525495dd",
   492 => x"3f80def8",
   493 => x"08841108",
   494 => x"70ffbfff",
   495 => x"0684130c",
   496 => x"53841108",
   497 => x"70e1ff06",
   498 => x"84130c53",
   499 => x"84110870",
   500 => x"82800784",
   501 => x"130c5384",
   502 => x"11087080",
   503 => x"c0800784",
   504 => x"130c5353",
   505 => x"735195a5",
   506 => x"3f80def8",
   507 => x"08841108",
   508 => x"ffbfff06",
   509 => x"84120c53",
   510 => x"aa519591",
   511 => x"3f825195",
   512 => x"b13f853d",
   513 => x"0d04fb3d",
   514 => x"0d777033",
   515 => x"53567180",
   516 => x"2e818f38",
   517 => x"71558116",
   518 => x"80def808",
   519 => x"84110881",
   520 => x"80800784",
   521 => x"120c8411",
   522 => x"08e1ff06",
   523 => x"84120c76",
   524 => x"842b9e80",
   525 => x"06841208",
   526 => x"70720784",
   527 => x"140c5584",
   528 => x"120880c0",
   529 => x"80078413",
   530 => x"0c565456",
   531 => x"815194bd",
   532 => x"3f80def8",
   533 => x"08841108",
   534 => x"ffbfff06",
   535 => x"84120c84",
   536 => x"1108e1ff",
   537 => x"0684120c",
   538 => x"75882b9e",
   539 => x"80068412",
   540 => x"08710784",
   541 => x"130c8412",
   542 => x"0880c080",
   543 => x"0784130c",
   544 => x"55538151",
   545 => x"94873f80",
   546 => x"def80884",
   547 => x"1108ffbf",
   548 => x"ff068412",
   549 => x"0c53ae51",
   550 => x"93f33f75",
   551 => x"335574fe",
   552 => x"f538873d",
   553 => x"0d04ff3d",
   554 => x"0d028f05",
   555 => x"33705252",
   556 => x"959f3f71",
   557 => x"51968e3f",
   558 => x"71800c83",
   559 => x"3d0d04ff",
   560 => x"3d0d800b",
   561 => x"80eefc08",
   562 => x"52527072",
   563 => x"2e098106",
   564 => x"83388152",
   565 => x"7180eefc",
   566 => x"0c80df80",
   567 => x"08528180",
   568 => x"0b8c130c",
   569 => x"833d0d04",
   570 => x"fa3d0d02",
   571 => x"a3053356",
   572 => x"758d2e80",
   573 => x"f3387588",
   574 => x"32703077",
   575 => x"80ff3270",
   576 => x"30728025",
   577 => x"71802507",
   578 => x"54515658",
   579 => x"55749438",
   580 => x"9f76278b",
   581 => x"3880f584",
   582 => x"33559e75",
   583 => x"27ae3888",
   584 => x"3d0d0480",
   585 => x"f5843356",
   586 => x"75802ef3",
   587 => x"38885190",
   588 => x"fd3fa051",
   589 => x"90f83f88",
   590 => x"5190f33f",
   591 => x"80f58433",
   592 => x"ff055776",
   593 => x"80f58434",
   594 => x"883d0d04",
   595 => x"755190de",
   596 => x"3f80f584",
   597 => x"33811155",
   598 => x"577380f5",
   599 => x"84347580",
   600 => x"f4e01834",
   601 => x"883d0d04",
   602 => x"8a5190c2",
   603 => x"3f80f584",
   604 => x"33811156",
   605 => x"547480f5",
   606 => x"8434800b",
   607 => x"80f4e015",
   608 => x"34805680",
   609 => x"0b80f4e0",
   610 => x"17335654",
   611 => x"74a02e83",
   612 => x"38815474",
   613 => x"802e9038",
   614 => x"73802e8b",
   615 => x"38811670",
   616 => x"81ff0657",
   617 => x"57dd3975",
   618 => x"802ebf38",
   619 => x"800b80f5",
   620 => x"80335555",
   621 => x"747427ab",
   622 => x"38735774",
   623 => x"10101075",
   624 => x"10057654",
   625 => x"80f4e053",
   626 => x"80ef8005",
   627 => x"51a0a63f",
   628 => x"8008802e",
   629 => x"a6388115",
   630 => x"7081ff06",
   631 => x"56547675",
   632 => x"26d93880",
   633 => x"ce84518f",
   634 => x"df3f80ce",
   635 => x"80518fd8",
   636 => x"3f800b80",
   637 => x"f5843488",
   638 => x"3d0d0474",
   639 => x"101080f4",
   640 => x"a0057008",
   641 => x"80f5880c",
   642 => x"56800b80",
   643 => x"f58434e7",
   644 => x"39fd3d0d",
   645 => x"8a518f96",
   646 => x"3f800b80",
   647 => x"f5843480",
   648 => x"0b80f580",
   649 => x"34800b80",
   650 => x"f5880c80",
   651 => x"ce985280",
   652 => x"ef80519d",
   653 => x"f43f80ce",
   654 => x"9c5280f5",
   655 => x"803370a0",
   656 => x"2980f0a0",
   657 => x"0552549d",
   658 => x"e03f80f5",
   659 => x"80337010",
   660 => x"1080f4a0",
   661 => x"0599c871",
   662 => x"0c548105",
   663 => x"537280f5",
   664 => x"803480ce",
   665 => x"a4527281",
   666 => x"ff06708a",
   667 => x"2980ef80",
   668 => x"0552539d",
   669 => x"b43f80ce",
   670 => x"ac5280f5",
   671 => x"803370a0",
   672 => x"2980f0a0",
   673 => x"0552549d",
   674 => x"a03f80f5",
   675 => x"80337010",
   676 => x"1080f4a0",
   677 => x"059d8a71",
   678 => x"0c548105",
   679 => x"537280f5",
   680 => x"803480cf",
   681 => x"d8527281",
   682 => x"ff06708a",
   683 => x"2980ef80",
   684 => x"0552539c",
   685 => x"f43f80ce",
   686 => x"b85280f5",
   687 => x"803370a0",
   688 => x"2980f0a0",
   689 => x"0552549c",
   690 => x"e03f80f5",
   691 => x"80337010",
   692 => x"1080f4a0",
   693 => x"0599c871",
   694 => x"0c548105",
   695 => x"537280f5",
   696 => x"803480ce",
   697 => x"c8527281",
   698 => x"ff06708a",
   699 => x"2980ef80",
   700 => x"0552539c",
   701 => x"b43f80ce",
   702 => x"d05280f5",
   703 => x"803370a0",
   704 => x"2980f0a0",
   705 => x"0552549c",
   706 => x"a03f80f5",
   707 => x"80337010",
   708 => x"1080f4a0",
   709 => x"059fda71",
   710 => x"0c548105",
   711 => x"537280f5",
   712 => x"803480ce",
   713 => x"e0527281",
   714 => x"ff06708a",
   715 => x"2980ef80",
   716 => x"0552539b",
   717 => x"f43f80ce",
   718 => x"e45280f5",
   719 => x"803370a0",
   720 => x"2980f0a0",
   721 => x"0552549b",
   722 => x"e03f80f5",
   723 => x"80337010",
   724 => x"1080f4a0",
   725 => x"059fe671",
   726 => x"0c548105",
   727 => x"537280f5",
   728 => x"803480ce",
   729 => x"f4527281",
   730 => x"ff06708a",
   731 => x"2980ef80",
   732 => x"0552539b",
   733 => x"b43f80dc",
   734 => x"885280f5",
   735 => x"803370a0",
   736 => x"2980f0a0",
   737 => x"0552549b",
   738 => x"a03f80f5",
   739 => x"80337010",
   740 => x"1080f4a0",
   741 => x"0598b271",
   742 => x"0c548105",
   743 => x"537280f5",
   744 => x"803480cd",
   745 => x"f8527281",
   746 => x"ff06708a",
   747 => x"2980ef80",
   748 => x"0552539a",
   749 => x"f43f80dc",
   750 => x"885280f5",
   751 => x"803370a0",
   752 => x"2980f0a0",
   753 => x"0552549a",
   754 => x"e03f80f5",
   755 => x"80337010",
   756 => x"1080f4a0",
   757 => x"0598b971",
   758 => x"0c548105",
   759 => x"537280f5",
   760 => x"803480ce",
   761 => x"80518be0",
   762 => x"3f810b80",
   763 => x"f58c348e",
   764 => x"ab3f8008",
   765 => x"ae3880f5",
   766 => x"88085372",
   767 => x"8d3880f5",
   768 => x"8c335372",
   769 => x"ea38853d",
   770 => x"0d04722d",
   771 => x"800b80f5",
   772 => x"880c80ce",
   773 => x"80518bb0",
   774 => x"3f80f58c",
   775 => x"335372cf",
   776 => x"38e4398e",
   777 => x"8a3f8008",
   778 => x"81ff0651",
   779 => x"f9ba3fff",
   780 => x"be39800b",
   781 => x"80f58c34",
   782 => x"04fc3d0d",
   783 => x"8a518aee",
   784 => x"3f80cefc",
   785 => x"518b813f",
   786 => x"800b80f5",
   787 => x"80335354",
   788 => x"73722780",
   789 => x"ea387310",
   790 => x"10107410",
   791 => x"0580ef80",
   792 => x"05705253",
   793 => x"8ae23f73",
   794 => x"852b80f0",
   795 => x"a0113353",
   796 => x"5571802e",
   797 => x"b2387251",
   798 => x"9a9c3f80",
   799 => x"0881ff06",
   800 => x"52718926",
   801 => x"9338a051",
   802 => x"8aa43f81",
   803 => x"127081ff",
   804 => x"06535389",
   805 => x"7227ef38",
   806 => x"80cf9451",
   807 => x"8aaa3f80",
   808 => x"f0a01551",
   809 => x"8aa23f8a",
   810 => x"518a833f",
   811 => x"81147081",
   812 => x"ff0680f5",
   813 => x"80335255",
   814 => x"52717426",
   815 => x"ff98388a",
   816 => x"5189eb3f",
   817 => x"863d0d04",
   818 => x"f63d0d80",
   819 => x"0b80f4e0",
   820 => x"3380f4e0",
   821 => x"59555673",
   822 => x"a02e0981",
   823 => x"06963881",
   824 => x"167081ff",
   825 => x"0680f4e0",
   826 => x"11703353",
   827 => x"59575473",
   828 => x"a02eec38",
   829 => x"80588077",
   830 => x"33565474",
   831 => x"742e8338",
   832 => x"815474a0",
   833 => x"2e81ce38",
   834 => x"7381fb38",
   835 => x"74a02e81",
   836 => x"c4388118",
   837 => x"7081ff06",
   838 => x"59548178",
   839 => x"26d83890",
   840 => x"538c3dfc",
   841 => x"05527651",
   842 => x"9e9a3f80",
   843 => x"0859800b",
   844 => x"80f4e033",
   845 => x"80f4e059",
   846 => x"555673a0",
   847 => x"2e098106",
   848 => x"96388116",
   849 => x"7081ff06",
   850 => x"80f4e011",
   851 => x"70335759",
   852 => x"575873a0",
   853 => x"2eec3880",
   854 => x"58807733",
   855 => x"56547474",
   856 => x"2e833881",
   857 => x"5474a02e",
   858 => x"81ac3873",
   859 => x"828c3874",
   860 => x"a02e81a2",
   861 => x"38811870",
   862 => x"81ff0659",
   863 => x"55827826",
   864 => x"d8389053",
   865 => x"8c3df805",
   866 => x"5276519d",
   867 => x"b73f8008",
   868 => x"57800883",
   869 => x"38905778",
   870 => x"fc065580",
   871 => x"56757727",
   872 => x"ab387583",
   873 => x"06597880",
   874 => x"2e819c38",
   875 => x"80d1d851",
   876 => x"88963f74",
   877 => x"70840556",
   878 => x"0852a051",
   879 => x"88ad3fa0",
   880 => x"5187eb3f",
   881 => x"81165676",
   882 => x"7626d738",
   883 => x"8a5187de",
   884 => x"3f8c3d0d",
   885 => x"04811670",
   886 => x"81ff0680",
   887 => x"f4e01170",
   888 => x"335c5257",
   889 => x"5778a02e",
   890 => x"098106fe",
   891 => x"a5388116",
   892 => x"7081ff06",
   893 => x"80f4e011",
   894 => x"70335c52",
   895 => x"575778a0",
   896 => x"2ed338fe",
   897 => x"8d398116",
   898 => x"7081ff06",
   899 => x"80f4e011",
   900 => x"595755fd",
   901 => x"e1398116",
   902 => x"7081ff06",
   903 => x"80f4e011",
   904 => x"70335752",
   905 => x"575773a0",
   906 => x"2e098106",
   907 => x"fec73881",
   908 => x"167081ff",
   909 => x"0680f4e0",
   910 => x"11703357",
   911 => x"52575773",
   912 => x"a02ed338",
   913 => x"feaf3980",
   914 => x"cf985186",
   915 => x"fb3f7452",
   916 => x"a0518797",
   917 => x"3f80cf9c",
   918 => x"5186ed3f",
   919 => x"80d1d851",
   920 => x"86e63f74",
   921 => x"70840556",
   922 => x"0852a051",
   923 => x"86fd3fa0",
   924 => x"5186bb3f",
   925 => x"811656fe",
   926 => x"ce398116",
   927 => x"7081ff06",
   928 => x"80f4e011",
   929 => x"595755fd",
   930 => x"d039f63d",
   931 => x"0d800b80",
   932 => x"f4e03380",
   933 => x"f4e05955",
   934 => x"5673a02e",
   935 => x"09810696",
   936 => x"38811670",
   937 => x"81ff0680",
   938 => x"f4e01170",
   939 => x"33535957",
   940 => x"5473a02e",
   941 => x"ec388058",
   942 => x"80773356",
   943 => x"5474742e",
   944 => x"83388154",
   945 => x"74a02e81",
   946 => x"8f387381",
   947 => x"bc3874a0",
   948 => x"2e818538",
   949 => x"81187081",
   950 => x"ff065954",
   951 => x"817826d8",
   952 => x"3890538c",
   953 => x"3dfc0552",
   954 => x"76519ad8",
   955 => x"3f800859",
   956 => x"800b80f4",
   957 => x"e03380f4",
   958 => x"e0595556",
   959 => x"73a02e09",
   960 => x"81069638",
   961 => x"81167081",
   962 => x"ff0680f4",
   963 => x"e0117033",
   964 => x"57595758",
   965 => x"73a02eec",
   966 => x"38805880",
   967 => x"77335654",
   968 => x"74742e83",
   969 => x"38815474",
   970 => x"a02e80ed",
   971 => x"3873819a",
   972 => x"3874a02e",
   973 => x"80e33881",
   974 => x"187081ff",
   975 => x"06595582",
   976 => x"7826d838",
   977 => x"90538c3d",
   978 => x"f8055276",
   979 => x"5199f53f",
   980 => x"8008790c",
   981 => x"8c3d0d04",
   982 => x"81167081",
   983 => x"ff0680f4",
   984 => x"e0117033",
   985 => x"5c525757",
   986 => x"78a02e09",
   987 => x"8106fee4",
   988 => x"38811670",
   989 => x"81ff0680",
   990 => x"f4e01170",
   991 => x"335c5257",
   992 => x"5778a02e",
   993 => x"d338fecc",
   994 => x"39811670",
   995 => x"81ff0680",
   996 => x"f4e01159",
   997 => x"5755fea0",
   998 => x"39811670",
   999 => x"81ff0680",
  1000 => x"f4e01170",
  1001 => x"33575257",
  1002 => x"5773a02e",
  1003 => x"098106ff",
  1004 => x"86388116",
  1005 => x"7081ff06",
  1006 => x"80f4e011",
  1007 => x"70335752",
  1008 => x"575773a0",
  1009 => x"2ed338fe",
  1010 => x"ee398116",
  1011 => x"7081ff06",
  1012 => x"80f4e011",
  1013 => x"595755fe",
  1014 => x"c239803d",
  1015 => x"0d8c5183",
  1016 => x"cd3f823d",
  1017 => x"0d04fc3d",
  1018 => x"0df881c0",
  1019 => x"8e80539f",
  1020 => x"0b80def8",
  1021 => x"087481ff",
  1022 => x"0684120c",
  1023 => x"80eefc08",
  1024 => x"54565471",
  1025 => x"802e9f38",
  1026 => x"729f2a73",
  1027 => x"10075373",
  1028 => x"802e9f38",
  1029 => x"ff147381",
  1030 => x"ff068417",
  1031 => x"0c80eefc",
  1032 => x"08535471",
  1033 => x"e338720a",
  1034 => x"100a739f",
  1035 => x"2b075373",
  1036 => x"e338863d",
  1037 => x"0d04f73d",
  1038 => x"0d80def8",
  1039 => x"08700881",
  1040 => x"0a0680ee",
  1041 => x"f80c5385",
  1042 => x"8c3f85ba",
  1043 => x"3fa39852",
  1044 => x"80eef808",
  1045 => x"843891a6",
  1046 => x"527180f5",
  1047 => x"900ce9d2",
  1048 => x"3f86be3f",
  1049 => x"80def008",
  1050 => x"53fac98e",
  1051 => x"868c730c",
  1052 => x"72087084",
  1053 => x"2a810651",
  1054 => x"5473f538",
  1055 => x"80def808",
  1056 => x"88110881",
  1057 => x"ff078812",
  1058 => x"0c7480ee",
  1059 => x"fc0c9411",
  1060 => x"08818007",
  1061 => x"94120c8c",
  1062 => x"11088180",
  1063 => x"078c120c",
  1064 => x"5380df80",
  1065 => x"08528180",
  1066 => x"0b80c013",
  1067 => x"0c80d294",
  1068 => x"5182953f",
  1069 => x"8c5181f6",
  1070 => x"3f80dbb8",
  1071 => x"5182893f",
  1072 => x"80eef808",
  1073 => x"802e81a0",
  1074 => x"3880dbc0",
  1075 => x"5181f93f",
  1076 => x"80dbcc51",
  1077 => x"eeb03ff2",
  1078 => x"b83ff881",
  1079 => x"c08e8053",
  1080 => x"9f0b80de",
  1081 => x"f8085555",
  1082 => x"80eef808",
  1083 => x"802e80d3",
  1084 => x"387281ff",
  1085 => x"0684150c",
  1086 => x"80eefc08",
  1087 => x"5271802e",
  1088 => x"9f38729f",
  1089 => x"2a731007",
  1090 => x"5374802e",
  1091 => x"9f38ff15",
  1092 => x"7381ff06",
  1093 => x"84160c80",
  1094 => x"eefc0853",
  1095 => x"5571e338",
  1096 => x"720a100a",
  1097 => x"739f2b07",
  1098 => x"5374e338",
  1099 => x"8ae03f72",
  1100 => x"0a100a73",
  1101 => x"9f2b0753",
  1102 => x"80fd5182",
  1103 => x"f53f80de",
  1104 => x"f8085472",
  1105 => x"81ff0684",
  1106 => x"150c80ee",
  1107 => x"fc085473",
  1108 => x"802edc38",
  1109 => x"729f2a73",
  1110 => x"10075380",
  1111 => x"fd5182d2",
  1112 => x"3f80def8",
  1113 => x"0854dc39",
  1114 => x"80dbd851",
  1115 => x"80da3f80",
  1116 => x"dbe85180",
  1117 => x"d33f80db",
  1118 => x"cc51ed8a",
  1119 => x"3ff1923f",
  1120 => x"f881c08e",
  1121 => x"80539f0b",
  1122 => x"80def808",
  1123 => x"555580ee",
  1124 => x"f808fedd",
  1125 => x"38ffac39",
  1126 => x"ff3d0d02",
  1127 => x"8f053380",
  1128 => x"def40852",
  1129 => x"710c800b",
  1130 => x"800c833d",
  1131 => x"0d04ff3d",
  1132 => x"0d028f05",
  1133 => x"335180f5",
  1134 => x"90085271",
  1135 => x"2d800881",
  1136 => x"ff06800c",
  1137 => x"833d0d04",
  1138 => x"fe3d0d74",
  1139 => x"70335353",
  1140 => x"71802e93",
  1141 => x"38811372",
  1142 => x"5280f590",
  1143 => x"08535371",
  1144 => x"2d723352",
  1145 => x"71ef3884",
  1146 => x"3d0d04f4",
  1147 => x"3d0d7f02",
  1148 => x"8405bb05",
  1149 => x"33555788",
  1150 => x"0b8c3d5a",
  1151 => x"5a895380",
  1152 => x"dcb05278",
  1153 => x"5189943f",
  1154 => x"737a2e80",
  1155 => x"fa387956",
  1156 => x"73902e80",
  1157 => x"e73802a7",
  1158 => x"0558768f",
  1159 => x"06547389",
  1160 => x"26bf3875",
  1161 => x"18b01555",
  1162 => x"55737534",
  1163 => x"76842aff",
  1164 => x"177081ff",
  1165 => x"06585557",
  1166 => x"75e03879",
  1167 => x"19557575",
  1168 => x"34787033",
  1169 => x"55557380",
  1170 => x"2e933881",
  1171 => x"15745280",
  1172 => x"f5900857",
  1173 => x"55752d74",
  1174 => x"335473ef",
  1175 => x"388e3d0d",
  1176 => x"047518b7",
  1177 => x"15555573",
  1178 => x"75347684",
  1179 => x"2aff1770",
  1180 => x"81ff0658",
  1181 => x"555775ff",
  1182 => x"a138c039",
  1183 => x"8470575a",
  1184 => x"02a70558",
  1185 => x"ff943982",
  1186 => x"70575af4",
  1187 => x"39ff3d0d",
  1188 => x"80df8408",
  1189 => x"74101075",
  1190 => x"10059412",
  1191 => x"0c52850b",
  1192 => x"98130c98",
  1193 => x"12087081",
  1194 => x"06515170",
  1195 => x"f638833d",
  1196 => x"0d04fd3d",
  1197 => x"0d80df84",
  1198 => x"0876b0ea",
  1199 => x"2994120c",
  1200 => x"54850b98",
  1201 => x"150c9814",
  1202 => x"08708106",
  1203 => x"515372f6",
  1204 => x"38853d0d",
  1205 => x"04803d0d",
  1206 => x"80df8408",
  1207 => x"51870b84",
  1208 => x"120cff0b",
  1209 => x"b4120ca7",
  1210 => x"0bb8120c",
  1211 => x"87e80ba4",
  1212 => x"120ca70b",
  1213 => x"a8120cb0",
  1214 => x"ea0b9412",
  1215 => x"0c870b98",
  1216 => x"120c823d",
  1217 => x"0d04803d",
  1218 => x"0d80df88",
  1219 => x"0851b60b",
  1220 => x"8c120c83",
  1221 => x"0b88120c",
  1222 => x"823d0d04",
  1223 => x"803d0d80",
  1224 => x"df880884",
  1225 => x"11088106",
  1226 => x"800c5182",
  1227 => x"3d0d04ff",
  1228 => x"3d0d80df",
  1229 => x"88085284",
  1230 => x"12087081",
  1231 => x"06515170",
  1232 => x"802ef438",
  1233 => x"71087081",
  1234 => x"ff06800c",
  1235 => x"51833d0d",
  1236 => x"04fe3d0d",
  1237 => x"02930533",
  1238 => x"53728a2e",
  1239 => x"9c3880df",
  1240 => x"88085284",
  1241 => x"12087089",
  1242 => x"2a708106",
  1243 => x"51515170",
  1244 => x"f2387272",
  1245 => x"0c843d0d",
  1246 => x"0480df88",
  1247 => x"08528412",
  1248 => x"0870892a",
  1249 => x"70810651",
  1250 => x"515170f2",
  1251 => x"388d720c",
  1252 => x"84120870",
  1253 => x"892a7081",
  1254 => x"06515151",
  1255 => x"70c538d2",
  1256 => x"39803d0d",
  1257 => x"80defc08",
  1258 => x"51800b84",
  1259 => x"120c83fe",
  1260 => x"800b8812",
  1261 => x"0c800b80",
  1262 => x"f5943480",
  1263 => x"0b80f598",
  1264 => x"34823d0d",
  1265 => x"04fa3d0d",
  1266 => x"02a30533",
  1267 => x"80defc08",
  1268 => x"80f59433",
  1269 => x"7081ff06",
  1270 => x"70101011",
  1271 => x"80f59833",
  1272 => x"7081ff06",
  1273 => x"72902911",
  1274 => x"70882b78",
  1275 => x"07770c53",
  1276 => x"5b5b5555",
  1277 => x"59545473",
  1278 => x"8a2e9838",
  1279 => x"7480cf2e",
  1280 => x"9238738c",
  1281 => x"2ea43881",
  1282 => x"16537280",
  1283 => x"f5983488",
  1284 => x"3d0d0471",
  1285 => x"a326a338",
  1286 => x"81175271",
  1287 => x"80f59434",
  1288 => x"800b80f5",
  1289 => x"9834883d",
  1290 => x"0d048052",
  1291 => x"71882b73",
  1292 => x"0c811252",
  1293 => x"97907226",
  1294 => x"f338800b",
  1295 => x"80f59434",
  1296 => x"800b80f5",
  1297 => x"9834df39",
  1298 => x"8c08028c",
  1299 => x"0cfd3d0d",
  1300 => x"80538c08",
  1301 => x"8c050852",
  1302 => x"8c088805",
  1303 => x"085182de",
  1304 => x"3f800870",
  1305 => x"800c5485",
  1306 => x"3d0d8c0c",
  1307 => x"048c0802",
  1308 => x"8c0cfd3d",
  1309 => x"0d81538c",
  1310 => x"088c0508",
  1311 => x"528c0888",
  1312 => x"05085182",
  1313 => x"b93f8008",
  1314 => x"70800c54",
  1315 => x"853d0d8c",
  1316 => x"0c048c08",
  1317 => x"028c0cf9",
  1318 => x"3d0d800b",
  1319 => x"8c08fc05",
  1320 => x"0c8c0888",
  1321 => x"05088025",
  1322 => x"ab388c08",
  1323 => x"88050830",
  1324 => x"8c088805",
  1325 => x"0c800b8c",
  1326 => x"08f4050c",
  1327 => x"8c08fc05",
  1328 => x"08883881",
  1329 => x"0b8c08f4",
  1330 => x"050c8c08",
  1331 => x"f405088c",
  1332 => x"08fc050c",
  1333 => x"8c088c05",
  1334 => x"088025ab",
  1335 => x"388c088c",
  1336 => x"0508308c",
  1337 => x"088c050c",
  1338 => x"800b8c08",
  1339 => x"f0050c8c",
  1340 => x"08fc0508",
  1341 => x"8838810b",
  1342 => x"8c08f005",
  1343 => x"0c8c08f0",
  1344 => x"05088c08",
  1345 => x"fc050c80",
  1346 => x"538c088c",
  1347 => x"0508528c",
  1348 => x"08880508",
  1349 => x"5181a73f",
  1350 => x"8008708c",
  1351 => x"08f8050c",
  1352 => x"548c08fc",
  1353 => x"0508802e",
  1354 => x"8c388c08",
  1355 => x"f8050830",
  1356 => x"8c08f805",
  1357 => x"0c8c08f8",
  1358 => x"05087080",
  1359 => x"0c54893d",
  1360 => x"0d8c0c04",
  1361 => x"8c08028c",
  1362 => x"0cfb3d0d",
  1363 => x"800b8c08",
  1364 => x"fc050c8c",
  1365 => x"08880508",
  1366 => x"80259338",
  1367 => x"8c088805",
  1368 => x"08308c08",
  1369 => x"88050c81",
  1370 => x"0b8c08fc",
  1371 => x"050c8c08",
  1372 => x"8c050880",
  1373 => x"258c388c",
  1374 => x"088c0508",
  1375 => x"308c088c",
  1376 => x"050c8153",
  1377 => x"8c088c05",
  1378 => x"08528c08",
  1379 => x"88050851",
  1380 => x"ad3f8008",
  1381 => x"708c08f8",
  1382 => x"050c548c",
  1383 => x"08fc0508",
  1384 => x"802e8c38",
  1385 => x"8c08f805",
  1386 => x"08308c08",
  1387 => x"f8050c8c",
  1388 => x"08f80508",
  1389 => x"70800c54",
  1390 => x"873d0d8c",
  1391 => x"0c048c08",
  1392 => x"028c0cfd",
  1393 => x"3d0d810b",
  1394 => x"8c08fc05",
  1395 => x"0c800b8c",
  1396 => x"08f8050c",
  1397 => x"8c088c05",
  1398 => x"088c0888",
  1399 => x"050827ac",
  1400 => x"388c08fc",
  1401 => x"0508802e",
  1402 => x"a338800b",
  1403 => x"8c088c05",
  1404 => x"08249938",
  1405 => x"8c088c05",
  1406 => x"08108c08",
  1407 => x"8c050c8c",
  1408 => x"08fc0508",
  1409 => x"108c08fc",
  1410 => x"050cc939",
  1411 => x"8c08fc05",
  1412 => x"08802e80",
  1413 => x"c9388c08",
  1414 => x"8c05088c",
  1415 => x"08880508",
  1416 => x"26a1388c",
  1417 => x"08880508",
  1418 => x"8c088c05",
  1419 => x"08318c08",
  1420 => x"88050c8c",
  1421 => x"08f80508",
  1422 => x"8c08fc05",
  1423 => x"08078c08",
  1424 => x"f8050c8c",
  1425 => x"08fc0508",
  1426 => x"812a8c08",
  1427 => x"fc050c8c",
  1428 => x"088c0508",
  1429 => x"812a8c08",
  1430 => x"8c050cff",
  1431 => x"af398c08",
  1432 => x"90050880",
  1433 => x"2e8f388c",
  1434 => x"08880508",
  1435 => x"708c08f4",
  1436 => x"050c518d",
  1437 => x"398c08f8",
  1438 => x"0508708c",
  1439 => x"08f4050c",
  1440 => x"518c08f4",
  1441 => x"0508800c",
  1442 => x"853d0d8c",
  1443 => x"0c04803d",
  1444 => x"0d865184",
  1445 => x"963f8151",
  1446 => x"9f873ffc",
  1447 => x"3d0d7670",
  1448 => x"797b5555",
  1449 => x"55558f72",
  1450 => x"278c3872",
  1451 => x"75078306",
  1452 => x"5170802e",
  1453 => x"a738ff12",
  1454 => x"5271ff2e",
  1455 => x"98387270",
  1456 => x"81055433",
  1457 => x"74708105",
  1458 => x"5634ff12",
  1459 => x"5271ff2e",
  1460 => x"098106ea",
  1461 => x"3874800c",
  1462 => x"863d0d04",
  1463 => x"74517270",
  1464 => x"84055408",
  1465 => x"71708405",
  1466 => x"530c7270",
  1467 => x"84055408",
  1468 => x"71708405",
  1469 => x"530c7270",
  1470 => x"84055408",
  1471 => x"71708405",
  1472 => x"530c7270",
  1473 => x"84055408",
  1474 => x"71708405",
  1475 => x"530cf012",
  1476 => x"52718f26",
  1477 => x"c9388372",
  1478 => x"27953872",
  1479 => x"70840554",
  1480 => x"08717084",
  1481 => x"05530cfc",
  1482 => x"12527183",
  1483 => x"26ed3870",
  1484 => x"54ff8339",
  1485 => x"fd3d0d75",
  1486 => x"5384d813",
  1487 => x"08802e8a",
  1488 => x"38805372",
  1489 => x"800c853d",
  1490 => x"0d048180",
  1491 => x"5272518a",
  1492 => x"883f8008",
  1493 => x"84d8140c",
  1494 => x"ff538008",
  1495 => x"802ee438",
  1496 => x"8008549f",
  1497 => x"53807470",
  1498 => x"8405560c",
  1499 => x"ff135380",
  1500 => x"7324ce38",
  1501 => x"80747084",
  1502 => x"05560cff",
  1503 => x"13537280",
  1504 => x"25e338ff",
  1505 => x"bc39fd3d",
  1506 => x"0d757755",
  1507 => x"539f7427",
  1508 => x"8d389673",
  1509 => x"0cff5271",
  1510 => x"800c853d",
  1511 => x"0d0484d8",
  1512 => x"13085271",
  1513 => x"802e9338",
  1514 => x"73101012",
  1515 => x"70087972",
  1516 => x"0c515271",
  1517 => x"800c853d",
  1518 => x"0d047251",
  1519 => x"fef63fff",
  1520 => x"528008d3",
  1521 => x"3884d813",
  1522 => x"08741010",
  1523 => x"1170087a",
  1524 => x"720c5151",
  1525 => x"52dd39f9",
  1526 => x"3d0d797b",
  1527 => x"5856769f",
  1528 => x"2680e838",
  1529 => x"84d81608",
  1530 => x"5473802e",
  1531 => x"aa387610",
  1532 => x"10147008",
  1533 => x"55557380",
  1534 => x"2eba3880",
  1535 => x"5873812e",
  1536 => x"8f3873ff",
  1537 => x"2ea33880",
  1538 => x"750c7651",
  1539 => x"732d8058",
  1540 => x"77800c89",
  1541 => x"3d0d0475",
  1542 => x"51fe993f",
  1543 => x"ff588008",
  1544 => x"ef3884d8",
  1545 => x"160854c6",
  1546 => x"3996760c",
  1547 => x"810b800c",
  1548 => x"893d0d04",
  1549 => x"755181ed",
  1550 => x"3f765380",
  1551 => x"08527551",
  1552 => x"81ad3f80",
  1553 => x"08800c89",
  1554 => x"3d0d0496",
  1555 => x"760cff0b",
  1556 => x"800c893d",
  1557 => x"0d04fc3d",
  1558 => x"0d767856",
  1559 => x"53ff5474",
  1560 => x"9f26b138",
  1561 => x"84d81308",
  1562 => x"5271802e",
  1563 => x"ae387410",
  1564 => x"10127008",
  1565 => x"53538154",
  1566 => x"71802e98",
  1567 => x"38825471",
  1568 => x"ff2e9138",
  1569 => x"83547181",
  1570 => x"2e8a3880",
  1571 => x"730c7451",
  1572 => x"712d8054",
  1573 => x"73800c86",
  1574 => x"3d0d0472",
  1575 => x"51fd953f",
  1576 => x"8008f138",
  1577 => x"84d81308",
  1578 => x"52c439ff",
  1579 => x"3d0d7352",
  1580 => x"80df8c08",
  1581 => x"51fea03f",
  1582 => x"833d0d04",
  1583 => x"fe3d0d75",
  1584 => x"53745280",
  1585 => x"df8c0851",
  1586 => x"fdbc3f84",
  1587 => x"3d0d0480",
  1588 => x"3d0d80df",
  1589 => x"8c0851fc",
  1590 => x"db3f823d",
  1591 => x"0d04ff3d",
  1592 => x"0d735280",
  1593 => x"df8c0851",
  1594 => x"feec3f83",
  1595 => x"3d0d04fc",
  1596 => x"3d0d800b",
  1597 => x"80f5a40c",
  1598 => x"78527751",
  1599 => x"99973f80",
  1600 => x"08548008",
  1601 => x"ff2e8838",
  1602 => x"73800c86",
  1603 => x"3d0d0480",
  1604 => x"f5a40855",
  1605 => x"74802ef0",
  1606 => x"38767571",
  1607 => x"0c537380",
  1608 => x"0c863d0d",
  1609 => x"0498e93f",
  1610 => x"04fc3d0d",
  1611 => x"76707970",
  1612 => x"73078306",
  1613 => x"54545455",
  1614 => x"7080c338",
  1615 => x"71700870",
  1616 => x"0970f7fb",
  1617 => x"fdff1306",
  1618 => x"70f88482",
  1619 => x"81800651",
  1620 => x"51535354",
  1621 => x"70a63884",
  1622 => x"14727470",
  1623 => x"8405560c",
  1624 => x"70087009",
  1625 => x"70f7fbfd",
  1626 => x"ff130670",
  1627 => x"f8848281",
  1628 => x"80065151",
  1629 => x"53535470",
  1630 => x"802edc38",
  1631 => x"73527170",
  1632 => x"81055333",
  1633 => x"51707370",
  1634 => x"81055534",
  1635 => x"70f03874",
  1636 => x"800c863d",
  1637 => x"0d04fd3d",
  1638 => x"0d757071",
  1639 => x"83065355",
  1640 => x"5270b838",
  1641 => x"71700870",
  1642 => x"09f7fbfd",
  1643 => x"ff120670",
  1644 => x"f8848281",
  1645 => x"80065151",
  1646 => x"5253709d",
  1647 => x"38841370",
  1648 => x"087009f7",
  1649 => x"fbfdff12",
  1650 => x"0670f884",
  1651 => x"82818006",
  1652 => x"51515253",
  1653 => x"70802ee5",
  1654 => x"38725271",
  1655 => x"33517080",
  1656 => x"2e8a3881",
  1657 => x"12703352",
  1658 => x"5270f838",
  1659 => x"71743180",
  1660 => x"0c853d0d",
  1661 => x"04fa3d0d",
  1662 => x"787a7c70",
  1663 => x"54555552",
  1664 => x"72802e80",
  1665 => x"d9387174",
  1666 => x"07830651",
  1667 => x"70802e80",
  1668 => x"d438ff13",
  1669 => x"5372ff2e",
  1670 => x"b1387133",
  1671 => x"74335651",
  1672 => x"74712e09",
  1673 => x"8106a938",
  1674 => x"72802e81",
  1675 => x"87387081",
  1676 => x"ff065170",
  1677 => x"802e80fc",
  1678 => x"38811281",
  1679 => x"15ff1555",
  1680 => x"555272ff",
  1681 => x"2e098106",
  1682 => x"d1387133",
  1683 => x"74335651",
  1684 => x"7081ff06",
  1685 => x"7581ff06",
  1686 => x"71713151",
  1687 => x"52527080",
  1688 => x"0c883d0d",
  1689 => x"04717457",
  1690 => x"55837327",
  1691 => x"88387108",
  1692 => x"74082e88",
  1693 => x"38747655",
  1694 => x"52ff9739",
  1695 => x"fc135372",
  1696 => x"802eb138",
  1697 => x"74087009",
  1698 => x"f7fbfdff",
  1699 => x"120670f8",
  1700 => x"84828180",
  1701 => x"06515151",
  1702 => x"709a3884",
  1703 => x"15841757",
  1704 => x"55837327",
  1705 => x"d0387408",
  1706 => x"76082ed0",
  1707 => x"38747655",
  1708 => x"52fedf39",
  1709 => x"800b800c",
  1710 => x"883d0d04",
  1711 => x"f33d0d60",
  1712 => x"6264725a",
  1713 => x"5a5d5d80",
  1714 => x"5e767081",
  1715 => x"05583380",
  1716 => x"dcbd1133",
  1717 => x"70832a70",
  1718 => x"81065155",
  1719 => x"555672e9",
  1720 => x"3875ad2e",
  1721 => x"81ff3875",
  1722 => x"ab2e81fb",
  1723 => x"38773070",
  1724 => x"79078025",
  1725 => x"79903270",
  1726 => x"30707207",
  1727 => x"80257307",
  1728 => x"53575751",
  1729 => x"5372802e",
  1730 => x"873875b0",
  1731 => x"2e81e238",
  1732 => x"778a3888",
  1733 => x"5875b02e",
  1734 => x"83388a58",
  1735 => x"7752ff51",
  1736 => x"f2a63f80",
  1737 => x"0878535a",
  1738 => x"ff51f2c1",
  1739 => x"3f80085b",
  1740 => x"80705a55",
  1741 => x"80dcbd16",
  1742 => x"3370822a",
  1743 => x"70810651",
  1744 => x"54547280",
  1745 => x"2e80c138",
  1746 => x"d0165675",
  1747 => x"782580d7",
  1748 => x"38807924",
  1749 => x"757b2607",
  1750 => x"53729338",
  1751 => x"747a2e80",
  1752 => x"eb387a76",
  1753 => x"2580ed38",
  1754 => x"72802e80",
  1755 => x"e738ff77",
  1756 => x"70810559",
  1757 => x"33575980",
  1758 => x"dcbd1633",
  1759 => x"70822a70",
  1760 => x"81065154",
  1761 => x"5472c138",
  1762 => x"73830653",
  1763 => x"72802e97",
  1764 => x"38738106",
  1765 => x"c9175553",
  1766 => x"728538ff",
  1767 => x"a9165473",
  1768 => x"56777624",
  1769 => x"ffab3880",
  1770 => x"79248189",
  1771 => x"387d802e",
  1772 => x"84387430",
  1773 => x"557b802e",
  1774 => x"8c38ff17",
  1775 => x"53788338",
  1776 => x"7c53727c",
  1777 => x"0c74800c",
  1778 => x"8f3d0d04",
  1779 => x"8153757b",
  1780 => x"24ff9538",
  1781 => x"81757929",
  1782 => x"17787081",
  1783 => x"055a3358",
  1784 => x"5659ff93",
  1785 => x"39815e76",
  1786 => x"70810558",
  1787 => x"3356fdfd",
  1788 => x"39807733",
  1789 => x"54547280",
  1790 => x"f82e80c3",
  1791 => x"387280d8",
  1792 => x"32703070",
  1793 => x"80257607",
  1794 => x"51515372",
  1795 => x"802efe80",
  1796 => x"38811733",
  1797 => x"82185856",
  1798 => x"90705358",
  1799 => x"ff51f0a8",
  1800 => x"3f800878",
  1801 => x"535aff51",
  1802 => x"f0c33f80",
  1803 => x"085b8070",
  1804 => x"5a55fe80",
  1805 => x"39ff6054",
  1806 => x"55a2730c",
  1807 => x"fef73981",
  1808 => x"54ffba39",
  1809 => x"fd3d0d77",
  1810 => x"54765375",
  1811 => x"5280df8c",
  1812 => x"0851fce8",
  1813 => x"3f853d0d",
  1814 => x"04f33d0d",
  1815 => x"7f618b11",
  1816 => x"70f8065c",
  1817 => x"55555e72",
  1818 => x"96268338",
  1819 => x"90598079",
  1820 => x"24747a26",
  1821 => x"07538054",
  1822 => x"72742e09",
  1823 => x"810680cb",
  1824 => x"387d518b",
  1825 => x"ca3f7883",
  1826 => x"f72680c6",
  1827 => x"3878832a",
  1828 => x"70101010",
  1829 => x"80e6c805",
  1830 => x"8c110859",
  1831 => x"595a7678",
  1832 => x"2e83b038",
  1833 => x"841708fc",
  1834 => x"06568c17",
  1835 => x"08881808",
  1836 => x"718c120c",
  1837 => x"88120c58",
  1838 => x"75178411",
  1839 => x"08810784",
  1840 => x"120c537d",
  1841 => x"518b893f",
  1842 => x"88175473",
  1843 => x"800c8f3d",
  1844 => x"0d047889",
  1845 => x"2a79832a",
  1846 => x"5b537280",
  1847 => x"2ebf3878",
  1848 => x"862ab805",
  1849 => x"5a847327",
  1850 => x"b43880db",
  1851 => x"135a9473",
  1852 => x"27ab3878",
  1853 => x"8c2a80ee",
  1854 => x"055a80d4",
  1855 => x"73279e38",
  1856 => x"788f2a80",
  1857 => x"f7055a82",
  1858 => x"d4732791",
  1859 => x"3878922a",
  1860 => x"80fc055a",
  1861 => x"8ad47327",
  1862 => x"843880fe",
  1863 => x"5a791010",
  1864 => x"1080e6c8",
  1865 => x"058c1108",
  1866 => x"58557675",
  1867 => x"2ea33884",
  1868 => x"1708fc06",
  1869 => x"707a3155",
  1870 => x"56738f24",
  1871 => x"88d53873",
  1872 => x"8025fee6",
  1873 => x"388c1708",
  1874 => x"5776752e",
  1875 => x"098106df",
  1876 => x"38811a5a",
  1877 => x"80e6d808",
  1878 => x"577680e6",
  1879 => x"d02e82c0",
  1880 => x"38841708",
  1881 => x"fc06707a",
  1882 => x"31555673",
  1883 => x"8f2481f9",
  1884 => x"3880e6d0",
  1885 => x"0b80e6dc",
  1886 => x"0c80e6d0",
  1887 => x"0b80e6d8",
  1888 => x"0c738025",
  1889 => x"feb23883",
  1890 => x"ff762783",
  1891 => x"df387589",
  1892 => x"2a76832a",
  1893 => x"55537280",
  1894 => x"2ebf3875",
  1895 => x"862ab805",
  1896 => x"54847327",
  1897 => x"b43880db",
  1898 => x"13549473",
  1899 => x"27ab3875",
  1900 => x"8c2a80ee",
  1901 => x"055480d4",
  1902 => x"73279e38",
  1903 => x"758f2a80",
  1904 => x"f7055482",
  1905 => x"d4732791",
  1906 => x"3875922a",
  1907 => x"80fc0554",
  1908 => x"8ad47327",
  1909 => x"843880fe",
  1910 => x"54731010",
  1911 => x"1080e6c8",
  1912 => x"05881108",
  1913 => x"56587478",
  1914 => x"2e86cf38",
  1915 => x"841508fc",
  1916 => x"06537573",
  1917 => x"278d3888",
  1918 => x"15085574",
  1919 => x"782e0981",
  1920 => x"06ea388c",
  1921 => x"150880e6",
  1922 => x"c80b8405",
  1923 => x"08718c1a",
  1924 => x"0c76881a",
  1925 => x"0c788813",
  1926 => x"0c788c18",
  1927 => x"0c5d5879",
  1928 => x"53807a24",
  1929 => x"83e63872",
  1930 => x"822c8171",
  1931 => x"2b5c537a",
  1932 => x"7c268198",
  1933 => x"387b7b06",
  1934 => x"537282f1",
  1935 => x"3879fc06",
  1936 => x"84055a7a",
  1937 => x"10707d06",
  1938 => x"545b7282",
  1939 => x"e038841a",
  1940 => x"5af13988",
  1941 => x"178c1108",
  1942 => x"58587678",
  1943 => x"2e098106",
  1944 => x"fcc23882",
  1945 => x"1a5afdec",
  1946 => x"39781779",
  1947 => x"81078419",
  1948 => x"0c7080e6",
  1949 => x"dc0c7080",
  1950 => x"e6d80c80",
  1951 => x"e6d00b8c",
  1952 => x"120c8c11",
  1953 => x"0888120c",
  1954 => x"74810784",
  1955 => x"120c7411",
  1956 => x"75710c51",
  1957 => x"537d5187",
  1958 => x"b73f8817",
  1959 => x"54fcac39",
  1960 => x"80e6c80b",
  1961 => x"8405087a",
  1962 => x"545c7980",
  1963 => x"25fef838",
  1964 => x"82da397a",
  1965 => x"097c0670",
  1966 => x"80e6c80b",
  1967 => x"84050c5c",
  1968 => x"7a105b7a",
  1969 => x"7c268538",
  1970 => x"7a85b838",
  1971 => x"80e6c80b",
  1972 => x"88050870",
  1973 => x"841208fc",
  1974 => x"06707c31",
  1975 => x"7c72268f",
  1976 => x"72250757",
  1977 => x"575c5d55",
  1978 => x"72802e80",
  1979 => x"db38797a",
  1980 => x"1680e6c0",
  1981 => x"081b9011",
  1982 => x"5a55575b",
  1983 => x"80e6bc08",
  1984 => x"ff2e8838",
  1985 => x"a08f13e0",
  1986 => x"80065776",
  1987 => x"527d5186",
  1988 => x"c03f8008",
  1989 => x"548008ff",
  1990 => x"2e903880",
  1991 => x"08762782",
  1992 => x"99387480",
  1993 => x"e6c82e82",
  1994 => x"913880e6",
  1995 => x"c80b8805",
  1996 => x"08558415",
  1997 => x"08fc0670",
  1998 => x"7a317a72",
  1999 => x"268f7225",
  2000 => x"07525553",
  2001 => x"7283e638",
  2002 => x"74798107",
  2003 => x"84170c79",
  2004 => x"167080e6",
  2005 => x"c80b8805",
  2006 => x"0c758107",
  2007 => x"84120c54",
  2008 => x"7e525785",
  2009 => x"eb3f8817",
  2010 => x"54fae039",
  2011 => x"75832a70",
  2012 => x"54548074",
  2013 => x"24819b38",
  2014 => x"72822c81",
  2015 => x"712b80e6",
  2016 => x"cc080770",
  2017 => x"80e6c80b",
  2018 => x"84050c75",
  2019 => x"10101080",
  2020 => x"e6c80588",
  2021 => x"1108585a",
  2022 => x"5d53778c",
  2023 => x"180c7488",
  2024 => x"180c7688",
  2025 => x"190c768c",
  2026 => x"160cfcf3",
  2027 => x"39797a10",
  2028 => x"101080e6",
  2029 => x"c8057057",
  2030 => x"595d8c15",
  2031 => x"08577675",
  2032 => x"2ea33884",
  2033 => x"1708fc06",
  2034 => x"707a3155",
  2035 => x"56738f24",
  2036 => x"83ca3873",
  2037 => x"80258481",
  2038 => x"388c1708",
  2039 => x"5776752e",
  2040 => x"098106df",
  2041 => x"38881581",
  2042 => x"1b708306",
  2043 => x"555b5572",
  2044 => x"c9387c83",
  2045 => x"06537280",
  2046 => x"2efdb838",
  2047 => x"ff1df819",
  2048 => x"595d8818",
  2049 => x"08782eea",
  2050 => x"38fdb539",
  2051 => x"831a53fc",
  2052 => x"96398314",
  2053 => x"70822c81",
  2054 => x"712b80e6",
  2055 => x"cc080770",
  2056 => x"80e6c80b",
  2057 => x"84050c76",
  2058 => x"10101080",
  2059 => x"e6c80588",
  2060 => x"1108595b",
  2061 => x"5e5153fe",
  2062 => x"e13980e6",
  2063 => x"8c081758",
  2064 => x"8008762e",
  2065 => x"818d3880",
  2066 => x"e6bc08ff",
  2067 => x"2e83ec38",
  2068 => x"73763118",
  2069 => x"80e68c0c",
  2070 => x"73870670",
  2071 => x"57537280",
  2072 => x"2e883888",
  2073 => x"73317015",
  2074 => x"55567614",
  2075 => x"9fff06a0",
  2076 => x"80713117",
  2077 => x"70547f53",
  2078 => x"575383d5",
  2079 => x"3f800853",
  2080 => x"8008ff2e",
  2081 => x"81a03880",
  2082 => x"e68c0816",
  2083 => x"7080e68c",
  2084 => x"0c747580",
  2085 => x"e6c80b88",
  2086 => x"050c7476",
  2087 => x"31187081",
  2088 => x"07515556",
  2089 => x"587b80e6",
  2090 => x"c82e839c",
  2091 => x"38798f26",
  2092 => x"82cb3881",
  2093 => x"0b84150c",
  2094 => x"841508fc",
  2095 => x"06707a31",
  2096 => x"7a72268f",
  2097 => x"72250752",
  2098 => x"55537280",
  2099 => x"2efcf938",
  2100 => x"80db3980",
  2101 => x"089fff06",
  2102 => x"5372feeb",
  2103 => x"387780e6",
  2104 => x"8c0c80e6",
  2105 => x"c80b8805",
  2106 => x"087b1881",
  2107 => x"0784120c",
  2108 => x"5580e6b8",
  2109 => x"08782786",
  2110 => x"387780e6",
  2111 => x"b80c80e6",
  2112 => x"b4087827",
  2113 => x"fcac3877",
  2114 => x"80e6b40c",
  2115 => x"841508fc",
  2116 => x"06707a31",
  2117 => x"7a72268f",
  2118 => x"72250752",
  2119 => x"55537280",
  2120 => x"2efca538",
  2121 => x"88398074",
  2122 => x"5456fedb",
  2123 => x"397d5182",
  2124 => x"9f3f800b",
  2125 => x"800c8f3d",
  2126 => x"0d047353",
  2127 => x"807424a9",
  2128 => x"3872822c",
  2129 => x"81712b80",
  2130 => x"e6cc0807",
  2131 => x"7080e6c8",
  2132 => x"0b84050c",
  2133 => x"5d53778c",
  2134 => x"180c7488",
  2135 => x"180c7688",
  2136 => x"190c768c",
  2137 => x"160cf9b7",
  2138 => x"39831470",
  2139 => x"822c8171",
  2140 => x"2b80e6cc",
  2141 => x"08077080",
  2142 => x"e6c80b84",
  2143 => x"050c5e51",
  2144 => x"53d4397b",
  2145 => x"7b065372",
  2146 => x"fca33884",
  2147 => x"1a7b105c",
  2148 => x"5af139ff",
  2149 => x"1a811151",
  2150 => x"5af7b939",
  2151 => x"78177981",
  2152 => x"0784190c",
  2153 => x"8c180888",
  2154 => x"1908718c",
  2155 => x"120c8812",
  2156 => x"0c597080",
  2157 => x"e6dc0c70",
  2158 => x"80e6d80c",
  2159 => x"80e6d00b",
  2160 => x"8c120c8c",
  2161 => x"11088812",
  2162 => x"0c748107",
  2163 => x"84120c74",
  2164 => x"1175710c",
  2165 => x"5153f9bd",
  2166 => x"39751784",
  2167 => x"11088107",
  2168 => x"84120c53",
  2169 => x"8c170888",
  2170 => x"1808718c",
  2171 => x"120c8812",
  2172 => x"0c587d51",
  2173 => x"80da3f88",
  2174 => x"1754f5cf",
  2175 => x"39728415",
  2176 => x"0cf41af8",
  2177 => x"0670841e",
  2178 => x"08810607",
  2179 => x"841e0c70",
  2180 => x"1d545b85",
  2181 => x"0b84140c",
  2182 => x"850b8814",
  2183 => x"0c8f7b27",
  2184 => x"fdcf3888",
  2185 => x"1c527d51",
  2186 => x"82903f80",
  2187 => x"e6c80b88",
  2188 => x"050880e6",
  2189 => x"8c085955",
  2190 => x"fdb73977",
  2191 => x"80e68c0c",
  2192 => x"7380e6bc",
  2193 => x"0cfc9139",
  2194 => x"7284150c",
  2195 => x"fda33904",
  2196 => x"04fd3d0d",
  2197 => x"800b80f5",
  2198 => x"a40c7651",
  2199 => x"86cc3f80",
  2200 => x"08538008",
  2201 => x"ff2e8838",
  2202 => x"72800c85",
  2203 => x"3d0d0480",
  2204 => x"f5a40854",
  2205 => x"73802ef0",
  2206 => x"38757471",
  2207 => x"0c527280",
  2208 => x"0c853d0d",
  2209 => x"04fb3d0d",
  2210 => x"77705256",
  2211 => x"c23f80e6",
  2212 => x"c80b8805",
  2213 => x"08841108",
  2214 => x"fc06707b",
  2215 => x"319fef05",
  2216 => x"e08006e0",
  2217 => x"80055656",
  2218 => x"53a08074",
  2219 => x"24943880",
  2220 => x"527551ff",
  2221 => x"9c3f80e6",
  2222 => x"d0081553",
  2223 => x"7280082e",
  2224 => x"8f387551",
  2225 => x"ff8a3f80",
  2226 => x"5372800c",
  2227 => x"873d0d04",
  2228 => x"73305275",
  2229 => x"51fefa3f",
  2230 => x"8008ff2e",
  2231 => x"a83880e6",
  2232 => x"c80b8805",
  2233 => x"08757531",
  2234 => x"81078412",
  2235 => x"0c5380e6",
  2236 => x"8c087431",
  2237 => x"80e68c0c",
  2238 => x"7551fed4",
  2239 => x"3f810b80",
  2240 => x"0c873d0d",
  2241 => x"04805275",
  2242 => x"51fec63f",
  2243 => x"80e6c80b",
  2244 => x"88050880",
  2245 => x"08713156",
  2246 => x"538f7525",
  2247 => x"ffa43880",
  2248 => x"0880e6bc",
  2249 => x"083180e6",
  2250 => x"8c0c7481",
  2251 => x"0784140c",
  2252 => x"7551fe9c",
  2253 => x"3f8053ff",
  2254 => x"9039f63d",
  2255 => x"0d7c7e54",
  2256 => x"5b72802e",
  2257 => x"8283387a",
  2258 => x"51fe843f",
  2259 => x"f8138411",
  2260 => x"0870fe06",
  2261 => x"70138411",
  2262 => x"08fc065d",
  2263 => x"58595458",
  2264 => x"80e6d008",
  2265 => x"752e82de",
  2266 => x"38788416",
  2267 => x"0c807381",
  2268 => x"06545a72",
  2269 => x"7a2e81d5",
  2270 => x"38781584",
  2271 => x"11088106",
  2272 => x"515372a0",
  2273 => x"38781757",
  2274 => x"7981e638",
  2275 => x"88150853",
  2276 => x"7280e6d0",
  2277 => x"2e82f938",
  2278 => x"8c150870",
  2279 => x"8c150c73",
  2280 => x"88120c56",
  2281 => x"76810784",
  2282 => x"190c7618",
  2283 => x"77710c53",
  2284 => x"79819138",
  2285 => x"83ff7727",
  2286 => x"81c83876",
  2287 => x"892a7783",
  2288 => x"2a565372",
  2289 => x"802ebf38",
  2290 => x"76862ab8",
  2291 => x"05558473",
  2292 => x"27b43880",
  2293 => x"db135594",
  2294 => x"7327ab38",
  2295 => x"768c2a80",
  2296 => x"ee055580",
  2297 => x"d473279e",
  2298 => x"38768f2a",
  2299 => x"80f70555",
  2300 => x"82d47327",
  2301 => x"91387692",
  2302 => x"2a80fc05",
  2303 => x"558ad473",
  2304 => x"27843880",
  2305 => x"fe557410",
  2306 => x"101080e6",
  2307 => x"c8058811",
  2308 => x"08555673",
  2309 => x"762e82b3",
  2310 => x"38841408",
  2311 => x"fc065376",
  2312 => x"73278d38",
  2313 => x"88140854",
  2314 => x"73762e09",
  2315 => x"8106ea38",
  2316 => x"8c140870",
  2317 => x"8c1a0c74",
  2318 => x"881a0c78",
  2319 => x"88120c56",
  2320 => x"778c150c",
  2321 => x"7a51fc88",
  2322 => x"3f8c3d0d",
  2323 => x"04770878",
  2324 => x"71315977",
  2325 => x"05881908",
  2326 => x"54577280",
  2327 => x"e6d02e80",
  2328 => x"e0388c18",
  2329 => x"08708c15",
  2330 => x"0c738812",
  2331 => x"0c56fe89",
  2332 => x"39881508",
  2333 => x"8c160870",
  2334 => x"8c130c57",
  2335 => x"88170cfe",
  2336 => x"a3397683",
  2337 => x"2a705455",
  2338 => x"80752481",
  2339 => x"98387282",
  2340 => x"2c81712b",
  2341 => x"80e6cc08",
  2342 => x"0780e6c8",
  2343 => x"0b84050c",
  2344 => x"53741010",
  2345 => x"1080e6c8",
  2346 => x"05881108",
  2347 => x"5556758c",
  2348 => x"190c7388",
  2349 => x"190c7788",
  2350 => x"170c778c",
  2351 => x"150cff84",
  2352 => x"39815afd",
  2353 => x"b4397817",
  2354 => x"73810654",
  2355 => x"57729838",
  2356 => x"77087871",
  2357 => x"31597705",
  2358 => x"8c190888",
  2359 => x"1a08718c",
  2360 => x"120c8812",
  2361 => x"0c575776",
  2362 => x"81078419",
  2363 => x"0c7780e6",
  2364 => x"c80b8805",
  2365 => x"0c80e6c4",
  2366 => x"087726fe",
  2367 => x"c73880e6",
  2368 => x"c008527a",
  2369 => x"51fafe3f",
  2370 => x"7a51fac4",
  2371 => x"3ffeba39",
  2372 => x"81788c15",
  2373 => x"0c788815",
  2374 => x"0c738c1a",
  2375 => x"0c73881a",
  2376 => x"0c5afd80",
  2377 => x"39831570",
  2378 => x"822c8171",
  2379 => x"2b80e6cc",
  2380 => x"080780e6",
  2381 => x"c80b8405",
  2382 => x"0c515374",
  2383 => x"10101080",
  2384 => x"e6c80588",
  2385 => x"11085556",
  2386 => x"fee43974",
  2387 => x"53807524",
  2388 => x"a7387282",
  2389 => x"2c81712b",
  2390 => x"80e6cc08",
  2391 => x"0780e6c8",
  2392 => x"0b84050c",
  2393 => x"53758c19",
  2394 => x"0c738819",
  2395 => x"0c778817",
  2396 => x"0c778c15",
  2397 => x"0cfdcd39",
  2398 => x"83157082",
  2399 => x"2c81712b",
  2400 => x"80e6cc08",
  2401 => x"0780e6c8",
  2402 => x"0b84050c",
  2403 => x"5153d639",
  2404 => x"810b800c",
  2405 => x"04803d0d",
  2406 => x"72812e89",
  2407 => x"38800b80",
  2408 => x"0c823d0d",
  2409 => x"04735180",
  2410 => x"f83ffe3d",
  2411 => x"0d80f59c",
  2412 => x"0851708a",
  2413 => x"3880f5a8",
  2414 => x"7080f59c",
  2415 => x"0c517075",
  2416 => x"125252ff",
  2417 => x"537087fb",
  2418 => x"80802688",
  2419 => x"387080f5",
  2420 => x"9c0c7153",
  2421 => x"72800c84",
  2422 => x"3d0d04fd",
  2423 => x"3d0d800b",
  2424 => x"80dee408",
  2425 => x"54547281",
  2426 => x"2e9c3873",
  2427 => x"80f5a00c",
  2428 => x"ffbced3f",
  2429 => x"ffbc893f",
  2430 => x"80eed052",
  2431 => x"8151d4b6",
  2432 => x"3f800851",
  2433 => x"9f3f7280",
  2434 => x"f5a00cff",
  2435 => x"bcd23fff",
  2436 => x"bbee3f80",
  2437 => x"eed05281",
  2438 => x"51d49b3f",
  2439 => x"80085184",
  2440 => x"3f00ff39",
  2441 => x"f73d0d7b",
  2442 => x"80df8c08",
  2443 => x"82c81108",
  2444 => x"5a545a77",
  2445 => x"802e80da",
  2446 => x"38818818",
  2447 => x"841908ff",
  2448 => x"0581712b",
  2449 => x"59555980",
  2450 => x"742480ea",
  2451 => x"38807424",
  2452 => x"b5387382",
  2453 => x"2b781188",
  2454 => x"05565681",
  2455 => x"80190877",
  2456 => x"06537280",
  2457 => x"2eb63878",
  2458 => x"16700853",
  2459 => x"53795174",
  2460 => x"0853722d",
  2461 => x"ff14fc17",
  2462 => x"fc177981",
  2463 => x"2c5a5757",
  2464 => x"54738025",
  2465 => x"d6387708",
  2466 => x"5877ffad",
  2467 => x"3880df8c",
  2468 => x"0853bc13",
  2469 => x"08a53879",
  2470 => x"51ff863f",
  2471 => x"74085372",
  2472 => x"2dff14fc",
  2473 => x"17fc1779",
  2474 => x"812c5a57",
  2475 => x"57547380",
  2476 => x"25ffa838",
  2477 => x"d1398057",
  2478 => x"ff933972",
  2479 => x"51bc1308",
  2480 => x"53722d79",
  2481 => x"51feda3f",
  2482 => x"ff3d0d80",
  2483 => x"eed80bfc",
  2484 => x"05700852",
  2485 => x"5270ff2e",
  2486 => x"9138702d",
  2487 => x"fc127008",
  2488 => x"525270ff",
  2489 => x"2e098106",
  2490 => x"f138833d",
  2491 => x"0d0404ff",
  2492 => x"bbdb3f04",
  2493 => x"00000040",
  2494 => x"68656c70",
  2495 => x"00000000",
  2496 => x"3e200000",
  2497 => x"636f6d6d",
  2498 => x"616e6420",
  2499 => x"6e6f7420",
  2500 => x"666f756e",
  2501 => x"642e0a00",
  2502 => x"6d656d00",
  2503 => x"6c696b65",
  2504 => x"20780000",
  2505 => x"776d656d",
  2506 => x"00000000",
  2507 => x"77726974",
  2508 => x"6520776f",
  2509 => x"72640000",
  2510 => x"6558616d",
  2511 => x"696e6520",
  2512 => x"6d656d6f",
  2513 => x"72790000",
  2514 => x"636c6561",
  2515 => x"72000000",
  2516 => x"636c6561",
  2517 => x"72207363",
  2518 => x"7265656e",
  2519 => x"00000000",
  2520 => x"6c656400",
  2521 => x"73746172",
  2522 => x"74204c45",
  2523 => x"44207465",
  2524 => x"73740000",
  2525 => x"71756974",
  2526 => x"00000000",
  2527 => x"73757070",
  2528 => x"6f727465",
  2529 => x"6420636f",
  2530 => x"6d6d616e",
  2531 => x"64733a0a",
  2532 => x"0a000000",
  2533 => x"202d2000",
  2534 => x"0a307800",
  2535 => x"203a2000",
  2536 => x"0a677265",
  2537 => x"74682072",
  2538 => x"65676973",
  2539 => x"74657273",
  2540 => x"3a000000",
  2541 => x"0a636f6e",
  2542 => x"74726f6c",
  2543 => x"3a202020",
  2544 => x"20202030",
  2545 => x"78000000",
  2546 => x"0a737461",
  2547 => x"7475733a",
  2548 => x"20202020",
  2549 => x"20202030",
  2550 => x"78000000",
  2551 => x"0a6d6163",
  2552 => x"5f6d7362",
  2553 => x"3a202020",
  2554 => x"20202030",
  2555 => x"78000000",
  2556 => x"0a6d6163",
  2557 => x"5f6c7362",
  2558 => x"3a202020",
  2559 => x"20202030",
  2560 => x"78000000",
  2561 => x"0a6d6469",
  2562 => x"6f5f636f",
  2563 => x"6e74726f",
  2564 => x"6c3a2030",
  2565 => x"78000000",
  2566 => x"0a74785f",
  2567 => x"706f696e",
  2568 => x"7465723a",
  2569 => x"20202030",
  2570 => x"78000000",
  2571 => x"0a72785f",
  2572 => x"706f696e",
  2573 => x"7465723a",
  2574 => x"20202030",
  2575 => x"78000000",
  2576 => x"0a656463",
  2577 => x"6c5f6970",
  2578 => x"3a202020",
  2579 => x"20202030",
  2580 => x"78000000",
  2581 => x"0a686173",
  2582 => x"685f6d73",
  2583 => x"623a2020",
  2584 => x"20202030",
  2585 => x"78000000",
  2586 => x"0a686173",
  2587 => x"685f6c73",
  2588 => x"623a2020",
  2589 => x"20202030",
  2590 => x"78000000",
  2591 => x"0a6d6469",
  2592 => x"6f207068",
  2593 => x"79207265",
  2594 => x"67697374",
  2595 => x"65727300",
  2596 => x"0a206d64",
  2597 => x"696f2070",
  2598 => x"68793a20",
  2599 => x"30780000",
  2600 => x"0a202072",
  2601 => x"65673a20",
  2602 => x"00000000",
  2603 => x"2d3e2030",
  2604 => x"78000000",
  2605 => x"67726574",
  2606 => x"682d3e63",
  2607 => x"6f6e7472",
  2608 => x"6f6c3a20",
  2609 => x"30780000",
  2610 => x"67726574",
  2611 => x"682d3e73",
  2612 => x"74617475",
  2613 => x"73203a20",
  2614 => x"30780000",
  2615 => x"64657363",
  2616 => x"722d3e63",
  2617 => x"6f6e7472",
  2618 => x"6f6c3a20",
  2619 => x"30780000",
  2620 => x"77726974",
  2621 => x"65206164",
  2622 => x"64726573",
  2623 => x"733a2030",
  2624 => x"78000000",
  2625 => x"20206c65",
  2626 => x"6e677468",
  2627 => x"3a203078",
  2628 => x"00000000",
  2629 => x"0a0a0000",
  2630 => x"72656164",
  2631 => x"20206164",
  2632 => x"64726573",
  2633 => x"733a2030",
  2634 => x"78000000",
  2635 => x"20206578",
  2636 => x"70656374",
  2637 => x"3a203078",
  2638 => x"00000000",
  2639 => x"2020676f",
  2640 => x"743a2030",
  2641 => x"78000000",
  2642 => x"20657272",
  2643 => x"6f720000",
  2644 => x"206f6b00",
  2645 => x"6d656d6f",
  2646 => x"72792074",
  2647 => x"65737420",
  2648 => x"696e6974",
  2649 => x"00000000",
  2650 => x"70686173",
  2651 => x"65207368",
  2652 => x"69667420",
  2653 => x"202d2020",
  2654 => x"76616c75",
  2655 => x"653a2000",
  2656 => x"20207374",
  2657 => x"61747573",
  2658 => x"3a203078",
  2659 => x"00000000",
  2660 => x"20202020",
  2661 => x"20000000",
  2662 => x"6f6b2020",
  2663 => x"00000000",
  2664 => x"4641494c",
  2665 => x"00000000",
  2666 => x"44445220",
  2667 => x"6d656d6f",
  2668 => x"72792069",
  2669 => x"6e666f00",
  2670 => x"0a0a6175",
  2671 => x"746f2074",
  2672 => x"5f524552",
  2673 => x"45534820",
  2674 => x"3a000000",
  2675 => x"0a636c6f",
  2676 => x"636b2065",
  2677 => x"6e61626c",
  2678 => x"6520203a",
  2679 => x"30780000",
  2680 => x"0a696e69",
  2681 => x"74616c69",
  2682 => x"7a652020",
  2683 => x"2020203a",
  2684 => x"30780000",
  2685 => x"0a636f6c",
  2686 => x"756d6e20",
  2687 => x"73697a65",
  2688 => x"2020203a",
  2689 => x"00000000",
  2690 => x"0a62616e",
  2691 => x"6b73697a",
  2692 => x"65202020",
  2693 => x"2020203a",
  2694 => x"00000000",
  2695 => x"4d627974",
  2696 => x"65000000",
  2697 => x"0a745f52",
  2698 => x"43442020",
  2699 => x"20202020",
  2700 => x"2020203a",
  2701 => x"00000000",
  2702 => x"0a745f52",
  2703 => x"46432020",
  2704 => x"20202020",
  2705 => x"2020203a",
  2706 => x"00000000",
  2707 => x"0a745f52",
  2708 => x"50202020",
  2709 => x"20202020",
  2710 => x"2020203a",
  2711 => x"00000000",
  2712 => x"0a726566",
  2713 => x"72657368",
  2714 => x"20656e2e",
  2715 => x"2020203a",
  2716 => x"30780000",
  2717 => x"0a0a4444",
  2718 => x"52206672",
  2719 => x"65717565",
  2720 => x"6e637920",
  2721 => x"3a000000",
  2722 => x"0a444452",
  2723 => x"20646174",
  2724 => x"61207769",
  2725 => x"6474683a",
  2726 => x"00000000",
  2727 => x"0a6d6f62",
  2728 => x"696c6520",
  2729 => x"73757070",
  2730 => x"6f72743a",
  2731 => x"30780000",
  2732 => x"0a0a7374",
  2733 => x"61747573",
  2734 => x"20726561",
  2735 => x"64202020",
  2736 => x"3a307800",
  2737 => x"0a0a7365",
  2738 => x"6c662072",
  2739 => x"65667265",
  2740 => x"73682020",
  2741 => x"3a000000",
  2742 => x"20353132",
  2743 => x"00000000",
  2744 => x"34303639",
  2745 => x"00000000",
  2746 => x"312f3800",
  2747 => x"20617272",
  2748 => x"61790000",
  2749 => x"0a74656d",
  2750 => x"702d636f",
  2751 => x"6d702072",
  2752 => x"6566723a",
  2753 => x"00000000",
  2754 => x"c2b04300",
  2755 => x"0a647269",
  2756 => x"76652073",
  2757 => x"7472656e",
  2758 => x"6774683a",
  2759 => x"00000000",
  2760 => x"0a706f77",
  2761 => x"65722073",
  2762 => x"6176696e",
  2763 => x"6720203a",
  2764 => x"00000000",
  2765 => x"756e6b6e",
  2766 => x"6f776e00",
  2767 => x"0a745f58",
  2768 => x"50202020",
  2769 => x"20202020",
  2770 => x"2020203a",
  2771 => x"00000000",
  2772 => x"0a745f58",
  2773 => x"53522020",
  2774 => x"20202020",
  2775 => x"2020203a",
  2776 => x"00000000",
  2777 => x"0a745f43",
  2778 => x"4b452020",
  2779 => x"20202020",
  2780 => x"2020203a",
  2781 => x"00000000",
  2782 => x"0a434153",
  2783 => x"206c6174",
  2784 => x"656e6379",
  2785 => x"2020203a",
  2786 => x"00000000",
  2787 => x"0a6d6f62",
  2788 => x"696c6520",
  2789 => x"656e6162",
  2790 => x"6c65643a",
  2791 => x"30780000",
  2792 => x"0a0a7068",
  2793 => x"7920636f",
  2794 => x"6e666967",
  2795 => x"20302020",
  2796 => x"3a307800",
  2797 => x"0a0a7068",
  2798 => x"7920636f",
  2799 => x"6e666967",
  2800 => x"20312020",
  2801 => x"3a307800",
  2802 => x"31303234",
  2803 => x"00000000",
  2804 => x"32303438",
  2805 => x"00000000",
  2806 => x"66756c6c",
  2807 => x"00000000",
  2808 => x"37300000",
  2809 => x"64656570",
  2810 => x"20706f77",
  2811 => x"65722064",
  2812 => x"6f776e00",
  2813 => x"636c6f63",
  2814 => x"6b207374",
  2815 => x"6f700000",
  2816 => x"73656c66",
  2817 => x"20726566",
  2818 => x"72657368",
  2819 => x"00000000",
  2820 => x"706f7765",
  2821 => x"7220646f",
  2822 => x"776e0000",
  2823 => x"6e6f6e65",
  2824 => x"00000000",
  2825 => x"312f3200",
  2826 => x"312f3400",
  2827 => x"312f3100",
  2828 => x"332f3400",
  2829 => x"38350000",
  2830 => x"34350000",
  2831 => x"68616c66",
  2832 => x"00000000",
  2833 => x"31350000",
  2834 => x"61646472",
  2835 => x"6573733a",
  2836 => x"20307800",
  2837 => x"20646174",
  2838 => x"613a2030",
  2839 => x"78000000",
  2840 => x"0a0a4443",
  2841 => x"4d207068",
  2842 => x"61736520",
  2843 => x"73686966",
  2844 => x"74207465",
  2845 => x"7374696e",
  2846 => x"67000000",
  2847 => x"0a696e69",
  2848 => x"7469616c",
  2849 => x"3a200000",
  2850 => x"676f2064",
  2851 => x"6f776e00",
  2852 => x"7363616e",
  2853 => x"2072616e",
  2854 => x"67650000",
  2855 => x"09000000",
  2856 => x"676f2074",
  2857 => x"6f206579",
  2858 => x"65000000",
  2859 => x"6c6f7720",
  2860 => x"666f756e",
  2861 => x"64000000",
  2862 => x"68696768",
  2863 => x"20666f75",
  2864 => x"6e640000",
  2865 => x"0a6c6f77",
  2866 => x"3a202020",
  2867 => x"20202020",
  2868 => x"20200000",
  2869 => x"0a686967",
  2870 => x"683a2020",
  2871 => x"20202020",
  2872 => x"20200000",
  2873 => x"0a646966",
  2874 => x"663a2020",
  2875 => x"20202020",
  2876 => x"20200000",
  2877 => x"0a6d696e",
  2878 => x"5f657272",
  2879 => x"3a202020",
  2880 => x"20200000",
  2881 => x"0a6d696e",
  2882 => x"5f657272",
  2883 => x"5f706f73",
  2884 => x"3a200000",
  2885 => x"676f206d",
  2886 => x"696e5f65",
  2887 => x"72726f72",
  2888 => x"00000000",
  2889 => x"0a66696e",
  2890 => x"616c3a20",
  2891 => x"20202020",
  2892 => x"20200000",
  2893 => x"64636d5f",
  2894 => x"74657374",
  2895 => x"5f707320",
  2896 => x"646f6e65",
  2897 => x"00000000",
  2898 => x"6c6f7720",
  2899 => x"4e4f5420",
  2900 => x"666f756e",
  2901 => x"64000000",
  2902 => x"68696768",
  2903 => x"204e4f54",
  2904 => x"20666f75",
  2905 => x"6e640000",
  2906 => x"676f207a",
  2907 => x"65726f00",
  2908 => x"64617461",
  2909 => x"2076616c",
  2910 => x"69640000",
  2911 => x"6c6f7720",
  2912 => x"20666f75",
  2913 => x"6e640000",
  2914 => x"0a646966",
  2915 => x"662f323a",
  2916 => x"20202020",
  2917 => x"20200000",
  2918 => x"6c6f7720",
  2919 => x"204e4f54",
  2920 => x"20666f75",
  2921 => x"6e640000",
  2922 => x"64617461",
  2923 => x"204e4f54",
  2924 => x"2076616c",
  2925 => x"69640000",
  2926 => x"74657374",
  2927 => x"2e632000",
  2928 => x"286f6e20",
  2929 => x"73696d29",
  2930 => x"0a000000",
  2931 => x"696e6974",
  2932 => x"20646f6e",
  2933 => x"652e0000",
  2934 => x"286f6e20",
  2935 => x"68617264",
  2936 => x"77617265",
  2937 => x"290a0000",
  2938 => x"636f6d70",
  2939 => x"696c6564",
  2940 => x"3a204a61",
  2941 => x"6e203234",
  2942 => x"20323031",
  2943 => x"31202031",
  2944 => x"333a3535",
  2945 => x"3a33330a",
  2946 => x"00000000",
  2947 => x"30622020",
  2948 => x"20202020",
  2949 => x"20202020",
  2950 => x"20202020",
  2951 => x"20202020",
  2952 => x"20202020",
  2953 => x"20202020",
  2954 => x"20202020",
  2955 => x"20200000",
  2956 => x"20202020",
  2957 => x"20202020",
  2958 => x"00000000",
  2959 => x"00202020",
  2960 => x"20202020",
  2961 => x"20202828",
  2962 => x"28282820",
  2963 => x"20202020",
  2964 => x"20202020",
  2965 => x"20202020",
  2966 => x"20202020",
  2967 => x"20881010",
  2968 => x"10101010",
  2969 => x"10101010",
  2970 => x"10101010",
  2971 => x"10040404",
  2972 => x"04040404",
  2973 => x"04040410",
  2974 => x"10101010",
  2975 => x"10104141",
  2976 => x"41414141",
  2977 => x"01010101",
  2978 => x"01010101",
  2979 => x"01010101",
  2980 => x"01010101",
  2981 => x"01010101",
  2982 => x"10101010",
  2983 => x"10104242",
  2984 => x"42424242",
  2985 => x"02020202",
  2986 => x"02020202",
  2987 => x"02020202",
  2988 => x"02020202",
  2989 => x"02020202",
  2990 => x"10101010",
  2991 => x"20000000",
  2992 => x"00000000",
  2993 => x"00000000",
  2994 => x"00000000",
  2995 => x"00000000",
  2996 => x"00000000",
  2997 => x"00000000",
  2998 => x"00000000",
  2999 => x"00000000",
  3000 => x"00000000",
  3001 => x"00000000",
  3002 => x"00000000",
  3003 => x"00000000",
  3004 => x"00000000",
  3005 => x"00000000",
  3006 => x"00000000",
  3007 => x"00000000",
  3008 => x"00000000",
  3009 => x"00000000",
  3010 => x"00000000",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"00000000",
  3015 => x"00000000",
  3016 => x"00000000",
  3017 => x"00000000",
  3018 => x"00000000",
  3019 => x"00000000",
  3020 => x"00000000",
  3021 => x"00000000",
  3022 => x"00000000",
  3023 => x"00000000",
  3024 => x"43000000",
  3025 => x"64756d6d",
  3026 => x"792e6578",
  3027 => x"65000000",
  3028 => x"00ffffff",
  3029 => x"ff00ffff",
  3030 => x"ffff00ff",
  3031 => x"ffffff00",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00003760",
  3036 => x"fff00000",
  3037 => x"80000d00",
  3038 => x"80000800",
  3039 => x"80000600",
  3040 => x"80000300",
  3041 => x"80000200",
  3042 => x"80000100",
  3043 => x"00002f90",
  3044 => x"00000000",
  3045 => x"000031f8",
  3046 => x"00003254",
  3047 => x"000032b0",
  3048 => x"00000000",
  3049 => x"00000000",
  3050 => x"00000000",
  3051 => x"00000000",
  3052 => x"00000000",
  3053 => x"00000000",
  3054 => x"00000000",
  3055 => x"00000000",
  3056 => x"00000000",
  3057 => x"00002f40",
  3058 => x"00000000",
  3059 => x"00000000",
  3060 => x"00000000",
  3061 => x"00000000",
  3062 => x"00000000",
  3063 => x"00000000",
  3064 => x"00000000",
  3065 => x"00000000",
  3066 => x"00000000",
  3067 => x"00000000",
  3068 => x"00000000",
  3069 => x"00000000",
  3070 => x"00000000",
  3071 => x"00000000",
  3072 => x"00000000",
  3073 => x"00000000",
  3074 => x"00000000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000000",
  3084 => x"00000000",
  3085 => x"00000000",
  3086 => x"00000001",
  3087 => x"330eabcd",
  3088 => x"1234e66d",
  3089 => x"deec0005",
  3090 => x"000b0000",
  3091 => x"00000000",
  3092 => x"00000000",
  3093 => x"00000000",
  3094 => x"00000000",
  3095 => x"00000000",
  3096 => x"00000000",
  3097 => x"00000000",
  3098 => x"00000000",
  3099 => x"00000000",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00000000",
  3103 => x"00000000",
  3104 => x"00000000",
  3105 => x"00000000",
  3106 => x"00000000",
  3107 => x"00000000",
  3108 => x"00000000",
  3109 => x"00000000",
  3110 => x"00000000",
  3111 => x"00000000",
  3112 => x"00000000",
  3113 => x"00000000",
  3114 => x"00000000",
  3115 => x"00000000",
  3116 => x"00000000",
  3117 => x"00000000",
  3118 => x"00000000",
  3119 => x"00000000",
  3120 => x"00000000",
  3121 => x"00000000",
  3122 => x"00000000",
  3123 => x"00000000",
  3124 => x"00000000",
  3125 => x"00000000",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000000",
  3151 => x"00000000",
  3152 => x"00000000",
  3153 => x"00000000",
  3154 => x"00000000",
  3155 => x"00000000",
  3156 => x"00000000",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"00000000",
  3161 => x"00000000",
  3162 => x"00000000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"00000000",
  3166 => x"00000000",
  3167 => x"00000000",
  3168 => x"00000000",
  3169 => x"00000000",
  3170 => x"00000000",
  3171 => x"00000000",
  3172 => x"00000000",
  3173 => x"00000000",
  3174 => x"00000000",
  3175 => x"00000000",
  3176 => x"00000000",
  3177 => x"00000000",
  3178 => x"00000000",
  3179 => x"00000000",
  3180 => x"00000000",
  3181 => x"00000000",
  3182 => x"00000000",
  3183 => x"00000000",
  3184 => x"00000000",
  3185 => x"00000000",
  3186 => x"00000000",
  3187 => x"00000000",
  3188 => x"00000000",
  3189 => x"00000000",
  3190 => x"00000000",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00000000",
  3195 => x"00000000",
  3196 => x"00000000",
  3197 => x"00000000",
  3198 => x"00000000",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"00000000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000000",
  3246 => x"00000000",
  3247 => x"00000000",
  3248 => x"00000000",
  3249 => x"00000000",
  3250 => x"00000000",
  3251 => x"00000000",
  3252 => x"00000000",
  3253 => x"00000000",
  3254 => x"00000000",
  3255 => x"00000000",
  3256 => x"00000000",
  3257 => x"00000000",
  3258 => x"00000000",
  3259 => x"00000000",
  3260 => x"00000000",
  3261 => x"00000000",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00000000",
  3265 => x"00000000",
  3266 => x"00000000",
  3267 => x"00000000",
  3268 => x"00000000",
  3269 => x"00000000",
  3270 => x"00000000",
  3271 => x"00000000",
  3272 => x"00000000",
  3273 => x"00000000",
  3274 => x"00000000",
  3275 => x"00000000",
  3276 => x"00000000",
  3277 => x"00000000",
  3278 => x"00000000",
  3279 => x"ffffffff",
  3280 => x"00000000",
  3281 => x"00020000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"00003348",
  3285 => x"00003348",
  3286 => x"00003350",
  3287 => x"00003350",
  3288 => x"00003358",
  3289 => x"00003358",
  3290 => x"00003360",
  3291 => x"00003360",
  3292 => x"00003368",
  3293 => x"00003368",
  3294 => x"00003370",
  3295 => x"00003370",
  3296 => x"00003378",
  3297 => x"00003378",
  3298 => x"00003380",
  3299 => x"00003380",
  3300 => x"00003388",
  3301 => x"00003388",
  3302 => x"00003390",
  3303 => x"00003390",
  3304 => x"00003398",
  3305 => x"00003398",
  3306 => x"000033a0",
  3307 => x"000033a0",
  3308 => x"000033a8",
  3309 => x"000033a8",
  3310 => x"000033b0",
  3311 => x"000033b0",
  3312 => x"000033b8",
  3313 => x"000033b8",
  3314 => x"000033c0",
  3315 => x"000033c0",
  3316 => x"000033c8",
  3317 => x"000033c8",
  3318 => x"000033d0",
  3319 => x"000033d0",
  3320 => x"000033d8",
  3321 => x"000033d8",
  3322 => x"000033e0",
  3323 => x"000033e0",
  3324 => x"000033e8",
  3325 => x"000033e8",
  3326 => x"000033f0",
  3327 => x"000033f0",
  3328 => x"000033f8",
  3329 => x"000033f8",
  3330 => x"00003400",
  3331 => x"00003400",
  3332 => x"00003408",
  3333 => x"00003408",
  3334 => x"00003410",
  3335 => x"00003410",
  3336 => x"00003418",
  3337 => x"00003418",
  3338 => x"00003420",
  3339 => x"00003420",
  3340 => x"00003428",
  3341 => x"00003428",
  3342 => x"00003430",
  3343 => x"00003430",
  3344 => x"00003438",
  3345 => x"00003438",
  3346 => x"00003440",
  3347 => x"00003440",
  3348 => x"00003448",
  3349 => x"00003448",
  3350 => x"00003450",
  3351 => x"00003450",
  3352 => x"00003458",
  3353 => x"00003458",
  3354 => x"00003460",
  3355 => x"00003460",
  3356 => x"00003468",
  3357 => x"00003468",
  3358 => x"00003470",
  3359 => x"00003470",
  3360 => x"00003478",
  3361 => x"00003478",
  3362 => x"00003480",
  3363 => x"00003480",
  3364 => x"00003488",
  3365 => x"00003488",
  3366 => x"00003490",
  3367 => x"00003490",
  3368 => x"00003498",
  3369 => x"00003498",
  3370 => x"000034a0",
  3371 => x"000034a0",
  3372 => x"000034a8",
  3373 => x"000034a8",
  3374 => x"000034b0",
  3375 => x"000034b0",
  3376 => x"000034b8",
  3377 => x"000034b8",
  3378 => x"000034c0",
  3379 => x"000034c0",
  3380 => x"000034c8",
  3381 => x"000034c8",
  3382 => x"000034d0",
  3383 => x"000034d0",
  3384 => x"000034d8",
  3385 => x"000034d8",
  3386 => x"000034e0",
  3387 => x"000034e0",
  3388 => x"000034e8",
  3389 => x"000034e8",
  3390 => x"000034f0",
  3391 => x"000034f0",
  3392 => x"000034f8",
  3393 => x"000034f8",
  3394 => x"00003500",
  3395 => x"00003500",
  3396 => x"00003508",
  3397 => x"00003508",
  3398 => x"00003510",
  3399 => x"00003510",
  3400 => x"00003518",
  3401 => x"00003518",
  3402 => x"00003520",
  3403 => x"00003520",
  3404 => x"00003528",
  3405 => x"00003528",
  3406 => x"00003530",
  3407 => x"00003530",
  3408 => x"00003538",
  3409 => x"00003538",
  3410 => x"00003540",
  3411 => x"00003540",
  3412 => x"00003548",
  3413 => x"00003548",
  3414 => x"00003550",
  3415 => x"00003550",
  3416 => x"00003558",
  3417 => x"00003558",
  3418 => x"00003560",
  3419 => x"00003560",
  3420 => x"00003568",
  3421 => x"00003568",
  3422 => x"00003570",
  3423 => x"00003570",
  3424 => x"00003578",
  3425 => x"00003578",
  3426 => x"00003580",
  3427 => x"00003580",
  3428 => x"00003588",
  3429 => x"00003588",
  3430 => x"00003590",
  3431 => x"00003590",
  3432 => x"00003598",
  3433 => x"00003598",
  3434 => x"000035a0",
  3435 => x"000035a0",
  3436 => x"000035a8",
  3437 => x"000035a8",
  3438 => x"000035b0",
  3439 => x"000035b0",
  3440 => x"000035b8",
  3441 => x"000035b8",
  3442 => x"000035c0",
  3443 => x"000035c0",
  3444 => x"000035c8",
  3445 => x"000035c8",
  3446 => x"000035d0",
  3447 => x"000035d0",
  3448 => x"000035d8",
  3449 => x"000035d8",
  3450 => x"000035e0",
  3451 => x"000035e0",
  3452 => x"000035e8",
  3453 => x"000035e8",
  3454 => x"000035f0",
  3455 => x"000035f0",
  3456 => x"000035f8",
  3457 => x"000035f8",
  3458 => x"00003600",
  3459 => x"00003600",
  3460 => x"00003608",
  3461 => x"00003608",
  3462 => x"00003610",
  3463 => x"00003610",
  3464 => x"00003618",
  3465 => x"00003618",
  3466 => x"00003620",
  3467 => x"00003620",
  3468 => x"00003628",
  3469 => x"00003628",
  3470 => x"00003630",
  3471 => x"00003630",
  3472 => x"00003638",
  3473 => x"00003638",
  3474 => x"00003640",
  3475 => x"00003640",
  3476 => x"00003648",
  3477 => x"00003648",
  3478 => x"00003650",
  3479 => x"00003650",
  3480 => x"00003658",
  3481 => x"00003658",
  3482 => x"00003660",
  3483 => x"00003660",
  3484 => x"00003668",
  3485 => x"00003668",
  3486 => x"00003670",
  3487 => x"00003670",
  3488 => x"00003678",
  3489 => x"00003678",
  3490 => x"00003680",
  3491 => x"00003680",
  3492 => x"00003688",
  3493 => x"00003688",
  3494 => x"00003690",
  3495 => x"00003690",
  3496 => x"00003698",
  3497 => x"00003698",
  3498 => x"000036a0",
  3499 => x"000036a0",
  3500 => x"000036a8",
  3501 => x"000036a8",
  3502 => x"000036b0",
  3503 => x"000036b0",
  3504 => x"000036b8",
  3505 => x"000036b8",
  3506 => x"000036c0",
  3507 => x"000036c0",
  3508 => x"000036c8",
  3509 => x"000036c8",
  3510 => x"000036d0",
  3511 => x"000036d0",
  3512 => x"000036d8",
  3513 => x"000036d8",
  3514 => x"000036e0",
  3515 => x"000036e0",
  3516 => x"000036e8",
  3517 => x"000036e8",
  3518 => x"000036f0",
  3519 => x"000036f0",
  3520 => x"000036f8",
  3521 => x"000036f8",
  3522 => x"00003700",
  3523 => x"00003700",
  3524 => x"00003708",
  3525 => x"00003708",
  3526 => x"00003710",
  3527 => x"00003710",
  3528 => x"00003718",
  3529 => x"00003718",
  3530 => x"00003720",
  3531 => x"00003720",
  3532 => x"00003728",
  3533 => x"00003728",
  3534 => x"00003730",
  3535 => x"00003730",
  3536 => x"00003738",
  3537 => x"00003738",
  3538 => x"00003740",
  3539 => x"00003740",
  3540 => x"00002f44",
  3541 => x"ffffffff",
  3542 => x"00000000",
  3543 => x"ffffffff",
  3544 => x"00000000",
  3545 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
