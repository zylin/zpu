-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"82cb940c",
     3 => x"3a0b0b82",
     4 => x"a5be0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"82a68b2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b82cb",
   162 => x"80738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80dc",
   171 => x"c62d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80dd",
   179 => x"f82d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"82cb900c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82c73f82",
   257 => x"babe3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"fe3d0d0b",
   281 => x"0b82dbb8",
   282 => x"08538413",
   283 => x"0870882a",
   284 => x"70810651",
   285 => x"52527080",
   286 => x"2ef03871",
   287 => x"81ff0680",
   288 => x"0c843d0d",
   289 => x"04ff3d0d",
   290 => x"0b0b82db",
   291 => x"b8085271",
   292 => x"0870882a",
   293 => x"81327081",
   294 => x"06515151",
   295 => x"70f13873",
   296 => x"720c833d",
   297 => x"0d0482cb",
   298 => x"9008802e",
   299 => x"a43882cb",
   300 => x"9408822e",
   301 => x"bd388380",
   302 => x"800b0b0b",
   303 => x"82dbb80c",
   304 => x"82a0800b",
   305 => x"82dbbc0c",
   306 => x"8290800b",
   307 => x"82dbc00c",
   308 => x"04f88080",
   309 => x"80a40b0b",
   310 => x"0b82dbb8",
   311 => x"0cf88080",
   312 => x"82800b82",
   313 => x"dbbc0cf8",
   314 => x"80808480",
   315 => x"0b82dbc0",
   316 => x"0c0480c0",
   317 => x"a8808c0b",
   318 => x"0b0b82db",
   319 => x"b80c80c0",
   320 => x"a880940b",
   321 => x"82dbbc0c",
   322 => x"0b0b82c2",
   323 => x"f00b82db",
   324 => x"c00c04ff",
   325 => x"3d0d82db",
   326 => x"c4335170",
   327 => x"a73882cb",
   328 => x"9c087008",
   329 => x"52527080",
   330 => x"2e943884",
   331 => x"1282cb9c",
   332 => x"0c702d82",
   333 => x"cb9c0870",
   334 => x"08525270",
   335 => x"ee38810b",
   336 => x"82dbc434",
   337 => x"833d0d04",
   338 => x"04803d0d",
   339 => x"0b0b82db",
   340 => x"b408802e",
   341 => x"8e380b0b",
   342 => x"0b0b800b",
   343 => x"802e0981",
   344 => x"06853882",
   345 => x"3d0d040b",
   346 => x"0b82dbb4",
   347 => x"510b0b0b",
   348 => x"f58e3f82",
   349 => x"3d0d0404",
   350 => x"f63d0d7c",
   351 => x"729b2a81",
   352 => x"068c120c",
   353 => x"739f2a70",
   354 => x"94130c53",
   355 => x"55719138",
   356 => x"74085880",
   357 => x"c0780c72",
   358 => x"862a8106",
   359 => x"5271fe38",
   360 => x"728b2a9f",
   361 => x"0690160c",
   362 => x"90805180",
   363 => x"f0a63f80",
   364 => x"08888005",
   365 => x"f8800670",
   366 => x"535480ff",
   367 => x"5380720c",
   368 => x"8812ff14",
   369 => x"54527280",
   370 => x"25f33873",
   371 => x"98160c90",
   372 => x"805180ef",
   373 => x"ff3f8008",
   374 => x"888005f8",
   375 => x"80067053",
   376 => x"5480ff53",
   377 => x"80720c88",
   378 => x"12ff1454",
   379 => x"52728025",
   380 => x"f338739c",
   381 => x"160c7408",
   382 => x"94119817",
   383 => x"08710c59",
   384 => x"98117571",
   385 => x"0c545680",
   386 => x"0ba0160c",
   387 => x"800ba416",
   388 => x"0c800ba8",
   389 => x"160c800b",
   390 => x"ac160c94",
   391 => x"150882ff",
   392 => x"38901508",
   393 => x"77832a81",
   394 => x"06535371",
   395 => x"fe38728b",
   396 => x"2bf88080",
   397 => x"80810790",
   398 => x"1759780c",
   399 => x"76832a81",
   400 => x"065271fe",
   401 => x"3876832a",
   402 => x"707a842a",
   403 => x"56585890",
   404 => x"15087881",
   405 => x"06535371",
   406 => x"fe38728b",
   407 => x"2b820790",
   408 => x"1753720c",
   409 => x"76810652",
   410 => x"71fe3873",
   411 => x"81067990",
   412 => x"2a545271",
   413 => x"802e8338",
   414 => x"ff53728f",
   415 => x"2a708106",
   416 => x"515271cb",
   417 => x"3871738c",
   418 => x"2a810658",
   419 => x"5476802e",
   420 => x"80cc3878",
   421 => x"832a7a83",
   422 => x"2a7b842a",
   423 => x"59595990",
   424 => x"15087981",
   425 => x"06535371",
   426 => x"fe38728b",
   427 => x"2b80c207",
   428 => x"90175372",
   429 => x"0c778106",
   430 => x"5271fe38",
   431 => x"7681067a",
   432 => x"902a5452",
   433 => x"71802e83",
   434 => x"38ff5372",
   435 => x"852a8106",
   436 => x"53728b38",
   437 => x"81145483",
   438 => x"86d07425",
   439 => x"c2389015",
   440 => x"087a832a",
   441 => x"81065353",
   442 => x"71fe3872",
   443 => x"8b2b8207",
   444 => x"90175877",
   445 => x"0c79832a",
   446 => x"81065271",
   447 => x"fe387984",
   448 => x"2a81067a",
   449 => x"902a5452",
   450 => x"71802e83",
   451 => x"38ff5372",
   452 => x"8d2a548c",
   453 => x"1508802e",
   454 => x"81ab3873",
   455 => x"81065776",
   456 => x"81a33872",
   457 => x"862a8106",
   458 => x"5978802e",
   459 => x"81973881",
   460 => x"775b5b72",
   461 => x"842a9006",
   462 => x"7a872b07",
   463 => x"7b882b07",
   464 => x"760c8415",
   465 => x"5a811a33",
   466 => x"85163482",
   467 => x"1a338616",
   468 => x"34831a33",
   469 => x"87163484",
   470 => x"1a338816",
   471 => x"34851a33",
   472 => x"89163488",
   473 => x"167a3381",
   474 => x"1c337188",
   475 => x"2b07720c",
   476 => x"8c18821d",
   477 => x"33831e33",
   478 => x"71982b71",
   479 => x"902b077f",
   480 => x"84053370",
   481 => x"882b7207",
   482 => x"61850533",
   483 => x"71077077",
   484 => x"0c800c5d",
   485 => x"59595c5e",
   486 => x"5256598c",
   487 => x"3d0d0480",
   488 => x"77832a81",
   489 => x"065c537a",
   490 => x"732e0981",
   491 => x"06953881",
   492 => x"13537282",
   493 => x"24ff8b38",
   494 => x"81135382",
   495 => x"7325f038",
   496 => x"ff8039ff",
   497 => x"39738106",
   498 => x"5776802e",
   499 => x"a2387286",
   500 => x"2a708106",
   501 => x"51527197",
   502 => x"38715b81",
   503 => x"73842a90",
   504 => x"0671872b",
   505 => x"077c882b",
   506 => x"07770c5a",
   507 => x"fed43973",
   508 => x"81065978",
   509 => x"febd3872",
   510 => x"862a8106",
   511 => x"5271feb3",
   512 => x"38717274",
   513 => x"842a9006",
   514 => x"71872b07",
   515 => x"72882b07",
   516 => x"780c5b5b",
   517 => x"feac39fb",
   518 => x"3d0d777a",
   519 => x"728b2c81",
   520 => x"06565455",
   521 => x"80517371",
   522 => x"2e098106",
   523 => x"b9389813",
   524 => x"08a01408",
   525 => x"10101011",
   526 => x"7a84120c",
   527 => x"52a01408",
   528 => x"52527080",
   529 => x"ff2ea638",
   530 => x"70101010",
   531 => x"12759080",
   532 => x"07710c54",
   533 => x"a0130881",
   534 => x"05a0140c",
   535 => x"72087681",
   536 => x"07710c55",
   537 => x"81517080",
   538 => x"0c873d0d",
   539 => x"0487f812",
   540 => x"75b08007",
   541 => x"710c5273",
   542 => x"a0140c72",
   543 => x"08768107",
   544 => x"710c5581",
   545 => x"51e039fc",
   546 => x"ee3d0df8",
   547 => x"80809680",
   548 => x"0b82dbc8",
   549 => x"0c800b9a",
   550 => x"3d349302",
   551 => x"840580e1",
   552 => x"053480f2",
   553 => x"02840580",
   554 => x"e20534ff",
   555 => x"ae028405",
   556 => x"80e30534",
   557 => x"80f20b9b",
   558 => x"3d34a102",
   559 => x"840580e5",
   560 => x"0534de02",
   561 => x"840580e6",
   562 => x"0534ffad",
   563 => x"02840580",
   564 => x"e70534ff",
   565 => x"be0b9c3d",
   566 => x"34ef0284",
   567 => x"0580e905",
   568 => x"34800284",
   569 => x"0580ea05",
   570 => x"34a00284",
   571 => x"0580eb05",
   572 => x"34850b9d",
   573 => x"3d34dc02",
   574 => x"840580ed",
   575 => x"05348653",
   576 => x"83943df4",
   577 => x"9a055282",
   578 => x"dbcc5180",
   579 => x"f5df3f80",
   580 => x"5b8e0b9a",
   581 => x"3d5e5c7b",
   582 => x"1d5a7b7a",
   583 => x"34811c7c",
   584 => x"71267c05",
   585 => x"70725f5d",
   586 => x"5a5a7880",
   587 => x"268a3878",
   588 => x"e6388be9",
   589 => x"7a27e038",
   590 => x"82dbc851",
   591 => x"f8ba3f02",
   592 => x"80e50533",
   593 => x"579a3d33",
   594 => x"560280e3",
   595 => x"05335502",
   596 => x"80e20533",
   597 => x"540280e1",
   598 => x"05335399",
   599 => x"3d335282",
   600 => x"c2f45180",
   601 => x"f6b93f84",
   602 => x"d53f8008",
   603 => x"40805d80",
   604 => x"0b9a3d40",
   605 => x"5e82dbc8",
   606 => x"537e528b",
   607 => x"ea51fd97",
   608 => x"3f80089f",
   609 => x"2c80081f",
   610 => x"7f71265b",
   611 => x"5d7d0570",
   612 => x"1a707e41",
   613 => x"5f515b7a",
   614 => x"80268b38",
   615 => x"7ad738bf",
   616 => x"ffff7c27",
   617 => x"d0388496",
   618 => x"3f800860",
   619 => x"31705383",
   620 => x"953df48c",
   621 => x"05525c80",
   622 => x"c7913f66",
   623 => x"685c5a80",
   624 => x"7c2480f8",
   625 => x"388be282",
   626 => x"0a5e807e",
   627 => x"55557952",
   628 => x"7a538394",
   629 => x"3df3fc05",
   630 => x"51b6c13f",
   631 => x"62647154",
   632 => x"705582c3",
   633 => x"b8535c5a",
   634 => x"80f5b43f",
   635 => x"80588078",
   636 => x"5454825c",
   637 => x"80f70a7c",
   638 => x"525285fa",
   639 => x"3f913d7a",
   640 => x"557b565c",
   641 => x"bbc0c20a",
   642 => x"5e807e53",
   643 => x"537b51b6",
   644 => x"8b3f9afc",
   645 => x"0a5f807f",
   646 => x"55556062",
   647 => x"5b527953",
   648 => x"7b5198e9",
   649 => x"3f60625c",
   650 => x"527a5382",
   651 => x"c3c45180",
   652 => x"f4ed3f80",
   653 => x"0b800c83",
   654 => x"943d0d04",
   655 => x"9f820a5e",
   656 => x"807e5555",
   657 => x"79527a53",
   658 => x"83943df4",
   659 => x"84055195",
   660 => x"f63f6466",
   661 => x"5c5a8be2",
   662 => x"820a5e80",
   663 => x"7e555579",
   664 => x"527a5383",
   665 => x"943df3fc",
   666 => x"0551b5b0",
   667 => x"3f626471",
   668 => x"54705582",
   669 => x"c3b8535c",
   670 => x"5a80f4a3",
   671 => x"3f805880",
   672 => x"78545482",
   673 => x"5c80f70a",
   674 => x"7c525284",
   675 => x"e93f913d",
   676 => x"7a557b56",
   677 => x"5cbbc0c2",
   678 => x"0a5e807e",
   679 => x"53537b51",
   680 => x"b4fa3f9a",
   681 => x"fc0a5f80",
   682 => x"7f555560",
   683 => x"625b5279",
   684 => x"537b5197",
   685 => x"d83f6062",
   686 => x"5c527a53",
   687 => x"82c3c451",
   688 => x"80f3dc3f",
   689 => x"800b800c",
   690 => x"83943d0d",
   691 => x"04ff3d0d",
   692 => x"82cbb408",
   693 => x"74101075",
   694 => x"10059412",
   695 => x"0c52850b",
   696 => x"98130c98",
   697 => x"12087081",
   698 => x"06515170",
   699 => x"f638833d",
   700 => x"0d04fd3d",
   701 => x"0d82cbb4",
   702 => x"0876b0ea",
   703 => x"2994120c",
   704 => x"54850b98",
   705 => x"150c9814",
   706 => x"08708106",
   707 => x"515372f6",
   708 => x"38853d0d",
   709 => x"04fb3d0d",
   710 => x"77568055",
   711 => x"74762781",
   712 => x"993882cb",
   713 => x"b40854bf",
   714 => x"a9bc0b94",
   715 => x"150c850b",
   716 => x"98150c98",
   717 => x"14087081",
   718 => x"06515372",
   719 => x"f638bfa9",
   720 => x"bc0b9415",
   721 => x"0c850b98",
   722 => x"150c9814",
   723 => x"08708106",
   724 => x"515372f6",
   725 => x"38bfa9bc",
   726 => x"0b94150c",
   727 => x"850b9815",
   728 => x"0c981408",
   729 => x"70810651",
   730 => x"5372f638",
   731 => x"bfa9bc0b",
   732 => x"94150c85",
   733 => x"0b98150c",
   734 => x"98140870",
   735 => x"81065153",
   736 => x"72f638bf",
   737 => x"a9bc0b94",
   738 => x"150c850b",
   739 => x"98150c98",
   740 => x"14087081",
   741 => x"06515372",
   742 => x"f638bfa9",
   743 => x"bc0b9415",
   744 => x"0c850b98",
   745 => x"150c9814",
   746 => x"08708106",
   747 => x"515372f6",
   748 => x"38811555",
   749 => x"757526fe",
   750 => x"ee38873d",
   751 => x"0d04803d",
   752 => x"0d82cbb4",
   753 => x"08a01108",
   754 => x"800c5182",
   755 => x"3d0d0480",
   756 => x"3d0d7251",
   757 => x"80712787",
   758 => x"38ff1151",
   759 => x"70fb3882",
   760 => x"3d0d0480",
   761 => x"3d0d82cb",
   762 => x"b4085187",
   763 => x"0b84120c",
   764 => x"b0ea0ba4",
   765 => x"120c870b",
   766 => x"a8120c82",
   767 => x"3d0d048c",
   768 => x"08028c0c",
   769 => x"f53d0d8c",
   770 => x"08940508",
   771 => x"9d388c08",
   772 => x"8c05088c",
   773 => x"08900508",
   774 => x"8c088805",
   775 => x"08585654",
   776 => x"73760c74",
   777 => x"84170c81",
   778 => x"c039800b",
   779 => x"8c08f005",
   780 => x"0c800b8c",
   781 => x"08f4050c",
   782 => x"8c088c05",
   783 => x"088c0890",
   784 => x"05085654",
   785 => x"738c08f0",
   786 => x"050c748c",
   787 => x"08f4050c",
   788 => x"8c08f805",
   789 => x"8c08f005",
   790 => x"56568870",
   791 => x"54755376",
   792 => x"525480ef",
   793 => x"883fa00b",
   794 => x"8c089405",
   795 => x"08318c08",
   796 => x"ec050c8c",
   797 => x"08ec0508",
   798 => x"80249d38",
   799 => x"800b8c08",
   800 => x"f4050c8c",
   801 => x"08ec0508",
   802 => x"308c08fc",
   803 => x"0508712b",
   804 => x"8c08f005",
   805 => x"0c54b939",
   806 => x"8c08fc05",
   807 => x"088c08ec",
   808 => x"05082a8c",
   809 => x"08e8050c",
   810 => x"8c08fc05",
   811 => x"088c0894",
   812 => x"05082b8c",
   813 => x"08f4050c",
   814 => x"8c08f805",
   815 => x"088c0894",
   816 => x"05082b70",
   817 => x"8c08e805",
   818 => x"08078c08",
   819 => x"f0050c54",
   820 => x"8c08f005",
   821 => x"088c08f4",
   822 => x"05088c08",
   823 => x"88050858",
   824 => x"56547376",
   825 => x"0c748417",
   826 => x"0c8c0888",
   827 => x"0508800c",
   828 => x"8d3d0d8c",
   829 => x"0c048c08",
   830 => x"028c0cf4",
   831 => x"3d0d800b",
   832 => x"8c08f005",
   833 => x"0c800b8c",
   834 => x"08f4050c",
   835 => x"8c088805",
   836 => x"088c088c",
   837 => x"05085654",
   838 => x"738c08f0",
   839 => x"050c748c",
   840 => x"08f4050c",
   841 => x"8c08f805",
   842 => x"8c08f005",
   843 => x"56568870",
   844 => x"54755376",
   845 => x"525480ed",
   846 => x"b43f800b",
   847 => x"8c08e805",
   848 => x"0c800b8c",
   849 => x"08ec050c",
   850 => x"8c089005",
   851 => x"088c0894",
   852 => x"05085654",
   853 => x"738c08e8",
   854 => x"050c748c",
   855 => x"08ec050c",
   856 => x"8c08f005",
   857 => x"8c08e805",
   858 => x"56568870",
   859 => x"54755376",
   860 => x"525480ec",
   861 => x"f83f8c08",
   862 => x"f805088c",
   863 => x"08f00508",
   864 => x"258b3880",
   865 => x"0b8c08e4",
   866 => x"050c80ca",
   867 => x"398c08f0",
   868 => x"05088c08",
   869 => x"f8050825",
   870 => x"8a38820b",
   871 => x"8c08e405",
   872 => x"0cb4398c",
   873 => x"08fc0508",
   874 => x"8c08f405",
   875 => x"08278a38",
   876 => x"800b8c08",
   877 => x"e4050c9e",
   878 => x"398c08f4",
   879 => x"05088c08",
   880 => x"fc050827",
   881 => x"8a38820b",
   882 => x"8c08e405",
   883 => x"0c883981",
   884 => x"0b8c08e4",
   885 => x"050c8c08",
   886 => x"e4050880",
   887 => x"0c8e3d0d",
   888 => x"8c0c048c",
   889 => x"08028c0c",
   890 => x"d43d0d8c",
   891 => x"08880508",
   892 => x"518e953f",
   893 => x"80085473",
   894 => x"802e9038",
   895 => x"8c088805",
   896 => x"08708c08",
   897 => x"d0050c54",
   898 => x"8cf4398c",
   899 => x"088c0508",
   900 => x"518df53f",
   901 => x"80085473",
   902 => x"802e9038",
   903 => x"8c088c05",
   904 => x"08708c08",
   905 => x"d0050c54",
   906 => x"8cd4398c",
   907 => x"08880508",
   908 => x"518da13f",
   909 => x"80085473",
   910 => x"802e80c5",
   911 => x"388c088c",
   912 => x"0508518d",
   913 => x"8f3f8008",
   914 => x"5473802e",
   915 => x"a5388c08",
   916 => x"8805088c",
   917 => x"088c0508",
   918 => x"55558415",
   919 => x"08841508",
   920 => x"2e90388c",
   921 => x"da3f8008",
   922 => x"708c08d0",
   923 => x"050c548c",
   924 => x"8d398c08",
   925 => x"88050870",
   926 => x"8c08d005",
   927 => x"0c548bfe",
   928 => x"398c088c",
   929 => x"0508518c",
   930 => x"cb3f8008",
   931 => x"5473802e",
   932 => x"90388c08",
   933 => x"8c050870",
   934 => x"8c08d005",
   935 => x"0c548bde",
   936 => x"398c088c",
   937 => x"0508518b",
   938 => x"e23f8008",
   939 => x"5473802e",
   940 => x"80e7388c",
   941 => x"08880508",
   942 => x"518bd03f",
   943 => x"80085473",
   944 => x"802e80c6",
   945 => x"388c0890",
   946 => x"05088c08",
   947 => x"88050871",
   948 => x"58565494",
   949 => x"70547553",
   950 => x"76525480",
   951 => x"ea8f3f8c",
   952 => x"08900508",
   953 => x"8c088805",
   954 => x"088c088c",
   955 => x"05088412",
   956 => x"08841208",
   957 => x"0684140c",
   958 => x"8c089005",
   959 => x"08708c08",
   960 => x"d0050c51",
   961 => x"5656568a",
   962 => x"f5398c08",
   963 => x"88050870",
   964 => x"8c08d005",
   965 => x"0c548ae6",
   966 => x"398c0888",
   967 => x"0508518a",
   968 => x"ea3f8008",
   969 => x"5473802e",
   970 => x"90388c08",
   971 => x"8c050870",
   972 => x"8c08d005",
   973 => x"0c548ac6",
   974 => x"398c0888",
   975 => x"05088811",
   976 => x"088c08f4",
   977 => x"050c8c08",
   978 => x"8c050888",
   979 => x"11088c08",
   980 => x"f0050c8c",
   981 => x"08880508",
   982 => x"51515490",
   983 => x"14088c15",
   984 => x"08555573",
   985 => x"8c08e805",
   986 => x"0c748c08",
   987 => x"ec050c8c",
   988 => x"088c0508",
   989 => x"54901408",
   990 => x"8c150855",
   991 => x"55738c08",
   992 => x"e0050c74",
   993 => x"8c08e405",
   994 => x"0c8c08f4",
   995 => x"05088c08",
   996 => x"f0050831",
   997 => x"8c08dc05",
   998 => x"0c8c08dc",
   999 => x"05088025",
  1000 => x"8c388c08",
  1001 => x"dc050830",
  1002 => x"8c08dc05",
  1003 => x"0c8c08dc",
  1004 => x"0508bf24",
  1005 => x"81b3388c",
  1006 => x"08f00508",
  1007 => x"8c08f405",
  1008 => x"082580cc",
  1009 => x"388c08f0",
  1010 => x"05088105",
  1011 => x"8c08f005",
  1012 => x"0c8c08e0",
  1013 => x"05088006",
  1014 => x"8c08e405",
  1015 => x"0881068c",
  1016 => x"08e00508",
  1017 => x"9f2b8c08",
  1018 => x"e4050881",
  1019 => x"2a707207",
  1020 => x"8c08e005",
  1021 => x"08812a70",
  1022 => x"76078c08",
  1023 => x"e0050c74",
  1024 => x"72078c08",
  1025 => x"e4050c59",
  1026 => x"595b5b58",
  1027 => x"56ffa839",
  1028 => x"8c08f405",
  1029 => x"088c08f0",
  1030 => x"05082581",
  1031 => x"8f388c08",
  1032 => x"f4050881",
  1033 => x"058c08f4",
  1034 => x"050c8c08",
  1035 => x"e8050880",
  1036 => x"068c08ec",
  1037 => x"05088106",
  1038 => x"8c08e805",
  1039 => x"089f2b8c",
  1040 => x"08ec0508",
  1041 => x"812a7072",
  1042 => x"078c08e8",
  1043 => x"0508812a",
  1044 => x"7076078c",
  1045 => x"08e8050c",
  1046 => x"7472078c",
  1047 => x"08ec050c",
  1048 => x"59595b5b",
  1049 => x"5856ffa8",
  1050 => x"398c08f0",
  1051 => x"05088c08",
  1052 => x"f4050825",
  1053 => x"9d388c08",
  1054 => x"f405088c",
  1055 => x"08f0050c",
  1056 => x"80548055",
  1057 => x"738c08e0",
  1058 => x"050c748c",
  1059 => x"08e4050c",
  1060 => x"9b398c08",
  1061 => x"f005088c",
  1062 => x"08f4050c",
  1063 => x"80548055",
  1064 => x"738c08e8",
  1065 => x"050c748c",
  1066 => x"08ec050c",
  1067 => x"8c088805",
  1068 => x"088c088c",
  1069 => x"05085555",
  1070 => x"84150884",
  1071 => x"15082e84",
  1072 => x"e4388c08",
  1073 => x"88050854",
  1074 => x"84140880",
  1075 => x"2e81b538",
  1076 => x"8c08e005",
  1077 => x"088c08e4",
  1078 => x"05085654",
  1079 => x"738c08c8",
  1080 => x"050c748c",
  1081 => x"08cc050c",
  1082 => x"8c08e805",
  1083 => x"088c08ec",
  1084 => x"05085755",
  1085 => x"748c08c0",
  1086 => x"050c758c",
  1087 => x"08c4050c",
  1088 => x"8c08cc05",
  1089 => x"088c08c4",
  1090 => x"05087171",
  1091 => x"31708c08",
  1092 => x"ffbc050c",
  1093 => x"52555681",
  1094 => x"0b8c08ff",
  1095 => x"b4050c8c",
  1096 => x"08ffbc05",
  1097 => x"088c08cc",
  1098 => x"05085755",
  1099 => x"74762689",
  1100 => x"38800b8c",
  1101 => x"08ffb405",
  1102 => x"0c8c08c8",
  1103 => x"05088c08",
  1104 => x"c0050871",
  1105 => x"7131708c",
  1106 => x"08ffb805",
  1107 => x"0c8c08ff",
  1108 => x"b8050870",
  1109 => x"8c08ffb4",
  1110 => x"05083170",
  1111 => x"8c08ffb8",
  1112 => x"050c5259",
  1113 => x"5256548c",
  1114 => x"08ffb805",
  1115 => x"088c08ff",
  1116 => x"bc050856",
  1117 => x"54738c08",
  1118 => x"f8050c74",
  1119 => x"8c08fc05",
  1120 => x"0c81bb39",
  1121 => x"8c08e805",
  1122 => x"088c08ec",
  1123 => x"05085755",
  1124 => x"748c08ff",
  1125 => x"ac050c75",
  1126 => x"8c08ffb0",
  1127 => x"050c8c08",
  1128 => x"e005088c",
  1129 => x"08e40508",
  1130 => x"5654738c",
  1131 => x"08ffa405",
  1132 => x"0c748c08",
  1133 => x"ffa8050c",
  1134 => x"8c08ffb0",
  1135 => x"05088c08",
  1136 => x"ffa80508",
  1137 => x"71713170",
  1138 => x"8c08ffa0",
  1139 => x"050c5257",
  1140 => x"55810b8c",
  1141 => x"08ff9805",
  1142 => x"0c8c08ff",
  1143 => x"a005088c",
  1144 => x"08ffb005",
  1145 => x"08565473",
  1146 => x"75268938",
  1147 => x"800b8c08",
  1148 => x"ff98050c",
  1149 => x"8c08ffac",
  1150 => x"05088c08",
  1151 => x"ffa40508",
  1152 => x"71713170",
  1153 => x"8c08ff9c",
  1154 => x"050c8c08",
  1155 => x"ff9c0508",
  1156 => x"708c08ff",
  1157 => x"98050831",
  1158 => x"708c08ff",
  1159 => x"9c050c53",
  1160 => x"58525556",
  1161 => x"8c08ff9c",
  1162 => x"05088c08",
  1163 => x"ffa00508",
  1164 => x"5654738c",
  1165 => x"08f8050c",
  1166 => x"748c08fc",
  1167 => x"050c800b",
  1168 => x"8c08f805",
  1169 => x"0824b738",
  1170 => x"8c089005",
  1171 => x"0854800b",
  1172 => x"84150c8c",
  1173 => x"08900508",
  1174 => x"8c08f405",
  1175 => x"0888120c",
  1176 => x"8c089005",
  1177 => x"0857548c",
  1178 => x"08f80508",
  1179 => x"8c08fc05",
  1180 => x"08565473",
  1181 => x"8c170c74",
  1182 => x"90170c80",
  1183 => x"ce398c08",
  1184 => x"90050854",
  1185 => x"810b8415",
  1186 => x"0c8c0890",
  1187 => x"05088c08",
  1188 => x"f4050888",
  1189 => x"120c8c08",
  1190 => x"9005088c",
  1191 => x"08d40558",
  1192 => x"58548c08",
  1193 => x"f805088c",
  1194 => x"08fc0508",
  1195 => x"56547352",
  1196 => x"74537551",
  1197 => x"bee83f8c",
  1198 => x"08d40508",
  1199 => x"8c08d805",
  1200 => x"08565473",
  1201 => x"8c180c74",
  1202 => x"90180c8c",
  1203 => x"08900508",
  1204 => x"548c1408",
  1205 => x"f00a2682",
  1206 => x"b1388c08",
  1207 => x"9005088c",
  1208 => x"11087090",
  1209 => x"13080751",
  1210 => x"55557380",
  1211 => x"2e829b38",
  1212 => x"8c089005",
  1213 => x"088c0890",
  1214 => x"05089011",
  1215 => x"089f2a8c",
  1216 => x"12081070",
  1217 => x"72078c15",
  1218 => x"0c901308",
  1219 => x"1090150c",
  1220 => x"8c089005",
  1221 => x"08881108",
  1222 => x"ff058812",
  1223 => x"0c535858",
  1224 => x"5557ffa7",
  1225 => x"398c0890",
  1226 => x"05088c08",
  1227 => x"88050884",
  1228 => x"11088413",
  1229 => x"0c8c0890",
  1230 => x"05088c08",
  1231 => x"f4050888",
  1232 => x"120c8c08",
  1233 => x"9005088c",
  1234 => x"08ff9405",
  1235 => x"0c525654",
  1236 => x"8c08e805",
  1237 => x"088c08ec",
  1238 => x"05085755",
  1239 => x"748c08ff",
  1240 => x"8c050c75",
  1241 => x"8c08ff90",
  1242 => x"050c8c08",
  1243 => x"e005088c",
  1244 => x"08e40508",
  1245 => x"5654738c",
  1246 => x"08ff8405",
  1247 => x"0c748c08",
  1248 => x"ff88050c",
  1249 => x"8c08ff90",
  1250 => x"05088c08",
  1251 => x"ff880508",
  1252 => x"7012708c",
  1253 => x"08ff8005",
  1254 => x"0c525755",
  1255 => x"810b8c08",
  1256 => x"fef8050c",
  1257 => x"8c08ff80",
  1258 => x"05088c08",
  1259 => x"ff900508",
  1260 => x"56547474",
  1261 => x"26893880",
  1262 => x"0b8c08fe",
  1263 => x"f8050c8c",
  1264 => x"08ff8c05",
  1265 => x"088c08ff",
  1266 => x"84050870",
  1267 => x"12708c08",
  1268 => x"fefc050c",
  1269 => x"8c08fefc",
  1270 => x"05088c08",
  1271 => x"fef80508",
  1272 => x"11708c08",
  1273 => x"fefc050c",
  1274 => x"53585255",
  1275 => x"568c08fe",
  1276 => x"fc05088c",
  1277 => x"08ff8005",
  1278 => x"088c08ff",
  1279 => x"94050858",
  1280 => x"5654738c",
  1281 => x"170c7490",
  1282 => x"170c8c08",
  1283 => x"90050854",
  1284 => x"83740c8c",
  1285 => x"08900508",
  1286 => x"548c1408",
  1287 => x"f80a2684",
  1288 => x"3880cf39",
  1289 => x"8c089005",
  1290 => x"088c0890",
  1291 => x"05088c11",
  1292 => x"08800690",
  1293 => x"12088106",
  1294 => x"8c089005",
  1295 => x"088c1108",
  1296 => x"9f2b9012",
  1297 => x"08812a70",
  1298 => x"72078c14",
  1299 => x"08812a70",
  1300 => x"77078c1a",
  1301 => x"0c757207",
  1302 => x"901a0c8c",
  1303 => x"08900508",
  1304 => x"88110881",
  1305 => x"0588120c",
  1306 => x"51575c5f",
  1307 => x"5f5c5a58",
  1308 => x"555b8c08",
  1309 => x"90050870",
  1310 => x"8c08d005",
  1311 => x"0c548c08",
  1312 => x"d0050880",
  1313 => x"0cae3d0d",
  1314 => x"8c0c048c",
  1315 => x"08028c0c",
  1316 => x"ff3d0d80",
  1317 => x"0b8c08fc",
  1318 => x"050c8c08",
  1319 => x"88050851",
  1320 => x"7008822e",
  1321 => x"09810688",
  1322 => x"38810b8c",
  1323 => x"08fc050c",
  1324 => x"8c08fc05",
  1325 => x"0870800c",
  1326 => x"51833d0d",
  1327 => x"8c0c048c",
  1328 => x"08028c0c",
  1329 => x"803d0d82",
  1330 => x"c3d87080",
  1331 => x"0c51823d",
  1332 => x"0d8c0c04",
  1333 => x"8c08028c",
  1334 => x"0cff3d0d",
  1335 => x"800b8c08",
  1336 => x"fc050c8c",
  1337 => x"08880508",
  1338 => x"51700884",
  1339 => x"2e098106",
  1340 => x"8838810b",
  1341 => x"8c08fc05",
  1342 => x"0c8c08fc",
  1343 => x"05087080",
  1344 => x"0c51833d",
  1345 => x"0d8c0c04",
  1346 => x"8c08028c",
  1347 => x"0cff3d0d",
  1348 => x"800b8c08",
  1349 => x"fc050c8c",
  1350 => x"08880508",
  1351 => x"51700880",
  1352 => x"2e8f388c",
  1353 => x"08880508",
  1354 => x"51700881",
  1355 => x"2e833888",
  1356 => x"39810b8c",
  1357 => x"08fc050c",
  1358 => x"8c08fc05",
  1359 => x"0870800c",
  1360 => x"51833d0d",
  1361 => x"8c0c048c",
  1362 => x"08028c0c",
  1363 => x"e73d0d8c",
  1364 => x"08880508",
  1365 => x"568c088c",
  1366 => x"05088c08",
  1367 => x"90050856",
  1368 => x"54738c08",
  1369 => x"ffb8050c",
  1370 => x"748c08ff",
  1371 => x"bc050c8c",
  1372 => x"08940508",
  1373 => x"8c089805",
  1374 => x"08565473",
  1375 => x"8c08ffb0",
  1376 => x"050c748c",
  1377 => x"08ffb405",
  1378 => x"0c8c08ec",
  1379 => x"0570538c",
  1380 => x"08ffb805",
  1381 => x"70535154",
  1382 => x"80cae53f",
  1383 => x"8c08d805",
  1384 => x"70538c08",
  1385 => x"ffb00570",
  1386 => x"53515480",
  1387 => x"cad23f8c",
  1388 => x"08c40570",
  1389 => x"548c08d8",
  1390 => x"0570548c",
  1391 => x"08ec0570",
  1392 => x"54515154",
  1393 => x"f09d3f80",
  1394 => x"08708c08",
  1395 => x"c0050c8c",
  1396 => x"08c00508",
  1397 => x"53765254",
  1398 => x"b9f03f75",
  1399 => x"800c9b3d",
  1400 => x"0d8c0c04",
  1401 => x"8c08028c",
  1402 => x"0ce73d0d",
  1403 => x"8c088805",
  1404 => x"08568c08",
  1405 => x"8c05088c",
  1406 => x"08900508",
  1407 => x"5654738c",
  1408 => x"08ffb805",
  1409 => x"0c748c08",
  1410 => x"ffbc050c",
  1411 => x"8c089405",
  1412 => x"088c0898",
  1413 => x"05085654",
  1414 => x"738c08ff",
  1415 => x"b0050c74",
  1416 => x"8c08ffb4",
  1417 => x"050c8c08",
  1418 => x"ec057053",
  1419 => x"8c08ffb8",
  1420 => x"05705351",
  1421 => x"5480c9c8",
  1422 => x"3f8c08d8",
  1423 => x"0570538c",
  1424 => x"08ffb005",
  1425 => x"70535154",
  1426 => x"80c9b53f",
  1427 => x"8c08dc05",
  1428 => x"0881328c",
  1429 => x"08dc050c",
  1430 => x"8c08c405",
  1431 => x"70548c08",
  1432 => x"d8057054",
  1433 => x"8c08ec05",
  1434 => x"70545151",
  1435 => x"54eef43f",
  1436 => x"8008708c",
  1437 => x"08c0050c",
  1438 => x"8c08c005",
  1439 => x"08537652",
  1440 => x"54b8c73f",
  1441 => x"75800c9b",
  1442 => x"3d0d8c0c",
  1443 => x"048c0802",
  1444 => x"8c0cff83",
  1445 => x"3d0d8c08",
  1446 => x"8c05088c",
  1447 => x"08900508",
  1448 => x"5856758c",
  1449 => x"08ffb805",
  1450 => x"0c768c08",
  1451 => x"ffbc050c",
  1452 => x"8c089405",
  1453 => x"088c0898",
  1454 => x"05085856",
  1455 => x"758c08ff",
  1456 => x"b0050c76",
  1457 => x"8c08ffb4",
  1458 => x"050c8c08",
  1459 => x"ec057053",
  1460 => x"8c08ffb8",
  1461 => x"05705351",
  1462 => x"5680c8a4",
  1463 => x"3f8c08d8",
  1464 => x"0570538c",
  1465 => x"08ffb005",
  1466 => x"70535156",
  1467 => x"80c8913f",
  1468 => x"8c08ec05",
  1469 => x"8c08ffac",
  1470 => x"050c8c08",
  1471 => x"d8058c08",
  1472 => x"ffa8050c",
  1473 => x"8c08c405",
  1474 => x"8c08ffa4",
  1475 => x"050c8056",
  1476 => x"8057758c",
  1477 => x"08ff9805",
  1478 => x"0c768c08",
  1479 => x"ff9c050c",
  1480 => x"80568057",
  1481 => x"758c08ff",
  1482 => x"90050c76",
  1483 => x"8c08ff94",
  1484 => x"050c8c08",
  1485 => x"ffac0508",
  1486 => x"519ba23f",
  1487 => x"80085675",
  1488 => x"802e80d3",
  1489 => x"388c08ff",
  1490 => x"ac05088c",
  1491 => x"08fec405",
  1492 => x"0c800b8c",
  1493 => x"08fec005",
  1494 => x"0c8c08ff",
  1495 => x"ac05088c",
  1496 => x"08ffa805",
  1497 => x"08575784",
  1498 => x"17088417",
  1499 => x"082e8938",
  1500 => x"810b8c08",
  1501 => x"fec0050c",
  1502 => x"8c08fec4",
  1503 => x"05088c08",
  1504 => x"fec00508",
  1505 => x"84120c8c",
  1506 => x"08ffac05",
  1507 => x"088c08ff",
  1508 => x"a0050c56",
  1509 => x"99a0398c",
  1510 => x"08ffa805",
  1511 => x"08519abd",
  1512 => x"3f800856",
  1513 => x"75802e80",
  1514 => x"d3388c08",
  1515 => x"ffa80508",
  1516 => x"8c08febc",
  1517 => x"050c800b",
  1518 => x"8c08feb8",
  1519 => x"050c8c08",
  1520 => x"ffac0508",
  1521 => x"8c08ffa8",
  1522 => x"05085757",
  1523 => x"84170884",
  1524 => x"17082e89",
  1525 => x"38810b8c",
  1526 => x"08feb805",
  1527 => x"0c8c08fe",
  1528 => x"bc05088c",
  1529 => x"08feb805",
  1530 => x"0884120c",
  1531 => x"8c08ffa8",
  1532 => x"05088c08",
  1533 => x"ffa0050c",
  1534 => x"5798bb39",
  1535 => x"8c08ffac",
  1536 => x"05085199",
  1537 => x"a43f8008",
  1538 => x"5675802e",
  1539 => x"80f5388c",
  1540 => x"08ffa805",
  1541 => x"085198dd",
  1542 => x"3f800856",
  1543 => x"75802e91",
  1544 => x"3898bd3f",
  1545 => x"8008708c",
  1546 => x"08ffa005",
  1547 => x"0c569886",
  1548 => x"398c08ff",
  1549 => x"ac05088c",
  1550 => x"08feb405",
  1551 => x"0c800b8c",
  1552 => x"08feb005",
  1553 => x"0c8c08ff",
  1554 => x"ac05088c",
  1555 => x"08ffa805",
  1556 => x"08575784",
  1557 => x"17088417",
  1558 => x"082e8938",
  1559 => x"810b8c08",
  1560 => x"feb0050c",
  1561 => x"8c08feb4",
  1562 => x"05088c08",
  1563 => x"feb00508",
  1564 => x"84120c8c",
  1565 => x"08ffac05",
  1566 => x"088c08ff",
  1567 => x"a0050c56",
  1568 => x"97b4398c",
  1569 => x"08ffa805",
  1570 => x"0851989d",
  1571 => x"3f800856",
  1572 => x"75802e80",
  1573 => x"f5388c08",
  1574 => x"ffac0508",
  1575 => x"5197d63f",
  1576 => x"80085675",
  1577 => x"802e9138",
  1578 => x"97b63f80",
  1579 => x"08708c08",
  1580 => x"ffa0050c",
  1581 => x"5696ff39",
  1582 => x"8c08ffa8",
  1583 => x"05088c08",
  1584 => x"feac050c",
  1585 => x"800b8c08",
  1586 => x"fea8050c",
  1587 => x"8c08ffac",
  1588 => x"05088c08",
  1589 => x"ffa80508",
  1590 => x"57578417",
  1591 => x"08841708",
  1592 => x"2e893881",
  1593 => x"0b8c08fe",
  1594 => x"a8050c8c",
  1595 => x"08feac05",
  1596 => x"088c08fe",
  1597 => x"a8050884",
  1598 => x"120c8c08",
  1599 => x"ffa80508",
  1600 => x"8c08ffa0",
  1601 => x"050c5796",
  1602 => x"ad398c08",
  1603 => x"ffac0508",
  1604 => x"5196e23f",
  1605 => x"80085675",
  1606 => x"802e80d3",
  1607 => x"388c08ff",
  1608 => x"ac05088c",
  1609 => x"08fea405",
  1610 => x"0c800b8c",
  1611 => x"08fea005",
  1612 => x"0c8c08ff",
  1613 => x"ac05088c",
  1614 => x"08ffa805",
  1615 => x"08575784",
  1616 => x"17088417",
  1617 => x"082e8938",
  1618 => x"810b8c08",
  1619 => x"fea0050c",
  1620 => x"8c08fea4",
  1621 => x"05088c08",
  1622 => x"fea00508",
  1623 => x"84120c8c",
  1624 => x"08ffac05",
  1625 => x"088c08ff",
  1626 => x"a0050c56",
  1627 => x"95c8398c",
  1628 => x"08ffa805",
  1629 => x"085195fd",
  1630 => x"3f800856",
  1631 => x"75802e80",
  1632 => x"d3388c08",
  1633 => x"ffa80508",
  1634 => x"8c08fe9c",
  1635 => x"050c800b",
  1636 => x"8c08fe98",
  1637 => x"050c8c08",
  1638 => x"ffac0508",
  1639 => x"8c08ffa8",
  1640 => x"05085757",
  1641 => x"84170884",
  1642 => x"17082e89",
  1643 => x"38810b8c",
  1644 => x"08fe9805",
  1645 => x"0c8c08fe",
  1646 => x"9c05088c",
  1647 => x"08fe9805",
  1648 => x"0884120c",
  1649 => x"8c08ffa8",
  1650 => x"05088c08",
  1651 => x"ffa0050c",
  1652 => x"5794e339",
  1653 => x"8c08ffac",
  1654 => x"05089011",
  1655 => x"088c08ff",
  1656 => x"8c050c8c",
  1657 => x"08ffac05",
  1658 => x"088c1108",
  1659 => x"802a5959",
  1660 => x"5680778c",
  1661 => x"08ff8805",
  1662 => x"0c8c08ff",
  1663 => x"a8050890",
  1664 => x"11088c08",
  1665 => x"ff84050c",
  1666 => x"8c08ffa8",
  1667 => x"05088c11",
  1668 => x"08802a5a",
  1669 => x"5a515680",
  1670 => x"778c08ff",
  1671 => x"80050c8c",
  1672 => x"08ff8405",
  1673 => x"085a5680",
  1674 => x"0b8c08ff",
  1675 => x"8c050858",
  1676 => x"58800b8c",
  1677 => x"08fef005",
  1678 => x"5b567554",
  1679 => x"76557752",
  1680 => x"78537951",
  1681 => x"abfc3f8c",
  1682 => x"08fef005",
  1683 => x"088c08fe",
  1684 => x"f4050858",
  1685 => x"56758c08",
  1686 => x"fef8050c",
  1687 => x"768c08fe",
  1688 => x"fc050c8c",
  1689 => x"08ff8005",
  1690 => x"0859800b",
  1691 => x"8c08ff8c",
  1692 => x"05085858",
  1693 => x"800b8c08",
  1694 => x"fee8055b",
  1695 => x"56755476",
  1696 => x"55775278",
  1697 => x"537951ab",
  1698 => x"b93f8c08",
  1699 => x"fee80508",
  1700 => x"8c08feec",
  1701 => x"05085856",
  1702 => x"758c08fe",
  1703 => x"f0050c76",
  1704 => x"8c08fef4",
  1705 => x"050c8c08",
  1706 => x"ff840508",
  1707 => x"59800b8c",
  1708 => x"08ff8805",
  1709 => x"08585880",
  1710 => x"0b8c08fe",
  1711 => x"e0055b56",
  1712 => x"75547655",
  1713 => x"77527853",
  1714 => x"7951aaf6",
  1715 => x"3f8c08fe",
  1716 => x"e005088c",
  1717 => x"08fee405",
  1718 => x"08585675",
  1719 => x"8c08fee8",
  1720 => x"050c768c",
  1721 => x"08feec05",
  1722 => x"0c8c08ff",
  1723 => x"80050859",
  1724 => x"800b8c08",
  1725 => x"ff880508",
  1726 => x"5858800b",
  1727 => x"8c08fed8",
  1728 => x"055b5675",
  1729 => x"54765577",
  1730 => x"52785379",
  1731 => x"51aab33f",
  1732 => x"8c08fed8",
  1733 => x"05088c08",
  1734 => x"fedc0508",
  1735 => x"5856758c",
  1736 => x"08fee005",
  1737 => x"0c768c08",
  1738 => x"fee4050c",
  1739 => x"80568057",
  1740 => x"758c08fe",
  1741 => x"d8050c76",
  1742 => x"8c08fedc",
  1743 => x"050c8056",
  1744 => x"8057758c",
  1745 => x"08fed005",
  1746 => x"0c768c08",
  1747 => x"fed4050c",
  1748 => x"8c08fef0",
  1749 => x"05088c08",
  1750 => x"fef40508",
  1751 => x"5856758c",
  1752 => x"08fe9005",
  1753 => x"0c768c08",
  1754 => x"fe94050c",
  1755 => x"8c08fee8",
  1756 => x"05088c08",
  1757 => x"feec0508",
  1758 => x"5856758c",
  1759 => x"08fe8805",
  1760 => x"0c768c08",
  1761 => x"fe8c050c",
  1762 => x"8c08fe94",
  1763 => x"05088c08",
  1764 => x"fe8c0508",
  1765 => x"7012708c",
  1766 => x"08fe8405",
  1767 => x"0c525757",
  1768 => x"810b8c08",
  1769 => x"fdfc050c",
  1770 => x"8c08fe84",
  1771 => x"05088c08",
  1772 => x"fe940508",
  1773 => x"57577577",
  1774 => x"26893880",
  1775 => x"0b8c08fd",
  1776 => x"fc050c8c",
  1777 => x"08fe9005",
  1778 => x"088c08fe",
  1779 => x"88050870",
  1780 => x"12708c08",
  1781 => x"fe80050c",
  1782 => x"8c08fe80",
  1783 => x"05088c08",
  1784 => x"fdfc0508",
  1785 => x"11708c08",
  1786 => x"fe80050c",
  1787 => x"53515257",
  1788 => x"578c08fe",
  1789 => x"8005088c",
  1790 => x"08fe8405",
  1791 => x"08585675",
  1792 => x"8c08fec8",
  1793 => x"050c768c",
  1794 => x"08fecc05",
  1795 => x"0c8c08fe",
  1796 => x"f005088c",
  1797 => x"08fec805",
  1798 => x"0826a638",
  1799 => x"8c08fef0",
  1800 => x"05088c08",
  1801 => x"fec80508",
  1802 => x"2e098106",
  1803 => x"81c6388c",
  1804 => x"08fef405",
  1805 => x"088c08fe",
  1806 => x"cc050826",
  1807 => x"843881b4",
  1808 => x"398c08fe",
  1809 => x"d805088c",
  1810 => x"08fedc05",
  1811 => x"08585675",
  1812 => x"8c08fdf4",
  1813 => x"050c768c",
  1814 => x"08fdf805",
  1815 => x"0c815680",
  1816 => x"57758c08",
  1817 => x"fdec050c",
  1818 => x"768c08fd",
  1819 => x"f0050c8c",
  1820 => x"08fdf805",
  1821 => x"088c08fd",
  1822 => x"f0050870",
  1823 => x"12708c08",
  1824 => x"fde8050c",
  1825 => x"52575781",
  1826 => x"0b8c08fd",
  1827 => x"e0050c8c",
  1828 => x"08fde805",
  1829 => x"088c08fd",
  1830 => x"f8050857",
  1831 => x"57757726",
  1832 => x"8938800b",
  1833 => x"8c08fde0",
  1834 => x"050c8c08",
  1835 => x"fdf40508",
  1836 => x"8c08fdec",
  1837 => x"05087012",
  1838 => x"708c08fd",
  1839 => x"e4050c8c",
  1840 => x"08fde405",
  1841 => x"088c08fd",
  1842 => x"e0050811",
  1843 => x"708c08fd",
  1844 => x"e4050c53",
  1845 => x"51525757",
  1846 => x"8c08fde4",
  1847 => x"05088c08",
  1848 => x"fde80508",
  1849 => x"5856758c",
  1850 => x"08fed805",
  1851 => x"0c768c08",
  1852 => x"fedc050c",
  1853 => x"8c08fecc",
  1854 => x"05085780",
  1855 => x"77802b8c",
  1856 => x"08fef005",
  1857 => x"0c56800b",
  1858 => x"8c08fef4",
  1859 => x"050c8c08",
  1860 => x"fef80508",
  1861 => x"8c08fefc",
  1862 => x"05085856",
  1863 => x"758c08fd",
  1864 => x"d8050c76",
  1865 => x"8c08fddc",
  1866 => x"050c8c08",
  1867 => x"fef00508",
  1868 => x"8c08fef4",
  1869 => x"05085856",
  1870 => x"758c08fd",
  1871 => x"d0050c76",
  1872 => x"8c08fdd4",
  1873 => x"050c8c08",
  1874 => x"fddc0508",
  1875 => x"8c08fdd4",
  1876 => x"05087012",
  1877 => x"708c08fd",
  1878 => x"cc050c52",
  1879 => x"5757810b",
  1880 => x"8c08fdc4",
  1881 => x"050c8c08",
  1882 => x"fdcc0508",
  1883 => x"8c08fddc",
  1884 => x"05085757",
  1885 => x"75772689",
  1886 => x"38800b8c",
  1887 => x"08fdc405",
  1888 => x"0c8c08fd",
  1889 => x"d805088c",
  1890 => x"08fdd005",
  1891 => x"08701270",
  1892 => x"8c08fdc8",
  1893 => x"050c8c08",
  1894 => x"fdc80508",
  1895 => x"8c08fdc4",
  1896 => x"05081170",
  1897 => x"8c08fdc8",
  1898 => x"050c5351",
  1899 => x"5257578c",
  1900 => x"08fdc805",
  1901 => x"088c08fd",
  1902 => x"cc050858",
  1903 => x"56758c08",
  1904 => x"fed0050c",
  1905 => x"768c08fe",
  1906 => x"d4050c8c",
  1907 => x"08fef805",
  1908 => x"088c08fe",
  1909 => x"d0050826",
  1910 => x"a6388c08",
  1911 => x"fef80508",
  1912 => x"8c08fed0",
  1913 => x"05082e09",
  1914 => x"810681c6",
  1915 => x"388c08fe",
  1916 => x"fc05088c",
  1917 => x"08fed405",
  1918 => x"08268438",
  1919 => x"81b4398c",
  1920 => x"08fed805",
  1921 => x"088c08fe",
  1922 => x"dc050858",
  1923 => x"56758c08",
  1924 => x"fdbc050c",
  1925 => x"768c08fd",
  1926 => x"c0050c80",
  1927 => x"56815775",
  1928 => x"8c08fdb4",
  1929 => x"050c768c",
  1930 => x"08fdb805",
  1931 => x"0c8c08fd",
  1932 => x"c005088c",
  1933 => x"08fdb805",
  1934 => x"08701270",
  1935 => x"8c08fdb0",
  1936 => x"050c5257",
  1937 => x"57810b8c",
  1938 => x"08fda805",
  1939 => x"0c8c08fd",
  1940 => x"b005088c",
  1941 => x"08fdc005",
  1942 => x"08575775",
  1943 => x"77268938",
  1944 => x"800b8c08",
  1945 => x"fda8050c",
  1946 => x"8c08fdbc",
  1947 => x"05088c08",
  1948 => x"fdb40508",
  1949 => x"7012708c",
  1950 => x"08fdac05",
  1951 => x"0c8c08fd",
  1952 => x"ac05088c",
  1953 => x"08fda805",
  1954 => x"0811708c",
  1955 => x"08fdac05",
  1956 => x"0c535152",
  1957 => x"57578c08",
  1958 => x"fdac0508",
  1959 => x"8c08fdb0",
  1960 => x"05085856",
  1961 => x"758c08fe",
  1962 => x"d8050c76",
  1963 => x"8c08fedc",
  1964 => x"050c8c08",
  1965 => x"fec80508",
  1966 => x"802a708c",
  1967 => x"08fda405",
  1968 => x"0c578070",
  1969 => x"8c08fda0",
  1970 => x"050c568c",
  1971 => x"08fda005",
  1972 => x"088c08fd",
  1973 => x"a4050858",
  1974 => x"56758c08",
  1975 => x"fda0050c",
  1976 => x"768c08fd",
  1977 => x"a4050c8c",
  1978 => x"08fee005",
  1979 => x"088c08fe",
  1980 => x"e4050858",
  1981 => x"56758c08",
  1982 => x"fd98050c",
  1983 => x"768c08fd",
  1984 => x"9c050c8c",
  1985 => x"08fda405",
  1986 => x"088c08fd",
  1987 => x"9c050870",
  1988 => x"12708c08",
  1989 => x"fd94050c",
  1990 => x"52575781",
  1991 => x"0b8c08fd",
  1992 => x"8c050c8c",
  1993 => x"08fd9405",
  1994 => x"088c08fd",
  1995 => x"a4050857",
  1996 => x"57757726",
  1997 => x"8938800b",
  1998 => x"8c08fd8c",
  1999 => x"050c8c08",
  2000 => x"fda00508",
  2001 => x"8c08fd98",
  2002 => x"05087012",
  2003 => x"708c08fd",
  2004 => x"90050c8c",
  2005 => x"08fd9005",
  2006 => x"088c08fd",
  2007 => x"8c050811",
  2008 => x"708c08fd",
  2009 => x"90050c53",
  2010 => x"51525757",
  2011 => x"8c08fed8",
  2012 => x"05088c08",
  2013 => x"fedc0508",
  2014 => x"5856758c",
  2015 => x"08fd8405",
  2016 => x"0c768c08",
  2017 => x"fd88050c",
  2018 => x"8c08fd88",
  2019 => x"05088c08",
  2020 => x"fd940508",
  2021 => x"7012708c",
  2022 => x"08fd8005",
  2023 => x"0c525757",
  2024 => x"810b8c08",
  2025 => x"fcf8050c",
  2026 => x"8c08fd80",
  2027 => x"05088c08",
  2028 => x"fd880508",
  2029 => x"57577577",
  2030 => x"26893880",
  2031 => x"0b8c08fc",
  2032 => x"f8050c8c",
  2033 => x"08fd8405",
  2034 => x"088c08fd",
  2035 => x"90050870",
  2036 => x"12708c08",
  2037 => x"fcfc050c",
  2038 => x"8c08fcfc",
  2039 => x"05088c08",
  2040 => x"fcf80508",
  2041 => x"11708c08",
  2042 => x"fcfc050c",
  2043 => x"53515257",
  2044 => x"578c08fc",
  2045 => x"fc05088c",
  2046 => x"08fd8005",
  2047 => x"08585675",
  2048 => x"8c08fed8",
  2049 => x"050c768c",
  2050 => x"08fedc05",
  2051 => x"0c8c08fe",
  2052 => x"d805088c",
  2053 => x"08fedc05",
  2054 => x"08585675",
  2055 => x"8c08ff90",
  2056 => x"050c768c",
  2057 => x"08ff9405",
  2058 => x"0c8c08fe",
  2059 => x"d005088c",
  2060 => x"08fed405",
  2061 => x"08585675",
  2062 => x"8c08ff98",
  2063 => x"050c768c",
  2064 => x"08ff9c05",
  2065 => x"0c8c08ff",
  2066 => x"a405088c",
  2067 => x"08ffac05",
  2068 => x"088c08ff",
  2069 => x"a8050888",
  2070 => x"12088812",
  2071 => x"08058411",
  2072 => x"88150c8c",
  2073 => x"08ffa405",
  2074 => x"088c08fc",
  2075 => x"f4050c51",
  2076 => x"58585880",
  2077 => x"0b8c08fc",
  2078 => x"f0050c8c",
  2079 => x"08ffac05",
  2080 => x"088c08ff",
  2081 => x"a8050857",
  2082 => x"57841708",
  2083 => x"8417082e",
  2084 => x"8938810b",
  2085 => x"8c08fcf0",
  2086 => x"050c8c08",
  2087 => x"fcf40508",
  2088 => x"8c08fcf0",
  2089 => x"05088412",
  2090 => x"0c578c08",
  2091 => x"ff900508",
  2092 => x"f80a2684",
  2093 => x"3881a839",
  2094 => x"8c08ffa4",
  2095 => x"05088811",
  2096 => x"08810588",
  2097 => x"120c8c08",
  2098 => x"ff900508",
  2099 => x"80068c08",
  2100 => x"ff940508",
  2101 => x"81067052",
  2102 => x"59515675",
  2103 => x"802e80cf",
  2104 => x"388c08ff",
  2105 => x"9805089f",
  2106 => x"2b8c08ff",
  2107 => x"9c050881",
  2108 => x"2a707207",
  2109 => x"8c08ff98",
  2110 => x"0508812a",
  2111 => x"59595959",
  2112 => x"758c08ff",
  2113 => x"98050c76",
  2114 => x"8c08ff9c",
  2115 => x"050c8c08",
  2116 => x"ff980508",
  2117 => x"810a078c",
  2118 => x"08ff9c05",
  2119 => x"08800758",
  2120 => x"56758c08",
  2121 => x"ff98050c",
  2122 => x"768c08ff",
  2123 => x"9c050c8c",
  2124 => x"08ff9005",
  2125 => x"089f2b8c",
  2126 => x"08ff9405",
  2127 => x"08812a70",
  2128 => x"72078c08",
  2129 => x"ff900508",
  2130 => x"812a5959",
  2131 => x"5959758c",
  2132 => x"08ff9005",
  2133 => x"0c768c08",
  2134 => x"ff94050c",
  2135 => x"fecc398c",
  2136 => x"08ff9005",
  2137 => x"08f00a26",
  2138 => x"8196388c",
  2139 => x"08ffa405",
  2140 => x"08881108",
  2141 => x"ff058812",
  2142 => x"0c8c08ff",
  2143 => x"9405089f",
  2144 => x"2a8c08ff",
  2145 => x"90050810",
  2146 => x"7072078c",
  2147 => x"08ff9405",
  2148 => x"08105b53",
  2149 => x"5a5a5675",
  2150 => x"8c08ff90",
  2151 => x"050c768c",
  2152 => x"08ff9405",
  2153 => x"0c800b8c",
  2154 => x"08ff9805",
  2155 => x"08248338",
  2156 => x"a1398c08",
  2157 => x"ff900508",
  2158 => x"80078c08",
  2159 => x"ff940508",
  2160 => x"81075856",
  2161 => x"758c08ff",
  2162 => x"90050c76",
  2163 => x"8c08ff94",
  2164 => x"050c8c08",
  2165 => x"ff9c0508",
  2166 => x"9f2a8c08",
  2167 => x"ff980508",
  2168 => x"10707207",
  2169 => x"8c08ff9c",
  2170 => x"0508105a",
  2171 => x"58595975",
  2172 => x"8c08ff98",
  2173 => x"050c768c",
  2174 => x"08ff9c05",
  2175 => x"0cfee039",
  2176 => x"8c08ff90",
  2177 => x"05088006",
  2178 => x"708c08fc",
  2179 => x"e8050c8c",
  2180 => x"08ff9405",
  2181 => x"0881ff06",
  2182 => x"708c08fc",
  2183 => x"ec050c58",
  2184 => x"568c08fc",
  2185 => x"e805088c",
  2186 => x"08fcec05",
  2187 => x"08585675",
  2188 => x"8c08fce8",
  2189 => x"050c768c",
  2190 => x"08fcec05",
  2191 => x"0c8c08fc",
  2192 => x"e8050857",
  2193 => x"7683bc38",
  2194 => x"8c08fcec",
  2195 => x"05085675",
  2196 => x"81802e09",
  2197 => x"810683ab",
  2198 => x"388c08ff",
  2199 => x"90050898",
  2200 => x"2b8c08ff",
  2201 => x"94050888",
  2202 => x"2a707207",
  2203 => x"8c08ff90",
  2204 => x"0508882a",
  2205 => x"71810651",
  2206 => x"59595959",
  2207 => x"75802e81",
  2208 => x"b8388c08",
  2209 => x"ff900508",
  2210 => x"8c08ff94",
  2211 => x"05085856",
  2212 => x"758c08fc",
  2213 => x"e0050c76",
  2214 => x"8c08fce4",
  2215 => x"050c8056",
  2216 => x"81805775",
  2217 => x"8c08fcd8",
  2218 => x"050c768c",
  2219 => x"08fcdc05",
  2220 => x"0c8c08fc",
  2221 => x"e405088c",
  2222 => x"08fcdc05",
  2223 => x"08701270",
  2224 => x"8c08fcd4",
  2225 => x"050c5257",
  2226 => x"57810b8c",
  2227 => x"08fccc05",
  2228 => x"0c8c08fc",
  2229 => x"d405088c",
  2230 => x"08fce405",
  2231 => x"08575775",
  2232 => x"77268938",
  2233 => x"800b8c08",
  2234 => x"fccc050c",
  2235 => x"8c08fce0",
  2236 => x"05088c08",
  2237 => x"fcd80508",
  2238 => x"7012708c",
  2239 => x"08fcd005",
  2240 => x"0c8c08fc",
  2241 => x"d005088c",
  2242 => x"08fccc05",
  2243 => x"0811708c",
  2244 => x"08fcd005",
  2245 => x"0c535152",
  2246 => x"57578c08",
  2247 => x"fcd00508",
  2248 => x"8c08fcd4",
  2249 => x"05085856",
  2250 => x"758c08ff",
  2251 => x"90050c76",
  2252 => x"8c08ff94",
  2253 => x"050c81cb",
  2254 => x"398c08ff",
  2255 => x"98050870",
  2256 => x"8c08ff9c",
  2257 => x"05080751",
  2258 => x"5675802e",
  2259 => x"81b5388c",
  2260 => x"08ff9005",
  2261 => x"088c08ff",
  2262 => x"94050858",
  2263 => x"56758c08",
  2264 => x"fcc4050c",
  2265 => x"768c08fc",
  2266 => x"c8050c80",
  2267 => x"56818057",
  2268 => x"758c08fc",
  2269 => x"bc050c76",
  2270 => x"8c08fcc0",
  2271 => x"050c8c08",
  2272 => x"fcc80508",
  2273 => x"8c08fcc0",
  2274 => x"05087012",
  2275 => x"708c08fc",
  2276 => x"b8050c52",
  2277 => x"5757810b",
  2278 => x"8c08fcb0",
  2279 => x"050c8c08",
  2280 => x"fcb80508",
  2281 => x"8c08fcc8",
  2282 => x"05085757",
  2283 => x"75772689",
  2284 => x"38800b8c",
  2285 => x"08fcb005",
  2286 => x"0c8c08fc",
  2287 => x"c405088c",
  2288 => x"08fcbc05",
  2289 => x"08701270",
  2290 => x"8c08fcb4",
  2291 => x"050c8c08",
  2292 => x"fcb40508",
  2293 => x"8c08fcb0",
  2294 => x"05081170",
  2295 => x"8c08fcb4",
  2296 => x"050c5351",
  2297 => x"5257578c",
  2298 => x"08fcb405",
  2299 => x"088c08fc",
  2300 => x"b8050858",
  2301 => x"56758c08",
  2302 => x"ff90050c",
  2303 => x"768c08ff",
  2304 => x"94050c8c",
  2305 => x"08ffa405",
  2306 => x"08568c08",
  2307 => x"ff900508",
  2308 => x"8c08ff94",
  2309 => x"05085957",
  2310 => x"768c170c",
  2311 => x"7790170c",
  2312 => x"8c08ffa4",
  2313 => x"05085683",
  2314 => x"760c8c08",
  2315 => x"ffa40508",
  2316 => x"8c08ffa0",
  2317 => x"050c8c08",
  2318 => x"ffa00508",
  2319 => x"708c08c0",
  2320 => x"050c8c08",
  2321 => x"c0050853",
  2322 => x"8c088805",
  2323 => x"0852569c",
  2324 => x"f93f8c08",
  2325 => x"88050880",
  2326 => x"0c80ff3d",
  2327 => x"0d8c0c04",
  2328 => x"8c08028c",
  2329 => x"0c803d0d",
  2330 => x"82c3d870",
  2331 => x"800c5182",
  2332 => x"3d0d8c0c",
  2333 => x"048c0802",
  2334 => x"8c0cff3d",
  2335 => x"0d800b8c",
  2336 => x"08fc050c",
  2337 => x"8c088805",
  2338 => x"08517008",
  2339 => x"822e0981",
  2340 => x"06883881",
  2341 => x"0b8c08fc",
  2342 => x"050c8c08",
  2343 => x"fc050870",
  2344 => x"800c5183",
  2345 => x"3d0d8c0c",
  2346 => x"048c0802",
  2347 => x"8c0cff3d",
  2348 => x"0d800b8c",
  2349 => x"08fc050c",
  2350 => x"8c088805",
  2351 => x"08517008",
  2352 => x"842e0981",
  2353 => x"06883881",
  2354 => x"0b8c08fc",
  2355 => x"050c8c08",
  2356 => x"fc050870",
  2357 => x"800c5183",
  2358 => x"3d0d8c0c",
  2359 => x"048c0802",
  2360 => x"8c0cff3d",
  2361 => x"0d800b8c",
  2362 => x"08fc050c",
  2363 => x"8c088805",
  2364 => x"08517008",
  2365 => x"802e8f38",
  2366 => x"8c088805",
  2367 => x"08517008",
  2368 => x"812e8338",
  2369 => x"8839810b",
  2370 => x"8c08fc05",
  2371 => x"0c8c08fc",
  2372 => x"05087080",
  2373 => x"0c51833d",
  2374 => x"0d8c0c04",
  2375 => x"8c08028c",
  2376 => x"0cffbc3d",
  2377 => x"0d8c088c",
  2378 => x"05088c08",
  2379 => x"90050855",
  2380 => x"53728c08",
  2381 => x"cc050c73",
  2382 => x"8c08d005",
  2383 => x"0c8c0894",
  2384 => x"05088c08",
  2385 => x"98050855",
  2386 => x"53728c08",
  2387 => x"c4050c73",
  2388 => x"8c08c805",
  2389 => x"0c8c08ec",
  2390 => x"0570538c",
  2391 => x"08cc0570",
  2392 => x"535153ab",
  2393 => x"9b3f8c08",
  2394 => x"d8057053",
  2395 => x"8c08c405",
  2396 => x"70535153",
  2397 => x"ab8a3f8c",
  2398 => x"08ec058c",
  2399 => x"08c0050c",
  2400 => x"8c08d805",
  2401 => x"8c08ffbc",
  2402 => x"050c8c08",
  2403 => x"c0050851",
  2404 => x"8efa3f80",
  2405 => x"08537280",
  2406 => x"2e8f388c",
  2407 => x"08c00508",
  2408 => x"8c08ffb8",
  2409 => x"050c8dbd",
  2410 => x"398c08ff",
  2411 => x"bc050851",
  2412 => x"8eda3f80",
  2413 => x"08537280",
  2414 => x"2e90388c",
  2415 => x"08ffbc05",
  2416 => x"088c08ff",
  2417 => x"b8050c8d",
  2418 => x"9c398c08",
  2419 => x"c005088c",
  2420 => x"08c00508",
  2421 => x"8c08ffbc",
  2422 => x"05088412",
  2423 => x"08841208",
  2424 => x"3284140c",
  2425 => x"8c08c005",
  2426 => x"08545555",
  2427 => x"558de93f",
  2428 => x"80085372",
  2429 => x"92388c08",
  2430 => x"c0050851",
  2431 => x"8da63f80",
  2432 => x"08537283",
  2433 => x"38b6398c",
  2434 => x"08c00508",
  2435 => x"8c08ffbc",
  2436 => x"05085454",
  2437 => x"73087308",
  2438 => x"2e098106",
  2439 => x"91388cef",
  2440 => x"3f800870",
  2441 => x"8c08ffb8",
  2442 => x"050c538c",
  2443 => x"b8398c08",
  2444 => x"c005088c",
  2445 => x"08ffb805",
  2446 => x"0c8caa39",
  2447 => x"8c08ffbc",
  2448 => x"0508518d",
  2449 => x"933f8008",
  2450 => x"5372802e",
  2451 => x"ac388c08",
  2452 => x"c0050853",
  2453 => x"80548055",
  2454 => x"738c140c",
  2455 => x"7490140c",
  2456 => x"8c08c005",
  2457 => x"0853800b",
  2458 => x"88140c8c",
  2459 => x"08c00508",
  2460 => x"8c08ffb8",
  2461 => x"050c8bed",
  2462 => x"398c08ff",
  2463 => x"bc050851",
  2464 => x"8ca23f80",
  2465 => x"08537280",
  2466 => x"2e98388c",
  2467 => x"08c00508",
  2468 => x"5384730c",
  2469 => x"8c08c005",
  2470 => x"088c08ff",
  2471 => x"b8050c8b",
  2472 => x"c4398c08",
  2473 => x"c005088c",
  2474 => x"08c00508",
  2475 => x"8c08ffbc",
  2476 => x"05088812",
  2477 => x"08881208",
  2478 => x"3188140c",
  2479 => x"8c08c005",
  2480 => x"08515555",
  2481 => x"55901308",
  2482 => x"8c140854",
  2483 => x"54728c08",
  2484 => x"ffa8050c",
  2485 => x"738c08ff",
  2486 => x"ac050c8c",
  2487 => x"08ffbc05",
  2488 => x"08539013",
  2489 => x"088c1408",
  2490 => x"5454728c",
  2491 => x"08ffa005",
  2492 => x"0c738c08",
  2493 => x"ffa4050c",
  2494 => x"8c08ffa0",
  2495 => x"05088c08",
  2496 => x"ffa80508",
  2497 => x"26a6388c",
  2498 => x"08ffa005",
  2499 => x"088c08ff",
  2500 => x"a805082e",
  2501 => x"09810681",
  2502 => x"de388c08",
  2503 => x"ffa40508",
  2504 => x"8c08ffac",
  2505 => x"05082684",
  2506 => x"3881cc39",
  2507 => x"8c08ffa8",
  2508 => x"05088c08",
  2509 => x"ffac0508",
  2510 => x"5553728c",
  2511 => x"08ff9005",
  2512 => x"0c738c08",
  2513 => x"ff94050c",
  2514 => x"8c08ff90",
  2515 => x"05088c08",
  2516 => x"ff940508",
  2517 => x"5553728c",
  2518 => x"08ff8805",
  2519 => x"0c738c08",
  2520 => x"ff8c050c",
  2521 => x"8c08ff8c",
  2522 => x"05088c08",
  2523 => x"ff940508",
  2524 => x"7012708c",
  2525 => x"08ff8405",
  2526 => x"0c525454",
  2527 => x"810b8c08",
  2528 => x"fefc050c",
  2529 => x"8c08ff84",
  2530 => x"05088c08",
  2531 => x"ff8c0508",
  2532 => x"54547274",
  2533 => x"26893880",
  2534 => x"0b8c08fe",
  2535 => x"fc050c8c",
  2536 => x"08ff8805",
  2537 => x"088c08ff",
  2538 => x"90050870",
  2539 => x"12708c08",
  2540 => x"ff80050c",
  2541 => x"8c08ff80",
  2542 => x"05088c08",
  2543 => x"fefc0508",
  2544 => x"11708c08",
  2545 => x"ff80050c",
  2546 => x"53515254",
  2547 => x"548c08ff",
  2548 => x"8005088c",
  2549 => x"08ff8405",
  2550 => x"08555372",
  2551 => x"8c08ffa8",
  2552 => x"050c738c",
  2553 => x"08ffac05",
  2554 => x"0c8c08c0",
  2555 => x"05088811",
  2556 => x"08ff0588",
  2557 => x"120c5388",
  2558 => x"0a538054",
  2559 => x"728c08ff",
  2560 => x"b0050c73",
  2561 => x"8c08ffb4",
  2562 => x"050c8053",
  2563 => x"8054728c",
  2564 => x"08ff9805",
  2565 => x"0c738c08",
  2566 => x"ff9c050c",
  2567 => x"8c08ffb0",
  2568 => x"0508708c",
  2569 => x"08ffb405",
  2570 => x"08075153",
  2571 => x"72802e84",
  2572 => x"8a388c08",
  2573 => x"ffa00508",
  2574 => x"8c08ffa8",
  2575 => x"05082682",
  2576 => x"8d388c08",
  2577 => x"ffa00508",
  2578 => x"8c08ffa8",
  2579 => x"05082e09",
  2580 => x"81069138",
  2581 => x"8c08ffa4",
  2582 => x"05088c08",
  2583 => x"ffac0508",
  2584 => x"2681eb38",
  2585 => x"8c08ff98",
  2586 => x"05088c08",
  2587 => x"ffb00508",
  2588 => x"078c08ff",
  2589 => x"9c05088c",
  2590 => x"08ffb405",
  2591 => x"08075553",
  2592 => x"728c08ff",
  2593 => x"98050c73",
  2594 => x"8c08ff9c",
  2595 => x"050c8c08",
  2596 => x"ffa80508",
  2597 => x"8c08ffac",
  2598 => x"05085553",
  2599 => x"728c08fe",
  2600 => x"f4050c73",
  2601 => x"8c08fef8",
  2602 => x"050c8c08",
  2603 => x"ffa00508",
  2604 => x"8c08ffa4",
  2605 => x"05085553",
  2606 => x"728c08fe",
  2607 => x"ec050c73",
  2608 => x"8c08fef0",
  2609 => x"050c8c08",
  2610 => x"fef80508",
  2611 => x"8c08fef0",
  2612 => x"05087171",
  2613 => x"31708c08",
  2614 => x"fee8050c",
  2615 => x"52545481",
  2616 => x"0b8c08fe",
  2617 => x"e0050c8c",
  2618 => x"08fee805",
  2619 => x"088c08fe",
  2620 => x"f8050854",
  2621 => x"54737326",
  2622 => x"8938800b",
  2623 => x"8c08fee0",
  2624 => x"050c8c08",
  2625 => x"fef40508",
  2626 => x"8c08feec",
  2627 => x"05087171",
  2628 => x"31708c08",
  2629 => x"fee4050c",
  2630 => x"8c08fee4",
  2631 => x"0508708c",
  2632 => x"08fee005",
  2633 => x"0831708c",
  2634 => x"08fee405",
  2635 => x"0c535152",
  2636 => x"54548c08",
  2637 => x"fee40508",
  2638 => x"8c08fee8",
  2639 => x"05085553",
  2640 => x"728c08ff",
  2641 => x"a8050c73",
  2642 => x"8c08ffac",
  2643 => x"050c8c08",
  2644 => x"ffb00508",
  2645 => x"9f2b8c08",
  2646 => x"ffb40508",
  2647 => x"812a7072",
  2648 => x"078c08ff",
  2649 => x"b0050881",
  2650 => x"2a565656",
  2651 => x"56728c08",
  2652 => x"ffb0050c",
  2653 => x"738c08ff",
  2654 => x"b4050c8c",
  2655 => x"08ffa805",
  2656 => x"088c08ff",
  2657 => x"ac050855",
  2658 => x"53728c08",
  2659 => x"fed8050c",
  2660 => x"738c08fe",
  2661 => x"dc050c8c",
  2662 => x"08fed805",
  2663 => x"088c08fe",
  2664 => x"dc050855",
  2665 => x"53728c08",
  2666 => x"fed0050c",
  2667 => x"738c08fe",
  2668 => x"d4050c8c",
  2669 => x"08fed405",
  2670 => x"088c08fe",
  2671 => x"dc050870",
  2672 => x"12708c08",
  2673 => x"fecc050c",
  2674 => x"52545481",
  2675 => x"0b8c08fe",
  2676 => x"c4050c8c",
  2677 => x"08fecc05",
  2678 => x"088c08fe",
  2679 => x"d4050854",
  2680 => x"54727426",
  2681 => x"8938800b",
  2682 => x"8c08fec4",
  2683 => x"050c8c08",
  2684 => x"fed00508",
  2685 => x"8c08fed8",
  2686 => x"05087012",
  2687 => x"708c08fe",
  2688 => x"c8050c8c",
  2689 => x"08fec805",
  2690 => x"088c08fe",
  2691 => x"c4050811",
  2692 => x"708c08fe",
  2693 => x"c8050c53",
  2694 => x"51525454",
  2695 => x"8c08fec8",
  2696 => x"05088c08",
  2697 => x"fecc0508",
  2698 => x"5553728c",
  2699 => x"08ffa805",
  2700 => x"0c738c08",
  2701 => x"ffac050c",
  2702 => x"fbe2398c",
  2703 => x"08ff9805",
  2704 => x"08800670",
  2705 => x"8c08febc",
  2706 => x"050c8c08",
  2707 => x"ff9c0508",
  2708 => x"81ff0670",
  2709 => x"8c08fec0",
  2710 => x"050c5454",
  2711 => x"8c08febc",
  2712 => x"05088c08",
  2713 => x"fec00508",
  2714 => x"5553728c",
  2715 => x"08febc05",
  2716 => x"0c738c08",
  2717 => x"fec0050c",
  2718 => x"8c08febc",
  2719 => x"05085473",
  2720 => x"83bc388c",
  2721 => x"08fec005",
  2722 => x"08537281",
  2723 => x"802e0981",
  2724 => x"0683ab38",
  2725 => x"8c08ff98",
  2726 => x"0508982b",
  2727 => x"8c08ff9c",
  2728 => x"0508882a",
  2729 => x"7072078c",
  2730 => x"08ff9805",
  2731 => x"08882a71",
  2732 => x"81065156",
  2733 => x"56565672",
  2734 => x"802e81b8",
  2735 => x"388c08ff",
  2736 => x"9805088c",
  2737 => x"08ff9c05",
  2738 => x"08555372",
  2739 => x"8c08feb4",
  2740 => x"050c738c",
  2741 => x"08feb805",
  2742 => x"0c805381",
  2743 => x"8054728c",
  2744 => x"08feac05",
  2745 => x"0c738c08",
  2746 => x"feb0050c",
  2747 => x"8c08feb8",
  2748 => x"05088c08",
  2749 => x"feb00508",
  2750 => x"7012708c",
  2751 => x"08fea805",
  2752 => x"0c525454",
  2753 => x"810b8c08",
  2754 => x"fea0050c",
  2755 => x"8c08fea8",
  2756 => x"05088c08",
  2757 => x"feb80508",
  2758 => x"54547274",
  2759 => x"26893880",
  2760 => x"0b8c08fe",
  2761 => x"a0050c8c",
  2762 => x"08feb405",
  2763 => x"088c08fe",
  2764 => x"ac050870",
  2765 => x"12708c08",
  2766 => x"fea4050c",
  2767 => x"8c08fea4",
  2768 => x"05088c08",
  2769 => x"fea00508",
  2770 => x"11708c08",
  2771 => x"fea4050c",
  2772 => x"53515254",
  2773 => x"548c08fe",
  2774 => x"a405088c",
  2775 => x"08fea805",
  2776 => x"08555372",
  2777 => x"8c08ff98",
  2778 => x"050c738c",
  2779 => x"08ff9c05",
  2780 => x"0c81cb39",
  2781 => x"8c08ffa8",
  2782 => x"0508708c",
  2783 => x"08ffac05",
  2784 => x"08075153",
  2785 => x"72802e81",
  2786 => x"b5388c08",
  2787 => x"ff980508",
  2788 => x"8c08ff9c",
  2789 => x"05085553",
  2790 => x"728c08fe",
  2791 => x"98050c73",
  2792 => x"8c08fe9c",
  2793 => x"050c8053",
  2794 => x"81805472",
  2795 => x"8c08fe90",
  2796 => x"050c738c",
  2797 => x"08fe9405",
  2798 => x"0c8c08fe",
  2799 => x"9c05088c",
  2800 => x"08fe9405",
  2801 => x"08701270",
  2802 => x"8c08fe8c",
  2803 => x"050c5254",
  2804 => x"54810b8c",
  2805 => x"08fe8405",
  2806 => x"0c8c08fe",
  2807 => x"8c05088c",
  2808 => x"08fe9c05",
  2809 => x"08545472",
  2810 => x"74268938",
  2811 => x"800b8c08",
  2812 => x"fe84050c",
  2813 => x"8c08fe98",
  2814 => x"05088c08",
  2815 => x"fe900508",
  2816 => x"7012708c",
  2817 => x"08fe8805",
  2818 => x"0c8c08fe",
  2819 => x"8805088c",
  2820 => x"08fe8405",
  2821 => x"0811708c",
  2822 => x"08fe8805",
  2823 => x"0c535152",
  2824 => x"54548c08",
  2825 => x"fe880508",
  2826 => x"8c08fe8c",
  2827 => x"05085553",
  2828 => x"728c08ff",
  2829 => x"98050c73",
  2830 => x"8c08ff9c",
  2831 => x"050c8c08",
  2832 => x"c0050855",
  2833 => x"8c08ff98",
  2834 => x"05088c08",
  2835 => x"ff9c0508",
  2836 => x"5553728c",
  2837 => x"160c7390",
  2838 => x"160c8c08",
  2839 => x"c005088c",
  2840 => x"08ffb805",
  2841 => x"0c8c08ff",
  2842 => x"b8050870",
  2843 => x"8c08d405",
  2844 => x"0c8c08d4",
  2845 => x"0508538c",
  2846 => x"08880508",
  2847 => x"52538cca",
  2848 => x"3f8c0888",
  2849 => x"0508800c",
  2850 => x"80c63d0d",
  2851 => x"8c0c048c",
  2852 => x"08028c0c",
  2853 => x"803d0d82",
  2854 => x"c3d87080",
  2855 => x"0c51823d",
  2856 => x"0d8c0c04",
  2857 => x"8c08028c",
  2858 => x"0cff3d0d",
  2859 => x"800b8c08",
  2860 => x"fc050c8c",
  2861 => x"08880508",
  2862 => x"51700882",
  2863 => x"2e098106",
  2864 => x"8838810b",
  2865 => x"8c08fc05",
  2866 => x"0c8c08fc",
  2867 => x"05087080",
  2868 => x"0c51833d",
  2869 => x"0d8c0c04",
  2870 => x"8c08028c",
  2871 => x"0cff3d0d",
  2872 => x"800b8c08",
  2873 => x"fc050c8c",
  2874 => x"08880508",
  2875 => x"51700884",
  2876 => x"2e098106",
  2877 => x"8838810b",
  2878 => x"8c08fc05",
  2879 => x"0c8c08fc",
  2880 => x"05087080",
  2881 => x"0c51833d",
  2882 => x"0d8c0c04",
  2883 => x"8c08028c",
  2884 => x"0cff3d0d",
  2885 => x"800b8c08",
  2886 => x"fc050c8c",
  2887 => x"08880508",
  2888 => x"51700880",
  2889 => x"2e8f388c",
  2890 => x"08880508",
  2891 => x"51700881",
  2892 => x"2e833888",
  2893 => x"39810b8c",
  2894 => x"08fc050c",
  2895 => x"8c08fc05",
  2896 => x"0870800c",
  2897 => x"51833d0d",
  2898 => x"8c0c048c",
  2899 => x"08028c0c",
  2900 => x"f63d0d83",
  2901 => x"0b8c08ec",
  2902 => x"050c800b",
  2903 => x"8c08e805",
  2904 => x"0c8c088c",
  2905 => x"05088025",
  2906 => x"8838810b",
  2907 => x"8c08e805",
  2908 => x"0c8c08e8",
  2909 => x"05088c08",
  2910 => x"f0050c8c",
  2911 => x"088c0508",
  2912 => x"8b38820b",
  2913 => x"8c08ec05",
  2914 => x"0c819e39",
  2915 => x"bc0b8c08",
  2916 => x"f4050c8c",
  2917 => x"08f00508",
  2918 => x"802ebe38",
  2919 => x"8c088c05",
  2920 => x"08810a2e",
  2921 => x"09810698",
  2922 => x"388f830a",
  2923 => x"53800b8c",
  2924 => x"08880508",
  2925 => x"56547275",
  2926 => x"0c738416",
  2927 => x"0c80fa39",
  2928 => x"8c088c05",
  2929 => x"0830708c",
  2930 => x"08fc050c",
  2931 => x"709f2c70",
  2932 => x"8c08f805",
  2933 => x"0c515397",
  2934 => x"398c088c",
  2935 => x"0508708c",
  2936 => x"08fc050c",
  2937 => x"709f2c70",
  2938 => x"8c08f805",
  2939 => x"0c51538c",
  2940 => x"08f80508",
  2941 => x"f00a26b1",
  2942 => x"388c08fc",
  2943 => x"05089f2a",
  2944 => x"8c08f805",
  2945 => x"08107072",
  2946 => x"078c08f8",
  2947 => x"050c8c08",
  2948 => x"fc050810",
  2949 => x"8c08fc05",
  2950 => x"0c8c08f4",
  2951 => x"0508ff05",
  2952 => x"8c08f405",
  2953 => x"0c5454c7",
  2954 => x"398c08ec",
  2955 => x"0570538c",
  2956 => x"08880508",
  2957 => x"52538992",
  2958 => x"3f8c0888",
  2959 => x"0508800c",
  2960 => x"8c3d0d8c",
  2961 => x"0c048c08",
  2962 => x"028c0cf9",
  2963 => x"3d0d800b",
  2964 => x"8c08fc05",
  2965 => x"0c8c0888",
  2966 => x"05088025",
  2967 => x"ab388c08",
  2968 => x"88050830",
  2969 => x"8c088805",
  2970 => x"0c800b8c",
  2971 => x"08f4050c",
  2972 => x"8c08fc05",
  2973 => x"08883881",
  2974 => x"0b8c08f4",
  2975 => x"050c8c08",
  2976 => x"f405088c",
  2977 => x"08fc050c",
  2978 => x"8c088c05",
  2979 => x"088025ab",
  2980 => x"388c088c",
  2981 => x"0508308c",
  2982 => x"088c050c",
  2983 => x"800b8c08",
  2984 => x"f0050c8c",
  2985 => x"08fc0508",
  2986 => x"8838810b",
  2987 => x"8c08f005",
  2988 => x"0c8c08f0",
  2989 => x"05088c08",
  2990 => x"fc050c80",
  2991 => x"538c088c",
  2992 => x"0508528c",
  2993 => x"08880508",
  2994 => x"5181a73f",
  2995 => x"8008708c",
  2996 => x"08f8050c",
  2997 => x"548c08fc",
  2998 => x"0508802e",
  2999 => x"8c388c08",
  3000 => x"f8050830",
  3001 => x"8c08f805",
  3002 => x"0c8c08f8",
  3003 => x"05087080",
  3004 => x"0c54893d",
  3005 => x"0d8c0c04",
  3006 => x"8c08028c",
  3007 => x"0cfb3d0d",
  3008 => x"800b8c08",
  3009 => x"fc050c8c",
  3010 => x"08880508",
  3011 => x"80259338",
  3012 => x"8c088805",
  3013 => x"08308c08",
  3014 => x"88050c81",
  3015 => x"0b8c08fc",
  3016 => x"050c8c08",
  3017 => x"8c050880",
  3018 => x"258c388c",
  3019 => x"088c0508",
  3020 => x"308c088c",
  3021 => x"050c8153",
  3022 => x"8c088c05",
  3023 => x"08528c08",
  3024 => x"88050851",
  3025 => x"ad3f8008",
  3026 => x"708c08f8",
  3027 => x"050c548c",
  3028 => x"08fc0508",
  3029 => x"802e8c38",
  3030 => x"8c08f805",
  3031 => x"08308c08",
  3032 => x"f8050c8c",
  3033 => x"08f80508",
  3034 => x"70800c54",
  3035 => x"873d0d8c",
  3036 => x"0c048c08",
  3037 => x"028c0cfd",
  3038 => x"3d0d810b",
  3039 => x"8c08fc05",
  3040 => x"0c800b8c",
  3041 => x"08f8050c",
  3042 => x"8c088c05",
  3043 => x"088c0888",
  3044 => x"050827ac",
  3045 => x"388c08fc",
  3046 => x"0508802e",
  3047 => x"a338800b",
  3048 => x"8c088c05",
  3049 => x"08249938",
  3050 => x"8c088c05",
  3051 => x"08108c08",
  3052 => x"8c050c8c",
  3053 => x"08fc0508",
  3054 => x"108c08fc",
  3055 => x"050cc939",
  3056 => x"8c08fc05",
  3057 => x"08802e80",
  3058 => x"c9388c08",
  3059 => x"8c05088c",
  3060 => x"08880508",
  3061 => x"26a1388c",
  3062 => x"08880508",
  3063 => x"8c088c05",
  3064 => x"08318c08",
  3065 => x"88050c8c",
  3066 => x"08f80508",
  3067 => x"8c08fc05",
  3068 => x"08078c08",
  3069 => x"f8050c8c",
  3070 => x"08fc0508",
  3071 => x"812a8c08",
  3072 => x"fc050c8c",
  3073 => x"088c0508",
  3074 => x"812a8c08",
  3075 => x"8c050cff",
  3076 => x"af398c08",
  3077 => x"90050880",
  3078 => x"2e8f388c",
  3079 => x"08880508",
  3080 => x"708c08f4",
  3081 => x"050c518d",
  3082 => x"398c08f8",
  3083 => x"0508708c",
  3084 => x"08f4050c",
  3085 => x"518c08f4",
  3086 => x"0508800c",
  3087 => x"853d0d8c",
  3088 => x"0c048c08",
  3089 => x"028c0ceb",
  3090 => x"3d0d800b",
  3091 => x"8c08f005",
  3092 => x"0c800b8c",
  3093 => x"08f4050c",
  3094 => x"8c088c05",
  3095 => x"088c0890",
  3096 => x"05085654",
  3097 => x"738c08f0",
  3098 => x"050c748c",
  3099 => x"08f4050c",
  3100 => x"8c08f805",
  3101 => x"8c08f005",
  3102 => x"56568870",
  3103 => x"54755376",
  3104 => x"5254a6e9",
  3105 => x"3f800b8c",
  3106 => x"08e8050c",
  3107 => x"800b8c08",
  3108 => x"ec050c8c",
  3109 => x"08940508",
  3110 => x"8c089805",
  3111 => x"08565473",
  3112 => x"8c08e805",
  3113 => x"0c748c08",
  3114 => x"ec050c8c",
  3115 => x"08f0058c",
  3116 => x"08e80556",
  3117 => x"56887054",
  3118 => x"75537652",
  3119 => x"54a6ae3f",
  3120 => x"800b8c08",
  3121 => x"e8050c80",
  3122 => x"0b8c08ec",
  3123 => x"050c8c08",
  3124 => x"fc050883",
  3125 => x"ffff068c",
  3126 => x"08cc050c",
  3127 => x"8c08fc05",
  3128 => x"08902a8c",
  3129 => x"08c4050c",
  3130 => x"8c08f405",
  3131 => x"0883ffff",
  3132 => x"068c08c8",
  3133 => x"050c8c08",
  3134 => x"f4050890",
  3135 => x"2a8c08c0",
  3136 => x"050c8c08",
  3137 => x"cc05088c",
  3138 => x"08c80508",
  3139 => x"29708c08",
  3140 => x"dc050c8c",
  3141 => x"08cc0508",
  3142 => x"8c08c005",
  3143 => x"0829708c",
  3144 => x"08d8050c",
  3145 => x"8c08c405",
  3146 => x"088c08c8",
  3147 => x"05082970",
  3148 => x"8c08d405",
  3149 => x"0c8c08c4",
  3150 => x"05088c08",
  3151 => x"c0050829",
  3152 => x"708c08d0",
  3153 => x"050c8c08",
  3154 => x"dc050890",
  3155 => x"2a8c08d8",
  3156 => x"0508118c",
  3157 => x"08d8050c",
  3158 => x"8c08d805",
  3159 => x"088c08d4",
  3160 => x"0508058c",
  3161 => x"08d8050c",
  3162 => x"51515151",
  3163 => x"548c08d8",
  3164 => x"05088c08",
  3165 => x"d4050827",
  3166 => x"8f388c08",
  3167 => x"d0050884",
  3168 => x"8080058c",
  3169 => x"08d0050c",
  3170 => x"8c08d805",
  3171 => x"08902a8c",
  3172 => x"08d00508",
  3173 => x"118c08e0",
  3174 => x"050c8c08",
  3175 => x"d8050883",
  3176 => x"ffff0670",
  3177 => x"902b8c08",
  3178 => x"dc050883",
  3179 => x"ffff0670",
  3180 => x"128c08e4",
  3181 => x"050c5257",
  3182 => x"51548c08",
  3183 => x"e005088c",
  3184 => x"08e40508",
  3185 => x"5654738c",
  3186 => x"08e8050c",
  3187 => x"748c08ec",
  3188 => x"050c8c08",
  3189 => x"fc05088c",
  3190 => x"08f00508",
  3191 => x"298c08f8",
  3192 => x"05088c08",
  3193 => x"f4050829",
  3194 => x"70128c08",
  3195 => x"e8050811",
  3196 => x"8c08e805",
  3197 => x"0c515555",
  3198 => x"8c08e805",
  3199 => x"088c08ec",
  3200 => x"05088c08",
  3201 => x"88050858",
  3202 => x"56547376",
  3203 => x"0c748417",
  3204 => x"0c8c0888",
  3205 => x"0508800c",
  3206 => x"973d0d8c",
  3207 => x"0c048c08",
  3208 => x"028c0cf6",
  3209 => x"3d0d800b",
  3210 => x"8c08f005",
  3211 => x"0c800b8c",
  3212 => x"08f4050c",
  3213 => x"8c088c05",
  3214 => x"088c0890",
  3215 => x"05085654",
  3216 => x"738c08f0",
  3217 => x"050c748c",
  3218 => x"08f4050c",
  3219 => x"8c08f805",
  3220 => x"8c08f005",
  3221 => x"56568870",
  3222 => x"54755376",
  3223 => x"5254a38d",
  3224 => x"3f800b8c",
  3225 => x"08f0050c",
  3226 => x"800b8c08",
  3227 => x"f4050c8c",
  3228 => x"08f80508",
  3229 => x"308c08ec",
  3230 => x"050c8c08",
  3231 => x"fc050880",
  3232 => x"2e8d388c",
  3233 => x"08ec0508",
  3234 => x"ff058c08",
  3235 => x"ec050c8c",
  3236 => x"08ec0508",
  3237 => x"8c08f005",
  3238 => x"0c8c08fc",
  3239 => x"0508308c",
  3240 => x"08f4050c",
  3241 => x"8c08f005",
  3242 => x"088c08f4",
  3243 => x"05088c08",
  3244 => x"88050858",
  3245 => x"56547376",
  3246 => x"0c748417",
  3247 => x"0c8c0888",
  3248 => x"0508800c",
  3249 => x"8c3d0d8c",
  3250 => x"0c048c08",
  3251 => x"028c0cc7",
  3252 => x"3d0d8c08",
  3253 => x"8c050855",
  3254 => x"9015088c",
  3255 => x"16085656",
  3256 => x"748c08f0",
  3257 => x"050c758c",
  3258 => x"08f4050c",
  3259 => x"8c088c05",
  3260 => x"08841108",
  3261 => x"8c08ec05",
  3262 => x"0c55800b",
  3263 => x"8c08e805",
  3264 => x"0c8c088c",
  3265 => x"0508518f",
  3266 => x"b83f8008",
  3267 => x"5574802e",
  3268 => x"aa388fff",
  3269 => x"0b8c08e8",
  3270 => x"050c8c08",
  3271 => x"f00508a0",
  3272 => x"8080078c",
  3273 => x"08f40508",
  3274 => x"80075755",
  3275 => x"748c08f0",
  3276 => x"050c758c",
  3277 => x"08f4050c",
  3278 => x"8d80398c",
  3279 => x"088c0508",
  3280 => x"518eca3f",
  3281 => x"80085574",
  3282 => x"802e9c38",
  3283 => x"8fff0b8c",
  3284 => x"08e8050c",
  3285 => x"80558056",
  3286 => x"748c08f0",
  3287 => x"050c758c",
  3288 => x"08f4050c",
  3289 => x"8cd4398c",
  3290 => x"088c0508",
  3291 => x"518dea3f",
  3292 => x"80085574",
  3293 => x"802e9b38",
  3294 => x"800b8c08",
  3295 => x"e8050c80",
  3296 => x"55805674",
  3297 => x"8c08f005",
  3298 => x"0c758c08",
  3299 => x"f4050c8c",
  3300 => x"a9398c08",
  3301 => x"f0050870",
  3302 => x"8c08f405",
  3303 => x"08075155",
  3304 => x"748b3880",
  3305 => x"0b8c08e8",
  3306 => x"050c8c8e",
  3307 => x"398c088c",
  3308 => x"05085588",
  3309 => x"1508f882",
  3310 => x"2586fc38",
  3311 => x"8c088c05",
  3312 => x"08f8820b",
  3313 => x"88120831",
  3314 => x"8c08e405",
  3315 => x"0c55800b",
  3316 => x"8c08e805",
  3317 => x"0cb80b8c",
  3318 => x"08e40508",
  3319 => x"25943880",
  3320 => x"55805674",
  3321 => x"8c08f005",
  3322 => x"0c758c08",
  3323 => x"f4050c82",
  3324 => x"a339800b",
  3325 => x"8c08e005",
  3326 => x"0c8c08d8",
  3327 => x"05578055",
  3328 => x"810b8c08",
  3329 => x"e4050855",
  3330 => x"56745275",
  3331 => x"537651ff",
  3332 => x"afed3f8c",
  3333 => x"08d80508",
  3334 => x"8c08dc05",
  3335 => x"08575574",
  3336 => x"8c08d005",
  3337 => x"0c758c08",
  3338 => x"d4050cff",
  3339 => x"56ff5775",
  3340 => x"8c08c805",
  3341 => x"0c768c08",
  3342 => x"cc050c8c",
  3343 => x"08d40508",
  3344 => x"8c08cc05",
  3345 => x"08701270",
  3346 => x"8c08c405",
  3347 => x"0c525657",
  3348 => x"810b8c08",
  3349 => x"ffbc050c",
  3350 => x"8c08c405",
  3351 => x"088c08d4",
  3352 => x"05085856",
  3353 => x"76762689",
  3354 => x"38800b8c",
  3355 => x"08ffbc05",
  3356 => x"0c8c08d0",
  3357 => x"05088c08",
  3358 => x"c8050870",
  3359 => x"12708c08",
  3360 => x"c0050c8c",
  3361 => x"08c00508",
  3362 => x"8c08ffbc",
  3363 => x"05081170",
  3364 => x"8c08c005",
  3365 => x"0c8c08c0",
  3366 => x"0508708c",
  3367 => x"08f00508",
  3368 => x"068c08c4",
  3369 => x"0508708c",
  3370 => x"08f40508",
  3371 => x"06727072",
  3372 => x"07515257",
  3373 => x"52525252",
  3374 => x"5a525755",
  3375 => x"76802e88",
  3376 => x"38810b8c",
  3377 => x"08e0050c",
  3378 => x"8c08d805",
  3379 => x"8c08e405",
  3380 => x"0855578c",
  3381 => x"08f00508",
  3382 => x"8c08f405",
  3383 => x"08575574",
  3384 => x"52755376",
  3385 => x"518ff73f",
  3386 => x"8c08d805",
  3387 => x"088c08dc",
  3388 => x"05088c08",
  3389 => x"e005089f",
  3390 => x"2c8c08e0",
  3391 => x"05087170",
  3392 => x"75078c08",
  3393 => x"f0050c73",
  3394 => x"72078c08",
  3395 => x"f4050c59",
  3396 => x"595b5957",
  3397 => x"8c08f005",
  3398 => x"08800670",
  3399 => x"8c08ffb4",
  3400 => x"050c8c08",
  3401 => x"f4050881",
  3402 => x"ff06708c",
  3403 => x"08ffb805",
  3404 => x"0c57558c",
  3405 => x"08ffb405",
  3406 => x"088c08ff",
  3407 => x"b8050857",
  3408 => x"55748c08",
  3409 => x"ffb4050c",
  3410 => x"758c08ff",
  3411 => x"b8050c8c",
  3412 => x"08ffb405",
  3413 => x"08567581",
  3414 => x"eb388c08",
  3415 => x"ffb80508",
  3416 => x"57768180",
  3417 => x"2e098106",
  3418 => x"81da388c",
  3419 => x"08f00508",
  3420 => x"982b8c08",
  3421 => x"f4050888",
  3422 => x"2a707207",
  3423 => x"8c08f005",
  3424 => x"08882a71",
  3425 => x"81065158",
  3426 => x"58585874",
  3427 => x"802e82e4",
  3428 => x"388c08f0",
  3429 => x"05088c08",
  3430 => x"f4050857",
  3431 => x"55748c08",
  3432 => x"ffac050c",
  3433 => x"758c08ff",
  3434 => x"b0050c80",
  3435 => x"56818057",
  3436 => x"758c08ff",
  3437 => x"a4050c76",
  3438 => x"8c08ffa8",
  3439 => x"050c8c08",
  3440 => x"ffb00508",
  3441 => x"8c08ffa8",
  3442 => x"05087012",
  3443 => x"708c08ff",
  3444 => x"a0050c52",
  3445 => x"5657810b",
  3446 => x"8c08ff98",
  3447 => x"050c8c08",
  3448 => x"ffa00508",
  3449 => x"8c08ffb0",
  3450 => x"05085856",
  3451 => x"76762689",
  3452 => x"38800b8c",
  3453 => x"08ff9805",
  3454 => x"0c8c08ff",
  3455 => x"ac05088c",
  3456 => x"08ffa405",
  3457 => x"08701270",
  3458 => x"8c08ff9c",
  3459 => x"050c8c08",
  3460 => x"ff9c0508",
  3461 => x"8c08ff98",
  3462 => x"05081170",
  3463 => x"8c08ff9c",
  3464 => x"050c525a",
  3465 => x"5257558c",
  3466 => x"08ff9c05",
  3467 => x"088c08ff",
  3468 => x"a0050857",
  3469 => x"55748c08",
  3470 => x"f0050c75",
  3471 => x"8c08f405",
  3472 => x"0c81b139",
  3473 => x"8c08f005",
  3474 => x"088c08f4",
  3475 => x"05085856",
  3476 => x"758c08ff",
  3477 => x"90050c76",
  3478 => x"8c08ff94",
  3479 => x"050c8055",
  3480 => x"80ff5674",
  3481 => x"8c08ff88",
  3482 => x"050c758c",
  3483 => x"08ff8c05",
  3484 => x"0c8c08ff",
  3485 => x"9405088c",
  3486 => x"08ff8c05",
  3487 => x"08701270",
  3488 => x"8c08ff84",
  3489 => x"050c5258",
  3490 => x"56810b8c",
  3491 => x"08fefc05",
  3492 => x"0c8c08ff",
  3493 => x"8405088c",
  3494 => x"08ff9405",
  3495 => x"08575575",
  3496 => x"75268938",
  3497 => x"800b8c08",
  3498 => x"fefc050c",
  3499 => x"8c08ff90",
  3500 => x"05088c08",
  3501 => x"ff880508",
  3502 => x"7012708c",
  3503 => x"08ff8005",
  3504 => x"0c8c08ff",
  3505 => x"8005088c",
  3506 => x"08fefc05",
  3507 => x"0811708c",
  3508 => x"08ff8005",
  3509 => x"0c535952",
  3510 => x"56578c08",
  3511 => x"ff800508",
  3512 => x"8c08ff84",
  3513 => x"05085755",
  3514 => x"748c08f0",
  3515 => x"050c758c",
  3516 => x"08f4050c",
  3517 => x"8c08f005",
  3518 => x"08f00a26",
  3519 => x"83388d39",
  3520 => x"8c08e805",
  3521 => x"0881058c",
  3522 => x"08e8050c",
  3523 => x"8c08f005",
  3524 => x"08982b8c",
  3525 => x"08f40508",
  3526 => x"882a7072",
  3527 => x"078c08f0",
  3528 => x"0508882a",
  3529 => x"58585858",
  3530 => x"748c08f0",
  3531 => x"050c758c",
  3532 => x"08f4050c",
  3533 => x"8584398c",
  3534 => x"088c0508",
  3535 => x"5587ff0b",
  3536 => x"88160825",
  3537 => x"9c388fff",
  3538 => x"0b8c08e8",
  3539 => x"050c8055",
  3540 => x"8056748c",
  3541 => x"08f0050c",
  3542 => x"758c08f4",
  3543 => x"050c84da",
  3544 => x"398c088c",
  3545 => x"05088811",
  3546 => x"0887ff05",
  3547 => x"8c08e805",
  3548 => x"0c8c08f0",
  3549 => x"05088006",
  3550 => x"708c08fe",
  3551 => x"f4050c8c",
  3552 => x"08f40508",
  3553 => x"81ff0670",
  3554 => x"8c08fef8",
  3555 => x"050c5957",
  3556 => x"558c08fe",
  3557 => x"f405088c",
  3558 => x"08fef805",
  3559 => x"08575574",
  3560 => x"8c08fef4",
  3561 => x"050c758c",
  3562 => x"08fef805",
  3563 => x"0c8c08fe",
  3564 => x"f4050856",
  3565 => x"7581eb38",
  3566 => x"8c08fef8",
  3567 => x"05085776",
  3568 => x"81802e09",
  3569 => x"810681da",
  3570 => x"388c08f0",
  3571 => x"0508982b",
  3572 => x"8c08f405",
  3573 => x"08882a70",
  3574 => x"72078c08",
  3575 => x"f0050888",
  3576 => x"2a718106",
  3577 => x"51585858",
  3578 => x"5874802e",
  3579 => x"82e4388c",
  3580 => x"08f00508",
  3581 => x"8c08f405",
  3582 => x"08575574",
  3583 => x"8c08feec",
  3584 => x"050c758c",
  3585 => x"08fef005",
  3586 => x"0c805681",
  3587 => x"8057758c",
  3588 => x"08fee405",
  3589 => x"0c768c08",
  3590 => x"fee8050c",
  3591 => x"8c08fef0",
  3592 => x"05088c08",
  3593 => x"fee80508",
  3594 => x"7012708c",
  3595 => x"08fee005",
  3596 => x"0c525657",
  3597 => x"810b8c08",
  3598 => x"fed8050c",
  3599 => x"8c08fee0",
  3600 => x"05088c08",
  3601 => x"fef00508",
  3602 => x"58567676",
  3603 => x"26893880",
  3604 => x"0b8c08fe",
  3605 => x"d8050c8c",
  3606 => x"08feec05",
  3607 => x"088c08fe",
  3608 => x"e4050870",
  3609 => x"12708c08",
  3610 => x"fedc050c",
  3611 => x"8c08fedc",
  3612 => x"05088c08",
  3613 => x"fed80508",
  3614 => x"11708c08",
  3615 => x"fedc050c",
  3616 => x"525a5257",
  3617 => x"558c08fe",
  3618 => x"dc05088c",
  3619 => x"08fee005",
  3620 => x"08575574",
  3621 => x"8c08f005",
  3622 => x"0c758c08",
  3623 => x"f4050c81",
  3624 => x"b1398c08",
  3625 => x"f005088c",
  3626 => x"08f40508",
  3627 => x"5856758c",
  3628 => x"08fed005",
  3629 => x"0c768c08",
  3630 => x"fed4050c",
  3631 => x"805580ff",
  3632 => x"56748c08",
  3633 => x"fec8050c",
  3634 => x"758c08fe",
  3635 => x"cc050c8c",
  3636 => x"08fed405",
  3637 => x"088c08fe",
  3638 => x"cc050870",
  3639 => x"12708c08",
  3640 => x"fec4050c",
  3641 => x"52585681",
  3642 => x"0b8c08fe",
  3643 => x"bc050c8c",
  3644 => x"08fec405",
  3645 => x"088c08fe",
  3646 => x"d4050857",
  3647 => x"55757526",
  3648 => x"8938800b",
  3649 => x"8c08febc",
  3650 => x"050c8c08",
  3651 => x"fed00508",
  3652 => x"8c08fec8",
  3653 => x"05087012",
  3654 => x"708c08fe",
  3655 => x"c0050c8c",
  3656 => x"08fec005",
  3657 => x"088c08fe",
  3658 => x"bc050811",
  3659 => x"708c08fe",
  3660 => x"c0050c53",
  3661 => x"59525657",
  3662 => x"8c08fec0",
  3663 => x"05088c08",
  3664 => x"fec40508",
  3665 => x"5755748c",
  3666 => x"08f0050c",
  3667 => x"758c08f4",
  3668 => x"050c8c08",
  3669 => x"f00508f8",
  3670 => x"0a268338",
  3671 => x"b5398c08",
  3672 => x"f005089f",
  3673 => x"2b8c08f4",
  3674 => x"0508812a",
  3675 => x"7072078c",
  3676 => x"08f00508",
  3677 => x"812a5858",
  3678 => x"5858748c",
  3679 => x"08f0050c",
  3680 => x"758c08f4",
  3681 => x"050c8c08",
  3682 => x"e8050881",
  3683 => x"058c08e8",
  3684 => x"050c8c08",
  3685 => x"f0050898",
  3686 => x"2b8c08f4",
  3687 => x"0508882a",
  3688 => x"7072078c",
  3689 => x"08f00508",
  3690 => x"882a5858",
  3691 => x"5858748c",
  3692 => x"08f0050c",
  3693 => x"758c08f4",
  3694 => x"050c8c08",
  3695 => x"f00508bf",
  3696 => x"ffff068c",
  3697 => x"08f8050c",
  3698 => x"8c08f405",
  3699 => x"08ff068c",
  3700 => x"08fc050c",
  3701 => x"8c08e805",
  3702 => x"08568070",
  3703 => x"8006778f",
  3704 => x"ff067094",
  3705 => x"2b535a58",
  3706 => x"55800b8c",
  3707 => x"08f80508",
  3708 => x"76078c08",
  3709 => x"f8050c70",
  3710 => x"8c08fc05",
  3711 => x"08078c08",
  3712 => x"fc050c8c",
  3713 => x"08ec0508",
  3714 => x"51568070",
  3715 => x"80067781",
  3716 => x"06709f2b",
  3717 => x"535a5855",
  3718 => x"800b8c08",
  3719 => x"f8050876",
  3720 => x"078c08f8",
  3721 => x"050c708c",
  3722 => x"08fc0508",
  3723 => x"078c08fc",
  3724 => x"050c568c",
  3725 => x"08f80508",
  3726 => x"8c08fc05",
  3727 => x"088c0888",
  3728 => x"05085957",
  3729 => x"5574770c",
  3730 => x"7584180c",
  3731 => x"8c088805",
  3732 => x"08800cbb",
  3733 => x"3d0d8c0c",
  3734 => x"048c0802",
  3735 => x"8c0cff3d",
  3736 => x"0d800b8c",
  3737 => x"08fc050c",
  3738 => x"8c088805",
  3739 => x"08517008",
  3740 => x"822e0981",
  3741 => x"06883881",
  3742 => x"0b8c08fc",
  3743 => x"050c8c08",
  3744 => x"fc050870",
  3745 => x"800c5183",
  3746 => x"3d0d8c0c",
  3747 => x"048c0802",
  3748 => x"8c0cff3d",
  3749 => x"0d800b8c",
  3750 => x"08fc050c",
  3751 => x"8c088805",
  3752 => x"08517008",
  3753 => x"842e0981",
  3754 => x"06883881",
  3755 => x"0b8c08fc",
  3756 => x"050c8c08",
  3757 => x"fc050870",
  3758 => x"800c5183",
  3759 => x"3d0d8c0c",
  3760 => x"048c0802",
  3761 => x"8c0cff3d",
  3762 => x"0d800b8c",
  3763 => x"08fc050c",
  3764 => x"8c088805",
  3765 => x"08517008",
  3766 => x"802e8f38",
  3767 => x"8c088805",
  3768 => x"08517008",
  3769 => x"812e8338",
  3770 => x"8839810b",
  3771 => x"8c08fc05",
  3772 => x"0c8c08fc",
  3773 => x"05087080",
  3774 => x"0c51833d",
  3775 => x"0d8c0c04",
  3776 => x"8c08028c",
  3777 => x"0cf83d0d",
  3778 => x"8c088805",
  3779 => x"087008bf",
  3780 => x"ffff068c",
  3781 => x"08f8050c",
  3782 => x"841108ff",
  3783 => x"068c08fc",
  3784 => x"050c8c08",
  3785 => x"88050870",
  3786 => x"08942a54",
  3787 => x"54518072",
  3788 => x"8fff068c",
  3789 => x"08f4050c",
  3790 => x"8c088805",
  3791 => x"0870089f",
  3792 => x"2a545451",
  3793 => x"80728106",
  3794 => x"8c08f005",
  3795 => x"0c8c088c",
  3796 => x"05088c08",
  3797 => x"f0050884",
  3798 => x"120c5151",
  3799 => x"8c08f405",
  3800 => x"0881bd38",
  3801 => x"8c08f805",
  3802 => x"08708c08",
  3803 => x"fc050807",
  3804 => x"5151708d",
  3805 => x"388c088c",
  3806 => x"05085182",
  3807 => x"710c82d8",
  3808 => x"398c088c",
  3809 => x"05088c08",
  3810 => x"f40508f8",
  3811 => x"82058812",
  3812 => x"0c8c08fc",
  3813 => x"0508982a",
  3814 => x"8c08f805",
  3815 => x"08882b70",
  3816 => x"72078c08",
  3817 => x"fc050888",
  3818 => x"2b565355",
  3819 => x"5551708c",
  3820 => x"08f8050c",
  3821 => x"718c08fc",
  3822 => x"050c8c08",
  3823 => x"8c050851",
  3824 => x"83710c8c",
  3825 => x"08f80508",
  3826 => x"f00a26b7",
  3827 => x"388c08fc",
  3828 => x"05089f2a",
  3829 => x"8c08f805",
  3830 => x"08107072",
  3831 => x"078c08fc",
  3832 => x"05081055",
  3833 => x"53545470",
  3834 => x"8c08f805",
  3835 => x"0c718c08",
  3836 => x"fc050c8c",
  3837 => x"088c0508",
  3838 => x"881108ff",
  3839 => x"0588120c",
  3840 => x"51c1398c",
  3841 => x"088c0508",
  3842 => x"538c08f8",
  3843 => x"05088c08",
  3844 => x"fc050853",
  3845 => x"51708c14",
  3846 => x"0c719014",
  3847 => x"0c81b939",
  3848 => x"8c08f405",
  3849 => x"088fff2e",
  3850 => x"09810680",
  3851 => x"e2388c08",
  3852 => x"f8050870",
  3853 => x"8c08fc05",
  3854 => x"08075151",
  3855 => x"708d388c",
  3856 => x"088c0508",
  3857 => x"5184710c",
  3858 => x"818e398c",
  3859 => x"08f80508",
  3860 => x"932a5280",
  3861 => x"72810651",
  3862 => x"5170802e",
  3863 => x"8c388c08",
  3864 => x"8c050851",
  3865 => x"81710c8a",
  3866 => x"398c088c",
  3867 => x"05085180",
  3868 => x"710c8c08",
  3869 => x"8c050853",
  3870 => x"8c08f805",
  3871 => x"088c08fc",
  3872 => x"05085351",
  3873 => x"708c140c",
  3874 => x"7190140c",
  3875 => x"80ca398c",
  3876 => x"088c0508",
  3877 => x"8c08f405",
  3878 => x"08f88105",
  3879 => x"88120c8c",
  3880 => x"088c0508",
  3881 => x"51518371",
  3882 => x"0c8c088c",
  3883 => x"05088c08",
  3884 => x"fc050898",
  3885 => x"2a8c08f8",
  3886 => x"0508882b",
  3887 => x"7072078c",
  3888 => x"08fc0508",
  3889 => x"882b7188",
  3890 => x"0a078c16",
  3891 => x"0c708007",
  3892 => x"90160c56",
  3893 => x"54555555",
  3894 => x"8a3d0d8c",
  3895 => x"0c048c08",
  3896 => x"028c0cf5",
  3897 => x"3d0d8c08",
  3898 => x"9405089d",
  3899 => x"388c088c",
  3900 => x"05088c08",
  3901 => x"9005088c",
  3902 => x"08880508",
  3903 => x"58565473",
  3904 => x"760c7484",
  3905 => x"170c81bf",
  3906 => x"39800b8c",
  3907 => x"08f0050c",
  3908 => x"800b8c08",
  3909 => x"f4050c8c",
  3910 => x"088c0508",
  3911 => x"8c089005",
  3912 => x"08565473",
  3913 => x"8c08f005",
  3914 => x"0c748c08",
  3915 => x"f4050c8c",
  3916 => x"08f8058c",
  3917 => x"08f00556",
  3918 => x"56887054",
  3919 => x"75537652",
  3920 => x"548daa3f",
  3921 => x"a00b8c08",
  3922 => x"94050831",
  3923 => x"8c08ec05",
  3924 => x"0c8c08ec",
  3925 => x"05088024",
  3926 => x"9d38800b",
  3927 => x"8c08f005",
  3928 => x"0c8c08ec",
  3929 => x"0508308c",
  3930 => x"08f80508",
  3931 => x"712a8c08",
  3932 => x"f4050c54",
  3933 => x"b9398c08",
  3934 => x"f805088c",
  3935 => x"08ec0508",
  3936 => x"2b8c08e8",
  3937 => x"050c8c08",
  3938 => x"f805088c",
  3939 => x"08940508",
  3940 => x"2a8c08f0",
  3941 => x"050c8c08",
  3942 => x"fc05088c",
  3943 => x"08940508",
  3944 => x"2a708c08",
  3945 => x"e8050807",
  3946 => x"8c08f405",
  3947 => x"0c548c08",
  3948 => x"f005088c",
  3949 => x"08f40508",
  3950 => x"8c088805",
  3951 => x"08585654",
  3952 => x"73760c74",
  3953 => x"84170c8c",
  3954 => x"08880508",
  3955 => x"800c8d3d",
  3956 => x"0d8c0c04",
  3957 => x"ff3d0d73",
  3958 => x"5282d480",
  3959 => x"0851973f",
  3960 => x"833d0d04",
  3961 => x"ff3d0d73",
  3962 => x"5282d480",
  3963 => x"085180f0",
  3964 => x"ee3f833d",
  3965 => x"0d04f33d",
  3966 => x"0d7f618b",
  3967 => x"1170f806",
  3968 => x"5c55555e",
  3969 => x"72962683",
  3970 => x"38905980",
  3971 => x"7924747a",
  3972 => x"26075380",
  3973 => x"5472742e",
  3974 => x"09810680",
  3975 => x"cb387d51",
  3976 => x"8ce43f78",
  3977 => x"83f72680",
  3978 => x"c6387883",
  3979 => x"2a701010",
  3980 => x"1082cbf8",
  3981 => x"058c1108",
  3982 => x"59595a76",
  3983 => x"782e83b0",
  3984 => x"38841708",
  3985 => x"fc06568c",
  3986 => x"17088818",
  3987 => x"08718c12",
  3988 => x"0c88120c",
  3989 => x"58751784",
  3990 => x"11088107",
  3991 => x"84120c53",
  3992 => x"7d518ca3",
  3993 => x"3f881754",
  3994 => x"73800c8f",
  3995 => x"3d0d0478",
  3996 => x"892a7983",
  3997 => x"2a5b5372",
  3998 => x"802ebf38",
  3999 => x"78862ab8",
  4000 => x"055a8473",
  4001 => x"27b43880",
  4002 => x"db135a94",
  4003 => x"7327ab38",
  4004 => x"788c2a80",
  4005 => x"ee055a80",
  4006 => x"d473279e",
  4007 => x"38788f2a",
  4008 => x"80f7055a",
  4009 => x"82d47327",
  4010 => x"91387892",
  4011 => x"2a80fc05",
  4012 => x"5a8ad473",
  4013 => x"27843880",
  4014 => x"fe5a7910",
  4015 => x"101082cb",
  4016 => x"f8058c11",
  4017 => x"08585576",
  4018 => x"752ea338",
  4019 => x"841708fc",
  4020 => x"06707a31",
  4021 => x"5556738f",
  4022 => x"2488d538",
  4023 => x"738025fe",
  4024 => x"e6388c17",
  4025 => x"08577675",
  4026 => x"2e098106",
  4027 => x"df38811a",
  4028 => x"5a82cc88",
  4029 => x"08577682",
  4030 => x"cc802e82",
  4031 => x"c0388417",
  4032 => x"08fc0670",
  4033 => x"7a315556",
  4034 => x"738f2481",
  4035 => x"f93882cc",
  4036 => x"800b82cc",
  4037 => x"8c0c82cc",
  4038 => x"800b82cc",
  4039 => x"880c7380",
  4040 => x"25feb238",
  4041 => x"83ff7627",
  4042 => x"83df3875",
  4043 => x"892a7683",
  4044 => x"2a555372",
  4045 => x"802ebf38",
  4046 => x"75862ab8",
  4047 => x"05548473",
  4048 => x"27b43880",
  4049 => x"db135494",
  4050 => x"7327ab38",
  4051 => x"758c2a80",
  4052 => x"ee055480",
  4053 => x"d473279e",
  4054 => x"38758f2a",
  4055 => x"80f70554",
  4056 => x"82d47327",
  4057 => x"91387592",
  4058 => x"2a80fc05",
  4059 => x"548ad473",
  4060 => x"27843880",
  4061 => x"fe547310",
  4062 => x"101082cb",
  4063 => x"f8058811",
  4064 => x"08565874",
  4065 => x"782e86cf",
  4066 => x"38841508",
  4067 => x"fc065375",
  4068 => x"73278d38",
  4069 => x"88150855",
  4070 => x"74782e09",
  4071 => x"8106ea38",
  4072 => x"8c150882",
  4073 => x"cbf80b84",
  4074 => x"0508718c",
  4075 => x"1a0c7688",
  4076 => x"1a0c7888",
  4077 => x"130c788c",
  4078 => x"180c5d58",
  4079 => x"7953807a",
  4080 => x"2483e638",
  4081 => x"72822c81",
  4082 => x"712b5c53",
  4083 => x"7a7c2681",
  4084 => x"98387b7b",
  4085 => x"06537282",
  4086 => x"f13879fc",
  4087 => x"0684055a",
  4088 => x"7a10707d",
  4089 => x"06545b72",
  4090 => x"82e03884",
  4091 => x"1a5af139",
  4092 => x"88178c11",
  4093 => x"08585876",
  4094 => x"782e0981",
  4095 => x"06fcc238",
  4096 => x"821a5afd",
  4097 => x"ec397817",
  4098 => x"79810784",
  4099 => x"190c7082",
  4100 => x"cc8c0c70",
  4101 => x"82cc880c",
  4102 => x"82cc800b",
  4103 => x"8c120c8c",
  4104 => x"11088812",
  4105 => x"0c748107",
  4106 => x"84120c74",
  4107 => x"1175710c",
  4108 => x"51537d51",
  4109 => x"88d13f88",
  4110 => x"1754fcac",
  4111 => x"3982cbf8",
  4112 => x"0b840508",
  4113 => x"7a545c79",
  4114 => x"8025fef8",
  4115 => x"3882da39",
  4116 => x"7a097c06",
  4117 => x"7082cbf8",
  4118 => x"0b84050c",
  4119 => x"5c7a105b",
  4120 => x"7a7c2685",
  4121 => x"387a85b8",
  4122 => x"3882cbf8",
  4123 => x"0b880508",
  4124 => x"70841208",
  4125 => x"fc06707c",
  4126 => x"317c7226",
  4127 => x"8f722507",
  4128 => x"57575c5d",
  4129 => x"5572802e",
  4130 => x"80db3879",
  4131 => x"7a1682cb",
  4132 => x"f0081b90",
  4133 => x"115a5557",
  4134 => x"5b82cbec",
  4135 => x"08ff2e88",
  4136 => x"38a08f13",
  4137 => x"e0800657",
  4138 => x"76527d51",
  4139 => x"88903f80",
  4140 => x"08548008",
  4141 => x"ff2e9038",
  4142 => x"80087627",
  4143 => x"82993874",
  4144 => x"82cbf82e",
  4145 => x"82913882",
  4146 => x"cbf80b88",
  4147 => x"05085584",
  4148 => x"1508fc06",
  4149 => x"707a317a",
  4150 => x"72268f72",
  4151 => x"25075255",
  4152 => x"537283e6",
  4153 => x"38747981",
  4154 => x"0784170c",
  4155 => x"79167082",
  4156 => x"cbf80b88",
  4157 => x"050c7581",
  4158 => x"0784120c",
  4159 => x"547e5257",
  4160 => x"87853f88",
  4161 => x"1754fae0",
  4162 => x"3975832a",
  4163 => x"70545480",
  4164 => x"7424819b",
  4165 => x"3872822c",
  4166 => x"81712b82",
  4167 => x"cbfc0807",
  4168 => x"7082cbf8",
  4169 => x"0b84050c",
  4170 => x"75101010",
  4171 => x"82cbf805",
  4172 => x"88110858",
  4173 => x"5a5d5377",
  4174 => x"8c180c74",
  4175 => x"88180c76",
  4176 => x"88190c76",
  4177 => x"8c160cfc",
  4178 => x"f339797a",
  4179 => x"10101082",
  4180 => x"cbf80570",
  4181 => x"57595d8c",
  4182 => x"15085776",
  4183 => x"752ea338",
  4184 => x"841708fc",
  4185 => x"06707a31",
  4186 => x"5556738f",
  4187 => x"2483ca38",
  4188 => x"73802584",
  4189 => x"81388c17",
  4190 => x"08577675",
  4191 => x"2e098106",
  4192 => x"df388815",
  4193 => x"811b7083",
  4194 => x"06555b55",
  4195 => x"72c9387c",
  4196 => x"83065372",
  4197 => x"802efdb8",
  4198 => x"38ff1df8",
  4199 => x"19595d88",
  4200 => x"1808782e",
  4201 => x"ea38fdb5",
  4202 => x"39831a53",
  4203 => x"fc963983",
  4204 => x"1470822c",
  4205 => x"81712b82",
  4206 => x"cbfc0807",
  4207 => x"7082cbf8",
  4208 => x"0b84050c",
  4209 => x"76101010",
  4210 => x"82cbf805",
  4211 => x"88110859",
  4212 => x"5b5e5153",
  4213 => x"fee13982",
  4214 => x"cbbc0817",
  4215 => x"58800876",
  4216 => x"2e818d38",
  4217 => x"82cbec08",
  4218 => x"ff2e83ed",
  4219 => x"38737631",
  4220 => x"1882cbbc",
  4221 => x"0c738706",
  4222 => x"70575372",
  4223 => x"802e8838",
  4224 => x"88733170",
  4225 => x"15555676",
  4226 => x"149fff06",
  4227 => x"a0807131",
  4228 => x"1770547f",
  4229 => x"53575385",
  4230 => x"a53f8008",
  4231 => x"538008ff",
  4232 => x"2e81a038",
  4233 => x"82cbbc08",
  4234 => x"167082cb",
  4235 => x"bc0c7475",
  4236 => x"82cbf80b",
  4237 => x"88050c74",
  4238 => x"76311870",
  4239 => x"81075155",
  4240 => x"56587b82",
  4241 => x"cbf82e83",
  4242 => x"9d38798f",
  4243 => x"2682cb38",
  4244 => x"810b8415",
  4245 => x"0c841508",
  4246 => x"fc06707a",
  4247 => x"317a7226",
  4248 => x"8f722507",
  4249 => x"52555372",
  4250 => x"802efcf9",
  4251 => x"3880db39",
  4252 => x"80089fff",
  4253 => x"065372fe",
  4254 => x"eb387782",
  4255 => x"cbbc0c82",
  4256 => x"cbf80b88",
  4257 => x"05087b18",
  4258 => x"81078412",
  4259 => x"0c5582cb",
  4260 => x"e8087827",
  4261 => x"86387782",
  4262 => x"cbe80c82",
  4263 => x"cbe40878",
  4264 => x"27fcac38",
  4265 => x"7782cbe4",
  4266 => x"0c841508",
  4267 => x"fc06707a",
  4268 => x"317a7226",
  4269 => x"8f722507",
  4270 => x"52555372",
  4271 => x"802efca5",
  4272 => x"38883980",
  4273 => x"745456fe",
  4274 => x"db397d51",
  4275 => x"83b93f80",
  4276 => x"0b800c8f",
  4277 => x"3d0d0473",
  4278 => x"53807424",
  4279 => x"a9387282",
  4280 => x"2c81712b",
  4281 => x"82cbfc08",
  4282 => x"077082cb",
  4283 => x"f80b8405",
  4284 => x"0c5d5377",
  4285 => x"8c180c74",
  4286 => x"88180c76",
  4287 => x"88190c76",
  4288 => x"8c160cf9",
  4289 => x"b7398314",
  4290 => x"70822c81",
  4291 => x"712b82cb",
  4292 => x"fc080770",
  4293 => x"82cbf80b",
  4294 => x"84050c5e",
  4295 => x"5153d439",
  4296 => x"7b7b0653",
  4297 => x"72fca338",
  4298 => x"841a7b10",
  4299 => x"5c5af139",
  4300 => x"ff1a8111",
  4301 => x"515af7b9",
  4302 => x"39781779",
  4303 => x"81078419",
  4304 => x"0c8c1808",
  4305 => x"88190871",
  4306 => x"8c120c88",
  4307 => x"120c5970",
  4308 => x"82cc8c0c",
  4309 => x"7082cc88",
  4310 => x"0c82cc80",
  4311 => x"0b8c120c",
  4312 => x"8c110888",
  4313 => x"120c7481",
  4314 => x"0784120c",
  4315 => x"74117571",
  4316 => x"0c5153f9",
  4317 => x"bd397517",
  4318 => x"84110881",
  4319 => x"0784120c",
  4320 => x"538c1708",
  4321 => x"88180871",
  4322 => x"8c120c88",
  4323 => x"120c587d",
  4324 => x"5181f43f",
  4325 => x"881754f5",
  4326 => x"cf397284",
  4327 => x"150cf41a",
  4328 => x"f8067084",
  4329 => x"1e088106",
  4330 => x"07841e0c",
  4331 => x"701d545b",
  4332 => x"850b8414",
  4333 => x"0c850b88",
  4334 => x"140c8f7b",
  4335 => x"27fdcf38",
  4336 => x"881c527d",
  4337 => x"5180e597",
  4338 => x"3f82cbf8",
  4339 => x"0b880508",
  4340 => x"82cbbc08",
  4341 => x"5955fdb6",
  4342 => x"397782cb",
  4343 => x"bc0c7382",
  4344 => x"cbec0cfc",
  4345 => x"90397284",
  4346 => x"150cfda2",
  4347 => x"39fc3d0d",
  4348 => x"7670797b",
  4349 => x"55555555",
  4350 => x"8f72278c",
  4351 => x"38727507",
  4352 => x"83065170",
  4353 => x"802ea738",
  4354 => x"ff125271",
  4355 => x"ff2e9838",
  4356 => x"72708105",
  4357 => x"54337470",
  4358 => x"81055634",
  4359 => x"ff125271",
  4360 => x"ff2e0981",
  4361 => x"06ea3874",
  4362 => x"800c863d",
  4363 => x"0d047451",
  4364 => x"72708405",
  4365 => x"54087170",
  4366 => x"8405530c",
  4367 => x"72708405",
  4368 => x"54087170",
  4369 => x"8405530c",
  4370 => x"72708405",
  4371 => x"54087170",
  4372 => x"8405530c",
  4373 => x"72708405",
  4374 => x"54087170",
  4375 => x"8405530c",
  4376 => x"f0125271",
  4377 => x"8f26c938",
  4378 => x"83722795",
  4379 => x"38727084",
  4380 => x"05540871",
  4381 => x"70840553",
  4382 => x"0cfc1252",
  4383 => x"718326ed",
  4384 => x"387054ff",
  4385 => x"83390404",
  4386 => x"fb3d0d77",
  4387 => x"893d8805",
  4388 => x"55795488",
  4389 => x"11085351",
  4390 => x"818a3f87",
  4391 => x"3d0d04fc",
  4392 => x"3d0d873d",
  4393 => x"70708405",
  4394 => x"52085653",
  4395 => x"745282d4",
  4396 => x"80088811",
  4397 => x"085254ab",
  4398 => x"973f863d",
  4399 => x"0d04fd3d",
  4400 => x"0d800b82",
  4401 => x"dc800c76",
  4402 => x"51819bc1",
  4403 => x"3f800853",
  4404 => x"8008ff2e",
  4405 => x"88387280",
  4406 => x"0c853d0d",
  4407 => x"0482dc80",
  4408 => x"08547380",
  4409 => x"2ef03875",
  4410 => x"74710c52",
  4411 => x"72800c85",
  4412 => x"3d0d04fd",
  4413 => x"3d0d7688",
  4414 => x"11085454",
  4415 => x"728c3872",
  4416 => x"84150c72",
  4417 => x"800c853d",
  4418 => x"0d047352",
  4419 => x"755180e7",
  4420 => x"a73f800b",
  4421 => x"88150c80",
  4422 => x"0b84150c",
  4423 => x"8008800c",
  4424 => x"853d0d04",
  4425 => x"fcc43d0d",
  4426 => x"83bf3d08",
  4427 => x"83c13d08",
  4428 => x"83c33d08",
  4429 => x"83c53d08",
  4430 => x"485e484b",
  4431 => x"80ef843f",
  4432 => x"8008084c",
  4433 => x"800b83bb",
  4434 => x"3d0c800b",
  4435 => x"83bc3d0c",
  4436 => x"80707169",
  4437 => x"8c052270",
  4438 => x"832a8132",
  4439 => x"70810651",
  4440 => x"5d5d4c4f",
  4441 => x"4d786d2e",
  4442 => x"0981068c",
  4443 => x"38669005",
  4444 => x"086d2e09",
  4445 => x"81069238",
  4446 => x"6651b49e",
  4447 => x"3fff5980",
  4448 => x"0881e438",
  4449 => x"668c0522",
  4450 => x"5a799a06",
  4451 => x"59788a2e",
  4452 => x"80c0387b",
  4453 => x"83a63d70",
  4454 => x"7183b93d",
  4455 => x"0c5e475d",
  4456 => x"800b83b8",
  4457 => x"3d0c800b",
  4458 => x"83b73d0c",
  4459 => x"80497c5e",
  4460 => x"807d3370",
  4461 => x"81ff065b",
  4462 => x"5b5b787b",
  4463 => x"2e833881",
  4464 => x"5b78a52e",
  4465 => x"81a9387a",
  4466 => x"802e81a3",
  4467 => x"38811d5d",
  4468 => x"df39668e",
  4469 => x"05227090",
  4470 => x"2b5a5b80",
  4471 => x"7924ffb3",
  4472 => x"3879fd06",
  4473 => x"597882ba",
  4474 => x"3d237a02",
  4475 => x"840589e2",
  4476 => x"0523669c",
  4477 => x"050882be",
  4478 => x"3d0c66a4",
  4479 => x"050882c0",
  4480 => x"3d0cb63d",
  4481 => x"7082b83d",
  4482 => x"0c82bb3d",
  4483 => x"0c88800b",
  4484 => x"82b93d0c",
  4485 => x"88800b82",
  4486 => x"bc3d0c80",
  4487 => x"0b82bd3d",
  4488 => x"0c64537b",
  4489 => x"5282b63d",
  4490 => x"705259a8",
  4491 => x"a33f8008",
  4492 => x"5a800b80",
  4493 => x"08248f38",
  4494 => x"785180d9",
  4495 => x"cf3f8008",
  4496 => x"802e8338",
  4497 => x"ff5a82b9",
  4498 => x"3d227086",
  4499 => x"2a708106",
  4500 => x"515a5b78",
  4501 => x"802e8e38",
  4502 => x"668c0522",
  4503 => x"80c00759",
  4504 => x"78678c05",
  4505 => x"23795978",
  4506 => x"800c83be",
  4507 => x"3d0d047c",
  4508 => x"7e315b7a",
  4509 => x"802eae38",
  4510 => x"7d7c0c7a",
  4511 => x"841d0c83",
  4512 => x"b73d081b",
  4513 => x"83b83d0c",
  4514 => x"881c83b7",
  4515 => x"3d088111",
  4516 => x"83b93d0c",
  4517 => x"8111515a",
  4518 => x"5c788724",
  4519 => x"80c33868",
  4520 => x"1b7d335b",
  4521 => x"497981ff",
  4522 => x"06597880",
  4523 => x"2ea69638",
  4524 => x"811d5d80",
  4525 => x"70714a45",
  4526 => x"43ff4162",
  4527 => x"83be3d34",
  4528 => x"7c335a79",
  4529 => x"81ff0681",
  4530 => x"1e5e407f",
  4531 => x"e0055978",
  4532 => x"80d82686",
  4533 => x"ec387810",
  4534 => x"1082c48c",
  4535 => x"05597808",
  4536 => x"0483be3d",
  4537 => x"dc055266",
  4538 => x"51fc883f",
  4539 => x"80088997",
  4540 => x"3865691c",
  4541 => x"7e335c4a",
  4542 => x"5cffaa39",
  4543 => x"62900743",
  4544 => x"62842a70",
  4545 => x"81065159",
  4546 => x"7898ba38",
  4547 => x"62862a70",
  4548 => x"81065159",
  4549 => x"78802e98",
  4550 => x"ac386465",
  4551 => x"84058212",
  4552 => x"225d4659",
  4553 => x"815f800b",
  4554 => x"83be3d34",
  4555 => x"60448061",
  4556 => x"24863862",
  4557 => x"feff0643",
  4558 => x"657b3070",
  4559 => x"7d079f2a",
  4560 => x"66307068",
  4561 => x"079f2a72",
  4562 => x"07525c51",
  4563 => x"5b5e7980",
  4564 => x"2e948938",
  4565 => x"7e812e89",
  4566 => x"d338817f",
  4567 => x"259ad438",
  4568 => x"7e822e8a",
  4569 => x"863882c6",
  4570 => x"f05e7d51",
  4571 => x"81929c3f",
  4572 => x"80085f7e",
  4573 => x"427e6425",
  4574 => x"83386342",
  4575 => x"83bd3d33",
  4576 => x"7081ff06",
  4577 => x"5a5b7880",
  4578 => x"2e908d38",
  4579 => x"61810542",
  4580 => x"62818406",
  4581 => x"416080f1",
  4582 => x"38676231",
  4583 => x"5a807a25",
  4584 => x"80e73890",
  4585 => x"7a25b438",
  4586 => x"82c3ec7c",
  4587 => x"0c900b84",
  4588 => x"1d0c83b7",
  4589 => x"3d089005",
  4590 => x"83b83d0c",
  4591 => x"881c83b7",
  4592 => x"3d088111",
  4593 => x"83b93d0c",
  4594 => x"8111515a",
  4595 => x"5c788724",
  4596 => x"858738f0",
  4597 => x"1a5a7990",
  4598 => x"24ce3882",
  4599 => x"c3ec7c0c",
  4600 => x"79841d0c",
  4601 => x"83b73d08",
  4602 => x"1a83b83d",
  4603 => x"0c881c83",
  4604 => x"b73d0881",
  4605 => x"1183b93d",
  4606 => x"0c811151",
  4607 => x"5a5c7887",
  4608 => x"2492bf38",
  4609 => x"83bd3d33",
  4610 => x"5b7a81ff",
  4611 => x"06597880",
  4612 => x"2e8f9b38",
  4613 => x"83be3dfc",
  4614 => x"057c0c81",
  4615 => x"0b841d0c",
  4616 => x"83b73d08",
  4617 => x"810583b8",
  4618 => x"3d0c881c",
  4619 => x"83b73d08",
  4620 => x"811183b9",
  4621 => x"3d0c8111",
  4622 => x"515a5c78",
  4623 => x"872485eb",
  4624 => x"38608180",
  4625 => x"2e84c238",
  4626 => x"637f315a",
  4627 => x"807a2580",
  4628 => x"f338907a",
  4629 => x"25b43882",
  4630 => x"c3fc7c0c",
  4631 => x"900b841d",
  4632 => x"0c83b73d",
  4633 => x"08900583",
  4634 => x"b83d0c88",
  4635 => x"1c83b73d",
  4636 => x"08811183",
  4637 => x"b93d0c81",
  4638 => x"11515a5c",
  4639 => x"78872483",
  4640 => x"f038f01a",
  4641 => x"5a799024",
  4642 => x"ce3882c3",
  4643 => x"fc7c0c79",
  4644 => x"841d0c83",
  4645 => x"b73d081a",
  4646 => x"83b83d0c",
  4647 => x"881c83b7",
  4648 => x"3d088111",
  4649 => x"83b93d0c",
  4650 => x"8111515a",
  4651 => x"5c877925",
  4652 => x"933883be",
  4653 => x"3ddc0552",
  4654 => x"6651f8b7",
  4655 => x"3f800885",
  4656 => x"c638655c",
  4657 => x"62882a81",
  4658 => x"32708106",
  4659 => x"51597880",
  4660 => x"2e8ea938",
  4661 => x"7d7c0c7e",
  4662 => x"841d0c83",
  4663 => x"b73d081f",
  4664 => x"83b83d0c",
  4665 => x"881c83b7",
  4666 => x"3d088111",
  4667 => x"83b93d0c",
  4668 => x"8111515a",
  4669 => x"5c788724",
  4670 => x"84e73862",
  4671 => x"822a7081",
  4672 => x"06515978",
  4673 => x"802e80f8",
  4674 => x"38676231",
  4675 => x"5a807a25",
  4676 => x"80ee3890",
  4677 => x"7a25b438",
  4678 => x"82c3ec7c",
  4679 => x"0c900b84",
  4680 => x"1d0c83b7",
  4681 => x"3d089005",
  4682 => x"83b83d0c",
  4683 => x"881c83b7",
  4684 => x"3d088111",
  4685 => x"83b93d0c",
  4686 => x"8111515a",
  4687 => x"5c788724",
  4688 => x"848838f0",
  4689 => x"1a5a7990",
  4690 => x"24ce3882",
  4691 => x"c3ec7c0c",
  4692 => x"79841d0c",
  4693 => x"83b73d08",
  4694 => x"1a83b83d",
  4695 => x"0c83b63d",
  4696 => x"08811183",
  4697 => x"b83d0c81",
  4698 => x"11515987",
  4699 => x"79259138",
  4700 => x"83be3ddc",
  4701 => x"05526651",
  4702 => x"f6f93f80",
  4703 => x"08848838",
  4704 => x"61596168",
  4705 => x"25833867",
  4706 => x"59681949",
  4707 => x"83b73d08",
  4708 => x"83e33880",
  4709 => x"0b83b73d",
  4710 => x"0c655c69",
  4711 => x"802ef88e",
  4712 => x"386951e8",
  4713 => x"bf3f807d",
  4714 => x"5f4af884",
  4715 => x"39629007",
  4716 => x"4362842a",
  4717 => x"70810651",
  4718 => x"59789397",
  4719 => x"3862862a",
  4720 => x"70810651",
  4721 => x"5978802e",
  4722 => x"93893864",
  4723 => x"65840582",
  4724 => x"12225d46",
  4725 => x"59805f80",
  4726 => x"0b83be3d",
  4727 => x"34facd39",
  4728 => x"62900743",
  4729 => x"62842a70",
  4730 => x"81065159",
  4731 => x"7892f238",
  4732 => x"62862a70",
  4733 => x"81065159",
  4734 => x"78802e92",
  4735 => x"e4386465",
  4736 => x"84057108",
  4737 => x"902b7090",
  4738 => x"2c515d46",
  4739 => x"59807b24",
  4740 => x"89a43881",
  4741 => x"5ffa9539",
  4742 => x"64658405",
  4743 => x"71084a46",
  4744 => x"59678025",
  4745 => x"f99a3867",
  4746 => x"30486284",
  4747 => x"077d335b",
  4748 => x"43f99039",
  4749 => x"811d5d62",
  4750 => x"90077d33",
  4751 => x"5b43f983",
  4752 => x"397f802e",
  4753 => x"9eff3882",
  4754 => x"ce3d5e7f",
  4755 => x"7e34815f",
  4756 => x"800b83be",
  4757 => x"3d34fa9b",
  4758 => x"3983be3d",
  4759 => x"dc055266",
  4760 => x"51f5903f",
  4761 => x"8008829f",
  4762 => x"3865f01b",
  4763 => x"5b5cfae6",
  4764 => x"3983be3d",
  4765 => x"dc055266",
  4766 => x"51f4f83f",
  4767 => x"80088287",
  4768 => x"3865f01b",
  4769 => x"5b5cfbfd",
  4770 => x"39676231",
  4771 => x"5a807a25",
  4772 => x"fbb63890",
  4773 => x"7a25b438",
  4774 => x"82c3fc7c",
  4775 => x"0c900b84",
  4776 => x"1d0c83b7",
  4777 => x"3d089005",
  4778 => x"83b83d0c",
  4779 => x"881c83b7",
  4780 => x"3d088111",
  4781 => x"83b93d0c",
  4782 => x"8111515a",
  4783 => x"5c788724",
  4784 => x"80d138f0",
  4785 => x"1a5a7990",
  4786 => x"24ce3882",
  4787 => x"c3fc7c0c",
  4788 => x"79841d0c",
  4789 => x"83b73d08",
  4790 => x"1a83b83d",
  4791 => x"0c881c83",
  4792 => x"b73d0881",
  4793 => x"1183b93d",
  4794 => x"0c811151",
  4795 => x"5a5c8779",
  4796 => x"25fad538",
  4797 => x"83be3ddc",
  4798 => x"05526651",
  4799 => x"f3f53f80",
  4800 => x"08818438",
  4801 => x"65646031",
  4802 => x"5b5c7980",
  4803 => x"24fac338",
  4804 => x"fbb23983",
  4805 => x"be3ddc05",
  4806 => x"526651f3",
  4807 => x"d63f8008",
  4808 => x"80e53865",
  4809 => x"f01b5b5c",
  4810 => x"ff9c3983",
  4811 => x"be3ddc05",
  4812 => x"526651f3",
  4813 => x"be3f8008",
  4814 => x"80cd3865",
  4815 => x"5c608180",
  4816 => x"2e098106",
  4817 => x"fa8238fe",
  4818 => x"c03983be",
  4819 => x"3ddc0552",
  4820 => x"6651f39f",
  4821 => x"3f8008af",
  4822 => x"3865f01b",
  4823 => x"5b5cfbe6",
  4824 => x"3983be3d",
  4825 => x"dc055266",
  4826 => x"51f3883f",
  4827 => x"80089838",
  4828 => x"655cfb87",
  4829 => x"3983be3d",
  4830 => x"dc055266",
  4831 => x"51f2f43f",
  4832 => x"8008802e",
  4833 => x"fc8d3869",
  4834 => x"802e8638",
  4835 => x"6951e4d4",
  4836 => x"3f668c05",
  4837 => x"2270862a",
  4838 => x"7081066b",
  4839 => x"5d515a47",
  4840 => x"78802ef5",
  4841 => x"c038ff59",
  4842 => x"f5bd397c",
  4843 => x"337081ff",
  4844 => x"065a5a78",
  4845 => x"80ec2efc",
  4846 => x"fb386290",
  4847 => x"077a81ff",
  4848 => x"06811f5f",
  4849 => x"4143f683",
  4850 => x"397c7081",
  4851 => x"055e3340",
  4852 => x"7faa2e9c",
  4853 => x"ce388060",
  4854 => x"d0057143",
  4855 => x"5a5a7889",
  4856 => x"26f5e838",
  4857 => x"79101010",
  4858 => x"7a100560",
  4859 => x"05d0057d",
  4860 => x"7081055f",
  4861 => x"33d0115b",
  4862 => x"415a8979",
  4863 => x"27e63879",
  4864 => x"4179ff25",
  4865 => x"f5c538ff",
  4866 => x"41f5c039",
  4867 => x"64658405",
  4868 => x"71085d46",
  4869 => x"59820b82",
  4870 => x"c78c6472",
  4871 => x"07454f5f",
  4872 => x"80f84080",
  4873 => x"0b83be3d",
  4874 => x"34f68139",
  4875 => x"897b27a4",
  4876 => x"38ff1e5e",
  4877 => x"8a527a51",
  4878 => x"81a1dd3f",
  4879 => x"8008b005",
  4880 => x"59787e34",
  4881 => x"8a527a51",
  4882 => x"81a1a73f",
  4883 => x"80085b7a",
  4884 => x"8926de38",
  4885 => x"ff1eb01c",
  4886 => x"5a5e787e",
  4887 => x"3483be3d",
  4888 => x"707f31ff",
  4889 => x"9c05405b",
  4890 => x"f68939ff",
  4891 => x"1e7b8f06",
  4892 => x"6f055a5e",
  4893 => x"78337e34",
  4894 => x"7a842a5b",
  4895 => x"7a802edd",
  4896 => x"38ff1e7b",
  4897 => x"8f066f05",
  4898 => x"5a5e7833",
  4899 => x"7e347a84",
  4900 => x"2a5b7ad7",
  4901 => x"38c73962",
  4902 => x"80c0077d",
  4903 => x"335b43f4",
  4904 => x"a23960ff",
  4905 => x"2e99e238",
  4906 => x"7f80e732",
  4907 => x"70307072",
  4908 => x"07802562",
  4909 => x"80c73270",
  4910 => x"30707207",
  4911 => x"80257307",
  4912 => x"53545e51",
  4913 => x"5b597980",
  4914 => x"2e863860",
  4915 => x"83388141",
  4916 => x"64658805",
  4917 => x"84120872",
  4918 => x"087083bf",
  4919 => x"3d0c7183",
  4920 => x"c03d0c54",
  4921 => x"54465981",
  4922 => x"82ff3f80",
  4923 => x"08802e91",
  4924 => x"ea388059",
  4925 => x"80795454",
  4926 => x"83ba3d08",
  4927 => x"83bc3d08",
  4928 => x"5b517952",
  4929 => x"8198963f",
  4930 => x"800b8008",
  4931 => x"2484d738",
  4932 => x"82c7a05e",
  4933 => x"835ff4db",
  4934 => x"3982ce3d",
  4935 => x"5e7f80c3",
  4936 => x"2e8f3862",
  4937 => x"842a7081",
  4938 => x"06515978",
  4939 => x"802e82f6",
  4940 => x"38885380",
  4941 => x"52b43d70",
  4942 => x"525980e3",
  4943 => x"fb3f7854",
  4944 => x"64658405",
  4945 => x"7108557f",
  4946 => x"546c5346",
  4947 => x"599ab93f",
  4948 => x"80085f80",
  4949 => x"08ff2efc",
  4950 => x"ae38800b",
  4951 => x"83be3d34",
  4952 => x"f4913982",
  4953 => x"c7a46384",
  4954 => x"2a708106",
  4955 => x"515a4e78",
  4956 => x"82893862",
  4957 => x"862a7081",
  4958 => x"06515978",
  4959 => x"802e81fb",
  4960 => x"38646584",
  4961 => x"05821222",
  4962 => x"5d465982",
  4963 => x"6381065a",
  4964 => x"5f7a802e",
  4965 => x"f3903878",
  4966 => x"802ef38a",
  4967 => x"38627f07",
  4968 => x"43800b83",
  4969 => x"be3d34f3",
  4970 => x"8339800b",
  4971 => x"83be3d34",
  4972 => x"64658405",
  4973 => x"71084046",
  4974 => x"597d802e",
  4975 => x"97d0387f",
  4976 => x"80d32e81",
  4977 => x"ff386284",
  4978 => x"2a708106",
  4979 => x"51597881",
  4980 => x"f3388061",
  4981 => x"24f39338",
  4982 => x"60537852",
  4983 => x"7d5180df",
  4984 => x"f53f605f",
  4985 => x"8008802e",
  4986 => x"f3893880",
  4987 => x"087e315f",
  4988 => x"607f25f2",
  4989 => x"fe38605f",
  4990 => x"f2f93962",
  4991 => x"842a7081",
  4992 => x"06515978",
  4993 => x"8d9c3862",
  4994 => x"862a7081",
  4995 => x"06515978",
  4996 => x"802e8d8e",
  4997 => x"38646584",
  4998 => x"05710852",
  4999 => x"46596879",
  5000 => x"237c5eef",
  5001 => x"8b39ab0b",
  5002 => x"83be3d34",
  5003 => x"7c335af1",
  5004 => x"9239805a",
  5005 => x"79101010",
  5006 => x"7a100560",
  5007 => x"05d0057d",
  5008 => x"7081055f",
  5009 => x"33d0115b",
  5010 => x"415a8979",
  5011 => x"27e63879",
  5012 => x"48f0f839",
  5013 => x"62818007",
  5014 => x"7d335b43",
  5015 => x"f0e53962",
  5016 => x"88077d33",
  5017 => x"5b43f0db",
  5018 => x"3982c78c",
  5019 => x"63842a70",
  5020 => x"8106515a",
  5021 => x"4e78802e",
  5022 => x"fdf93864",
  5023 => x"65840571",
  5024 => x"085d4659",
  5025 => x"fe853962",
  5026 => x"81077d33",
  5027 => x"5b43f0b3",
  5028 => x"3983bd3d",
  5029 => x"335978f0",
  5030 => x"a738a00b",
  5031 => x"83be3d34",
  5032 => x"7c335af0",
  5033 => x"9e396465",
  5034 => x"84054659",
  5035 => x"8319337e",
  5036 => x"34815ff7",
  5037 => x"9b397a30",
  5038 => x"5bad0b83",
  5039 => x"be3d3481",
  5040 => x"5ff0e939",
  5041 => x"7da23d0c",
  5042 => x"80705c5f",
  5043 => x"88537e52",
  5044 => x"a63d7052",
  5045 => x"5a80e0e0",
  5046 => x"3f7e6124",
  5047 => x"8197387a",
  5048 => x"1010a23d",
  5049 => x"08055978",
  5050 => x"08802eaf",
  5051 => x"38795478",
  5052 => x"085383be",
  5053 => x"3dfcc005",
  5054 => x"526a5197",
  5055 => x"8b3f8008",
  5056 => x"ff2ef983",
  5057 => x"3880081f",
  5058 => x"59786124",
  5059 => x"8e38811b",
  5060 => x"79405b78",
  5061 => x"612e0981",
  5062 => x"06c5387e",
  5063 => x"802ef0d3",
  5064 => x"38811f52",
  5065 => x"6a51ddce",
  5066 => x"3f80084a",
  5067 => x"8008802e",
  5068 => x"f8df3888",
  5069 => x"53805279",
  5070 => x"5180dffc",
  5071 => x"3f79557e",
  5072 => x"5483be3d",
  5073 => x"f38c0553",
  5074 => x"69526a51",
  5075 => x"97a23f80",
  5076 => x"087f2e09",
  5077 => x"8106f8af",
  5078 => x"38696a80",
  5079 => x"08055a5e",
  5080 => x"807934f0",
  5081 => x"8e39ad0b",
  5082 => x"83be3d34",
  5083 => x"82c7a05e",
  5084 => x"835fefff",
  5085 => x"3979557e",
  5086 => x"5483be3d",
  5087 => x"f38c0553",
  5088 => x"7e526a51",
  5089 => x"96ea3f80",
  5090 => x"085f8008",
  5091 => x"ff2ef7f7",
  5092 => x"387da23d",
  5093 => x"0cff8439",
  5094 => x"620a100a",
  5095 => x"70810651",
  5096 => x"5978802e",
  5097 => x"efea3861",
  5098 => x"820542ef",
  5099 => x"e339620a",
  5100 => x"100a7081",
  5101 => x"06515978",
  5102 => x"802ef185",
  5103 => x"38b00b82",
  5104 => x"ce3d347f",
  5105 => x"0284058a",
  5106 => x"b1053483",
  5107 => x"be3dfcbc",
  5108 => x"057c0c82",
  5109 => x"0b841d0c",
  5110 => x"83b73d08",
  5111 => x"820583b8",
  5112 => x"3d0c881c",
  5113 => x"83b73d08",
  5114 => x"811183b9",
  5115 => x"3d0c8111",
  5116 => x"515a5c87",
  5117 => x"7925f0c9",
  5118 => x"38f6b039",
  5119 => x"80e56025",
  5120 => x"82fe3880",
  5121 => x"59807954",
  5122 => x"5483ba3d",
  5123 => x"0883bc3d",
  5124 => x"085b5179",
  5125 => x"52818cc1",
  5126 => x"3f800886",
  5127 => x"d63882c7",
  5128 => x"b87c0c81",
  5129 => x"0b841d0c",
  5130 => x"83b73d08",
  5131 => x"810583b8",
  5132 => x"3d0c881c",
  5133 => x"83b73d08",
  5134 => x"811183b9",
  5135 => x"3d0c8111",
  5136 => x"515a5c78",
  5137 => x"872481ac",
  5138 => x"38a43d08",
  5139 => x"5b7aa63d",
  5140 => x"08248b38",
  5141 => x"62810659",
  5142 => x"78802ef1",
  5143 => x"9e386b7c",
  5144 => x"0c810b84",
  5145 => x"1d0c83b7",
  5146 => x"3d088105",
  5147 => x"83b83d0c",
  5148 => x"881c83b7",
  5149 => x"3d088111",
  5150 => x"83b93d0c",
  5151 => x"8111515a",
  5152 => x"5c788724",
  5153 => x"819b38ff",
  5154 => x"1b5a807a",
  5155 => x"25f0ec38",
  5156 => x"907a25b4",
  5157 => x"3882c3fc",
  5158 => x"7c0c900b",
  5159 => x"841d0c83",
  5160 => x"b73d0890",
  5161 => x"0583b83d",
  5162 => x"0c881c83",
  5163 => x"b73d0881",
  5164 => x"1183b93d",
  5165 => x"0c811151",
  5166 => x"5a5c7887",
  5167 => x"2480ca38",
  5168 => x"f01a5a79",
  5169 => x"9024ce38",
  5170 => x"82c3fc7c",
  5171 => x"0c79841d",
  5172 => x"0c83b73d",
  5173 => x"081a83b8",
  5174 => x"3d0c881c",
  5175 => x"83b73d08",
  5176 => x"811183b9",
  5177 => x"3d0c8111",
  5178 => x"515a5c87",
  5179 => x"7925f08b",
  5180 => x"38f4ee39",
  5181 => x"83be3ddc",
  5182 => x"05526651",
  5183 => x"e7f53f80",
  5184 => x"08f58438",
  5185 => x"655cfec1",
  5186 => x"3983be3d",
  5187 => x"dc055266",
  5188 => x"51e7e03f",
  5189 => x"8008f4ef",
  5190 => x"3865f01b",
  5191 => x"5b5cffa3",
  5192 => x"3983be3d",
  5193 => x"dc055266",
  5194 => x"51e7c83f",
  5195 => x"8008f4d7",
  5196 => x"3865a53d",
  5197 => x"08ff055b",
  5198 => x"5c798024",
  5199 => x"fed238ef",
  5200 => x"ba3983be",
  5201 => x"3ddc0552",
  5202 => x"6651e7a7",
  5203 => x"3f8008f4",
  5204 => x"b6386583",
  5205 => x"be3d335c",
  5206 => x"5cedae39",
  5207 => x"7ef5fe38",
  5208 => x"62810659",
  5209 => x"78802ef5",
  5210 => x"f438028d",
  5211 => x"8f055eb0",
  5212 => x"7e3483be",
  5213 => x"3d707f31",
  5214 => x"ff9c0540",
  5215 => x"5bebf439",
  5216 => x"a43d085b",
  5217 => x"817b2583",
  5218 => x"82387d70",
  5219 => x"81055f33",
  5220 => x"82ce3d34",
  5221 => x"ae028405",
  5222 => x"8ab10534",
  5223 => x"83be3dfc",
  5224 => x"bc057c0c",
  5225 => x"820b841d",
  5226 => x"0c83b73d",
  5227 => x"08820583",
  5228 => x"b83d0c88",
  5229 => x"1c83b73d",
  5230 => x"08811183",
  5231 => x"b93d0c81",
  5232 => x"11515a5c",
  5233 => x"78872480",
  5234 => x"fd388059",
  5235 => x"80795454",
  5236 => x"83ba3d08",
  5237 => x"83bc3d08",
  5238 => x"5b517952",
  5239 => x"818ae63f",
  5240 => x"8008802e",
  5241 => x"8191387d",
  5242 => x"7c0cff1b",
  5243 => x"841d0c83",
  5244 => x"b73d081b",
  5245 => x"ff0583b8",
  5246 => x"3d0c881c",
  5247 => x"83b73d08",
  5248 => x"811183b9",
  5249 => x"3d0c8111",
  5250 => x"515a5c78",
  5251 => x"872481d1",
  5252 => x"3883be3d",
  5253 => x"e8057c0c",
  5254 => x"6c841d0c",
  5255 => x"83b73d08",
  5256 => x"6d0583b8",
  5257 => x"3d0c881c",
  5258 => x"83b73d08",
  5259 => x"811183b9",
  5260 => x"3d0c8111",
  5261 => x"515a5c87",
  5262 => x"7925edbf",
  5263 => x"3883be3d",
  5264 => x"dc0552f2",
  5265 => x"a23983be",
  5266 => x"3ddc0552",
  5267 => x"6651e5a3",
  5268 => x"3f8008f2",
  5269 => x"b23865a5",
  5270 => x"3d085c5c",
  5271 => x"80598079",
  5272 => x"545483ba",
  5273 => x"3d0883bc",
  5274 => x"3d085b51",
  5275 => x"79528189",
  5276 => x"d43f8008",
  5277 => x"fef138ff",
  5278 => x"1b5a807a",
  5279 => x"25ff9238",
  5280 => x"907a25b4",
  5281 => x"3882c3fc",
  5282 => x"7c0c900b",
  5283 => x"841d0c83",
  5284 => x"b73d0890",
  5285 => x"0583b83d",
  5286 => x"0c881c83",
  5287 => x"b73d0881",
  5288 => x"1183b93d",
  5289 => x"0c811151",
  5290 => x"5a5c7887",
  5291 => x"2483db38",
  5292 => x"f01a5a79",
  5293 => x"9024ce38",
  5294 => x"82c3fc7c",
  5295 => x"0c79841d",
  5296 => x"0c83b73d",
  5297 => x"081a83b8",
  5298 => x"3d0c881c",
  5299 => x"83b73d08",
  5300 => x"811183b9",
  5301 => x"3d0c8111",
  5302 => x"515a5c87",
  5303 => x"7925feb1",
  5304 => x"3883be3d",
  5305 => x"dc055266",
  5306 => x"51e4883f",
  5307 => x"8008f197",
  5308 => x"386583bf",
  5309 => x"3de80571",
  5310 => x"0c6d8412",
  5311 => x"0c83b83d",
  5312 => x"086e0583",
  5313 => x"b93d0c5c",
  5314 => x"fe9c3962",
  5315 => x"81065978",
  5316 => x"fcf8387d",
  5317 => x"7c0c810b",
  5318 => x"841d0c83",
  5319 => x"b73d0881",
  5320 => x"0583b83d",
  5321 => x"0c881c83",
  5322 => x"b73d0881",
  5323 => x"1183b93d",
  5324 => x"0c811151",
  5325 => x"5a5c8779",
  5326 => x"25fdd638",
  5327 => x"83be3ddc",
  5328 => x"0552ffa3",
  5329 => x"39646584",
  5330 => x"0571085d",
  5331 => x"4659815f",
  5332 => x"e7d43964",
  5333 => x"65840571",
  5334 => x"085d4659",
  5335 => x"805fecf7",
  5336 => x"39646584",
  5337 => x"0571085d",
  5338 => x"46597a80",
  5339 => x"25eda438",
  5340 => x"f6c439a5",
  5341 => x"3d085a80",
  5342 => x"7a2589c8",
  5343 => x"38a43d08",
  5344 => x"5b7a7a24",
  5345 => x"82dd387d",
  5346 => x"7c0c7a84",
  5347 => x"1d0c83b7",
  5348 => x"3d081b83",
  5349 => x"b83d0c88",
  5350 => x"1c83b73d",
  5351 => x"08811183",
  5352 => x"b93d0c81",
  5353 => x"11515a5c",
  5354 => x"78872481",
  5355 => x"b638797b",
  5356 => x"315a807a",
  5357 => x"2580f338",
  5358 => x"907a25b4",
  5359 => x"3882c3fc",
  5360 => x"7c0c900b",
  5361 => x"841d0c83",
  5362 => x"b73d0890",
  5363 => x"0583b83d",
  5364 => x"0c881c83",
  5365 => x"b73d0881",
  5366 => x"1183b93d",
  5367 => x"0c811151",
  5368 => x"5a5c7887",
  5369 => x"2480e438",
  5370 => x"f01a5a79",
  5371 => x"9024ce38",
  5372 => x"82c3fc7c",
  5373 => x"0c79841d",
  5374 => x"0c83b73d",
  5375 => x"081a83b8",
  5376 => x"3d0c881c",
  5377 => x"83b73d08",
  5378 => x"811183b9",
  5379 => x"3d0c8111",
  5380 => x"515a5c87",
  5381 => x"79259338",
  5382 => x"83be3ddc",
  5383 => x"05526651",
  5384 => x"e1d13f80",
  5385 => x"08eee038",
  5386 => x"655c6281",
  5387 => x"06597880",
  5388 => x"2ee9c838",
  5389 => x"82c7bc7c",
  5390 => x"0c810b84",
  5391 => x"1d0c83b7",
  5392 => x"3d088105",
  5393 => x"83b83d0c",
  5394 => x"fbdc3983",
  5395 => x"be3ddc05",
  5396 => x"526651e1",
  5397 => x"9e3f8008",
  5398 => x"eead3865",
  5399 => x"f01b5b5c",
  5400 => x"ff893983",
  5401 => x"be3ddc05",
  5402 => x"526651e1",
  5403 => x"863f8008",
  5404 => x"ee953865",
  5405 => x"a63d08a6",
  5406 => x"3d087171",
  5407 => x"31525d5b",
  5408 => x"5c798024",
  5409 => x"feb238ff",
  5410 => x"a13983be",
  5411 => x"3ddc0552",
  5412 => x"6651e0df",
  5413 => x"3f8008ed",
  5414 => x"ee3865f0",
  5415 => x"1b5b5cfc",
  5416 => x"92396465",
  5417 => x"84057108",
  5418 => x"6b710c52",
  5419 => x"7e404659",
  5420 => x"e1fe397e",
  5421 => x"e5b038ff",
  5422 => x"1e7bb706",
  5423 => x"b0075b5e",
  5424 => x"797e347a",
  5425 => x"832a5b7a",
  5426 => x"ee386281",
  5427 => x"06597880",
  5428 => x"2eef8a38",
  5429 => x"79b02eef",
  5430 => x"8438ff1e",
  5431 => x"5eb07e34",
  5432 => x"f990397d",
  5433 => x"7c0c7984",
  5434 => x"1d0c83b7",
  5435 => x"3d081a83",
  5436 => x"b83d0c88",
  5437 => x"1c83b73d",
  5438 => x"08811183",
  5439 => x"b93d0c81",
  5440 => x"11515a5c",
  5441 => x"78872481",
  5442 => x"8b38791e",
  5443 => x"82c7bc7d",
  5444 => x"0c5e810b",
  5445 => x"841d0c83",
  5446 => x"b73d0881",
  5447 => x"0583b83d",
  5448 => x"0c881c83",
  5449 => x"b73d0881",
  5450 => x"1183b93d",
  5451 => x"0c811151",
  5452 => x"5a5c7887",
  5453 => x"24b0387d",
  5454 => x"7c0ca43d",
  5455 => x"087a3170",
  5456 => x"841e0c83",
  5457 => x"b83d0805",
  5458 => x"83b83d0c",
  5459 => x"881c83b7",
  5460 => x"3d088111",
  5461 => x"83b93d0c",
  5462 => x"8111515a",
  5463 => x"5c877925",
  5464 => x"e79938eb",
  5465 => x"fc3983be",
  5466 => x"3ddc0552",
  5467 => x"6651df83",
  5468 => x"3f8008ec",
  5469 => x"923865a6",
  5470 => x"3d087f72",
  5471 => x"0ca63d08",
  5472 => x"71317084",
  5473 => x"140c83ba",
  5474 => x"3d080583",
  5475 => x"ba3d0c5b",
  5476 => x"5cffb939",
  5477 => x"83be3ddc",
  5478 => x"05526651",
  5479 => x"ded53f80",
  5480 => x"08ebe438",
  5481 => x"65a63d08",
  5482 => x"7f1182c7",
  5483 => x"bc730c40",
  5484 => x"5b5c810b",
  5485 => x"841d0c83",
  5486 => x"b73d0881",
  5487 => x"0583b83d",
  5488 => x"0c881c83",
  5489 => x"b73d0881",
  5490 => x"1183b93d",
  5491 => x"0c811151",
  5492 => x"5a5c8779",
  5493 => x"25fee038",
  5494 => x"ff8c3983",
  5495 => x"ba3d0883",
  5496 => x"bc3d085b",
  5497 => x"51795280",
  5498 => x"f1b03f82",
  5499 => x"c7c05e83",
  5500 => x"5f8008e2",
  5501 => x"fe386282",
  5502 => x"800783bb",
  5503 => x"3d0883bd",
  5504 => x"3d086383",
  5505 => x"c03daa3d",
  5506 => x"a53d0c5f",
  5507 => x"45415f43",
  5508 => x"830ba13d",
  5509 => x"0c7f80e6",
  5510 => x"2ea73880",
  5511 => x"085a7f80",
  5512 => x"e52e83a9",
  5513 => x"38800859",
  5514 => x"7f80c52e",
  5515 => x"83af3879",
  5516 => x"79075978",
  5517 => x"802e8538",
  5518 => x"60810542",
  5519 => x"820ba13d",
  5520 => x"0c7db33d",
  5521 => x"0c7eb43d",
  5522 => x"0c800bb3",
  5523 => x"3d082487",
  5524 => x"9c38807b",
  5525 => x"3483be3d",
  5526 => x"f3941159",
  5527 => x"f3900557",
  5528 => x"6e566155",
  5529 => x"6f547d52",
  5530 => x"7e536a51",
  5531 => x"96d13f80",
  5532 => x"086080e7",
  5533 => x"32703070",
  5534 => x"72079f2a",
  5535 => x"515b5ba1",
  5536 => x"3d0c7f80",
  5537 => x"c72e8538",
  5538 => x"7881d038",
  5539 => x"62810659",
  5540 => x"7881c838",
  5541 => x"a33d0859",
  5542 => x"78a13d08",
  5543 => x"31a53d0c",
  5544 => x"6f6080e7",
  5545 => x"32703070",
  5546 => x"72078025",
  5547 => x"6380c732",
  5548 => x"70307072",
  5549 => x"07802573",
  5550 => x"0753545f",
  5551 => x"515c5a5e",
  5552 => x"79802e85",
  5553 => x"d238a53d",
  5554 => x"085afc7a",
  5555 => x"25873860",
  5556 => x"7a25829f",
  5557 => x"3880e559",
  5558 => x"7f80e72e",
  5559 => x"843880c5",
  5560 => x"5978407f",
  5561 => x"80e52485",
  5562 => x"b538ff1a",
  5563 => x"70a73d0c",
  5564 => x"83b93d71",
  5565 => x"5d435a7f",
  5566 => x"6234028d",
  5567 => x"dd055f80",
  5568 => x"7a248686",
  5569 => x"38ab7f34",
  5570 => x"028dde05",
  5571 => x"b33d705c",
  5572 => x"425f897b",
  5573 => x"2580fd38",
  5574 => x"ff1a5a8a",
  5575 => x"527a51ff",
  5576 => x"afd63f80",
  5577 => x"08b00559",
  5578 => x"787a348a",
  5579 => x"527a51ff",
  5580 => x"ae943f80",
  5581 => x"085b8008",
  5582 => x"8924dd38",
  5583 => x"ff1a8008",
  5584 => x"b0055a5a",
  5585 => x"787a3479",
  5586 => x"612780d9",
  5587 => x"38797081",
  5588 => x"055b337f",
  5589 => x"70810541",
  5590 => x"34ed3980",
  5591 => x"0862055b",
  5592 => x"7f80e62e",
  5593 => x"80fc3880",
  5594 => x"59807954",
  5595 => x"547d517e",
  5596 => x"5280fde5",
  5597 => x"3f800885",
  5598 => x"387aa43d",
  5599 => x"0ca33d08",
  5600 => x"59787b27",
  5601 => x"fe9238b0",
  5602 => x"7934a33d",
  5603 => x"088105a4",
  5604 => x"3d0cea39",
  5605 => x"b07f7081",
  5606 => x"054134b0",
  5607 => x"1b59787f",
  5608 => x"70810541",
  5609 => x"347e6231",
  5610 => x"a53d0870",
  5611 => x"12415a4d",
  5612 => x"81792580",
  5613 => x"ff38811f",
  5614 => x"5f83bc3d",
  5615 => x"33597880",
  5616 => x"2edfb038",
  5617 => x"ad0b83be",
  5618 => x"3d34dfa7",
  5619 => x"39810b80",
  5620 => x"085a5a7f",
  5621 => x"80c52e09",
  5622 => x"8106fcd3",
  5623 => x"388159fc",
  5624 => x"ce398008",
  5625 => x"335978b0",
  5626 => x"2ea8386e",
  5627 => x"087b055b",
  5628 => x"fef53980",
  5629 => x"e740a43d",
  5630 => x"0859787a",
  5631 => x"2483f938",
  5632 => x"79638106",
  5633 => x"5a5f7880",
  5634 => x"2effae38",
  5635 => x"811a5fff",
  5636 => x"a8398059",
  5637 => x"80795454",
  5638 => x"7d517e52",
  5639 => x"80fea63f",
  5640 => x"8008802e",
  5641 => x"c6388162",
  5642 => x"3170a13d",
  5643 => x"080c7b05",
  5644 => x"5bfeb439",
  5645 => x"62810659",
  5646 => x"78802efe",
  5647 => x"fc38811f",
  5648 => x"5ffef639",
  5649 => x"82c7b87c",
  5650 => x"0c810b84",
  5651 => x"1d0c83b7",
  5652 => x"3d088105",
  5653 => x"83b83d0c",
  5654 => x"881c83b7",
  5655 => x"3d088111",
  5656 => x"83b93d0c",
  5657 => x"8111515a",
  5658 => x"5c788724",
  5659 => x"81e03879",
  5660 => x"8938a43d",
  5661 => x"08802ee1",
  5662 => x"82386b7c",
  5663 => x"0c810b84",
  5664 => x"1d0c83b7",
  5665 => x"3d088105",
  5666 => x"83b83d0c",
  5667 => x"881c83b7",
  5668 => x"3d088111",
  5669 => x"83b93d0c",
  5670 => x"8111515a",
  5671 => x"5c788724",
  5672 => x"81c53879",
  5673 => x"305a807a",
  5674 => x"2580f338",
  5675 => x"907a25b4",
  5676 => x"3882c3fc",
  5677 => x"7c0c900b",
  5678 => x"841d0c83",
  5679 => x"b73d0890",
  5680 => x"0583b83d",
  5681 => x"0c881c83",
  5682 => x"b73d0881",
  5683 => x"1183b93d",
  5684 => x"0c811151",
  5685 => x"5a5c7887",
  5686 => x"2480db38",
  5687 => x"f01a5a79",
  5688 => x"9024ce38",
  5689 => x"82c3fc7c",
  5690 => x"0c79841d",
  5691 => x"0c83b73d",
  5692 => x"081a83b8",
  5693 => x"3d0c881c",
  5694 => x"83b73d08",
  5695 => x"811183b9",
  5696 => x"3d0c8111",
  5697 => x"515a5c87",
  5698 => x"79259338",
  5699 => x"83be3ddc",
  5700 => x"05526651",
  5701 => x"d7dd3f80",
  5702 => x"08e4ec38",
  5703 => x"655c7d7c",
  5704 => x"0ca43d08",
  5705 => x"841d0c83",
  5706 => x"b73d08a5",
  5707 => x"3d080583",
  5708 => x"b83d0cf1",
  5709 => x"f13983be",
  5710 => x"3ddc0552",
  5711 => x"6651d7b3",
  5712 => x"3f8008e4",
  5713 => x"c23865f0",
  5714 => x"1b5b5cff",
  5715 => x"923983be",
  5716 => x"3ddc0552",
  5717 => x"6651d79b",
  5718 => x"3f8008e4",
  5719 => x"aa3865a6",
  5720 => x"3d085b5c",
  5721 => x"fe893983",
  5722 => x"be3ddc05",
  5723 => x"526651d7",
  5724 => x"823f8008",
  5725 => x"e4913865",
  5726 => x"a63d0870",
  5727 => x"30515b5c",
  5728 => x"798024fe",
  5729 => x"a738ff96",
  5730 => x"398641e6",
  5731 => x"c33982c7",
  5732 => x"c45e865f",
  5733 => x"dbdd39a5",
  5734 => x"3d085afa",
  5735 => x"c6397f80",
  5736 => x"e62e0981",
  5737 => x"06fccf38",
  5738 => x"807a2581",
  5739 => x"8d38795f",
  5740 => x"608b3862",
  5741 => x"81065978",
  5742 => x"802efbfd",
  5743 => x"38601a81",
  5744 => x"055ffbf5",
  5745 => x"3983b73d",
  5746 => x"088a3880",
  5747 => x"0b83b73d",
  5748 => x"0ce3b439",
  5749 => x"83be3ddc",
  5750 => x"05526651",
  5751 => x"d6953f80",
  5752 => x"08e3a438",
  5753 => x"800b83b7",
  5754 => x"3d0ce39b",
  5755 => x"397d810a",
  5756 => x"325ead7b",
  5757 => x"34f8de39",
  5758 => x"787a3182",
  5759 => x"055f807a",
  5760 => x"25fbb638",
  5761 => x"81195ffb",
  5762 => x"b0397930",
  5763 => x"5bad7f34",
  5764 => x"028dde05",
  5765 => x"b33d705c",
  5766 => x"425f897b",
  5767 => x"25faf538",
  5768 => x"f9f63964",
  5769 => x"65840571",
  5770 => x"08434659",
  5771 => x"608025d9",
  5772 => x"8f38ff7d",
  5773 => x"335b41d9",
  5774 => x"8a39608d",
  5775 => x"38628106",
  5776 => x"59815f78",
  5777 => x"802efaf1",
  5778 => x"38608205",
  5779 => x"5ffaea39",
  5780 => x"fc3d0d82",
  5781 => x"d4800855",
  5782 => x"b8150880",
  5783 => x"2e933878",
  5784 => x"54775376",
  5785 => x"5282d480",
  5786 => x"0851d5b8",
  5787 => x"3f863d0d",
  5788 => x"047451b3",
  5789 => x"fb3f7854",
  5790 => x"77537652",
  5791 => x"82d48008",
  5792 => x"51d5a13f",
  5793 => x"863d0d04",
  5794 => x"f63d0d7c",
  5795 => x"7e615956",
  5796 => x"58805674",
  5797 => x"762e9c38",
  5798 => x"76547e53",
  5799 => x"74527751",
  5800 => x"82b73f80",
  5801 => x"08558008",
  5802 => x"ff2ea238",
  5803 => x"74800c8c",
  5804 => x"3d0d0476",
  5805 => x"5475538c",
  5806 => x"3df40552",
  5807 => x"77518299",
  5808 => x"3f800855",
  5809 => x"8008ff2e",
  5810 => x"098106e0",
  5811 => x"3880770c",
  5812 => x"818a780c",
  5813 => x"74800c8c",
  5814 => x"3d0d04fd",
  5815 => x"3d0d7754",
  5816 => x"76537552",
  5817 => x"82d48008",
  5818 => x"51ff9d3f",
  5819 => x"853d0d04",
  5820 => x"ec3d0d66",
  5821 => x"686a6c6e",
  5822 => x"735c405d",
  5823 => x"42424260",
  5824 => x"802e818c",
  5825 => x"38806008",
  5826 => x"5a5d7c7a",
  5827 => x"2780f838",
  5828 => x"933d5b7b",
  5829 => x"08841d08",
  5830 => x"7d567a08",
  5831 => x"557c5463",
  5832 => x"53405efe",
  5833 => x"e33f8008",
  5834 => x"588008ff",
  5835 => x"2e80f138",
  5836 => x"807a8008",
  5837 => x"3156567c",
  5838 => x"75268338",
  5839 => x"81568008",
  5840 => x"7a2780d1",
  5841 => x"3875802e",
  5842 => x"80cb3880",
  5843 => x"081d5d60",
  5844 => x"802ea238",
  5845 => x"80567580",
  5846 => x"08259438",
  5847 => x"751b5574",
  5848 => x"33777081",
  5849 => x"05593481",
  5850 => x"16567776",
  5851 => x"24ee387f",
  5852 => x"08840560",
  5853 => x"0c787084",
  5854 => x"055a0855",
  5855 => x"74802eaf",
  5856 => x"38797d26",
  5857 => x"ff8d387c",
  5858 => x"5574800c",
  5859 => x"963d0d04",
  5860 => x"ff5afef1",
  5861 => x"397d7c0c",
  5862 => x"7e841d0c",
  5863 => x"7c55ea39",
  5864 => x"818a620c",
  5865 => x"807c0c80",
  5866 => x"08800c96",
  5867 => x"3d0d0460",
  5868 => x"802e8438",
  5869 => x"74600c74",
  5870 => x"7c0cff1d",
  5871 => x"800c963d",
  5872 => x"0d04fc3d",
  5873 => x"0d795578",
  5874 => x"54775376",
  5875 => x"5282d480",
  5876 => x"0851fe9c",
  5877 => x"3f863d0d",
  5878 => x"04f83d0d",
  5879 => x"7b7d7f82",
  5880 => x"db805459",
  5881 => x"575580e9",
  5882 => x"a23f8008",
  5883 => x"81269438",
  5884 => x"74547480",
  5885 => x"2e863875",
  5886 => x"75348154",
  5887 => x"73800c8a",
  5888 => x"3d0d0482",
  5889 => x"c7cc5282",
  5890 => x"db805180",
  5891 => x"e7e83f80",
  5892 => x"0881c138",
  5893 => x"80085474",
  5894 => x"802ee138",
  5895 => x"80ff7625",
  5896 => x"d638ff80",
  5897 => x"16538eff",
  5898 => x"732784ef",
  5899 => x"38f08016",
  5900 => x"5383efff",
  5901 => x"732782a9",
  5902 => x"38fc8080",
  5903 => x"165380fb",
  5904 => x"ffff7327",
  5905 => x"84f7388f",
  5906 => x"ff0a1653",
  5907 => x"f7c00a73",
  5908 => x"2785b838",
  5909 => x"ff54c00a",
  5910 => x"7625ffa0",
  5911 => x"3875820a",
  5912 => x"06709e2c",
  5913 => x"70fc0751",
  5914 => x"51537275",
  5915 => x"70810557",
  5916 => x"347581fc",
  5917 => x"0a067098",
  5918 => x"2aff8007",
  5919 => x"51537275",
  5920 => x"70810557",
  5921 => x"347587f0",
  5922 => x"80800670",
  5923 => x"922aff80",
  5924 => x"07515372",
  5925 => x"75708105",
  5926 => x"5734758f",
  5927 => x"e0800670",
  5928 => x"8c2aff80",
  5929 => x"07515372",
  5930 => x"75708105",
  5931 => x"5734759f",
  5932 => x"c0067086",
  5933 => x"2aff8007",
  5934 => x"51537275",
  5935 => x"70810557",
  5936 => x"3475ffbf",
  5937 => x"06ff8007",
  5938 => x"53727534",
  5939 => x"860b800c",
  5940 => x"8a3d0d04",
  5941 => x"82c7d452",
  5942 => x"82db8051",
  5943 => x"80e6973f",
  5944 => x"800881d7",
  5945 => x"387581ff",
  5946 => x"0676882c",
  5947 => x"7081ff06",
  5948 => x"80085759",
  5949 => x"54587480",
  5950 => x"2efe8138",
  5951 => x"76802efd",
  5952 => x"ef388008",
  5953 => x"80ff1870",
  5954 => x"81ff0651",
  5955 => x"5456729e",
  5956 => x"26833881",
  5957 => x"568008a0",
  5958 => x"187081ff",
  5959 => x"06515454",
  5960 => x"728f2683",
  5961 => x"38815475",
  5962 => x"74075372",
  5963 => x"802eaa38",
  5964 => x"8008c019",
  5965 => x"545672be",
  5966 => x"26833881",
  5967 => x"568008ff",
  5968 => x"80197081",
  5969 => x"ff065154",
  5970 => x"547280fc",
  5971 => x"26833881",
  5972 => x"54757407",
  5973 => x"537280d0",
  5974 => x"38ff0b80",
  5975 => x"0c8a3d0d",
  5976 => x"04fcd080",
  5977 => x"1653ff54",
  5978 => x"8fff7327",
  5979 => x"fd8e3875",
  5980 => x"83e08006",
  5981 => x"708c2ae0",
  5982 => x"07515372",
  5983 => x"75708105",
  5984 => x"5734759f",
  5985 => x"c0067086",
  5986 => x"2aff8007",
  5987 => x"51537275",
  5988 => x"70810557",
  5989 => x"3475ffbf",
  5990 => x"06ff8007",
  5991 => x"53727534",
  5992 => x"830b800c",
  5993 => x"8a3d0d04",
  5994 => x"76757081",
  5995 => x"05573477",
  5996 => x"75348254",
  5997 => x"73800c8a",
  5998 => x"3d0d0482",
  5999 => x"c7dc5282",
  6000 => x"db805180",
  6001 => x"e4b03f80",
  6002 => x"0880db38",
  6003 => x"7581ff06",
  6004 => x"76882c70",
  6005 => x"81ff0680",
  6006 => x"08575954",
  6007 => x"5874802e",
  6008 => x"fc9a3876",
  6009 => x"802efc88",
  6010 => x"38800853",
  6011 => x"81a07727",
  6012 => x"83388153",
  6013 => x"7681ff2e",
  6014 => x"fedf3881",
  6015 => x"70740654",
  6016 => x"5472802e",
  6017 => x"fed33880",
  6018 => x"085381a0",
  6019 => x"78278338",
  6020 => x"73537781",
  6021 => x"ff2efec1",
  6022 => x"38727406",
  6023 => x"5372802e",
  6024 => x"feb738ff",
  6025 => x"833982c7",
  6026 => x"e45282db",
  6027 => x"805180e3",
  6028 => x"c53f8008",
  6029 => x"fbba3880",
  6030 => x"087681ff",
  6031 => x"0677882c",
  6032 => x"7081ff06",
  6033 => x"59555959",
  6034 => x"81547480",
  6035 => x"2efbad38",
  6036 => x"75802e82",
  6037 => x"9838df16",
  6038 => x"537280dd",
  6039 => x"26fdfa38",
  6040 => x"df185372",
  6041 => x"80dd26fd",
  6042 => x"f0387608",
  6043 => x"9c387377",
  6044 => x"0c9b7570",
  6045 => x"81055734",
  6046 => x"a4757081",
  6047 => x"05573480",
  6048 => x"c2757081",
  6049 => x"05573483",
  6050 => x"59757570",
  6051 => x"81055734",
  6052 => x"77753482",
  6053 => x"19800c8a",
  6054 => x"3d0d0475",
  6055 => x"8fc00670",
  6056 => x"862ac007",
  6057 => x"51537275",
  6058 => x"70810557",
  6059 => x"3475ffbf",
  6060 => x"06ff8007",
  6061 => x"53727534",
  6062 => x"8254fdf8",
  6063 => x"397580f0",
  6064 => x"80800670",
  6065 => x"922af007",
  6066 => x"51537275",
  6067 => x"70810557",
  6068 => x"34758fe0",
  6069 => x"8006708c",
  6070 => x"2aff8007",
  6071 => x"51537275",
  6072 => x"70810557",
  6073 => x"34759fc0",
  6074 => x"0670862a",
  6075 => x"ff800751",
  6076 => x"53727570",
  6077 => x"81055734",
  6078 => x"75ffbf06",
  6079 => x"ff800753",
  6080 => x"72753484",
  6081 => x"0b800c8a",
  6082 => x"3d0d0475",
  6083 => x"81c00a06",
  6084 => x"70982af8",
  6085 => x"07515372",
  6086 => x"75708105",
  6087 => x"57347587",
  6088 => x"f0808006",
  6089 => x"70922aff",
  6090 => x"80075153",
  6091 => x"72757081",
  6092 => x"05573475",
  6093 => x"8fe08006",
  6094 => x"708c2aff",
  6095 => x"80075153",
  6096 => x"72757081",
  6097 => x"05573475",
  6098 => x"9fc00670",
  6099 => x"862aff80",
  6100 => x"07515372",
  6101 => x"75708105",
  6102 => x"573475ff",
  6103 => x"bf06ff80",
  6104 => x"07537275",
  6105 => x"34850b80",
  6106 => x"0c8a3d0d",
  6107 => x"04760880",
  6108 => x"2e9d3880",
  6109 => x"08770c9b",
  6110 => x"75708105",
  6111 => x"5734a875",
  6112 => x"70810557",
  6113 => x"3480c275",
  6114 => x"70810557",
  6115 => x"34835977",
  6116 => x"75348119",
  6117 => x"800c8a3d",
  6118 => x"0d04fa3d",
  6119 => x"0d7882d4",
  6120 => x"80085455",
  6121 => x"b8130880",
  6122 => x"2e81b638",
  6123 => x"8c152270",
  6124 => x"83ffff06",
  6125 => x"70832a81",
  6126 => x"32708106",
  6127 => x"51555556",
  6128 => x"72802e80",
  6129 => x"dc387384",
  6130 => x"2a813281",
  6131 => x"0657ff53",
  6132 => x"7680f738",
  6133 => x"73822a70",
  6134 => x"81065153",
  6135 => x"72802eb9",
  6136 => x"38b01508",
  6137 => x"5473802e",
  6138 => x"9c3880c0",
  6139 => x"15537373",
  6140 => x"2e8f3873",
  6141 => x"5282d480",
  6142 => x"0851ace3",
  6143 => x"3f8c1522",
  6144 => x"5676b016",
  6145 => x"0c75db06",
  6146 => x"53728c16",
  6147 => x"23800b84",
  6148 => x"160c9015",
  6149 => x"08750c72",
  6150 => x"56758807",
  6151 => x"53728c16",
  6152 => x"23901508",
  6153 => x"802e80c1",
  6154 => x"388c1522",
  6155 => x"70810655",
  6156 => x"53739e38",
  6157 => x"720a100a",
  6158 => x"70810651",
  6159 => x"53728538",
  6160 => x"94150854",
  6161 => x"7388160c",
  6162 => x"80537280",
  6163 => x"0c883d0d",
  6164 => x"04800b88",
  6165 => x"160c9415",
  6166 => x"08309816",
  6167 => x"0c8053ea",
  6168 => x"397251a8",
  6169 => x"8b3ffec4",
  6170 => x"397451b8",
  6171 => x"e43f8c15",
  6172 => x"22708106",
  6173 => x"55537380",
  6174 => x"2effb938",
  6175 => x"d439ef3d",
  6176 => x"0d636590",
  6177 => x"11085e40",
  6178 => x"4080537b",
  6179 => x"60900508",
  6180 => x"2481b338",
  6181 => x"941f70ff",
  6182 => x"1e70822b",
  6183 => x"73116494",
  6184 => x"05705c43",
  6185 => x"5f610570",
  6186 => x"087f0881",
  6187 => x"0557555c",
  6188 => x"5e425780",
  6189 => x"f8bc3f80",
  6190 => x"085d8008",
  6191 => x"818f387e",
  6192 => x"527f5180",
  6193 => x"c9e53f80",
  6194 => x"0b800824",
  6195 => x"80f63881",
  6196 => x"1d5d8070",
  6197 => x"7f635a58",
  6198 => x"5b587670",
  6199 => x"84055808",
  6200 => x"7083ffff",
  6201 => x"067b0571",
  6202 => x"902a7190",
  6203 => x"2a057090",
  6204 => x"2a5d5283",
  6205 => x"ffff0682",
  6206 => x"18227072",
  6207 => x"311b585b",
  6208 => x"5483ffff",
  6209 => x"06762270",
  6210 => x"72317790",
  6211 => x"2c057090",
  6212 => x"2c5b5243",
  6213 => x"53727623",
  6214 => x"74821723",
  6215 => x"8416567a",
  6216 => x"7727ffb6",
  6217 => x"387b1010",
  6218 => x"1e597808",
  6219 => x"9738fc19",
  6220 => x"597d7927",
  6221 => x"8a387808",
  6222 => x"8638ff1c",
  6223 => x"5cf0397b",
  6224 => x"6090050c",
  6225 => x"7c537280",
  6226 => x"0c933d0d",
  6227 => x"0480705b",
  6228 => x"58767084",
  6229 => x"05580870",
  6230 => x"83ffff06",
  6231 => x"707f291c",
  6232 => x"72902a60",
  6233 => x"2971902a",
  6234 => x"0570902a",
  6235 => x"5e5283ff",
  6236 => x"ff068219",
  6237 => x"22707231",
  6238 => x"1c594552",
  6239 => x"83ffff06",
  6240 => x"77227072",
  6241 => x"3178902c",
  6242 => x"0570902c",
  6243 => x"5c525651",
  6244 => x"53727623",
  6245 => x"74821723",
  6246 => x"8416567a",
  6247 => x"7727ffb1",
  6248 => x"387808fe",
  6249 => x"9a38fc19",
  6250 => x"597d7927",
  6251 => x"8a387808",
  6252 => x"8638ff1c",
  6253 => x"5cf0397b",
  6254 => x"6090050c",
  6255 => x"fe81398c",
  6256 => x"08c83d0d",
  6257 => x"bc3d0880",
  6258 => x"c03d0880",
  6259 => x"c23d0880",
  6260 => x"c53d0880",
  6261 => x"c73d088c",
  6262 => x"0c5d4b43",
  6263 => x"40800bbe",
  6264 => x"3d0880c0",
  6265 => x"3d085bba",
  6266 => x"3d0c79bb",
  6267 => x"3d0c6080",
  6268 => x"c0050857",
  6269 => x"4875682e",
  6270 => x"09810680",
  6271 => x"d938b83d",
  6272 => x"08578077",
  6273 => x"2480f838",
  6274 => x"677a0c76",
  6275 => x"9ffe0a06",
  6276 => x"56759ffe",
  6277 => x"0a2e8184",
  6278 => x"38b83d08",
  6279 => x"ba3d085a",
  6280 => x"58805680",
  6281 => x"76545477",
  6282 => x"51785280",
  6283 => x"e8ab3f80",
  6284 => x"0881a538",
  6285 => x"80c13d08",
  6286 => x"5881780c",
  6287 => x"82c7b85f",
  6288 => x"8c08802e",
  6289 => x"8638811f",
  6290 => x"8c080c7e",
  6291 => x"5675800c",
  6292 => x"ba3d0d8c",
  6293 => x"0c047f80",
  6294 => x"c4050884",
  6295 => x"170c8160",
  6296 => x"80c40508",
  6297 => x"2b88170c",
  6298 => x"75527f51",
  6299 => x"bbe33f67",
  6300 => x"6080c005",
  6301 => x"0cb83d08",
  6302 => x"57768025",
  6303 => x"ff8a3881",
  6304 => x"7a0c76fe",
  6305 => x"0a0670ba",
  6306 => x"3d0c709f",
  6307 => x"fe0a0657",
  6308 => x"57759ffe",
  6309 => x"0a2e0981",
  6310 => x"06fefe38",
  6311 => x"80c13d08",
  6312 => x"5680ce8f",
  6313 => x"760cb93d",
  6314 => x"0883ff38",
  6315 => x"76bfffff",
  6316 => x"0682c7ec",
  6317 => x"40567583",
  6318 => x"f1388c08",
  6319 => x"802eff8b",
  6320 => x"38831f33",
  6321 => x"7f880558",
  6322 => x"56758438",
  6323 => x"831f5776",
  6324 => x"8c080c7e",
  6325 => x"56fef639",
  6326 => x"ba3dffb4",
  6327 => x"1156ffb0",
  6328 => x"05547752",
  6329 => x"78537f51",
  6330 => x"80cb843f",
  6331 => x"8008b93d",
  6332 => x"0870942a",
  6333 => x"8fff065e",
  6334 => x"59417b83",
  6335 => x"b438a73d",
  6336 => x"08a73d08",
  6337 => x"0588b211",
  6338 => x"5d56a07c",
  6339 => x"258e8138",
  6340 => x"80c07c31",
  6341 => x"88921779",
  6342 => x"722bbc3d",
  6343 => x"08722a07",
  6344 => x"b53d7156",
  6345 => x"70555d51",
  6346 => x"5757ff94",
  6347 => x"9e3fb23d",
  6348 => x"08b43d08",
  6349 => x"b23d5d5a",
  6350 => x"58807624",
  6351 => x"91a23877",
  6352 => x"b73d0c78",
  6353 => x"b83d0cb6",
  6354 => x"3d0890ff",
  6355 => x"0a05b73d",
  6356 => x"0cf7cd1c",
  6357 => x"5c814ebf",
  6358 => x"fc0a5680",
  6359 => x"765555b6",
  6360 => x"3d08b83d",
  6361 => x"08585276",
  6362 => x"537a51fe",
  6363 => x"e4f63f83",
  6364 => x"feca8fa7",
  6365 => x"56869bbd",
  6366 => x"86e17655",
  6367 => x"55b03d08",
  6368 => x"b23d0858",
  6369 => x"52765379",
  6370 => x"51fee681",
  6371 => x"3f83fe9a",
  6372 => x"94a856f8",
  6373 => x"db8391b3",
  6374 => x"765555b2",
  6375 => x"3d08b43d",
  6376 => x"08585276",
  6377 => x"53ba3dd0",
  6378 => x"0551fee3",
  6379 => x"9a3fae3d",
  6380 => x"08b03d08",
  6381 => x"7d54ae3d",
  6382 => x"535a58ff",
  6383 => x"938d3faa",
  6384 => x"3d4c83fe",
  6385 => x"cd889356",
  6386 => x"8584fdf3",
  6387 => x"fb765555",
  6388 => x"ac3d08ae",
  6389 => x"3d085852",
  6390 => x"76536b51",
  6391 => x"fee5ae3f",
  6392 => x"a83dab3d",
  6393 => x"08ad3d08",
  6394 => x"59557756",
  6395 => x"78537954",
  6396 => x"705245fe",
  6397 => x"e2d13fa8",
  6398 => x"3d08aa3d",
  6399 => x"08715370",
  6400 => x"545f5d80",
  6401 => x"edef3f80",
  6402 => x"08438056",
  6403 => x"80765454",
  6404 => x"7c517d52",
  6405 => x"80ea863f",
  6406 => x"800b8008",
  6407 => x"248cc338",
  6408 => x"810ba23d",
  6409 => x"0c629626",
  6410 => x"ae386210",
  6411 => x"101082c9",
  6412 => x"a0058411",
  6413 => x"08710855",
  6414 => x"55b93d08",
  6415 => x"bb3d0859",
  6416 => x"52567652",
  6417 => x"80e9d63f",
  6418 => x"800b8008",
  6419 => x"24637131",
  6420 => x"4456800b",
  6421 => x"a23d0ca7",
  6422 => x"3d087c31",
  6423 => x"ff055a80",
  6424 => x"7a454b6a",
  6425 => x"7a248bd1",
  6426 => x"38806324",
  6427 => x"9aad3880",
  6428 => x"0ba63d0c",
  6429 => x"624f6363",
  6430 => x"05448962",
  6431 => x"27833880",
  6432 => x"42815885",
  6433 => x"62258738",
  6434 => x"61fc0542",
  6435 => x"8058810b",
  6436 => x"a13d0cff",
  6437 => x"70a53d0c",
  6438 => x"46618526",
  6439 => x"829c3861",
  6440 => x"101082c7",
  6441 => x"f8055675",
  6442 => x"080482c7",
  6443 => x"c05ffc8a",
  6444 => x"39b83d08",
  6445 => x"ba3d0858",
  6446 => x"b73d0c76",
  6447 => x"b83d0cb6",
  6448 => x"3d08fc0a",
  6449 => x"069ffc0a",
  6450 => x"07b73d0c",
  6451 => x"f8811c5c",
  6452 => x"804eb23d",
  6453 => x"b13d5c5a",
  6454 => x"bffc0a56",
  6455 => x"80765555",
  6456 => x"b63d08b8",
  6457 => x"3d085852",
  6458 => x"76537a51",
  6459 => x"fee1f53f",
  6460 => x"83feca8f",
  6461 => x"a756869b",
  6462 => x"bd86e176",
  6463 => x"5555b03d",
  6464 => x"08b23d08",
  6465 => x"58527653",
  6466 => x"7951fee3",
  6467 => x"803f83fe",
  6468 => x"9a94a856",
  6469 => x"f8db8391",
  6470 => x"b3765555",
  6471 => x"b23d08b4",
  6472 => x"3d085852",
  6473 => x"7653ba3d",
  6474 => x"d00551fe",
  6475 => x"e0993fae",
  6476 => x"3d08b03d",
  6477 => x"087d54ae",
  6478 => x"3d535a58",
  6479 => x"ff908c3f",
  6480 => x"aa3d4c83",
  6481 => x"fecd8893",
  6482 => x"568584fd",
  6483 => x"f3fb7655",
  6484 => x"55ac3d08",
  6485 => x"ae3d0858",
  6486 => x"5276536b",
  6487 => x"51fee2ad",
  6488 => x"3fa83dab",
  6489 => x"3d08ad3d",
  6490 => x"08595577",
  6491 => x"56785379",
  6492 => x"54705245",
  6493 => x"fedfd03f",
  6494 => x"a83d08aa",
  6495 => x"3d087153",
  6496 => x"70545f5d",
  6497 => x"80eaee3f",
  6498 => x"80084380",
  6499 => x"56807654",
  6500 => x"547c517d",
  6501 => x"5280e785",
  6502 => x"3f800880",
  6503 => x"25fd8138",
  6504 => x"89c03980",
  6505 => x"0ba13d0c",
  6506 => x"68630581",
  6507 => x"1170485d",
  6508 => x"a43d0c7b",
  6509 => x"80248338",
  6510 => x"815c845a",
  6511 => x"806080c4",
  6512 => x"050c987c",
  6513 => x"26973880",
  6514 => x"5781177a",
  6515 => x"10941158",
  6516 => x"5b577b76",
  6517 => x"27f33876",
  6518 => x"6080c405",
  6519 => x"0c7f80c4",
  6520 => x"0508527f",
  6521 => x"51b3e03f",
  6522 => x"80086080",
  6523 => x"c0050c80",
  6524 => x"0880088e",
  6525 => x"68275840",
  6526 => x"4d77802e",
  6527 => x"86903875",
  6528 => x"802e868a",
  6529 => x"38b83d08",
  6530 => x"ba3d0871",
  6531 => x"b93d0c70",
  6532 => x"ba3d0c64",
  6533 => x"a53d0c67",
  6534 => x"a73d0c5a",
  6535 => x"58825c80",
  6536 => x"63258ad7",
  6537 => x"3862832b",
  6538 => x"80f80682",
  6539 => x"c9a01108",
  6540 => x"82c9a412",
  6541 => x"0865842c",
  6542 => x"70842a70",
  6543 => x"81065154",
  6544 => x"5d405e56",
  6545 => x"7588e438",
  6546 => x"79802e9f",
  6547 => x"3882c8f8",
  6548 => x"58798106",
  6549 => x"567587e9",
  6550 => x"3879812c",
  6551 => x"8819595a",
  6552 => x"79ef38b8",
  6553 => x"3d08ba3d",
  6554 => x"085a587c",
  6555 => x"547d5577",
  6556 => x"52785364",
  6557 => x"51fefda4",
  6558 => x"3fa83d08",
  6559 => x"aa3d0871",
  6560 => x"bb3d0c70",
  6561 => x"bc3d0c5a",
  6562 => x"58a13d08",
  6563 => x"802e80d9",
  6564 => x"38805a9f",
  6565 => x"fc0a5680",
  6566 => x"76545477",
  6567 => x"51785280",
  6568 => x"e4fb3f79",
  6569 => x"8008248b",
  6570 => x"f3388066",
  6571 => x"25bb3879",
  6572 => x"802eb638",
  6573 => x"800ba43d",
  6574 => x"082584ba",
  6575 => x"38a33d08",
  6576 => x"63ff0544",
  6577 => x"4680c882",
  6578 => x"0a568076",
  6579 => x"55557752",
  6580 => x"78536451",
  6581 => x"fedfb63f",
  6582 => x"a83d08aa",
  6583 => x"3d085ab9",
  6584 => x"3d0c78ba",
  6585 => x"3d0c811c",
  6586 => x"5c7b5264",
  6587 => x"51ff8cdb",
  6588 => x"3fb83d08",
  6589 => x"ba3d0858",
  6590 => x"547655a8",
  6591 => x"3d08aa3d",
  6592 => x"08585276",
  6593 => x"536b51fe",
  6594 => x"df833f80",
  6595 => x"f0820a56",
  6596 => x"80765555",
  6597 => x"aa3d08ac",
  6598 => x"3d085852",
  6599 => x"7653ac3d",
  6600 => x"51fedca3",
  6601 => x"3fac3d08",
  6602 => x"ae3d0858",
  6603 => x"b53d0c76",
  6604 => x"b63d0cb4",
  6605 => x"3d0886bf",
  6606 => x"0a05b53d",
  6607 => x"0c65802e",
  6608 => x"96bd386f",
  6609 => x"802e94f2",
  6610 => x"38651010",
  6611 => x"1082c998",
  6612 => x"05841108",
  6613 => x"71085656",
  6614 => x"568ffc0a",
  6615 => x"56807653",
  6616 => x"536451fe",
  6617 => x"fbb63fb4",
  6618 => x"3d08b63d",
  6619 => x"08585476",
  6620 => x"55a83d08",
  6621 => x"aa3d0858",
  6622 => x"5276536b",
  6623 => x"51fedce4",
  6624 => x"3faa3d08",
  6625 => x"ac3d0858",
  6626 => x"b53d0c76",
  6627 => x"b63d0c80",
  6628 => x"0bb93d08",
  6629 => x"bb3d085b",
  6630 => x"595c80c8",
  6631 => x"820a5d80",
  6632 => x"5e775178",
  6633 => x"5280e6cd",
  6634 => x"3f800880",
  6635 => x"08536552",
  6636 => x"5aff8b97",
  6637 => x"3fa83d08",
  6638 => x"aa3d0858",
  6639 => x"547655b8",
  6640 => x"3d08ba3d",
  6641 => x"08585276",
  6642 => x"536b51fe",
  6643 => x"dc963faa",
  6644 => x"3d08ac3d",
  6645 => x"085ab93d",
  6646 => x"0c78ba3d",
  6647 => x"0cb01a56",
  6648 => x"757f7081",
  6649 => x"054134b8",
  6650 => x"3d08ba3d",
  6651 => x"08b63d08",
  6652 => x"b83d085a",
  6653 => x"55785671",
  6654 => x"5370545a",
  6655 => x"5880e29d",
  6656 => x"3f800b80",
  6657 => x"082486cc",
  6658 => x"38775478",
  6659 => x"559ffc0a",
  6660 => x"56807653",
  6661 => x"536451fe",
  6662 => x"dbca3fb4",
  6663 => x"3d08b63d",
  6664 => x"08715570",
  6665 => x"56aa3d08",
  6666 => x"ac3d085a",
  6667 => x"5378545a",
  6668 => x"5880e1e9",
  6669 => x"3f800b80",
  6670 => x"082485ed",
  6671 => x"38811c5c",
  6672 => x"7b662581",
  6673 => x"b1387c54",
  6674 => x"7d557752",
  6675 => x"78536b51",
  6676 => x"fedcba3f",
  6677 => x"aa3d08ac",
  6678 => x"3d0858b5",
  6679 => x"3d0c76b6",
  6680 => x"3d0c7c54",
  6681 => x"7d55b83d",
  6682 => x"08ba3d08",
  6683 => x"58527653",
  6684 => x"6451fedc",
  6685 => x"983fa83d",
  6686 => x"08aa3d08",
  6687 => x"71bb3d0c",
  6688 => x"70bc3d0c",
  6689 => x"5a58fe99",
  6690 => x"398ffc0a",
  6691 => x"58807855",
  6692 => x"7056b53d",
  6693 => x"08b73d08",
  6694 => x"59537754",
  6695 => x"655259fe",
  6696 => x"d9a53fa8",
  6697 => x"3d08aa3d",
  6698 => x"08585376",
  6699 => x"54b83d08",
  6700 => x"ba3d0858",
  6701 => x"51765280",
  6702 => x"def73f80",
  6703 => x"08802484",
  6704 => x"e838b43d",
  6705 => x"08b63d08",
  6706 => x"58547655",
  6707 => x"77527853",
  6708 => x"6b51feda",
  6709 => x"8f3faa3d",
  6710 => x"08ac3d08",
  6711 => x"58537654",
  6712 => x"b83d08ba",
  6713 => x"3d085851",
  6714 => x"765280e0",
  6715 => x"b03f800b",
  6716 => x"80082492",
  6717 => x"f9386cb7",
  6718 => x"3d08b93d",
  6719 => x"085bba3d",
  6720 => x"0c79bb3d",
  6721 => x"0ca33d08",
  6722 => x"a63d0848",
  6723 => x"445f800b",
  6724 => x"a73d0857",
  6725 => x"58777624",
  6726 => x"83388158",
  6727 => x"80780657",
  6728 => x"628e2487",
  6729 => x"e5388170",
  6730 => x"79065859",
  6731 => x"76802e87",
  6732 => x"d9386210",
  6733 => x"101082c9",
  6734 => x"a0057008",
  6735 => x"84120880",
  6736 => x"6c245340",
  6737 => x"5e568066",
  6738 => x"2585c838",
  6739 => x"810bb93d",
  6740 => x"08bb3d08",
  6741 => x"5b595c7c",
  6742 => x"547d5577",
  6743 => x"52785364",
  6744 => x"51fef7b8",
  6745 => x"3fa83d08",
  6746 => x"aa3d0858",
  6747 => x"51765280",
  6748 => x"e3833f80",
  6749 => x"08800853",
  6750 => x"65525aff",
  6751 => x"87cd3f7c",
  6752 => x"547d55a8",
  6753 => x"3d08aa3d",
  6754 => x"08585276",
  6755 => x"536b51fe",
  6756 => x"d9fb3faa",
  6757 => x"3d08ac3d",
  6758 => x"08585476",
  6759 => x"55b83d08",
  6760 => x"ba3d0858",
  6761 => x"527653ac",
  6762 => x"3d51fed8",
  6763 => x"b73fac3d",
  6764 => x"08ae3d08",
  6765 => x"5ab93d0c",
  6766 => x"78ba3d0c",
  6767 => x"b01a5675",
  6768 => x"7f708105",
  6769 => x"41347b66",
  6770 => x"2e828f38",
  6771 => x"80c8820a",
  6772 => x"56807655",
  6773 => x"55b83d08",
  6774 => x"ba3d0858",
  6775 => x"52765364",
  6776 => x"51fed9a9",
  6777 => x"3fa83d08",
  6778 => x"aa3d0871",
  6779 => x"bb3d0c70",
  6780 => x"bc3d0c5a",
  6781 => x"58805680",
  6782 => x"76545477",
  6783 => x"51785280",
  6784 => x"d8d73f80",
  6785 => x"08802e82",
  6786 => x"cb38811c",
  6787 => x"5cfec839",
  6788 => x"a07c31ba",
  6789 => x"3d08712b",
  6790 => x"b43d7155",
  6791 => x"70545c51",
  6792 => x"56ff86a7",
  6793 => x"3fb23d08",
  6794 => x"b43d08b2",
  6795 => x"3d5d5a58",
  6796 => x"758025f2",
  6797 => x"8a3883a8",
  6798 => x"3979304b",
  6799 => x"8044f4a9",
  6800 => x"39811c78",
  6801 => x"08841a08",
  6802 => x"59557756",
  6803 => x"7d537e54",
  6804 => x"65525cfe",
  6805 => x"d8b73fa8",
  6806 => x"3d08aa3d",
  6807 => x"085f5df7",
  6808 => x"f8396252",
  6809 => x"6451ff85",
  6810 => x"e23f7c53",
  6811 => x"7d54a83d",
  6812 => x"08aa3d08",
  6813 => x"58517652",
  6814 => x"80d9ca3f",
  6815 => x"80083070",
  6816 => x"8008079f",
  6817 => x"2a647131",
  6818 => x"455156f3",
  6819 => x"9339800b",
  6820 => x"a13d0c80",
  6821 => x"692583f7",
  6822 => x"386869a5",
  6823 => x"3d0c6947",
  6824 => x"5cf69739",
  6825 => x"925c8049",
  6826 => x"f6903979",
  6827 => x"8f0682c9",
  6828 => x"980882c9",
  6829 => x"9c085955",
  6830 => x"77567853",
  6831 => x"79546552",
  6832 => x"5afef4d8",
  6833 => x"3fa83d08",
  6834 => x"aa3d0871",
  6835 => x"bb3d0c70",
  6836 => x"bc3d0c5a",
  6837 => x"58835cf6",
  6838 => x"ef39b83d",
  6839 => x"08ba3d08",
  6840 => x"71567057",
  6841 => x"58527653",
  6842 => x"6451fed4",
  6843 => x"da3fa83d",
  6844 => x"08aa3d08",
  6845 => x"71bb3d0c",
  6846 => x"70bc3d0c",
  6847 => x"7e557f56",
  6848 => x"71537054",
  6849 => x"5a5880da",
  6850 => x"a83f8008",
  6851 => x"80249a38",
  6852 => x"7c537d54",
  6853 => x"77517852",
  6854 => x"80d6be3f",
  6855 => x"8008b538",
  6856 => x"79810656",
  6857 => x"75802eac",
  6858 => x"38ff1f70",
  6859 => x"33575f75",
  6860 => x"b92e0981",
  6861 => x"0690387e",
  6862 => x"6d2e0981",
  6863 => x"06eb3862",
  6864 => x"810543b0",
  6865 => x"6d347e7f",
  6866 => x"81057133",
  6867 => x"81055840",
  6868 => x"57757734",
  6869 => x"60527f51",
  6870 => x"a9f73f80",
  6871 => x"7f3480c1",
  6872 => x"3d086381",
  6873 => x"05710c56",
  6874 => x"8c08802e",
  6875 => x"85387e8c",
  6876 => x"080c6c80",
  6877 => x"0cba3d0d",
  6878 => x"8c0c0462",
  6879 => x"305b7a80",
  6880 => x"2ef68638",
  6881 => x"7a832b80",
  6882 => x"f80682c9",
  6883 => x"a4110882",
  6884 => x"c9a01208",
  6885 => x"56567853",
  6886 => x"79546552",
  6887 => x"56fed5ed",
  6888 => x"3fa83d08",
  6889 => x"aa3d0871",
  6890 => x"bb3d0c70",
  6891 => x"bc3d0c7c",
  6892 => x"842c5c5a",
  6893 => x"5879802e",
  6894 => x"f5cf3882",
  6895 => x"c8f87a81",
  6896 => x"06575b75",
  6897 => x"81db3879",
  6898 => x"812c881c",
  6899 => x"5c5a7980",
  6900 => x"2ef5b638",
  6901 => x"79810656",
  6902 => x"75802eeb",
  6903 => x"3881c239",
  6904 => x"9f820a56",
  6905 => x"80765555",
  6906 => x"77527853",
  6907 => x"7a51fed2",
  6908 => x"d63fb03d",
  6909 => x"08b23d08",
  6910 => x"5ab73d0c",
  6911 => x"78b83d0c",
  6912 => x"b63d0890",
  6913 => x"ff0a05b7",
  6914 => x"3d0cf7cd",
  6915 => x"1c5c814e",
  6916 => x"eec53975",
  6917 => x"79065675",
  6918 => x"802efab0",
  6919 => x"38807048",
  6920 => x"4a696624",
  6921 => x"81de3880",
  6922 => x"d0820a56",
  6923 => x"80765555",
  6924 => x"7c527d53",
  6925 => x"6451fed4",
  6926 => x"d43fa83d",
  6927 => x"08aa3d08",
  6928 => x"58537654",
  6929 => x"b83d08ba",
  6930 => x"3d085851",
  6931 => x"765280db",
  6932 => x"b83f6980",
  6933 => x"082581ac",
  6934 => x"386c5fb1",
  6935 => x"7f708105",
  6936 => x"41346281",
  6937 => x"05436652",
  6938 => x"7f51a7e5",
  6939 => x"3f69802e",
  6940 => x"fde23867",
  6941 => x"30706907",
  6942 => x"9f2a5156",
  6943 => x"676a2e85",
  6944 => x"387580d1",
  6945 => x"3869527f",
  6946 => x"51a7c63f",
  6947 => x"fdc63981",
  6948 => x"7071a63d",
  6949 => x"0c71485d",
  6950 => x"49f29f39",
  6951 => x"815af48a",
  6952 => x"39811c7b",
  6953 => x"08841d08",
  6954 => x"59557756",
  6955 => x"78537954",
  6956 => x"65525cfe",
  6957 => x"d3d73fa8",
  6958 => x"3d08aa3d",
  6959 => x"0871bb3d",
  6960 => x"0c70bc3d",
  6961 => x"0c7b812c",
  6962 => x"881e5e5c",
  6963 => x"5a5879fe",
  6964 => x"8338f3b5",
  6965 => x"3967527f",
  6966 => x"51a6f63f",
  6967 => x"69527f51",
  6968 => x"a6ef3ffc",
  6969 => x"ef397781",
  6970 => x"0a325378",
  6971 => x"5479517a",
  6972 => x"5280d8a9",
  6973 => x"3f800880",
  6974 => x"25f7fb38",
  6975 => x"79b93d0c",
  6976 => x"7aba3d0c",
  6977 => x"680943fe",
  6978 => x"dd396aa6",
  6979 => x"3d087879",
  6980 => x"4b4c5959",
  6981 => x"6f802e80",
  6982 => x"c3388162",
  6983 => x"258bb938",
  6984 => x"65ff05a6",
  6985 => x"3d087131",
  6986 => x"595aa53d",
  6987 => x"087a2594",
  6988 => x"3879a63d",
  6989 => x"08316f11",
  6990 => x"a13d0ca6",
  6991 => x"3d0805a6",
  6992 => x"3d0c7658",
  6993 => x"655c8066",
  6994 => x"2483be38",
  6995 => x"6a1c641d",
  6996 => x"454b8152",
  6997 => x"7f51aaed",
  6998 => x"3f80084a",
  6999 => x"78802456",
  7000 => x"8064259b",
  7001 => x"3875802e",
  7002 => x"9638635c",
  7003 => x"78642583",
  7004 => x"38785c6a",
  7005 => x"7c31797d",
  7006 => x"31657e31",
  7007 => x"465a4b80",
  7008 => x"0ba63d08",
  7009 => x"25b8386f",
  7010 => x"802e889d",
  7011 => x"38807825",
  7012 => x"a3387753",
  7013 => x"69527f51",
  7014 => x"ad8d3f80",
  7015 => x"08615480",
  7016 => x"08536052",
  7017 => x"4aaab93f",
  7018 => x"80086153",
  7019 => x"605256a5",
  7020 => x"a03f7541",
  7021 => x"a53d0878",
  7022 => x"315a7982",
  7023 => x"bd388152",
  7024 => x"7f51aa81",
  7025 => x"3f800847",
  7026 => x"806f258e",
  7027 => x"386e5380",
  7028 => x"08527f51",
  7029 => x"acd13f80",
  7030 => x"08478058",
  7031 => x"81622581",
  7032 => x"d6386381",
  7033 => x"059f065c",
  7034 => x"6e81b238",
  7035 => x"7b802e85",
  7036 => x"38a07c31",
  7037 => x"5c847c25",
  7038 => x"86c438fc",
  7039 => x"1c6b1171",
  7040 => x"1b5b4c64",
  7041 => x"0544806b",
  7042 => x"258d386a",
  7043 => x"5360527f",
  7044 => x"51add43f",
  7045 => x"80084180",
  7046 => x"64258d38",
  7047 => x"63536652",
  7048 => x"7f51adc3",
  7049 => x"3f800847",
  7050 => x"a13d0880",
  7051 => x"c5388066",
  7052 => x"25568262",
  7053 => x"2581ff38",
  7054 => x"75802e81",
  7055 => x"f9388066",
  7056 => x"24fdc138",
  7057 => x"80548553",
  7058 => x"66527f51",
  7059 => x"a4a53f80",
  7060 => x"08800853",
  7061 => x"615247ae",
  7062 => x"d23f800b",
  7063 => x"800825fd",
  7064 => x"a3386c5f",
  7065 => x"b17f7081",
  7066 => x"05413462",
  7067 => x"810543fb",
  7068 => x"f5396652",
  7069 => x"6051aeb3",
  7070 => x"3f800880",
  7071 => x"25ffaf38",
  7072 => x"62ff0543",
  7073 => x"80548a53",
  7074 => x"60527f51",
  7075 => x"a3e53f80",
  7076 => x"08416f81",
  7077 => x"8c38a33d",
  7078 => x"0846ff92",
  7079 => x"39669005",
  7080 => x"08101067",
  7081 => x"05901108",
  7082 => x"5256a686",
  7083 => x"3f638008",
  7084 => x"319f065c",
  7085 => x"feb639b9",
  7086 => x"3d08782e",
  7087 => x"098106fe",
  7088 => x"a138b83d",
  7089 => x"0870bfff",
  7090 => x"ff065757",
  7091 => x"75782e09",
  7092 => x"8106fe8e",
  7093 => x"38769ffe",
  7094 => x"0a065675",
  7095 => x"782efe82",
  7096 => x"386a8105",
  7097 => x"64810545",
  7098 => x"4b816481",
  7099 => x"059f065d",
  7100 => x"586e802e",
  7101 => x"fdf638ff",
  7102 => x"a4397953",
  7103 => x"60527f51",
  7104 => x"aaa53f80",
  7105 => x"0841fdb6",
  7106 => x"396a6631",
  7107 => x"59806b11",
  7108 => x"4c640544",
  7109 => x"81527f51",
  7110 => x"a7ab3f80",
  7111 => x"084afcbc",
  7112 => x"3980548a",
  7113 => x"5369527f",
  7114 => x"51a2c83f",
  7115 => x"8008a43d",
  7116 => x"08474afd",
  7117 => x"f939815c",
  7118 => x"6f802e81",
  7119 => x"ef388079",
  7120 => x"258d3878",
  7121 => x"5369527f",
  7122 => x"51ab9c3f",
  7123 => x"80084a69",
  7124 => x"48778294",
  7125 => x"38815c66",
  7126 => x"526051e2",
  7127 => x"a13f8008",
  7128 => x"b0056853",
  7129 => x"615257ac",
  7130 => x"c23f8008",
  7131 => x"6a546753",
  7132 => x"60525aad",
  7133 => x"8d3f8008",
  7134 => x"56815b80",
  7135 => x"088c0508",
  7136 => x"802e81d6",
  7137 => x"3875527f",
  7138 => x"51a1c63f",
  7139 => x"7a620756",
  7140 => x"758d38b9",
  7141 => x"3d088106",
  7142 => x"5675802e",
  7143 => x"81fe3880",
  7144 => x"7a24828c",
  7145 => x"38796207",
  7146 => x"56758d38",
  7147 => x"b93d0881",
  7148 => x"06567580",
  7149 => x"2e81f938",
  7150 => x"7a802486",
  7151 => x"bc38767f",
  7152 => x"70810541",
  7153 => x"347b662e",
  7154 => x"83883880",
  7155 => x"548a5360",
  7156 => x"527f51a1",
  7157 => x"9e3f8008",
  7158 => x"41676a2e",
  7159 => x"82c93880",
  7160 => x"548a5367",
  7161 => x"527f51a1",
  7162 => x"8a3f8008",
  7163 => x"4880548a",
  7164 => x"5369527f",
  7165 => x"51a0fc3f",
  7166 => x"8008811d",
  7167 => x"5d4a6652",
  7168 => x"6051e0fa",
  7169 => x"3f8008b0",
  7170 => x"05685361",
  7171 => x"5257ab9b",
  7172 => x"3f80086a",
  7173 => x"54675360",
  7174 => x"525aabe6",
  7175 => x"3f800856",
  7176 => x"815b8008",
  7177 => x"8c0508fe",
  7178 => x"dc38af39",
  7179 => x"66527e7f",
  7180 => x"81056253",
  7181 => x"4056e0c6",
  7182 => x"3f8008b0",
  7183 => x"05577676",
  7184 => x"347b6625",
  7185 => x"828c3880",
  7186 => x"548a5360",
  7187 => x"527f51a0",
  7188 => x"a23f8008",
  7189 => x"811d5d41",
  7190 => x"d3398008",
  7191 => x"526051aa",
  7192 => x"ca3f8008",
  7193 => x"5bfe9e39",
  7194 => x"69840508",
  7195 => x"527f519e",
  7196 => x"d63f8008",
  7197 => x"68900508",
  7198 => x"10108805",
  7199 => x"54688c05",
  7200 => x"5380088c",
  7201 => x"05524aff",
  7202 => x"a6e33f81",
  7203 => x"5369527f",
  7204 => x"51a8d43f",
  7205 => x"80084a81",
  7206 => x"5cfdbc39",
  7207 => x"76b92ebb",
  7208 => x"38798024",
  7209 => x"1757767f",
  7210 => x"70810541",
  7211 => x"34f7b739",
  7212 => x"807b25f2",
  7213 => x"38815360",
  7214 => x"527f51a8",
  7215 => x"aa3f8008",
  7216 => x"67538008",
  7217 => x"5241a9e3",
  7218 => x"3f800b80",
  7219 => x"0825ba38",
  7220 => x"81175776",
  7221 => x"ba2e0981",
  7222 => x"06cc38b9",
  7223 => x"7f708105",
  7224 => x"4134ff1f",
  7225 => x"7033575f",
  7226 => x"75b92e09",
  7227 => x"8106819a",
  7228 => x"387e6d2e",
  7229 => x"098106ea",
  7230 => x"38628105",
  7231 => x"6d4043b1",
  7232 => x"7f708105",
  7233 => x"4134f6de",
  7234 => x"398008ff",
  7235 => x"99387681",
  7236 => x"06567580",
  7237 => x"2eff8f38",
  7238 => x"81175776",
  7239 => x"ba2e0981",
  7240 => x"06ff8338",
  7241 => x"ffb53980",
  7242 => x"548a5369",
  7243 => x"527f519e",
  7244 => x"c23f8008",
  7245 => x"8008811e",
  7246 => x"5e494afd",
  7247 => x"c1397b83",
  7248 => x"24f9c338",
  7249 => x"9c1c6b11",
  7250 => x"711b5b4c",
  7251 => x"640544f9",
  7252 => x"b5398153",
  7253 => x"60527f51",
  7254 => x"a78d3f80",
  7255 => x"08675380",
  7256 => x"085241a8",
  7257 => x"c63f8008",
  7258 => x"8024fef6",
  7259 => x"38800889",
  7260 => x"38768106",
  7261 => x"5675feea",
  7262 => x"38ff1f70",
  7263 => x"33575f75",
  7264 => x"b02ef638",
  7265 => x"811f5ff5",
  7266 => x"dd397e7f",
  7267 => x"81057133",
  7268 => x"81055840",
  7269 => x"57757734",
  7270 => x"f5cc396a",
  7271 => x"63316330",
  7272 => x"a73d0c4b",
  7273 => x"804fe5d2",
  7274 => x"39a53d08",
  7275 => x"5360527f",
  7276 => x"51a4f43f",
  7277 => x"800841f8",
  7278 => x"85396510",
  7279 => x"101082c9",
  7280 => x"98058411",
  7281 => x"08710856",
  7282 => x"56b53d08",
  7283 => x"b73d0859",
  7284 => x"53567653",
  7285 => x"6451fec9",
  7286 => x"b43fa83d",
  7287 => x"08aa3d08",
  7288 => x"58b53d0c",
  7289 => x"76b63d0c",
  7290 => x"810bb93d",
  7291 => x"08bb3d08",
  7292 => x"5b595c77",
  7293 => x"51785280",
  7294 => x"d1fb3f80",
  7295 => x"08800853",
  7296 => x"65525afe",
  7297 => x"f6c53fa8",
  7298 => x"3d08aa3d",
  7299 => x"08585476",
  7300 => x"55b83d08",
  7301 => x"ba3d0858",
  7302 => x"5276536b",
  7303 => x"51fec7c4",
  7304 => x"3faa3d08",
  7305 => x"ac3d085a",
  7306 => x"b93d0c78",
  7307 => x"ba3d0cb0",
  7308 => x"1a56757f",
  7309 => x"70810541",
  7310 => x"347b662e",
  7311 => x"eccb3881",
  7312 => x"1c5c80c8",
  7313 => x"820a5680",
  7314 => x"765555b8",
  7315 => x"3d08ba3d",
  7316 => x"08585276",
  7317 => x"536451fe",
  7318 => x"c8b33fa8",
  7319 => x"3d08aa3d",
  7320 => x"0871bb3d",
  7321 => x"0c70bc3d",
  7322 => x"0c5a58ff",
  7323 => x"8639ff1f",
  7324 => x"7033575f",
  7325 => x"75b02ef6",
  7326 => x"38811f5f",
  7327 => x"f1d63965",
  7328 => x"66484a80",
  7329 => x"d0820a56",
  7330 => x"80765555",
  7331 => x"b83d08ba",
  7332 => x"3d085852",
  7333 => x"76536451",
  7334 => x"fec6c93f",
  7335 => x"a83d08aa",
  7336 => x"3d08b63d",
  7337 => x"08b83d08",
  7338 => x"71577058",
  7339 => x"73557256",
  7340 => x"5c5a5c5a",
  7341 => x"80cafa3f",
  7342 => x"800b8008",
  7343 => x"25f4a738",
  7344 => x"79b93d0c",
  7345 => x"7aba3d0c",
  7346 => x"6c5fb17f",
  7347 => x"70810541",
  7348 => x"34628105",
  7349 => x"43f38f39",
  7350 => x"88b3165c",
  7351 => x"6df4ed38",
  7352 => x"b60ba83d",
  7353 => x"08316b11",
  7354 => x"4c640544",
  7355 => x"81527f51",
  7356 => x"9fd33f80",
  7357 => x"084af4e4",
  7358 => x"3976b92e",
  7359 => x"fbdd3881",
  7360 => x"1756757f",
  7361 => x"70810541",
  7362 => x"34f2db39",
  7363 => x"f83d0d7a",
  7364 => x"5877802e",
  7365 => x"81993882",
  7366 => x"d4800854",
  7367 => x"b8140880",
  7368 => x"2e80ed38",
  7369 => x"8c182270",
  7370 => x"902b7090",
  7371 => x"2c70832a",
  7372 => x"81328106",
  7373 => x"5c515754",
  7374 => x"7880cd38",
  7375 => x"90180857",
  7376 => x"76802e80",
  7377 => x"c3387708",
  7378 => x"77317779",
  7379 => x"0c768306",
  7380 => x"7a585555",
  7381 => x"73853894",
  7382 => x"18085675",
  7383 => x"88190c80",
  7384 => x"7525a538",
  7385 => x"74537652",
  7386 => x"9c180851",
  7387 => x"a4180854",
  7388 => x"732d800b",
  7389 => x"80082580",
  7390 => x"ca388008",
  7391 => x"17758008",
  7392 => x"31565774",
  7393 => x"8024dd38",
  7394 => x"800b800c",
  7395 => x"8a3d0d04",
  7396 => x"735181dc",
  7397 => x"3f8c1822",
  7398 => x"70902b70",
  7399 => x"902c7083",
  7400 => x"2a813281",
  7401 => x"065c5157",
  7402 => x"5478dd38",
  7403 => x"ff8e3981",
  7404 => x"e68c5282",
  7405 => x"d4800851",
  7406 => x"8fe53f80",
  7407 => x"08800c8a",
  7408 => x"3d0d048c",
  7409 => x"182280c0",
  7410 => x"0754738c",
  7411 => x"1923ff0b",
  7412 => x"800c8a3d",
  7413 => x"0d04803d",
  7414 => x"0d725180",
  7415 => x"710c800b",
  7416 => x"84120c80",
  7417 => x"0b88120c",
  7418 => x"028e0522",
  7419 => x"8c122302",
  7420 => x"9205228e",
  7421 => x"1223800b",
  7422 => x"90120c80",
  7423 => x"0b94120c",
  7424 => x"800b9812",
  7425 => x"0c709c12",
  7426 => x"0c829dc0",
  7427 => x"0ba0120c",
  7428 => x"829e8c0b",
  7429 => x"a4120c82",
  7430 => x"9f880ba8",
  7431 => x"120c829f",
  7432 => x"d90bac12",
  7433 => x"0c823d0d",
  7434 => x"04fa3d0d",
  7435 => x"797080dc",
  7436 => x"298c1154",
  7437 => x"7a535657",
  7438 => x"ff93bb3f",
  7439 => x"80088008",
  7440 => x"55568008",
  7441 => x"802ea238",
  7442 => x"80088c05",
  7443 => x"54800b80",
  7444 => x"080c7680",
  7445 => x"0884050c",
  7446 => x"73800888",
  7447 => x"050c7453",
  7448 => x"80527351",
  7449 => x"95d23f75",
  7450 => x"5473800c",
  7451 => x"883d0d04",
  7452 => x"fc3d0d76",
  7453 => x"81eb840b",
  7454 => x"bc120c55",
  7455 => x"810bb816",
  7456 => x"0c800b84",
  7457 => x"dc160c83",
  7458 => x"0b84e016",
  7459 => x"0c84e815",
  7460 => x"84e4160c",
  7461 => x"74548053",
  7462 => x"84528415",
  7463 => x"0851feb6",
  7464 => x"3f745481",
  7465 => x"53895288",
  7466 => x"150851fe",
  7467 => x"a93f7454",
  7468 => x"82538a52",
  7469 => x"8c150851",
  7470 => x"fe9c3f86",
  7471 => x"3d0d04f9",
  7472 => x"3d0d7982",
  7473 => x"d4800854",
  7474 => x"57b81308",
  7475 => x"802e80c8",
  7476 => x"3884dc13",
  7477 => x"56881608",
  7478 => x"841708ff",
  7479 => x"05555580",
  7480 => x"74249f38",
  7481 => x"8c152270",
  7482 => x"902b7090",
  7483 => x"2c515458",
  7484 => x"72802e80",
  7485 => x"ca3880dc",
  7486 => x"15ff1555",
  7487 => x"55738025",
  7488 => x"e3387508",
  7489 => x"5372802e",
  7490 => x"9f387256",
  7491 => x"88160884",
  7492 => x"1708ff05",
  7493 => x"5555c839",
  7494 => x"7251fed4",
  7495 => x"3f82d480",
  7496 => x"0884dc05",
  7497 => x"56ffae39",
  7498 => x"84527651",
  7499 => x"fdfb3f80",
  7500 => x"08760c80",
  7501 => x"08802e80",
  7502 => x"c0388008",
  7503 => x"56ce3981",
  7504 => x"0b8c1623",
  7505 => x"72750c72",
  7506 => x"88160c72",
  7507 => x"84160c72",
  7508 => x"90160c72",
  7509 => x"94160c72",
  7510 => x"98160cff",
  7511 => x"0b8e1623",
  7512 => x"72b0160c",
  7513 => x"72b4160c",
  7514 => x"7280c416",
  7515 => x"0c7280c8",
  7516 => x"160c7480",
  7517 => x"0c893d0d",
  7518 => x"048c770c",
  7519 => x"800b800c",
  7520 => x"893d0d04",
  7521 => x"ff3d0d81",
  7522 => x"e68c5273",
  7523 => x"518c903f",
  7524 => x"833d0d04",
  7525 => x"803d0d82",
  7526 => x"d4800851",
  7527 => x"e73f823d",
  7528 => x"0d04fb3d",
  7529 => x"0d777052",
  7530 => x"56ff9dda",
  7531 => x"3f82cbf8",
  7532 => x"0b880508",
  7533 => x"841108fc",
  7534 => x"06707b31",
  7535 => x"9fef05e0",
  7536 => x"8006e080",
  7537 => x"05565653",
  7538 => x"a0807424",
  7539 => x"95388052",
  7540 => x"7551ff9d",
  7541 => x"e93f82cc",
  7542 => x"80081553",
  7543 => x"7280082e",
  7544 => x"90387551",
  7545 => x"ff9da03f",
  7546 => x"80537280",
  7547 => x"0c873d0d",
  7548 => x"04733052",
  7549 => x"7551ff9d",
  7550 => x"c53f8008",
  7551 => x"ff2ea938",
  7552 => x"82cbf80b",
  7553 => x"88050875",
  7554 => x"75318107",
  7555 => x"84120c53",
  7556 => x"82cbbc08",
  7557 => x"743182cb",
  7558 => x"bc0c7551",
  7559 => x"ff9ce83f",
  7560 => x"810b800c",
  7561 => x"873d0d04",
  7562 => x"80527551",
  7563 => x"ff9d8f3f",
  7564 => x"82cbf80b",
  7565 => x"88050880",
  7566 => x"08713156",
  7567 => x"538f7525",
  7568 => x"ffa03880",
  7569 => x"0882cbec",
  7570 => x"083182cb",
  7571 => x"bc0c7481",
  7572 => x"0784140c",
  7573 => x"7551ff9c",
  7574 => x"ae3f8053",
  7575 => x"ff8c39f6",
  7576 => x"3d0d7c7e",
  7577 => x"545b7280",
  7578 => x"2e828538",
  7579 => x"7a51ff9c",
  7580 => x"953ff813",
  7581 => x"84110870",
  7582 => x"fe067013",
  7583 => x"841108fc",
  7584 => x"065d5859",
  7585 => x"545882cc",
  7586 => x"8008752e",
  7587 => x"82df3878",
  7588 => x"84160c80",
  7589 => x"73810654",
  7590 => x"5a727a2e",
  7591 => x"81d63878",
  7592 => x"15841108",
  7593 => x"81065153",
  7594 => x"72a03878",
  7595 => x"17577981",
  7596 => x"e7388815",
  7597 => x"08537282",
  7598 => x"cc802e82",
  7599 => x"fb388c15",
  7600 => x"08708c15",
  7601 => x"0c738812",
  7602 => x"0c567681",
  7603 => x"0784190c",
  7604 => x"76187771",
  7605 => x"0c537981",
  7606 => x"913883ff",
  7607 => x"772781c9",
  7608 => x"3876892a",
  7609 => x"77832a56",
  7610 => x"5372802e",
  7611 => x"bf387686",
  7612 => x"2ab80555",
  7613 => x"847327b4",
  7614 => x"3880db13",
  7615 => x"55947327",
  7616 => x"ab38768c",
  7617 => x"2a80ee05",
  7618 => x"5580d473",
  7619 => x"279e3876",
  7620 => x"8f2a80f7",
  7621 => x"055582d4",
  7622 => x"73279138",
  7623 => x"76922a80",
  7624 => x"fc05558a",
  7625 => x"d4732784",
  7626 => x"3880fe55",
  7627 => x"74101010",
  7628 => x"82cbf805",
  7629 => x"88110855",
  7630 => x"5673762e",
  7631 => x"82b53884",
  7632 => x"1408fc06",
  7633 => x"53767327",
  7634 => x"8d388814",
  7635 => x"08547376",
  7636 => x"2e098106",
  7637 => x"ea388c14",
  7638 => x"08708c1a",
  7639 => x"0c74881a",
  7640 => x"0c788812",
  7641 => x"0c56778c",
  7642 => x"150c7a51",
  7643 => x"ff9a983f",
  7644 => x"8c3d0d04",
  7645 => x"77087871",
  7646 => x"31597705",
  7647 => x"88190854",
  7648 => x"577282cc",
  7649 => x"802e80e0",
  7650 => x"388c1808",
  7651 => x"708c150c",
  7652 => x"7388120c",
  7653 => x"56fe8839",
  7654 => x"8815088c",
  7655 => x"1608708c",
  7656 => x"130c5788",
  7657 => x"170cfea2",
  7658 => x"3976832a",
  7659 => x"70545580",
  7660 => x"75248199",
  7661 => x"3872822c",
  7662 => x"81712b82",
  7663 => x"cbfc0807",
  7664 => x"82cbf80b",
  7665 => x"84050c53",
  7666 => x"74101010",
  7667 => x"82cbf805",
  7668 => x"88110855",
  7669 => x"56758c19",
  7670 => x"0c738819",
  7671 => x"0c778817",
  7672 => x"0c778c15",
  7673 => x"0cff8339",
  7674 => x"815afdb3",
  7675 => x"39781773",
  7676 => x"81065457",
  7677 => x"72983877",
  7678 => x"08787131",
  7679 => x"5977058c",
  7680 => x"1908881a",
  7681 => x"08718c12",
  7682 => x"0c88120c",
  7683 => x"57577681",
  7684 => x"0784190c",
  7685 => x"7782cbf8",
  7686 => x"0b88050c",
  7687 => x"82cbf408",
  7688 => x"7726fec6",
  7689 => x"3882cbf0",
  7690 => x"08527a51",
  7691 => x"faf43f7a",
  7692 => x"51ff98d3",
  7693 => x"3ffeb939",
  7694 => x"81788c15",
  7695 => x"0c788815",
  7696 => x"0c738c1a",
  7697 => x"0c73881a",
  7698 => x"0c5afcfe",
  7699 => x"39831570",
  7700 => x"822c8171",
  7701 => x"2b82cbfc",
  7702 => x"080782cb",
  7703 => x"f80b8405",
  7704 => x"0c515374",
  7705 => x"10101082",
  7706 => x"cbf80588",
  7707 => x"11085556",
  7708 => x"fee33974",
  7709 => x"53807524",
  7710 => x"a7387282",
  7711 => x"2c81712b",
  7712 => x"82cbfc08",
  7713 => x"0782cbf8",
  7714 => x"0b84050c",
  7715 => x"53758c19",
  7716 => x"0c738819",
  7717 => x"0c778817",
  7718 => x"0c778c15",
  7719 => x"0cfdcb39",
  7720 => x"83157082",
  7721 => x"2c81712b",
  7722 => x"82cbfc08",
  7723 => x"0782cbf8",
  7724 => x"0b84050c",
  7725 => x"5153d639",
  7726 => x"f23d0d60",
  7727 => x"62881108",
  7728 => x"7057575f",
  7729 => x"5a74802e",
  7730 => x"8190388c",
  7731 => x"1a227083",
  7732 => x"2a813270",
  7733 => x"81065155",
  7734 => x"58738638",
  7735 => x"901a0891",
  7736 => x"387951cd",
  7737 => x"b53fff54",
  7738 => x"800880ee",
  7739 => x"388c1a22",
  7740 => x"587d0857",
  7741 => x"807883ff",
  7742 => x"ff06700a",
  7743 => x"100a7081",
  7744 => x"06515657",
  7745 => x"5573752e",
  7746 => x"80d73874",
  7747 => x"90387608",
  7748 => x"84180888",
  7749 => x"19595659",
  7750 => x"74802ef2",
  7751 => x"38745488",
  7752 => x"80752784",
  7753 => x"38888054",
  7754 => x"73537852",
  7755 => x"9c1a0851",
  7756 => x"a41a0854",
  7757 => x"732d800b",
  7758 => x"80082582",
  7759 => x"e6388008",
  7760 => x"19758008",
  7761 => x"317f8805",
  7762 => x"08800831",
  7763 => x"70618805",
  7764 => x"0c565659",
  7765 => x"73ffb438",
  7766 => x"80547380",
  7767 => x"0c903d0d",
  7768 => x"04758132",
  7769 => x"70810676",
  7770 => x"41515473",
  7771 => x"802e81c1",
  7772 => x"38749038",
  7773 => x"76088418",
  7774 => x"08881959",
  7775 => x"56597480",
  7776 => x"2ef23888",
  7777 => x"1a087883",
  7778 => x"ffff0670",
  7779 => x"892a7081",
  7780 => x"06515659",
  7781 => x"5673802e",
  7782 => x"82fa3875",
  7783 => x"75278d38",
  7784 => x"77872a70",
  7785 => x"81065154",
  7786 => x"7382b538",
  7787 => x"74762783",
  7788 => x"38745675",
  7789 => x"53785279",
  7790 => x"085189b9",
  7791 => x"3f881a08",
  7792 => x"7631881b",
  7793 => x"0c790816",
  7794 => x"7a0c7456",
  7795 => x"75197577",
  7796 => x"317f8805",
  7797 => x"08783170",
  7798 => x"6188050c",
  7799 => x"56565973",
  7800 => x"802efef4",
  7801 => x"388c1a22",
  7802 => x"58ff8639",
  7803 => x"77785479",
  7804 => x"537b5256",
  7805 => x"88ff3f88",
  7806 => x"1a087831",
  7807 => x"881b0c79",
  7808 => x"08187a0c",
  7809 => x"7c76315d",
  7810 => x"7c8e3879",
  7811 => x"51f1fd3f",
  7812 => x"8008818f",
  7813 => x"3880085f",
  7814 => x"75197577",
  7815 => x"317f8805",
  7816 => x"08783170",
  7817 => x"6188050c",
  7818 => x"56565973",
  7819 => x"802efea8",
  7820 => x"38748183",
  7821 => x"38760884",
  7822 => x"18088819",
  7823 => x"59565974",
  7824 => x"802ef238",
  7825 => x"74538a52",
  7826 => x"7851878a",
  7827 => x"3f800879",
  7828 => x"3181055d",
  7829 => x"80088438",
  7830 => x"81155d81",
  7831 => x"5f7c5874",
  7832 => x"7d278338",
  7833 => x"7458941a",
  7834 => x"08881b08",
  7835 => x"11575c80",
  7836 => x"7a085c54",
  7837 => x"901a087b",
  7838 => x"27833881",
  7839 => x"54757825",
  7840 => x"843873ba",
  7841 => x"387b7824",
  7842 => x"fee2387b",
  7843 => x"5378529c",
  7844 => x"1a0851a4",
  7845 => x"1a085473",
  7846 => x"2d800856",
  7847 => x"80088024",
  7848 => x"fee2388c",
  7849 => x"1a2280c0",
  7850 => x"0754738c",
  7851 => x"1b23ff54",
  7852 => x"73800c90",
  7853 => x"3d0d047e",
  7854 => x"ffa338ff",
  7855 => x"87397553",
  7856 => x"78527a51",
  7857 => x"87af3f79",
  7858 => x"08167a0c",
  7859 => x"7951f0bc",
  7860 => x"3f8008cf",
  7861 => x"387c7631",
  7862 => x"5d7cfebc",
  7863 => x"38feac39",
  7864 => x"901a087a",
  7865 => x"08713176",
  7866 => x"1170565a",
  7867 => x"575282d4",
  7868 => x"8008519e",
  7869 => x"e33f8008",
  7870 => x"802effa7",
  7871 => x"38800890",
  7872 => x"1b0c8008",
  7873 => x"167a0c77",
  7874 => x"941b0c74",
  7875 => x"881b0c74",
  7876 => x"56fd9939",
  7877 => x"79085890",
  7878 => x"1a087827",
  7879 => x"83388154",
  7880 => x"75752784",
  7881 => x"3873b338",
  7882 => x"941a0856",
  7883 => x"75752680",
  7884 => x"d3387553",
  7885 => x"78529c1a",
  7886 => x"0851a41a",
  7887 => x"0854732d",
  7888 => x"80085680",
  7889 => x"088024fd",
  7890 => x"83388c1a",
  7891 => x"2280c007",
  7892 => x"54738c1b",
  7893 => x"23ff54fe",
  7894 => x"d7397553",
  7895 => x"78527751",
  7896 => x"86933f79",
  7897 => x"08167a0c",
  7898 => x"7951efa0",
  7899 => x"3f800880",
  7900 => x"2efcd938",
  7901 => x"8c1a2280",
  7902 => x"c0075473",
  7903 => x"8c1b23ff",
  7904 => x"54fead39",
  7905 => x"74755479",
  7906 => x"53785256",
  7907 => x"85e73f88",
  7908 => x"1a087531",
  7909 => x"881b0c79",
  7910 => x"08157a0c",
  7911 => x"fcae39f9",
  7912 => x"3d0d797b",
  7913 => x"5853800b",
  7914 => x"82d48008",
  7915 => x"53567272",
  7916 => x"2e80c038",
  7917 => x"84dc1355",
  7918 => x"74762eb7",
  7919 => x"38881508",
  7920 => x"841608ff",
  7921 => x"05545480",
  7922 => x"73249d38",
  7923 => x"8c142270",
  7924 => x"902b7090",
  7925 => x"2c515358",
  7926 => x"7180d838",
  7927 => x"80dc14ff",
  7928 => x"14545472",
  7929 => x"8025e538",
  7930 => x"74085574",
  7931 => x"d03882d4",
  7932 => x"80085284",
  7933 => x"dc125574",
  7934 => x"802eb138",
  7935 => x"88150884",
  7936 => x"1608ff05",
  7937 => x"54548073",
  7938 => x"249c388c",
  7939 => x"14227090",
  7940 => x"2b70902c",
  7941 => x"51535871",
  7942 => x"ad3880dc",
  7943 => x"14ff1454",
  7944 => x"54728025",
  7945 => x"e6387408",
  7946 => x"5574d138",
  7947 => x"75800c89",
  7948 => x"3d0d0473",
  7949 => x"51762d75",
  7950 => x"80080780",
  7951 => x"dc15ff15",
  7952 => x"555556ff",
  7953 => x"9e397351",
  7954 => x"762d7580",
  7955 => x"080780dc",
  7956 => x"15ff1555",
  7957 => x"5556ca39",
  7958 => x"fc3d0d76",
  7959 => x"79555573",
  7960 => x"802e9638",
  7961 => x"82c89052",
  7962 => x"7351a78a",
  7963 => x"3f800894",
  7964 => x"3877b016",
  7965 => x"0c73b416",
  7966 => x"0c82c890",
  7967 => x"5372800c",
  7968 => x"863d0d04",
  7969 => x"82c7b452",
  7970 => x"7351a6ea",
  7971 => x"3f805380",
  7972 => x"08732e09",
  7973 => x"8106e638",
  7974 => x"77b0160c",
  7975 => x"73b4160c",
  7976 => x"d83982db",
  7977 => x"9c08800c",
  7978 => x"0482c8a0",
  7979 => x"0b800c04",
  7980 => x"fe3d0d75",
  7981 => x"53745282",
  7982 => x"d4800851",
  7983 => x"ff9a3f84",
  7984 => x"3d0d0480",
  7985 => x"3d0d82d4",
  7986 => x"800851dd",
  7987 => x"3f823d0d",
  7988 => x"04ea3d0d",
  7989 => x"688c1122",
  7990 => x"700a100a",
  7991 => x"81065758",
  7992 => x"567480e5",
  7993 => x"388e1622",
  7994 => x"70902b70",
  7995 => x"902c5155",
  7996 => x"58807424",
  7997 => x"b138983d",
  7998 => x"c4055373",
  7999 => x"5282d480",
  8000 => x"0851a9e3",
  8001 => x"3f800b80",
  8002 => x"08249738",
  8003 => x"7983e080",
  8004 => x"06547380",
  8005 => x"c0802e81",
  8006 => x"91387382",
  8007 => x"80802e81",
  8008 => x"93388c16",
  8009 => x"22577690",
  8010 => x"80075473",
  8011 => x"8c172388",
  8012 => x"805282d4",
  8013 => x"800851ff",
  8014 => x"81bc3f80",
  8015 => x"089d388c",
  8016 => x"16228207",
  8017 => x"54738c17",
  8018 => x"2380c316",
  8019 => x"70770c90",
  8020 => x"170c810b",
  8021 => x"94170c98",
  8022 => x"3d0d0482",
  8023 => x"d4800881",
  8024 => x"eb840bbc",
  8025 => x"120c548c",
  8026 => x"16228180",
  8027 => x"0754738c",
  8028 => x"17238008",
  8029 => x"760c8008",
  8030 => x"90170c88",
  8031 => x"800b9417",
  8032 => x"0c74802e",
  8033 => x"d2388e16",
  8034 => x"2270902b",
  8035 => x"70902c53",
  8036 => x"5558afea",
  8037 => x"3f800880",
  8038 => x"2effbc38",
  8039 => x"8c162281",
  8040 => x"0754738c",
  8041 => x"1723983d",
  8042 => x"0d04810b",
  8043 => x"8c172258",
  8044 => x"55fef339",
  8045 => x"a8160882",
  8046 => x"9f882e09",
  8047 => x"8106fee2",
  8048 => x"388c1622",
  8049 => x"88800754",
  8050 => x"738c1723",
  8051 => x"88800b80",
  8052 => x"cc170cfe",
  8053 => x"da39fa3d",
  8054 => x"0d7a7902",
  8055 => x"8805a705",
  8056 => x"33565253",
  8057 => x"8373278a",
  8058 => x"38708306",
  8059 => x"5271802e",
  8060 => x"a838ff13",
  8061 => x"5372ff2e",
  8062 => x"97387033",
  8063 => x"5273722e",
  8064 => x"91388111",
  8065 => x"ff145451",
  8066 => x"72ff2e09",
  8067 => x"8106eb38",
  8068 => x"80517080",
  8069 => x"0c883d0d",
  8070 => x"04707257",
  8071 => x"55835175",
  8072 => x"82802914",
  8073 => x"ff125256",
  8074 => x"708025f3",
  8075 => x"38837327",
  8076 => x"bf387408",
  8077 => x"76327009",
  8078 => x"f7fbfdff",
  8079 => x"120670f8",
  8080 => x"84828180",
  8081 => x"06515151",
  8082 => x"70802e99",
  8083 => x"38745180",
  8084 => x"52703357",
  8085 => x"73772eff",
  8086 => x"b9388111",
  8087 => x"81135351",
  8088 => x"837227ed",
  8089 => x"38fc1384",
  8090 => x"16565372",
  8091 => x"8326c338",
  8092 => x"7451fefe",
  8093 => x"39fa3d0d",
  8094 => x"787a7c72",
  8095 => x"72725757",
  8096 => x"57595656",
  8097 => x"747627b2",
  8098 => x"38761551",
  8099 => x"757127aa",
  8100 => x"38707717",
  8101 => x"ff145455",
  8102 => x"5371ff2e",
  8103 => x"9638ff14",
  8104 => x"ff145454",
  8105 => x"72337434",
  8106 => x"ff125271",
  8107 => x"ff2e0981",
  8108 => x"06ec3875",
  8109 => x"800c883d",
  8110 => x"0d04768f",
  8111 => x"269738ff",
  8112 => x"125271ff",
  8113 => x"2eed3872",
  8114 => x"70810554",
  8115 => x"33747081",
  8116 => x"055634eb",
  8117 => x"39747607",
  8118 => x"83065170",
  8119 => x"e2387575",
  8120 => x"54517270",
  8121 => x"84055408",
  8122 => x"71708405",
  8123 => x"530c7270",
  8124 => x"84055408",
  8125 => x"71708405",
  8126 => x"530c7270",
  8127 => x"84055408",
  8128 => x"71708405",
  8129 => x"530c7270",
  8130 => x"84055408",
  8131 => x"71708405",
  8132 => x"530cf012",
  8133 => x"52718f26",
  8134 => x"c9388372",
  8135 => x"27953872",
  8136 => x"70840554",
  8137 => x"08717084",
  8138 => x"05530cfc",
  8139 => x"12527183",
  8140 => x"26ed3870",
  8141 => x"54ff8839",
  8142 => x"fc3d0d76",
  8143 => x"7971028c",
  8144 => x"059f0533",
  8145 => x"57555355",
  8146 => x"8372278a",
  8147 => x"38748306",
  8148 => x"5170802e",
  8149 => x"a238ff12",
  8150 => x"5271ff2e",
  8151 => x"93387373",
  8152 => x"70810555",
  8153 => x"34ff1252",
  8154 => x"71ff2e09",
  8155 => x"8106ef38",
  8156 => x"74800c86",
  8157 => x"3d0d0474",
  8158 => x"74882b75",
  8159 => x"07707190",
  8160 => x"2b075154",
  8161 => x"518f7227",
  8162 => x"a5387271",
  8163 => x"70840553",
  8164 => x"0c727170",
  8165 => x"8405530c",
  8166 => x"72717084",
  8167 => x"05530c72",
  8168 => x"71708405",
  8169 => x"530cf012",
  8170 => x"52718f26",
  8171 => x"dd388372",
  8172 => x"27903872",
  8173 => x"71708405",
  8174 => x"530cfc12",
  8175 => x"52718326",
  8176 => x"f2387053",
  8177 => x"ff9039f9",
  8178 => x"3d0d797b",
  8179 => x"80cc1208",
  8180 => x"56585673",
  8181 => x"802ea538",
  8182 => x"76101014",
  8183 => x"70085555",
  8184 => x"73802eb5",
  8185 => x"38730875",
  8186 => x"0c800b90",
  8187 => x"150c800b",
  8188 => x"8c150c73",
  8189 => x"5574800c",
  8190 => x"893d0d04",
  8191 => x"90538452",
  8192 => x"7551a29e",
  8193 => x"3f800880",
  8194 => x"cc170c80",
  8195 => x"08558008",
  8196 => x"802ee238",
  8197 => x"800854c0",
  8198 => x"3981772b",
  8199 => x"70101094",
  8200 => x"05545881",
  8201 => x"527551a1",
  8202 => x"f93f8008",
  8203 => x"80085654",
  8204 => x"8008802e",
  8205 => x"c0387680",
  8206 => x"0884050c",
  8207 => x"77800888",
  8208 => x"050c800b",
  8209 => x"90150c80",
  8210 => x"0b8c150c",
  8211 => x"7355ffa5",
  8212 => x"39ff3d0d",
  8213 => x"74527180",
  8214 => x"2e953873",
  8215 => x"84130810",
  8216 => x"1080cc12",
  8217 => x"08057008",
  8218 => x"740c7371",
  8219 => x"0c515183",
  8220 => x"3d0d04f5",
  8221 => x"3d0d7d7f",
  8222 => x"61639013",
  8223 => x"0894145b",
  8224 => x"5d5b5c5c",
  8225 => x"5c805782",
  8226 => x"16227a71",
  8227 => x"29197722",
  8228 => x"7c712972",
  8229 => x"902a0570",
  8230 => x"902a7383",
  8231 => x"ffff0672",
  8232 => x"84808029",
  8233 => x"057b7084",
  8234 => x"055d0c81",
  8235 => x"1c5c5253",
  8236 => x"5a555578",
  8237 => x"7724d038",
  8238 => x"77802e96",
  8239 => x"3878881c",
  8240 => x"08259638",
  8241 => x"7810101b",
  8242 => x"7894120c",
  8243 => x"54811990",
  8244 => x"1c0c7a80",
  8245 => x"0c8d3d0d",
  8246 => x"04841b08",
  8247 => x"8105527b",
  8248 => x"51fde43f",
  8249 => x"8008901c",
  8250 => x"08101088",
  8251 => x"05548c1c",
  8252 => x"5380088c",
  8253 => x"055254ff",
  8254 => x"85f33f7a",
  8255 => x"527b51fe",
  8256 => x"d03f7379",
  8257 => x"10101179",
  8258 => x"94120c55",
  8259 => x"811a9012",
  8260 => x"0c5bffbe",
  8261 => x"39f63d0d",
  8262 => x"7c7e6062",
  8263 => x"5e5c5959",
  8264 => x"8952881b",
  8265 => x"51feda9e",
  8266 => x"3f800857",
  8267 => x"80568155",
  8268 => x"7477258c",
  8269 => x"38741081",
  8270 => x"17575576",
  8271 => x"7524f638",
  8272 => x"75527851",
  8273 => x"fd813f80",
  8274 => x"08618008",
  8275 => x"94050c56",
  8276 => x"810b8008",
  8277 => x"90050c89",
  8278 => x"57767a25",
  8279 => x"80cf3876",
  8280 => x"18587770",
  8281 => x"81055933",
  8282 => x"d005548a",
  8283 => x"53755278",
  8284 => x"51fe803f",
  8285 => x"80088118",
  8286 => x"58567977",
  8287 => x"24e43881",
  8288 => x"1858767b",
  8289 => x"25a0387a",
  8290 => x"77315777",
  8291 => x"70810559",
  8292 => x"33d00554",
  8293 => x"8a537552",
  8294 => x"7851fdd7",
  8295 => x"3f8008ff",
  8296 => x"18585676",
  8297 => x"e6387580",
  8298 => x"0c8c3d0d",
  8299 => x"048a1858",
  8300 => x"d139fe3d",
  8301 => x"0d745280",
  8302 => x"72fc8080",
  8303 => x"06525370",
  8304 => x"732e0981",
  8305 => x"06873890",
  8306 => x"72712b53",
  8307 => x"537181ff",
  8308 => x"0a065170",
  8309 => x"88388813",
  8310 => x"72882b53",
  8311 => x"53718f0a",
  8312 => x"06517088",
  8313 => x"38841372",
  8314 => x"842b5353",
  8315 => x"71830a06",
  8316 => x"51708838",
  8317 => x"82137282",
  8318 => x"2b535380",
  8319 => x"72249338",
  8320 => x"8113729e",
  8321 => x"2a708106",
  8322 => x"515253a0",
  8323 => x"5270802e",
  8324 => x"83387252",
  8325 => x"71800c84",
  8326 => x"3d0d04fc",
  8327 => x"3d0d7670",
  8328 => x"08708706",
  8329 => x"53535570",
  8330 => x"802eaa38",
  8331 => x"71810651",
  8332 => x"80537073",
  8333 => x"2e098106",
  8334 => x"9538710a",
  8335 => x"100a7081",
  8336 => x"06525370",
  8337 => x"802e80f0",
  8338 => x"3872750c",
  8339 => x"81537280",
  8340 => x"0c863d0d",
  8341 => x"04707283",
  8342 => x"ffff0652",
  8343 => x"5470802e",
  8344 => x"80cd3871",
  8345 => x"81ff0651",
  8346 => x"70883888",
  8347 => x"1472882a",
  8348 => x"5354718f",
  8349 => x"06517088",
  8350 => x"38841472",
  8351 => x"842a5354",
  8352 => x"71830651",
  8353 => x"70883882",
  8354 => x"1472822a",
  8355 => x"53547181",
  8356 => x"06517091",
  8357 => x"38811472",
  8358 => x"0a100a53",
  8359 => x"54a05371",
  8360 => x"802effaa",
  8361 => x"3871750c",
  8362 => x"73800c86",
  8363 => x"3d0d0490",
  8364 => x"72712a53",
  8365 => x"54ffac39",
  8366 => x"71822a75",
  8367 => x"0c820b80",
  8368 => x"0c863d0d",
  8369 => x"04ff3d0d",
  8370 => x"81527351",
  8371 => x"f9f93f74",
  8372 => x"80089405",
  8373 => x"0c810b80",
  8374 => x"0890050c",
  8375 => x"833d0d04",
  8376 => x"ee3d0d65",
  8377 => x"67901208",
  8378 => x"90120858",
  8379 => x"56575373",
  8380 => x"75258d38",
  8381 => x"72767177",
  8382 => x"90140859",
  8383 => x"57585442",
  8384 => x"74147088",
  8385 => x"15082484",
  8386 => x"15080553",
  8387 => x"65525ef9",
  8388 => x"b63f8008",
  8389 => x"80089405",
  8390 => x"7060822b",
  8391 => x"72114346",
  8392 => x"5941427f",
  8393 => x"7f278d38",
  8394 => x"80777084",
  8395 => x"05590c7e",
  8396 => x"7726f538",
  8397 => x"94137410",
  8398 => x"10119418",
  8399 => x"77101011",
  8400 => x"6341445d",
  8401 => x"5d5f7a61",
  8402 => x"2781b838",
  8403 => x"7a087083",
  8404 => x"ffff0659",
  8405 => x"5377802e",
  8406 => x"80c7387e",
  8407 => x"7d575780",
  8408 => x"5a767084",
  8409 => x"05580870",
  8410 => x"83ffff06",
  8411 => x"82182271",
  8412 => x"7b29057c",
  8413 => x"1173902a",
  8414 => x"7c297a22",
  8415 => x"5e7d0571",
  8416 => x"902a0570",
  8417 => x"902a5f59",
  8418 => x"51515454",
  8419 => x"74762372",
  8420 => x"82172384",
  8421 => x"16567b77",
  8422 => x"26c73879",
  8423 => x"760c7a08",
  8424 => x"5372902a",
  8425 => x"5877802e",
  8426 => x"80cd387e",
  8427 => x"7d575780",
  8428 => x"7d08705b",
  8429 => x"565a7670",
  8430 => x"84055808",
  8431 => x"7083ffff",
  8432 => x"06707a29",
  8433 => x"7b902a05",
  8434 => x"7c115151",
  8435 => x"54547276",
  8436 => x"23748217",
  8437 => x"23841674",
  8438 => x"902a7929",
  8439 => x"71088213",
  8440 => x"225d5b7b",
  8441 => x"0574902a",
  8442 => x"0570902a",
  8443 => x"5c56567b",
  8444 => x"7726c338",
  8445 => x"74760c84",
  8446 => x"1b841e5e",
  8447 => x"5b607b26",
  8448 => x"feca3862",
  8449 => x"60055680",
  8450 => x"7e259038",
  8451 => x"fc165675",
  8452 => x"088938ff",
  8453 => x"1e5e7d80",
  8454 => x"24f2387d",
  8455 => x"6290050c",
  8456 => x"61800c94",
  8457 => x"3d0d04f7",
  8458 => x"3d0d7b7d",
  8459 => x"7f708306",
  8460 => x"58585a5a",
  8461 => x"7480dd38",
  8462 => x"75822c56",
  8463 => x"75802eb6",
  8464 => x"3880c81a",
  8465 => x"08705657",
  8466 => x"76802e80",
  8467 => x"f8387581",
  8468 => x"065574a9",
  8469 => x"3875812c",
  8470 => x"5675802e",
  8471 => x"99387608",
  8472 => x"70595574",
  8473 => x"802e80c6",
  8474 => x"38745775",
  8475 => x"81065574",
  8476 => x"802ee238",
  8477 => x"88397880",
  8478 => x"0c8b3d0d",
  8479 => x"04765378",
  8480 => x"527951fc",
  8481 => x"db3f8008",
  8482 => x"79537a52",
  8483 => x"55f7c23f",
  8484 => x"7459c239",
  8485 => x"80547410",
  8486 => x"1082cae4",
  8487 => x"05700854",
  8488 => x"55785279",
  8489 => x"51f7cc3f",
  8490 => x"800859ff",
  8491 => x"8b397653",
  8492 => x"76527951",
  8493 => x"fcaa3f80",
  8494 => x"08770c80",
  8495 => x"08788008",
  8496 => x"0c57ffa7",
  8497 => x"3984f152",
  8498 => x"7951fbf9",
  8499 => x"3f800880",
  8500 => x"c81b0c80",
  8501 => x"08758008",
  8502 => x"0c768106",
  8503 => x"56577480",
  8504 => x"2efef238",
  8505 => x"ff9739f5",
  8506 => x"3d0d7d7f",
  8507 => x"6170852c",
  8508 => x"84130890",
  8509 => x"14081281",
  8510 => x"05881508",
  8511 => x"595e5959",
  8512 => x"5a5c5c72",
  8513 => x"79258c38",
  8514 => x"81157310",
  8515 => x"54557873",
  8516 => x"24f63874",
  8517 => x"527b51f5",
  8518 => x"ae3f8008",
  8519 => x"80089405",
  8520 => x"555a8076",
  8521 => x"25903875",
  8522 => x"53807470",
  8523 => x"8405560c",
  8524 => x"ff135372",
  8525 => x"f438941b",
  8526 => x"901c0810",
  8527 => x"1011799f",
  8528 => x"065a5853",
  8529 => x"77802ebf",
  8530 => x"38a07831",
  8531 => x"55805672",
  8532 => x"08782b76",
  8533 => x"07747084",
  8534 => x"05560c72",
  8535 => x"70840554",
  8536 => x"08752a56",
  8537 => x"767326e7",
  8538 => x"3875740c",
  8539 => x"75802e84",
  8540 => x"38811959",
  8541 => x"ff19901b",
  8542 => x"0c7a527b",
  8543 => x"51f5d23f",
  8544 => x"79800c8d",
  8545 => x"3d0d0472",
  8546 => x"70840554",
  8547 => x"08747084",
  8548 => x"05560c72",
  8549 => x"7727dd38",
  8550 => x"72708405",
  8551 => x"54087470",
  8552 => x"8405560c",
  8553 => x"767326df",
  8554 => x"38ca39fb",
  8555 => x"3d0d7779",
  8556 => x"90110890",
  8557 => x"13087131",
  8558 => x"70565455",
  8559 => x"575470ab",
  8560 => x"38941473",
  8561 => x"822b7111",
  8562 => x"71199405",
  8563 => x"52545255",
  8564 => x"fc12fc12",
  8565 => x"71087108",
  8566 => x"56565252",
  8567 => x"73732e09",
  8568 => x"81068f38",
  8569 => x"717526e8",
  8570 => x"38805271",
  8571 => x"800c873d",
  8572 => x"0d04ff51",
  8573 => x"72742683",
  8574 => x"38815170",
  8575 => x"800c873d",
  8576 => x"0d04f33d",
  8577 => x"0d7f6163",
  8578 => x"70557154",
  8579 => x"575456ff",
  8580 => x"9a3f8008",
  8581 => x"54800880",
  8582 => x"2e81c638",
  8583 => x"80547380",
  8584 => x"082481dc",
  8585 => x"38841308",
  8586 => x"527551f3",
  8587 => x"9a3f8008",
  8588 => x"7480088c",
  8589 => x"050c9014",
  8590 => x"08941571",
  8591 => x"10101194",
  8592 => x"19901a08",
  8593 => x"10101180",
  8594 => x"0894055d",
  8595 => x"415d415a",
  8596 => x"5c5d805a",
  8597 => x"77708405",
  8598 => x"59087083",
  8599 => x"ffff067a",
  8600 => x"7084055c",
  8601 => x"087083ff",
  8602 => x"ff067271",
  8603 => x"311e7490",
  8604 => x"2a73902a",
  8605 => x"3171902c",
  8606 => x"1170902c",
  8607 => x"41515551",
  8608 => x"56575754",
  8609 => x"73772372",
  8610 => x"82182384",
  8611 => x"17577b79",
  8612 => x"26c23877",
  8613 => x"7e27ac38",
  8614 => x"77708405",
  8615 => x"59087083",
  8616 => x"ffff067b",
  8617 => x"1170902c",
  8618 => x"73902a05",
  8619 => x"70902c5e",
  8620 => x"53515454",
  8621 => x"73772372",
  8622 => x"82182384",
  8623 => x"17577d78",
  8624 => x"26d638fc",
  8625 => x"17577608",
  8626 => x"8d38ff1b",
  8627 => x"fc18585b",
  8628 => x"7608802e",
  8629 => x"f5387a90",
  8630 => x"1e0c7c80",
  8631 => x"0c8f3d0d",
  8632 => x"04800852",
  8633 => x"7551f1df",
  8634 => x"3f80085d",
  8635 => x"810b8008",
  8636 => x"90050c73",
  8637 => x"80089405",
  8638 => x"0c7c800c",
  8639 => x"8f3d0d04",
  8640 => x"72755455",
  8641 => x"810b8414",
  8642 => x"08537652",
  8643 => x"54f1b83f",
  8644 => x"80087480",
  8645 => x"088c050c",
  8646 => x"90140894",
  8647 => x"15711010",
  8648 => x"11941990",
  8649 => x"1a081010",
  8650 => x"11800894",
  8651 => x"055d415d",
  8652 => x"415a5c5d",
  8653 => x"805afe9c",
  8654 => x"39fa3d0d",
  8655 => x"787a7c54",
  8656 => x"57725876",
  8657 => x"9ffe0a06",
  8658 => x"86bf0a05",
  8659 => x"53538072",
  8660 => x"25953871",
  8661 => x"54805573",
  8662 => x"7553730c",
  8663 => x"7184140c",
  8664 => x"72800c88",
  8665 => x"3d0d0471",
  8666 => x"3070942c",
  8667 => x"53519372",
  8668 => x"25a73880",
  8669 => x"54ec129f",
  8670 => x"71318171",
  8671 => x"2b515252",
  8672 => x"9e722583",
  8673 => x"38815170",
  8674 => x"55737553",
  8675 => x"730c7184",
  8676 => x"140c7280",
  8677 => x"0c883d0d",
  8678 => x"04a08080",
  8679 => x"722c5480",
  8680 => x"55ffb439",
  8681 => x"f63d0d7c",
  8682 => x"7e941190",
  8683 => x"12081010",
  8684 => x"11fc1170",
  8685 => x"0870575a",
  8686 => x"51575853",
  8687 => x"59f3f33f",
  8688 => x"80087fa0",
  8689 => x"0b800831",
  8690 => x"710c5353",
  8691 => x"8a0b8008",
  8692 => x"2580e838",
  8693 => x"80577376",
  8694 => x"26bd38f5",
  8695 => x"13537280",
  8696 => x"2e80c038",
  8697 => x"a0733175",
  8698 => x"742b7872",
  8699 => x"2a079ffc",
  8700 => x"0a075b58",
  8701 => x"80557574",
  8702 => x"278538fc",
  8703 => x"14085576",
  8704 => x"732b7579",
  8705 => x"2a075b79",
  8706 => x"7b54790c",
  8707 => x"72841a0c",
  8708 => x"78800c8c",
  8709 => x"3d0d04fc",
  8710 => x"147008f5",
  8711 => x"15555854",
  8712 => x"72c23874",
  8713 => x"9ffc0a07",
  8714 => x"5a765b79",
  8715 => x"7b54790c",
  8716 => x"72841a0c",
  8717 => x"78800c8c",
  8718 => x"3d0d048b",
  8719 => x"0b800831",
  8720 => x"75712a9f",
  8721 => x"fc0a075b",
  8722 => x"57805875",
  8723 => x"74278538",
  8724 => x"fc140858",
  8725 => x"95137571",
  8726 => x"2b79792a",
  8727 => x"075c5279",
  8728 => x"7b54790c",
  8729 => x"72841a0c",
  8730 => x"78800c8c",
  8731 => x"3d0d04f3",
  8732 => x"3d0d6264",
  8733 => x"6264575f",
  8734 => x"75405b59",
  8735 => x"81527f51",
  8736 => x"eec53f80",
  8737 => x"08800894",
  8738 => x"057e70bf",
  8739 => x"ffff0670",
  8740 => x"5f71fe0a",
  8741 => x"06704270",
  8742 => x"942a5b52",
  8743 => x"57555957",
  8744 => x"75802e87",
  8745 => x"38739080",
  8746 => x"0a075b7d",
  8747 => x"5372802e",
  8748 => x"80d63872",
  8749 => x"5c8f3df4",
  8750 => x"0551f2df",
  8751 => x"3f800855",
  8752 => x"8008802e",
  8753 => x"80ff38a0",
  8754 => x"0b800831",
  8755 => x"7b712b7d",
  8756 => x"07790c53",
  8757 => x"7a80082a",
  8758 => x"5b7a7084",
  8759 => x"1a0c7030",
  8760 => x"70720780",
  8761 => x"25827131",
  8762 => x"70901c0c",
  8763 => x"51515454",
  8764 => x"75802eaf",
  8765 => x"387416f7",
  8766 => x"cd05790c",
  8767 => x"b575317a",
  8768 => x"0c76800c",
  8769 => x"8f3d0d04",
  8770 => x"8f3df005",
  8771 => x"51f28c3f",
  8772 => x"7a780c81",
  8773 => x"0b90180c",
  8774 => x"810b8008",
  8775 => x"a0055653",
  8776 => x"75d338f7",
  8777 => x"ce15790c",
  8778 => x"72852b73",
  8779 => x"101019fc",
  8780 => x"11085354",
  8781 => x"54f0fb3f",
  8782 => x"73800831",
  8783 => x"7a0c7680",
  8784 => x"0c8f3d0d",
  8785 => x"047b780c",
  8786 => x"7a70841a",
  8787 => x"0c703070",
  8788 => x"72078025",
  8789 => x"82713170",
  8790 => x"901c0c51",
  8791 => x"515454ff",
  8792 => x"8f39f03d",
  8793 => x"0d626466",
  8794 => x"953de411",
  8795 => x"577256f8",
  8796 => x"05545858",
  8797 => x"58fcad3f",
  8798 => x"923de011",
  8799 => x"547653f0",
  8800 => x"0551fca0",
  8801 => x"3f901708",
  8802 => x"90170831",
  8803 => x"852b7b7b",
  8804 => x"31115156",
  8805 => x"807625ae",
  8806 => x"38759080",
  8807 => x"0a296005",
  8808 => x"407d7f58",
  8809 => x"5476557f",
  8810 => x"61585276",
  8811 => x"53923de8",
  8812 => x"0551feb6",
  8813 => x"e73f7b7d",
  8814 => x"58780c76",
  8815 => x"84190c77",
  8816 => x"800c923d",
  8817 => x"0d047530",
  8818 => x"7090800a",
  8819 => x"291f5f56",
  8820 => x"7d7f5854",
  8821 => x"76557f61",
  8822 => x"58527653",
  8823 => x"923de805",
  8824 => x"51feb6b8",
  8825 => x"3f7b7d58",
  8826 => x"780c7684",
  8827 => x"190c7780",
  8828 => x"0c923d0d",
  8829 => x"04f33d0d",
  8830 => x"7f61575c",
  8831 => x"9ffc0a57",
  8832 => x"80587597",
  8833 => x"249b3875",
  8834 => x"10101082",
  8835 => x"c9a00584",
  8836 => x"11087108",
  8837 => x"7e0c841e",
  8838 => x"0c7c800c",
  8839 => x"568f3d0d",
  8840 => x"04807625",
  8841 => x"a5388d3d",
  8842 => x"5b80c882",
  8843 => x"0a59805a",
  8844 => x"78547955",
  8845 => x"76527753",
  8846 => x"7a51fe98",
  8847 => x"d03f7c7e",
  8848 => x"ff185859",
  8849 => x"57758024",
  8850 => x"e738767c",
  8851 => x"0c77841d",
  8852 => x"0c7b800c",
  8853 => x"8f3d0d04",
  8854 => x"ef3d0d63",
  8855 => x"6567405d",
  8856 => x"427b802e",
  8857 => x"84ff3861",
  8858 => x"51fef49a",
  8859 => x"3ff81c70",
  8860 => x"84120870",
  8861 => x"fc067062",
  8862 => x"8b0570f8",
  8863 => x"06415945",
  8864 => x"5b5c4157",
  8865 => x"96742782",
  8866 => x"c438807b",
  8867 => x"247e7c26",
  8868 => x"07598054",
  8869 => x"78742e09",
  8870 => x"810682aa",
  8871 => x"38777b25",
  8872 => x"81fc3877",
  8873 => x"1782cbf8",
  8874 => x"0b880508",
  8875 => x"5e567c76",
  8876 => x"2e84c238",
  8877 => x"84160870",
  8878 => x"fe061784",
  8879 => x"11088106",
  8880 => x"51555573",
  8881 => x"828c3874",
  8882 => x"fc06597c",
  8883 => x"762e84e3",
  8884 => x"3877195f",
  8885 => x"7e7b2581",
  8886 => x"fe387981",
  8887 => x"06547382",
  8888 => x"c1387677",
  8889 => x"08318411",
  8890 => x"08fc0656",
  8891 => x"5a75802e",
  8892 => x"91387c76",
  8893 => x"2e84f138",
  8894 => x"74191859",
  8895 => x"787b2584",
  8896 => x"8f387980",
  8897 => x"2e829b38",
  8898 => x"7715567a",
  8899 => x"76248292",
  8900 => x"388c1a08",
  8901 => x"881b0871",
  8902 => x"8c120c88",
  8903 => x"120c5579",
  8904 => x"76595788",
  8905 => x"1761fc05",
  8906 => x"575975a4",
  8907 => x"2685f738",
  8908 => x"7b795555",
  8909 => x"93762780",
  8910 => x"c9387b70",
  8911 => x"84055d08",
  8912 => x"7c56790c",
  8913 => x"74708405",
  8914 => x"56088c18",
  8915 => x"0c901754",
  8916 => x"9b7627ae",
  8917 => x"38747084",
  8918 => x"05560874",
  8919 => x"0c747084",
  8920 => x"05560894",
  8921 => x"180c9817",
  8922 => x"54a37627",
  8923 => x"95387470",
  8924 => x"84055608",
  8925 => x"740c7470",
  8926 => x"84055608",
  8927 => x"9c180ca0",
  8928 => x"17547470",
  8929 => x"84055608",
  8930 => x"74708405",
  8931 => x"560c7470",
  8932 => x"84055608",
  8933 => x"74708405",
  8934 => x"560c7408",
  8935 => x"740c777b",
  8936 => x"3156758f",
  8937 => x"2680ca38",
  8938 => x"84170881",
  8939 => x"06780784",
  8940 => x"180c7717",
  8941 => x"84110881",
  8942 => x"0784120c",
  8943 => x"546151fe",
  8944 => x"f1c53f88",
  8945 => x"17547380",
  8946 => x"0c933d0d",
  8947 => x"04905bfd",
  8948 => x"b9397856",
  8949 => x"fe84398c",
  8950 => x"16088817",
  8951 => x"08718c12",
  8952 => x"0c88120c",
  8953 => x"557e707c",
  8954 => x"3157588f",
  8955 => x"7627ffb8",
  8956 => x"387a1784",
  8957 => x"18088106",
  8958 => x"7c078419",
  8959 => x"0c768107",
  8960 => x"84120c76",
  8961 => x"11841108",
  8962 => x"81078412",
  8963 => x"0c558805",
  8964 => x"526151d4",
  8965 => x"ca3f6151",
  8966 => x"fef0ec3f",
  8967 => x"881754ff",
  8968 => x"a5397d52",
  8969 => x"6151fee3",
  8970 => x"cd3f8008",
  8971 => x"59800880",
  8972 => x"2e81a338",
  8973 => x"8008f805",
  8974 => x"60840508",
  8975 => x"fe066105",
  8976 => x"55577674",
  8977 => x"2e83ec38",
  8978 => x"fc185675",
  8979 => x"a42681ac",
  8980 => x"387b8008",
  8981 => x"55559376",
  8982 => x"2780d838",
  8983 => x"74708405",
  8984 => x"56088008",
  8985 => x"70840580",
  8986 => x"0c0c8008",
  8987 => x"75708405",
  8988 => x"57087170",
  8989 => x"8405530c",
  8990 => x"549b7627",
  8991 => x"b6387470",
  8992 => x"84055608",
  8993 => x"74708405",
  8994 => x"560c7470",
  8995 => x"84055608",
  8996 => x"74708405",
  8997 => x"560ca376",
  8998 => x"27993874",
  8999 => x"70840556",
  9000 => x"08747084",
  9001 => x"05560c74",
  9002 => x"70840556",
  9003 => x"08747084",
  9004 => x"05560c74",
  9005 => x"70840556",
  9006 => x"08747084",
  9007 => x"05560c74",
  9008 => x"70840556",
  9009 => x"08747084",
  9010 => x"05560c74",
  9011 => x"08740c7b",
  9012 => x"526151d3",
  9013 => x"8a3f6151",
  9014 => x"feefac3f",
  9015 => x"78547380",
  9016 => x"0c933d0d",
  9017 => x"047d5261",
  9018 => x"51fee28a",
  9019 => x"3f800880",
  9020 => x"0c933d0d",
  9021 => x"04841608",
  9022 => x"55fbcc39",
  9023 => x"75537b52",
  9024 => x"800851fe",
  9025 => x"ede73f7b",
  9026 => x"526151d2",
  9027 => x"d23fc739",
  9028 => x"8c160888",
  9029 => x"1708718c",
  9030 => x"120c8812",
  9031 => x"0c558c1a",
  9032 => x"08881b08",
  9033 => x"718c120c",
  9034 => x"88120c55",
  9035 => x"79795957",
  9036 => x"fbf13977",
  9037 => x"19901c55",
  9038 => x"55737524",
  9039 => x"fb9c387a",
  9040 => x"177082cb",
  9041 => x"f80b8805",
  9042 => x"0c757c31",
  9043 => x"81078412",
  9044 => x"0c5d8417",
  9045 => x"0881067b",
  9046 => x"0784180c",
  9047 => x"6151feee",
  9048 => x"a63f8817",
  9049 => x"54fcdf39",
  9050 => x"74191890",
  9051 => x"1c555d73",
  9052 => x"7d24fb8e",
  9053 => x"388c1a08",
  9054 => x"881b0871",
  9055 => x"8c120c88",
  9056 => x"120c5588",
  9057 => x"1a61fc05",
  9058 => x"575975a4",
  9059 => x"2681b038",
  9060 => x"7b795555",
  9061 => x"93762780",
  9062 => x"c9387b70",
  9063 => x"84055d08",
  9064 => x"7c56790c",
  9065 => x"74708405",
  9066 => x"56088c1b",
  9067 => x"0c901a54",
  9068 => x"9b7627ae",
  9069 => x"38747084",
  9070 => x"05560874",
  9071 => x"0c747084",
  9072 => x"05560894",
  9073 => x"1b0c981a",
  9074 => x"54a37627",
  9075 => x"95387470",
  9076 => x"84055608",
  9077 => x"740c7470",
  9078 => x"84055608",
  9079 => x"9c1b0ca0",
  9080 => x"1a547470",
  9081 => x"84055608",
  9082 => x"74708405",
  9083 => x"560c7470",
  9084 => x"84055608",
  9085 => x"74708405",
  9086 => x"560c7408",
  9087 => x"740c7a1a",
  9088 => x"7082cbf8",
  9089 => x"0b88050c",
  9090 => x"7d7c3181",
  9091 => x"0784120c",
  9092 => x"54841a08",
  9093 => x"81067b07",
  9094 => x"841b0c61",
  9095 => x"51feece7",
  9096 => x"3f7854fd",
  9097 => x"b9397553",
  9098 => x"7b527851",
  9099 => x"feebbe3f",
  9100 => x"faec3984",
  9101 => x"1708fc06",
  9102 => x"18605858",
  9103 => x"fae03975",
  9104 => x"537b5278",
  9105 => x"51feeba5",
  9106 => x"3f7a1a70",
  9107 => x"82cbf80b",
  9108 => x"88050c7d",
  9109 => x"7c318107",
  9110 => x"84120c54",
  9111 => x"841a0881",
  9112 => x"067b0784",
  9113 => x"1b0cffb3",
  9114 => x"39fd3d0d",
  9115 => x"75775353",
  9116 => x"71547330",
  9117 => x"7075079f",
  9118 => x"2a7075fe",
  9119 => x"0a060790",
  9120 => x"810a119f",
  9121 => x"fe0a7231",
  9122 => x"07709f2a",
  9123 => x"81713180",
  9124 => x"0c515151",
  9125 => x"5151853d",
  9126 => x"0d04fd3d",
  9127 => x"0d757753",
  9128 => x"53715473",
  9129 => x"30707507",
  9130 => x"9f2a7075",
  9131 => x"fe0a0607",
  9132 => x"9ffe0a71",
  9133 => x"319f2a80",
  9134 => x"0c515151",
  9135 => x"853d0d04",
  9136 => x"f93d0d79",
  9137 => x"7c557b54",
  9138 => x"8e112270",
  9139 => x"902b7090",
  9140 => x"2c555782",
  9141 => x"d4800853",
  9142 => x"585686f9",
  9143 => x"3f800857",
  9144 => x"800b8008",
  9145 => x"24933880",
  9146 => x"d0160880",
  9147 => x"080580d0",
  9148 => x"170c7680",
  9149 => x"0c893d0d",
  9150 => x"048c1622",
  9151 => x"83dfff06",
  9152 => x"55748c17",
  9153 => x"2376800c",
  9154 => x"893d0d04",
  9155 => x"fa3d0d78",
  9156 => x"8c112270",
  9157 => x"882a7081",
  9158 => x"06515758",
  9159 => x"5674a938",
  9160 => x"8c162283",
  9161 => x"dfff0655",
  9162 => x"748c1723",
  9163 => x"7a547953",
  9164 => x"8e162270",
  9165 => x"902b7090",
  9166 => x"2c545682",
  9167 => x"d4800852",
  9168 => x"5683a73f",
  9169 => x"883d0d04",
  9170 => x"82548053",
  9171 => x"8e162270",
  9172 => x"902b7090",
  9173 => x"2c545682",
  9174 => x"d4800852",
  9175 => x"5785be3f",
  9176 => x"8c162283",
  9177 => x"dfff0655",
  9178 => x"748c1723",
  9179 => x"7a547953",
  9180 => x"8e162270",
  9181 => x"902b7090",
  9182 => x"2c545682",
  9183 => x"d4800852",
  9184 => x"5682e73f",
  9185 => x"883d0d04",
  9186 => x"f93d0d79",
  9187 => x"7c557b54",
  9188 => x"8e112270",
  9189 => x"902b7090",
  9190 => x"2c555782",
  9191 => x"d4800853",
  9192 => x"585684f9",
  9193 => x"3f800857",
  9194 => x"8008ff2e",
  9195 => x"99388c16",
  9196 => x"22a08007",
  9197 => x"55748c17",
  9198 => x"23800880",
  9199 => x"d0170c76",
  9200 => x"800c893d",
  9201 => x"0d048c16",
  9202 => x"2283dfff",
  9203 => x"0655748c",
  9204 => x"17237680",
  9205 => x"0c893d0d",
  9206 => x"04fe3d0d",
  9207 => x"748e1122",
  9208 => x"70902b70",
  9209 => x"902c5551",
  9210 => x"515382d4",
  9211 => x"80085183",
  9212 => x"c23f843d",
  9213 => x"0d04fb3d",
  9214 => x"0d777970",
  9215 => x"72078306",
  9216 => x"53545270",
  9217 => x"93387173",
  9218 => x"73085456",
  9219 => x"54717308",
  9220 => x"2e80c438",
  9221 => x"73755452",
  9222 => x"71337081",
  9223 => x"ff065254",
  9224 => x"70802e9d",
  9225 => x"38723355",
  9226 => x"70752e09",
  9227 => x"81069538",
  9228 => x"81128114",
  9229 => x"71337081",
  9230 => x"ff065456",
  9231 => x"545270e5",
  9232 => x"38723355",
  9233 => x"7381ff06",
  9234 => x"7581ff06",
  9235 => x"71713180",
  9236 => x"0c525287",
  9237 => x"3d0d0471",
  9238 => x"0970f7fb",
  9239 => x"fdff1406",
  9240 => x"70f88482",
  9241 => x"81800651",
  9242 => x"51517097",
  9243 => x"38841484",
  9244 => x"16710854",
  9245 => x"56547175",
  9246 => x"082edc38",
  9247 => x"73755452",
  9248 => x"ff963980",
  9249 => x"0b800c87",
  9250 => x"3d0d04fd",
  9251 => x"3d0d7570",
  9252 => x"71830653",
  9253 => x"555270b8",
  9254 => x"38717008",
  9255 => x"7009f7fb",
  9256 => x"fdff1206",
  9257 => x"70f88482",
  9258 => x"81800651",
  9259 => x"51525370",
  9260 => x"9d388413",
  9261 => x"70087009",
  9262 => x"f7fbfdff",
  9263 => x"120670f8",
  9264 => x"84828180",
  9265 => x"06515152",
  9266 => x"5370802e",
  9267 => x"e5387252",
  9268 => x"71335170",
  9269 => x"802e8a38",
  9270 => x"81127033",
  9271 => x"525270f8",
  9272 => x"38717431",
  9273 => x"800c853d",
  9274 => x"0d04fb3d",
  9275 => x"0d800b82",
  9276 => x"dc800c7a",
  9277 => x"53795278",
  9278 => x"5184933f",
  9279 => x"80085580",
  9280 => x"08ff2e88",
  9281 => x"3874800c",
  9282 => x"873d0d04",
  9283 => x"82dc8008",
  9284 => x"5675802e",
  9285 => x"f0387776",
  9286 => x"710c5474",
  9287 => x"800c873d",
  9288 => x"0d04fb3d",
  9289 => x"0d787a29",
  9290 => x"527751fe",
  9291 => x"d9c83f80",
  9292 => x"08800855",
  9293 => x"56800880",
  9294 => x"2e80e338",
  9295 => x"8008fc05",
  9296 => x"08fc06fc",
  9297 => x"055574a4",
  9298 => x"2680da38",
  9299 => x"937527bb",
  9300 => x"38800b80",
  9301 => x"08708405",
  9302 => x"800c0c80",
  9303 => x"08548074",
  9304 => x"70840556",
  9305 => x"0c9b7527",
  9306 => x"a2388074",
  9307 => x"70840556",
  9308 => x"0c807470",
  9309 => x"8405560c",
  9310 => x"a375278f",
  9311 => x"38807470",
  9312 => x"8405560c",
  9313 => x"80747084",
  9314 => x"05560c80",
  9315 => x"74708405",
  9316 => x"560c8074",
  9317 => x"70840556",
  9318 => x"0c80740c",
  9319 => x"75547380",
  9320 => x"0c873d0d",
  9321 => x"04745380",
  9322 => x"52800851",
  9323 => x"db8a3f75",
  9324 => x"54ec39fd",
  9325 => x"3d0d800b",
  9326 => x"82dc800c",
  9327 => x"765184d7",
  9328 => x"3f800853",
  9329 => x"8008ff2e",
  9330 => x"88387280",
  9331 => x"0c853d0d",
  9332 => x"0482dc80",
  9333 => x"08547380",
  9334 => x"2ef03875",
  9335 => x"74710c52",
  9336 => x"72800c85",
  9337 => x"3d0d04fc",
  9338 => x"3d0d800b",
  9339 => x"82dc800c",
  9340 => x"78527751",
  9341 => x"86bf3f80",
  9342 => x"08548008",
  9343 => x"ff2e8838",
  9344 => x"73800c86",
  9345 => x"3d0d0482",
  9346 => x"dc800855",
  9347 => x"74802ef0",
  9348 => x"38767571",
  9349 => x"0c537380",
  9350 => x"0c863d0d",
  9351 => x"04fb3d0d",
  9352 => x"800b82dc",
  9353 => x"800c7a53",
  9354 => x"79527851",
  9355 => x"849b3f80",
  9356 => x"08558008",
  9357 => x"ff2e8838",
  9358 => x"74800c87",
  9359 => x"3d0d0482",
  9360 => x"dc800856",
  9361 => x"75802ef0",
  9362 => x"38777671",
  9363 => x"0c547480",
  9364 => x"0c873d0d",
  9365 => x"04fb3d0d",
  9366 => x"800b82dc",
  9367 => x"800c7a53",
  9368 => x"79527851",
  9369 => x"82a03f80",
  9370 => x"08558008",
  9371 => x"ff2e8838",
  9372 => x"74800c87",
  9373 => x"3d0d0482",
  9374 => x"dc800856",
  9375 => x"75802ef0",
  9376 => x"38777671",
  9377 => x"0c547480",
  9378 => x"0c873d0d",
  9379 => x"04fe3d0d",
  9380 => x"82dbf808",
  9381 => x"51708a38",
  9382 => x"82dc8470",
  9383 => x"82dbf80c",
  9384 => x"51707512",
  9385 => x"5252ff53",
  9386 => x"7087fb80",
  9387 => x"80268838",
  9388 => x"7082dbf8",
  9389 => x"0c715372",
  9390 => x"800c843d",
  9391 => x"0d04fd3d",
  9392 => x"0d800b82",
  9393 => x"cb940854",
  9394 => x"5472812e",
  9395 => x"9e387382",
  9396 => x"dbfc0cfd",
  9397 => x"e3d03ffd",
  9398 => x"e2a63f82",
  9399 => x"dba05281",
  9400 => x"51fdeba3",
  9401 => x"3f800851",
  9402 => x"85cb3f72",
  9403 => x"82dbfc0c",
  9404 => x"fde3b33f",
  9405 => x"fde2893f",
  9406 => x"82dba052",
  9407 => x"8151fdeb",
  9408 => x"863f8008",
  9409 => x"5185ae3f",
  9410 => x"00ff3900",
  9411 => x"ff39f53d",
  9412 => x"0d7e6082",
  9413 => x"dbfc0870",
  9414 => x"5b585b5b",
  9415 => x"7580c538",
  9416 => x"777a25a2",
  9417 => x"38771b70",
  9418 => x"337081ff",
  9419 => x"06585859",
  9420 => x"758a2e99",
  9421 => x"387681ff",
  9422 => x"0651fde2",
  9423 => x"c83f8118",
  9424 => x"58797824",
  9425 => x"e0387980",
  9426 => x"0c8d3d0d",
  9427 => x"048d51fd",
  9428 => x"e2b33f78",
  9429 => x"337081ff",
  9430 => x"065257fd",
  9431 => x"e2a73f81",
  9432 => x"1858de39",
  9433 => x"79557a54",
  9434 => x"7d538552",
  9435 => x"8d3dfc05",
  9436 => x"51fde1ce",
  9437 => x"3f800856",
  9438 => x"84b43f7b",
  9439 => x"80080c75",
  9440 => x"800c8d3d",
  9441 => x"0d04f63d",
  9442 => x"0d7d7f82",
  9443 => x"dbfc0870",
  9444 => x"5b585a5a",
  9445 => x"7580c438",
  9446 => x"777925b6",
  9447 => x"38fde1c0",
  9448 => x"3f800881",
  9449 => x"ff06708d",
  9450 => x"32703070",
  9451 => x"9f2a5151",
  9452 => x"5757768a",
  9453 => x"2e80c638",
  9454 => x"75802e80",
  9455 => x"c038771a",
  9456 => x"56767634",
  9457 => x"7651fde1",
  9458 => x"bc3f8118",
  9459 => x"58787824",
  9460 => x"cc387756",
  9461 => x"75800c8c",
  9462 => x"3d0d0478",
  9463 => x"5579547c",
  9464 => x"5384528c",
  9465 => x"3dfc0551",
  9466 => x"fde0d73f",
  9467 => x"80085683",
  9468 => x"bd3f7a80",
  9469 => x"080c7580",
  9470 => x"0c8c3d0d",
  9471 => x"04771a56",
  9472 => x"8a763481",
  9473 => x"18588d51",
  9474 => x"fde0fa3f",
  9475 => x"8a51fde0",
  9476 => x"f43f7756",
  9477 => x"ffbe39fb",
  9478 => x"3d0d82db",
  9479 => x"fc087056",
  9480 => x"54738838",
  9481 => x"74800c87",
  9482 => x"3d0d0477",
  9483 => x"53835287",
  9484 => x"3dfc0551",
  9485 => x"fde08b3f",
  9486 => x"80085482",
  9487 => x"f13f7580",
  9488 => x"080c7380",
  9489 => x"0c873d0d",
  9490 => x"04fa3d0d",
  9491 => x"82dbfc08",
  9492 => x"802ea338",
  9493 => x"7a557954",
  9494 => x"78538652",
  9495 => x"883dfc05",
  9496 => x"51fddfde",
  9497 => x"3f800856",
  9498 => x"82c43f76",
  9499 => x"80080c75",
  9500 => x"800c883d",
  9501 => x"0d0482b6",
  9502 => x"3f9d0b80",
  9503 => x"080cff0b",
  9504 => x"800c883d",
  9505 => x"0d04fb3d",
  9506 => x"0d777956",
  9507 => x"56807054",
  9508 => x"54737525",
  9509 => x"9f387410",
  9510 => x"1010f805",
  9511 => x"52721670",
  9512 => x"3370742b",
  9513 => x"76078116",
  9514 => x"f8165656",
  9515 => x"56515174",
  9516 => x"7324ea38",
  9517 => x"73800c87",
  9518 => x"3d0d04fc",
  9519 => x"3d0d7678",
  9520 => x"5555bc53",
  9521 => x"80527351",
  9522 => x"d4ee3f84",
  9523 => x"527451ff",
  9524 => x"b53f8008",
  9525 => x"74238452",
  9526 => x"841551ff",
  9527 => x"a93f8008",
  9528 => x"82152384",
  9529 => x"52881551",
  9530 => x"ff9c3f80",
  9531 => x"0884150c",
  9532 => x"84528c15",
  9533 => x"51ff8f3f",
  9534 => x"80088815",
  9535 => x"23845290",
  9536 => x"1551ff82",
  9537 => x"3f80088a",
  9538 => x"15238452",
  9539 => x"941551fe",
  9540 => x"f53f8008",
  9541 => x"8c152384",
  9542 => x"52981551",
  9543 => x"fee83f80",
  9544 => x"088e1523",
  9545 => x"88529c15",
  9546 => x"51fedb3f",
  9547 => x"80089015",
  9548 => x"0c863d0d",
  9549 => x"04e93d0d",
  9550 => x"6a82dbfc",
  9551 => x"08575775",
  9552 => x"933880c0",
  9553 => x"800b8418",
  9554 => x"0c75ac18",
  9555 => x"0c75800c",
  9556 => x"993d0d04",
  9557 => x"893d7055",
  9558 => x"6a54558a",
  9559 => x"52993dff",
  9560 => x"bc0551fd",
  9561 => x"dddc3f80",
  9562 => x"08775375",
  9563 => x"5256fecb",
  9564 => x"3fbc3f77",
  9565 => x"80080c75",
  9566 => x"800c993d",
  9567 => x"0d04fc3d",
  9568 => x"0d815482",
  9569 => x"dbfc0888",
  9570 => x"3873800c",
  9571 => x"863d0d04",
  9572 => x"765397b9",
  9573 => x"52863dfc",
  9574 => x"0551fddd",
  9575 => x"a53f8008",
  9576 => x"548c3f74",
  9577 => x"80080c73",
  9578 => x"800c863d",
  9579 => x"0d0482d4",
  9580 => x"8008800c",
  9581 => x"04f73d0d",
  9582 => x"7b82d480",
  9583 => x"0882c811",
  9584 => x"085a545a",
  9585 => x"77802e80",
  9586 => x"da388188",
  9587 => x"18841908",
  9588 => x"ff058171",
  9589 => x"2b595559",
  9590 => x"80742480",
  9591 => x"ea388074",
  9592 => x"24b53873",
  9593 => x"822b7811",
  9594 => x"88055656",
  9595 => x"81801908",
  9596 => x"77065372",
  9597 => x"802eb638",
  9598 => x"78167008",
  9599 => x"53537951",
  9600 => x"74085372",
  9601 => x"2dff14fc",
  9602 => x"17fc1779",
  9603 => x"812c5a57",
  9604 => x"57547380",
  9605 => x"25d63877",
  9606 => x"085877ff",
  9607 => x"ad3882d4",
  9608 => x"800853bc",
  9609 => x"1308a538",
  9610 => x"7951f9dc",
  9611 => x"3f740853",
  9612 => x"722dff14",
  9613 => x"fc17fc17",
  9614 => x"79812c5a",
  9615 => x"57575473",
  9616 => x"8025ffa8",
  9617 => x"38d13980",
  9618 => x"57ff9339",
  9619 => x"7251bc13",
  9620 => x"0853722d",
  9621 => x"7951f9b0",
  9622 => x"3f8c0802",
  9623 => x"8c0cee3d",
  9624 => x"0d8c0888",
  9625 => x"05088c08",
  9626 => x"8c050855",
  9627 => x"53728c08",
  9628 => x"d0050c73",
  9629 => x"8c08d405",
  9630 => x"0c8c0890",
  9631 => x"05088c08",
  9632 => x"94050855",
  9633 => x"53728c08",
  9634 => x"c8050c73",
  9635 => x"8c08cc05",
  9636 => x"0c8c08ec",
  9637 => x"0570538c",
  9638 => x"08d00570",
  9639 => x"535153fe",
  9640 => x"c8de3f8c",
  9641 => x"08d80570",
  9642 => x"538c08c8",
  9643 => x"05705351",
  9644 => x"53fec8cc",
  9645 => x"3f8c08ec",
  9646 => x"05705253",
  9647 => x"80c83f80",
  9648 => x"08537292",
  9649 => x"388c08d8",
  9650 => x"05705253",
  9651 => x"b93f8008",
  9652 => x"53728338",
  9653 => x"8a39810b",
  9654 => x"8c08c405",
  9655 => x"0c9b398c",
  9656 => x"08d80570",
  9657 => x"538c08ec",
  9658 => x"05705351",
  9659 => x"538ccf3f",
  9660 => x"8008708c",
  9661 => x"08c4050c",
  9662 => x"538c08c4",
  9663 => x"0508800c",
  9664 => x"943d0d8c",
  9665 => x"0c048c08",
  9666 => x"028c0cff",
  9667 => x"3d0d800b",
  9668 => x"8c08fc05",
  9669 => x"0c8c0888",
  9670 => x"05085170",
  9671 => x"08802e8f",
  9672 => x"388c0888",
  9673 => x"05085170",
  9674 => x"08812e83",
  9675 => x"38883981",
  9676 => x"0b8c08fc",
  9677 => x"050c8c08",
  9678 => x"fc050870",
  9679 => x"800c5183",
  9680 => x"3d0d8c0c",
  9681 => x"048c0802",
  9682 => x"8c0cee3d",
  9683 => x"0d8c0888",
  9684 => x"05088c08",
  9685 => x"8c050855",
  9686 => x"53728c08",
  9687 => x"d0050c73",
  9688 => x"8c08d405",
  9689 => x"0c8c0890",
  9690 => x"05088c08",
  9691 => x"94050855",
  9692 => x"53728c08",
  9693 => x"c8050c73",
  9694 => x"8c08cc05",
  9695 => x"0c8c08ec",
  9696 => x"0570538c",
  9697 => x"08d00570",
  9698 => x"535153fe",
  9699 => x"c6f23f8c",
  9700 => x"08d80570",
  9701 => x"538c08c8",
  9702 => x"05705351",
  9703 => x"53fec6e0",
  9704 => x"3f8c08ec",
  9705 => x"05705253",
  9706 => x"80c83f80",
  9707 => x"08537292",
  9708 => x"388c08d8",
  9709 => x"05705253",
  9710 => x"b93f8008",
  9711 => x"53728338",
  9712 => x"8a39810b",
  9713 => x"8c08c405",
  9714 => x"0c9b398c",
  9715 => x"08d80570",
  9716 => x"538c08ec",
  9717 => x"05705351",
  9718 => x"538ae33f",
  9719 => x"8008708c",
  9720 => x"08c4050c",
  9721 => x"538c08c4",
  9722 => x"0508800c",
  9723 => x"943d0d8c",
  9724 => x"0c048c08",
  9725 => x"028c0cff",
  9726 => x"3d0d800b",
  9727 => x"8c08fc05",
  9728 => x"0c8c0888",
  9729 => x"05085170",
  9730 => x"08802e8f",
  9731 => x"388c0888",
  9732 => x"05085170",
  9733 => x"08812e83",
  9734 => x"38883981",
  9735 => x"0b8c08fc",
  9736 => x"050c8c08",
  9737 => x"fc050870",
  9738 => x"800c5183",
  9739 => x"3d0d8c0c",
  9740 => x"048c0802",
  9741 => x"8c0cee3d",
  9742 => x"0d8c0888",
  9743 => x"05088c08",
  9744 => x"8c050855",
  9745 => x"53728c08",
  9746 => x"d0050c73",
  9747 => x"8c08d405",
  9748 => x"0c8c0890",
  9749 => x"05088c08",
  9750 => x"94050855",
  9751 => x"53728c08",
  9752 => x"c8050c73",
  9753 => x"8c08cc05",
  9754 => x"0c8c08ec",
  9755 => x"0570538c",
  9756 => x"08d00570",
  9757 => x"535153fe",
  9758 => x"c5863f8c",
  9759 => x"08d80570",
  9760 => x"538c08c8",
  9761 => x"05705351",
  9762 => x"53fec4f4",
  9763 => x"3f8c08ec",
  9764 => x"05705253",
  9765 => x"80c83f80",
  9766 => x"08537292",
  9767 => x"388c08d8",
  9768 => x"05705253",
  9769 => x"b93f8008",
  9770 => x"53728338",
  9771 => x"8a39ff0b",
  9772 => x"8c08c405",
  9773 => x"0c9b398c",
  9774 => x"08d80570",
  9775 => x"538c08ec",
  9776 => x"05705351",
  9777 => x"5388f73f",
  9778 => x"8008708c",
  9779 => x"08c4050c",
  9780 => x"538c08c4",
  9781 => x"0508800c",
  9782 => x"943d0d8c",
  9783 => x"0c048c08",
  9784 => x"028c0cff",
  9785 => x"3d0d800b",
  9786 => x"8c08fc05",
  9787 => x"0c8c0888",
  9788 => x"05085170",
  9789 => x"08802e8f",
  9790 => x"388c0888",
  9791 => x"05085170",
  9792 => x"08812e83",
  9793 => x"38883981",
  9794 => x"0b8c08fc",
  9795 => x"050c8c08",
  9796 => x"fc050870",
  9797 => x"800c5183",
  9798 => x"3d0d8c0c",
  9799 => x"048c0802",
  9800 => x"8c0cee3d",
  9801 => x"0d8c0888",
  9802 => x"05088c08",
  9803 => x"8c050855",
  9804 => x"53728c08",
  9805 => x"d0050c73",
  9806 => x"8c08d405",
  9807 => x"0c8c0890",
  9808 => x"05088c08",
  9809 => x"94050855",
  9810 => x"53728c08",
  9811 => x"c8050c73",
  9812 => x"8c08cc05",
  9813 => x"0c8c08ec",
  9814 => x"0570538c",
  9815 => x"08d00570",
  9816 => x"535153fe",
  9817 => x"c39a3f8c",
  9818 => x"08d80570",
  9819 => x"538c08c8",
  9820 => x"05705351",
  9821 => x"53fec388",
  9822 => x"3f8c08ec",
  9823 => x"05705253",
  9824 => x"80c83f80",
  9825 => x"08537292",
  9826 => x"388c08d8",
  9827 => x"05705253",
  9828 => x"b93f8008",
  9829 => x"53728338",
  9830 => x"8a39810b",
  9831 => x"8c08c405",
  9832 => x"0c9b398c",
  9833 => x"08d80570",
  9834 => x"538c08ec",
  9835 => x"05705351",
  9836 => x"53878b3f",
  9837 => x"8008708c",
  9838 => x"08c4050c",
  9839 => x"538c08c4",
  9840 => x"0508800c",
  9841 => x"943d0d8c",
  9842 => x"0c048c08",
  9843 => x"028c0cff",
  9844 => x"3d0d800b",
  9845 => x"8c08fc05",
  9846 => x"0c8c0888",
  9847 => x"05085170",
  9848 => x"08802e8f",
  9849 => x"388c0888",
  9850 => x"05085170",
  9851 => x"08812e83",
  9852 => x"38883981",
  9853 => x"0b8c08fc",
  9854 => x"050c8c08",
  9855 => x"fc050870",
  9856 => x"800c5183",
  9857 => x"3d0d8c0c",
  9858 => x"048c0802",
  9859 => x"8c0cee3d",
  9860 => x"0d8c0888",
  9861 => x"05088c08",
  9862 => x"8c050855",
  9863 => x"53728c08",
  9864 => x"d0050c73",
  9865 => x"8c08d405",
  9866 => x"0c8c0890",
  9867 => x"05088c08",
  9868 => x"94050855",
  9869 => x"53728c08",
  9870 => x"c8050c73",
  9871 => x"8c08cc05",
  9872 => x"0c8c08ec",
  9873 => x"0570538c",
  9874 => x"08d00570",
  9875 => x"535153fe",
  9876 => x"c1ae3f8c",
  9877 => x"08d80570",
  9878 => x"538c08c8",
  9879 => x"05705351",
  9880 => x"53fec19c",
  9881 => x"3f8c08ec",
  9882 => x"05705253",
  9883 => x"80c83f80",
  9884 => x"08537292",
  9885 => x"388c08d8",
  9886 => x"05705253",
  9887 => x"b93f8008",
  9888 => x"53728338",
  9889 => x"8a39810b",
  9890 => x"8c08c405",
  9891 => x"0c9b398c",
  9892 => x"08d80570",
  9893 => x"538c08ec",
  9894 => x"05705351",
  9895 => x"53859f3f",
  9896 => x"8008708c",
  9897 => x"08c4050c",
  9898 => x"538c08c4",
  9899 => x"0508800c",
  9900 => x"943d0d8c",
  9901 => x"0c048c08",
  9902 => x"028c0cff",
  9903 => x"3d0d800b",
  9904 => x"8c08fc05",
  9905 => x"0c8c0888",
  9906 => x"05085170",
  9907 => x"08802e8f",
  9908 => x"388c0888",
  9909 => x"05085170",
  9910 => x"08812e83",
  9911 => x"38883981",
  9912 => x"0b8c08fc",
  9913 => x"050c8c08",
  9914 => x"fc050870",
  9915 => x"800c5183",
  9916 => x"3d0d8c0c",
  9917 => x"048c0802",
  9918 => x"8c0cec3d",
  9919 => x"0d8c0888",
  9920 => x"05088c08",
  9921 => x"8c050857",
  9922 => x"55748c08",
  9923 => x"e0050c75",
  9924 => x"8c08e405",
  9925 => x"0c8c08ec",
  9926 => x"0570538c",
  9927 => x"08e00570",
  9928 => x"535155fe",
  9929 => x"bfda3f8c",
  9930 => x"08ec0570",
  9931 => x"5255838e",
  9932 => x"3f800855",
  9933 => x"74802e8b",
  9934 => x"38800b8c",
  9935 => x"08d4050c",
  9936 => x"81fc398c",
  9937 => x"08ec0570",
  9938 => x"525582b3",
  9939 => x"3f800855",
  9940 => x"74802e8b",
  9941 => x"38800b8c",
  9942 => x"08d4050c",
  9943 => x"81e0398c",
  9944 => x"08ec0570",
  9945 => x"525581e3",
  9946 => x"3f800855",
  9947 => x"74802ea9",
  9948 => x"388c08f0",
  9949 => x"0508802e",
  9950 => x"8b38810a",
  9951 => x"0b8c08d0",
  9952 => x"050c8939",
  9953 => x"fe0a0b8c",
  9954 => x"08d0050c",
  9955 => x"8c08d005",
  9956 => x"088c08d4",
  9957 => x"050c81a6",
  9958 => x"398c08f4",
  9959 => x"05088025",
  9960 => x"8b38800b",
  9961 => x"8c08d405",
  9962 => x"0c819339",
  9963 => x"9e0b8c08",
  9964 => x"f4050825",
  9965 => x"a9388c08",
  9966 => x"f0050880",
  9967 => x"2e8b3881",
  9968 => x"0a0b8c08",
  9969 => x"cc050c89",
  9970 => x"39fe0a0b",
  9971 => x"8c08cc05",
  9972 => x"0c8c08cc",
  9973 => x"05088c08",
  9974 => x"d4050c80",
  9975 => x"e139bc0b",
  9976 => x"8c08f405",
  9977 => x"08318c08",
  9978 => x"d8057156",
  9979 => x"58558c08",
  9980 => x"f805088c",
  9981 => x"08fc0508",
  9982 => x"57557452",
  9983 => x"75537651",
  9984 => x"fec1db3f",
  9985 => x"8c08d805",
  9986 => x"088c08dc",
  9987 => x"0508708c",
  9988 => x"08e8050c",
  9989 => x"8c08e805",
  9990 => x"088c08c8",
  9991 => x"050c5755",
  9992 => x"8c08f005",
  9993 => x"08802e8c",
  9994 => x"388c08c8",
  9995 => x"0508308c",
  9996 => x"08c8050c",
  9997 => x"8c08c805",
  9998 => x"088c08d4",
  9999 => x"050c8c08",
 10000 => x"d4050880",
 10001 => x"0c963d0d",
 10002 => x"8c0c048c",
 10003 => x"08028c0c",
 10004 => x"ff3d0d80",
 10005 => x"0b8c08fc",
 10006 => x"050c8c08",
 10007 => x"88050851",
 10008 => x"7008842e",
 10009 => x"09810688",
 10010 => x"38810b8c",
 10011 => x"08fc050c",
 10012 => x"8c08fc05",
 10013 => x"0870800c",
 10014 => x"51833d0d",
 10015 => x"8c0c048c",
 10016 => x"08028c0c",
 10017 => x"ff3d0d80",
 10018 => x"0b8c08fc",
 10019 => x"050c8c08",
 10020 => x"88050851",
 10021 => x"7008802e",
 10022 => x"8f388c08",
 10023 => x"88050851",
 10024 => x"7008812e",
 10025 => x"83388839",
 10026 => x"810b8c08",
 10027 => x"fc050c8c",
 10028 => x"08fc0508",
 10029 => x"70800c51",
 10030 => x"833d0d8c",
 10031 => x"0c048c08",
 10032 => x"028c0cff",
 10033 => x"3d0d800b",
 10034 => x"8c08fc05",
 10035 => x"0c8c0888",
 10036 => x"05085170",
 10037 => x"08822e09",
 10038 => x"81068838",
 10039 => x"810b8c08",
 10040 => x"fc050c8c",
 10041 => x"08fc0508",
 10042 => x"70800c51",
 10043 => x"833d0d8c",
 10044 => x"0c048c08",
 10045 => x"028c0cfd",
 10046 => x"3d0d8053",
 10047 => x"8c088c05",
 10048 => x"08528c08",
 10049 => x"88050851",
 10050 => x"fea4e73f",
 10051 => x"80087080",
 10052 => x"0c54853d",
 10053 => x"0d8c0c04",
 10054 => x"8c08028c",
 10055 => x"0cfd3d0d",
 10056 => x"81538c08",
 10057 => x"8c050852",
 10058 => x"8c088805",
 10059 => x"0851fea4",
 10060 => x"c13f8008",
 10061 => x"70800c54",
 10062 => x"853d0d8c",
 10063 => x"0c048c08",
 10064 => x"028c0cf0",
 10065 => x"3d0d8c08",
 10066 => x"88050851",
 10067 => x"87b73f80",
 10068 => x"08527192",
 10069 => x"388c088c",
 10070 => x"05085187",
 10071 => x"a83f8008",
 10072 => x"52718338",
 10073 => x"8b39810b",
 10074 => x"8c08fc05",
 10075 => x"0c86a139",
 10076 => x"8c088805",
 10077 => x"085186d9",
 10078 => x"3f800852",
 10079 => x"71802eaf",
 10080 => x"388c088c",
 10081 => x"05085186",
 10082 => x"c83f8008",
 10083 => x"5271802e",
 10084 => x"9e388c08",
 10085 => x"8c05088c",
 10086 => x"08880508",
 10087 => x"84120884",
 10088 => x"12083170",
 10089 => x"8c08fc05",
 10090 => x"0c525452",
 10091 => x"85e2398c",
 10092 => x"08880508",
 10093 => x"51869a3f",
 10094 => x"80085271",
 10095 => x"802eab38",
 10096 => x"8c088805",
 10097 => x"08528412",
 10098 => x"08802e8a",
 10099 => x"38ff0b8c",
 10100 => x"08f8050c",
 10101 => x"8839810b",
 10102 => x"8c08f805",
 10103 => x"0c8c08f8",
 10104 => x"05088c08",
 10105 => x"fc050c85",
 10106 => x"a7398c08",
 10107 => x"8c050851",
 10108 => x"85df3f80",
 10109 => x"08527180",
 10110 => x"2eab388c",
 10111 => x"088c0508",
 10112 => x"52841208",
 10113 => x"802e8a38",
 10114 => x"810b8c08",
 10115 => x"f4050c88",
 10116 => x"39ff0b8c",
 10117 => x"08f4050c",
 10118 => x"8c08f405",
 10119 => x"088c08fc",
 10120 => x"050c84ec",
 10121 => x"398c0888",
 10122 => x"05085184",
 10123 => x"f03f8008",
 10124 => x"5271802e",
 10125 => x"9c388c08",
 10126 => x"8c050851",
 10127 => x"84df3f80",
 10128 => x"08527180",
 10129 => x"2e8b3880",
 10130 => x"0b8c08fc",
 10131 => x"050c84c0",
 10132 => x"398c0888",
 10133 => x"05085184",
 10134 => x"c43f8008",
 10135 => x"5271802e",
 10136 => x"ab388c08",
 10137 => x"8c050852",
 10138 => x"84120880",
 10139 => x"2e8a3881",
 10140 => x"0b8c08f0",
 10141 => x"050c8839",
 10142 => x"ff0b8c08",
 10143 => x"f0050c8c",
 10144 => x"08f00508",
 10145 => x"8c08fc05",
 10146 => x"0c848539",
 10147 => x"8c088c05",
 10148 => x"08518489",
 10149 => x"3f800852",
 10150 => x"71802eab",
 10151 => x"388c0888",
 10152 => x"05085284",
 10153 => x"1208802e",
 10154 => x"8a38ff0b",
 10155 => x"8c08ec05",
 10156 => x"0c883981",
 10157 => x"0b8c08ec",
 10158 => x"050c8c08",
 10159 => x"ec05088c",
 10160 => x"08fc050c",
 10161 => x"83ca398c",
 10162 => x"08880508",
 10163 => x"8c088c05",
 10164 => x"08535384",
 10165 => x"13088413",
 10166 => x"082eab38",
 10167 => x"8c088805",
 10168 => x"08528412",
 10169 => x"08802e8a",
 10170 => x"38ff0b8c",
 10171 => x"08e8050c",
 10172 => x"8839810b",
 10173 => x"8c08e805",
 10174 => x"0c8c08e8",
 10175 => x"05088c08",
 10176 => x"fc050c83",
 10177 => x"8b398c08",
 10178 => x"8805088c",
 10179 => x"088c0508",
 10180 => x"53538812",
 10181 => x"08881408",
 10182 => x"25ab388c",
 10183 => x"08880508",
 10184 => x"52841208",
 10185 => x"802e8a38",
 10186 => x"ff0b8c08",
 10187 => x"e4050c88",
 10188 => x"39810b8c",
 10189 => x"08e4050c",
 10190 => x"8c08e405",
 10191 => x"088c08fc",
 10192 => x"050c82cc",
 10193 => x"398c0888",
 10194 => x"05088c08",
 10195 => x"8c050853",
 10196 => x"53881308",
 10197 => x"88130825",
 10198 => x"ab388c08",
 10199 => x"88050852",
 10200 => x"84120880",
 10201 => x"2e8a3881",
 10202 => x"0b8c08e0",
 10203 => x"050c8839",
 10204 => x"ff0b8c08",
 10205 => x"e0050c8c",
 10206 => x"08e00508",
 10207 => x"8c08fc05",
 10208 => x"0c828d39",
 10209 => x"8c088805",
 10210 => x"088c08dc",
 10211 => x"050c8c08",
 10212 => x"8c05088c",
 10213 => x"08d8050c",
 10214 => x"8c08dc05",
 10215 => x"088c08d8",
 10216 => x"05085452",
 10217 => x"8c12088c",
 10218 => x"140826b1",
 10219 => x"388c08dc",
 10220 => x"05088c08",
 10221 => x"d8050854",
 10222 => x"528c1208",
 10223 => x"8c14082e",
 10224 => x"09810680",
 10225 => x"c2388c08",
 10226 => x"dc05088c",
 10227 => x"08d80508",
 10228 => x"54529012",
 10229 => x"08901408",
 10230 => x"268338ab",
 10231 => x"398c0888",
 10232 => x"05085284",
 10233 => x"1208802e",
 10234 => x"8a38ff0b",
 10235 => x"8c08d405",
 10236 => x"0c883981",
 10237 => x"0b8c08d4",
 10238 => x"050c8c08",
 10239 => x"d405088c",
 10240 => x"08fc050c",
 10241 => x"818a398c",
 10242 => x"088c0508",
 10243 => x"8c08d005",
 10244 => x"0c8c0888",
 10245 => x"05088c08",
 10246 => x"cc050c8c",
 10247 => x"08d00508",
 10248 => x"8c08cc05",
 10249 => x"0854528c",
 10250 => x"12088c14",
 10251 => x"0826b138",
 10252 => x"8c08d005",
 10253 => x"088c08cc",
 10254 => x"05085452",
 10255 => x"8c12088c",
 10256 => x"14082e09",
 10257 => x"810680c1",
 10258 => x"388c08d0",
 10259 => x"05088c08",
 10260 => x"cc050854",
 10261 => x"52901208",
 10262 => x"90140826",
 10263 => x"8338aa39",
 10264 => x"8c088805",
 10265 => x"08528412",
 10266 => x"08802e8a",
 10267 => x"38810b8c",
 10268 => x"08c8050c",
 10269 => x"8839ff0b",
 10270 => x"8c08c805",
 10271 => x"0c8c08c8",
 10272 => x"05088c08",
 10273 => x"fc050c88",
 10274 => x"39800b8c",
 10275 => x"08fc050c",
 10276 => x"8c08fc05",
 10277 => x"08800c92",
 10278 => x"3d0d8c0c",
 10279 => x"048c0802",
 10280 => x"8c0cff3d",
 10281 => x"0d800b8c",
 10282 => x"08fc050c",
 10283 => x"8c088805",
 10284 => x"08517008",
 10285 => x"822e0981",
 10286 => x"06883881",
 10287 => x"0b8c08fc",
 10288 => x"050c8c08",
 10289 => x"fc050870",
 10290 => x"800c5183",
 10291 => x"3d0d8c0c",
 10292 => x"048c0802",
 10293 => x"8c0cff3d",
 10294 => x"0d800b8c",
 10295 => x"08fc050c",
 10296 => x"8c088805",
 10297 => x"08517008",
 10298 => x"842e0981",
 10299 => x"06883881",
 10300 => x"0b8c08fc",
 10301 => x"050c8c08",
 10302 => x"fc050870",
 10303 => x"800c5183",
 10304 => x"3d0d8c0c",
 10305 => x"048c0802",
 10306 => x"8c0cff3d",
 10307 => x"0d800b8c",
 10308 => x"08fc050c",
 10309 => x"8c088805",
 10310 => x"08517008",
 10311 => x"802e8f38",
 10312 => x"8c088805",
 10313 => x"08517008",
 10314 => x"812e8338",
 10315 => x"8839810b",
 10316 => x"8c08fc05",
 10317 => x"0c8c08fc",
 10318 => x"05087080",
 10319 => x"0c51833d",
 10320 => x"0d8c0c04",
 10321 => x"ff3d0d82",
 10322 => x"dba80bfc",
 10323 => x"05700852",
 10324 => x"5270ff2e",
 10325 => x"9138702d",
 10326 => x"fc127008",
 10327 => x"525270ff",
 10328 => x"2e098106",
 10329 => x"f138833d",
 10330 => x"0d0404fd",
 10331 => x"c7a53f04",
 10332 => x"00000040",
 10333 => x"0a53656e",
 10334 => x"64696e67",
 10335 => x"20313530",
 10336 => x"30204d62",
 10337 => x"79746520",
 10338 => x"6f662064",
 10339 => x"61746120",
 10340 => x"746f2025",
 10341 => x"2e303278",
 10342 => x"3a252e30",
 10343 => x"32783a25",
 10344 => x"2e303278",
 10345 => x"3a252e30",
 10346 => x"32783a25",
 10347 => x"2e303278",
 10348 => x"3a252e30",
 10349 => x"32780a00",
 10350 => x"0a54696d",
 10351 => x"653a2025",
 10352 => x"660a0000",
 10353 => x"42697472",
 10354 => x"6174653a",
 10355 => x"20256620",
 10356 => x"4d627073",
 10357 => x"0a000000",
 10358 => x"00000000",
 10359 => x"00000000",
 10360 => x"00000000",
 10361 => x"00000000",
 10362 => x"00000000",
 10363 => x"20202020",
 10364 => x"20202020",
 10365 => x"20202020",
 10366 => x"20202020",
 10367 => x"30303030",
 10368 => x"30303030",
 10369 => x"30303030",
 10370 => x"30303030",
 10371 => x"00004e91",
 10372 => x"00004a41",
 10373 => x"00004a41",
 10374 => x"00004e87",
 10375 => x"00004a41",
 10376 => x"00004a41",
 10377 => x"00004a41",
 10378 => x"00004a41",
 10379 => x"00004a41",
 10380 => x"00004a41",
 10381 => x"00004a18",
 10382 => x"00004e26",
 10383 => x"00004a41",
 10384 => x"00004a2a",
 10385 => x"00004bc9",
 10386 => x"00004a41",
 10387 => x"00004e54",
 10388 => x"00004e32",
 10389 => x"00004e32",
 10390 => x"00004e32",
 10391 => x"00004e32",
 10392 => x"00004e32",
 10393 => x"00004e32",
 10394 => x"00004e32",
 10395 => x"00004e32",
 10396 => x"00004e32",
 10397 => x"00004a41",
 10398 => x"00004a41",
 10399 => x"00004a41",
 10400 => x"00004a41",
 10401 => x"00004a41",
 10402 => x"00004a41",
 10403 => x"00004a41",
 10404 => x"00004a41",
 10405 => x"00004a41",
 10406 => x"00004d19",
 10407 => x"000049e0",
 10408 => x"00004ca2",
 10409 => x"00004a41",
 10410 => x"00004ca2",
 10411 => x"00004a41",
 10412 => x"00004a41",
 10413 => x"00004a41",
 10414 => x"00004a41",
 10415 => x"00004e5f",
 10416 => x"00004a41",
 10417 => x"00004a41",
 10418 => x"000049ad",
 10419 => x"00004a41",
 10420 => x"00004a41",
 10421 => x"00004a41",
 10422 => x"00004daa",
 10423 => x"00004a41",
 10424 => x"000046fc",
 10425 => x"00004a41",
 10426 => x"00004a41",
 10427 => x"00004d63",
 10428 => x"00004a41",
 10429 => x"00004a41",
 10430 => x"00004a41",
 10431 => x"00004a41",
 10432 => x"00004a41",
 10433 => x"00004a41",
 10434 => x"00004a41",
 10435 => x"00004a41",
 10436 => x"00004a41",
 10437 => x"00004a41",
 10438 => x"00004d19",
 10439 => x"000049e4",
 10440 => x"00004ca2",
 10441 => x"00004ca2",
 10442 => x"00004ca2",
 10443 => x"00004c97",
 10444 => x"000049e4",
 10445 => x"00004a41",
 10446 => x"00004a41",
 10447 => x"00004bab",
 10448 => x"00004a41",
 10449 => x"00004dfb",
 10450 => x"000049b1",
 10451 => x"00004c0c",
 10452 => x"00004a37",
 10453 => x"00004a41",
 10454 => x"00004daa",
 10455 => x"00004a41",
 10456 => x"00004700",
 10457 => x"00004a41",
 10458 => x"00004a41",
 10459 => x"00004e69",
 10460 => x"62756720",
 10461 => x"696e2076",
 10462 => x"66707269",
 10463 => x"6e74663a",
 10464 => x"20626164",
 10465 => x"20626173",
 10466 => x"65000000",
 10467 => x"30313233",
 10468 => x"34353637",
 10469 => x"38396162",
 10470 => x"63646566",
 10471 => x"00000000",
 10472 => x"496e6600",
 10473 => x"30313233",
 10474 => x"34353637",
 10475 => x"38394142",
 10476 => x"43444546",
 10477 => x"00000000",
 10478 => x"30000000",
 10479 => x"2e000000",
 10480 => x"4e614e00",
 10481 => x"286e756c",
 10482 => x"6c290000",
 10483 => x"432d5554",
 10484 => x"462d3800",
 10485 => x"432d534a",
 10486 => x"49530000",
 10487 => x"432d4555",
 10488 => x"434a5000",
 10489 => x"432d4a49",
 10490 => x"53000000",
 10491 => x"496e6669",
 10492 => x"6e697479",
 10493 => x"00000000",
 10494 => x"00006aa4",
 10495 => x"00006aa4",
 10496 => x"00006a8e",
 10497 => x"000065a3",
 10498 => x"00006a93",
 10499 => x"000065a8",
 10500 => x"43000000",
 10501 => x"49534f2d",
 10502 => x"38383539",
 10503 => x"2d310000",
 10504 => x"0000a3bc",
 10505 => x"0000a3b4",
 10506 => x"0000a3b4",
 10507 => x"0000a3b4",
 10508 => x"0000a3b4",
 10509 => x"0000a3b4",
 10510 => x"0000a3b4",
 10511 => x"0000a3b4",
 10512 => x"0000a3b4",
 10513 => x"0000a3b4",
 10514 => x"ffffffff",
 10515 => x"ffffffff",
 10516 => x"3c9cd2b2",
 10517 => x"97d889bc",
 10518 => x"3949f623",
 10519 => x"d5a8a733",
 10520 => x"32a50ffd",
 10521 => x"44f4a73d",
 10522 => x"255bba08",
 10523 => x"cf8c979d",
 10524 => x"0ac80628",
 10525 => x"64ac6f43",
 10526 => x"4341c379",
 10527 => x"37e08000",
 10528 => x"4693b8b5",
 10529 => x"b5056e17",
 10530 => x"4d384f03",
 10531 => x"e93ff9f5",
 10532 => x"5a827748",
 10533 => x"f9301d32",
 10534 => x"75154fdd",
 10535 => x"7f73bf3c",
 10536 => x"3ff00000",
 10537 => x"00000000",
 10538 => x"40240000",
 10539 => x"00000000",
 10540 => x"40590000",
 10541 => x"00000000",
 10542 => x"408f4000",
 10543 => x"00000000",
 10544 => x"40c38800",
 10545 => x"00000000",
 10546 => x"40f86a00",
 10547 => x"00000000",
 10548 => x"412e8480",
 10549 => x"00000000",
 10550 => x"416312d0",
 10551 => x"00000000",
 10552 => x"4197d784",
 10553 => x"00000000",
 10554 => x"41cdcd65",
 10555 => x"00000000",
 10556 => x"4202a05f",
 10557 => x"20000000",
 10558 => x"42374876",
 10559 => x"e8000000",
 10560 => x"426d1a94",
 10561 => x"a2000000",
 10562 => x"42a2309c",
 10563 => x"e5400000",
 10564 => x"42d6bcc4",
 10565 => x"1e900000",
 10566 => x"430c6bf5",
 10567 => x"26340000",
 10568 => x"4341c379",
 10569 => x"37e08000",
 10570 => x"43763457",
 10571 => x"85d8a000",
 10572 => x"43abc16d",
 10573 => x"674ec800",
 10574 => x"43e158e4",
 10575 => x"60913d00",
 10576 => x"4415af1d",
 10577 => x"78b58c40",
 10578 => x"444b1ae4",
 10579 => x"d6e2ef50",
 10580 => x"4480f0cf",
 10581 => x"064dd592",
 10582 => x"44b52d02",
 10583 => x"c7e14af6",
 10584 => x"44ea7843",
 10585 => x"79d99db4",
 10586 => x"00000005",
 10587 => x"00000019",
 10588 => x"0000007d",
 10589 => x"64756d6d",
 10590 => x"792e6578",
 10591 => x"65000000",
 10592 => x"00ffffff",
 10593 => x"ff00ffff",
 10594 => x"ffff00ff",
 10595 => x"ffffff00",
 10596 => x"00000000",
 10597 => x"00000000",
 10598 => x"00000000",
 10599 => x"0000adb0",
 10600 => x"fff00000",
 10601 => x"80000e00",
 10602 => x"80000c00",
 10603 => x"80000800",
 10604 => x"80000600",
 10605 => x"80000200",
 10606 => x"80000100",
 10607 => x"00000000",
 10608 => x"00000000",
 10609 => x"00000000",
 10610 => x"00000000",
 10611 => x"00000000",
 10612 => x"00000000",
 10613 => x"00000000",
 10614 => x"00000000",
 10615 => x"00000000",
 10616 => x"00000000",
 10617 => x"00000000",
 10618 => x"00000000",
 10619 => x"ffffffff",
 10620 => x"00000000",
 10621 => x"00020000",
 10622 => x"00000000",
 10623 => x"00000000",
 10624 => x"0000a5f8",
 10625 => x"0000a5f8",
 10626 => x"0000a600",
 10627 => x"0000a600",
 10628 => x"0000a608",
 10629 => x"0000a608",
 10630 => x"0000a610",
 10631 => x"0000a610",
 10632 => x"0000a618",
 10633 => x"0000a618",
 10634 => x"0000a620",
 10635 => x"0000a620",
 10636 => x"0000a628",
 10637 => x"0000a628",
 10638 => x"0000a630",
 10639 => x"0000a630",
 10640 => x"0000a638",
 10641 => x"0000a638",
 10642 => x"0000a640",
 10643 => x"0000a640",
 10644 => x"0000a648",
 10645 => x"0000a648",
 10646 => x"0000a650",
 10647 => x"0000a650",
 10648 => x"0000a658",
 10649 => x"0000a658",
 10650 => x"0000a660",
 10651 => x"0000a660",
 10652 => x"0000a668",
 10653 => x"0000a668",
 10654 => x"0000a670",
 10655 => x"0000a670",
 10656 => x"0000a678",
 10657 => x"0000a678",
 10658 => x"0000a680",
 10659 => x"0000a680",
 10660 => x"0000a688",
 10661 => x"0000a688",
 10662 => x"0000a690",
 10663 => x"0000a690",
 10664 => x"0000a698",
 10665 => x"0000a698",
 10666 => x"0000a6a0",
 10667 => x"0000a6a0",
 10668 => x"0000a6a8",
 10669 => x"0000a6a8",
 10670 => x"0000a6b0",
 10671 => x"0000a6b0",
 10672 => x"0000a6b8",
 10673 => x"0000a6b8",
 10674 => x"0000a6c0",
 10675 => x"0000a6c0",
 10676 => x"0000a6c8",
 10677 => x"0000a6c8",
 10678 => x"0000a6d0",
 10679 => x"0000a6d0",
 10680 => x"0000a6d8",
 10681 => x"0000a6d8",
 10682 => x"0000a6e0",
 10683 => x"0000a6e0",
 10684 => x"0000a6e8",
 10685 => x"0000a6e8",
 10686 => x"0000a6f0",
 10687 => x"0000a6f0",
 10688 => x"0000a6f8",
 10689 => x"0000a6f8",
 10690 => x"0000a700",
 10691 => x"0000a700",
 10692 => x"0000a708",
 10693 => x"0000a708",
 10694 => x"0000a710",
 10695 => x"0000a710",
 10696 => x"0000a718",
 10697 => x"0000a718",
 10698 => x"0000a720",
 10699 => x"0000a720",
 10700 => x"0000a728",
 10701 => x"0000a728",
 10702 => x"0000a730",
 10703 => x"0000a730",
 10704 => x"0000a738",
 10705 => x"0000a738",
 10706 => x"0000a740",
 10707 => x"0000a740",
 10708 => x"0000a748",
 10709 => x"0000a748",
 10710 => x"0000a750",
 10711 => x"0000a750",
 10712 => x"0000a758",
 10713 => x"0000a758",
 10714 => x"0000a760",
 10715 => x"0000a760",
 10716 => x"0000a768",
 10717 => x"0000a768",
 10718 => x"0000a770",
 10719 => x"0000a770",
 10720 => x"0000a778",
 10721 => x"0000a778",
 10722 => x"0000a780",
 10723 => x"0000a780",
 10724 => x"0000a788",
 10725 => x"0000a788",
 10726 => x"0000a790",
 10727 => x"0000a790",
 10728 => x"0000a798",
 10729 => x"0000a798",
 10730 => x"0000a7a0",
 10731 => x"0000a7a0",
 10732 => x"0000a7a8",
 10733 => x"0000a7a8",
 10734 => x"0000a7b0",
 10735 => x"0000a7b0",
 10736 => x"0000a7b8",
 10737 => x"0000a7b8",
 10738 => x"0000a7c0",
 10739 => x"0000a7c0",
 10740 => x"0000a7c8",
 10741 => x"0000a7c8",
 10742 => x"0000a7d0",
 10743 => x"0000a7d0",
 10744 => x"0000a7d8",
 10745 => x"0000a7d8",
 10746 => x"0000a7e0",
 10747 => x"0000a7e0",
 10748 => x"0000a7e8",
 10749 => x"0000a7e8",
 10750 => x"0000a7f0",
 10751 => x"0000a7f0",
 10752 => x"0000a7f8",
 10753 => x"0000a7f8",
 10754 => x"0000a800",
 10755 => x"0000a800",
 10756 => x"0000a808",
 10757 => x"0000a808",
 10758 => x"0000a810",
 10759 => x"0000a810",
 10760 => x"0000a818",
 10761 => x"0000a818",
 10762 => x"0000a820",
 10763 => x"0000a820",
 10764 => x"0000a828",
 10765 => x"0000a828",
 10766 => x"0000a830",
 10767 => x"0000a830",
 10768 => x"0000a838",
 10769 => x"0000a838",
 10770 => x"0000a840",
 10771 => x"0000a840",
 10772 => x"0000a848",
 10773 => x"0000a848",
 10774 => x"0000a850",
 10775 => x"0000a850",
 10776 => x"0000a858",
 10777 => x"0000a858",
 10778 => x"0000a860",
 10779 => x"0000a860",
 10780 => x"0000a868",
 10781 => x"0000a868",
 10782 => x"0000a870",
 10783 => x"0000a870",
 10784 => x"0000a878",
 10785 => x"0000a878",
 10786 => x"0000a880",
 10787 => x"0000a880",
 10788 => x"0000a888",
 10789 => x"0000a888",
 10790 => x"0000a890",
 10791 => x"0000a890",
 10792 => x"0000a898",
 10793 => x"0000a898",
 10794 => x"0000a8a0",
 10795 => x"0000a8a0",
 10796 => x"0000a8a8",
 10797 => x"0000a8a8",
 10798 => x"0000a8b0",
 10799 => x"0000a8b0",
 10800 => x"0000a8b8",
 10801 => x"0000a8b8",
 10802 => x"0000a8c0",
 10803 => x"0000a8c0",
 10804 => x"0000a8c8",
 10805 => x"0000a8c8",
 10806 => x"0000a8d0",
 10807 => x"0000a8d0",
 10808 => x"0000a8d8",
 10809 => x"0000a8d8",
 10810 => x"0000a8e0",
 10811 => x"0000a8e0",
 10812 => x"0000a8e8",
 10813 => x"0000a8e8",
 10814 => x"0000a8f0",
 10815 => x"0000a8f0",
 10816 => x"0000a8f8",
 10817 => x"0000a8f8",
 10818 => x"0000a900",
 10819 => x"0000a900",
 10820 => x"0000a908",
 10821 => x"0000a908",
 10822 => x"0000a910",
 10823 => x"0000a910",
 10824 => x"0000a918",
 10825 => x"0000a918",
 10826 => x"0000a920",
 10827 => x"0000a920",
 10828 => x"0000a928",
 10829 => x"0000a928",
 10830 => x"0000a930",
 10831 => x"0000a930",
 10832 => x"0000a938",
 10833 => x"0000a938",
 10834 => x"0000a940",
 10835 => x"0000a940",
 10836 => x"0000a948",
 10837 => x"0000a948",
 10838 => x"0000a950",
 10839 => x"0000a950",
 10840 => x"0000a958",
 10841 => x"0000a958",
 10842 => x"0000a960",
 10843 => x"0000a960",
 10844 => x"0000a968",
 10845 => x"0000a968",
 10846 => x"0000a970",
 10847 => x"0000a970",
 10848 => x"0000a978",
 10849 => x"0000a978",
 10850 => x"0000a980",
 10851 => x"0000a980",
 10852 => x"0000a988",
 10853 => x"0000a988",
 10854 => x"0000a990",
 10855 => x"0000a990",
 10856 => x"0000a998",
 10857 => x"0000a998",
 10858 => x"0000a9a0",
 10859 => x"0000a9a0",
 10860 => x"0000a9a8",
 10861 => x"0000a9a8",
 10862 => x"0000a9b0",
 10863 => x"0000a9b0",
 10864 => x"0000a9b8",
 10865 => x"0000a9b8",
 10866 => x"0000a9c0",
 10867 => x"0000a9c0",
 10868 => x"0000a9c8",
 10869 => x"0000a9c8",
 10870 => x"0000a9d0",
 10871 => x"0000a9d0",
 10872 => x"0000a9d8",
 10873 => x"0000a9d8",
 10874 => x"0000a9e0",
 10875 => x"0000a9e0",
 10876 => x"0000a9e8",
 10877 => x"0000a9e8",
 10878 => x"0000a9f0",
 10879 => x"0000a9f0",
 10880 => x"0000aa04",
 10881 => x"00000000",
 10882 => x"0000ac6c",
 10883 => x"0000acc8",
 10884 => x"0000ad24",
 10885 => x"00000000",
 10886 => x"00000000",
 10887 => x"00000000",
 10888 => x"00000000",
 10889 => x"00000000",
 10890 => x"00000000",
 10891 => x"00000000",
 10892 => x"00000000",
 10893 => x"00000000",
 10894 => x"0000a410",
 10895 => x"00000000",
 10896 => x"00000000",
 10897 => x"00000000",
 10898 => x"00000000",
 10899 => x"00000000",
 10900 => x"00000000",
 10901 => x"00000000",
 10902 => x"00000000",
 10903 => x"00000000",
 10904 => x"00000000",
 10905 => x"00000000",
 10906 => x"00000000",
 10907 => x"00000000",
 10908 => x"00000000",
 10909 => x"00000000",
 10910 => x"00000000",
 10911 => x"00000000",
 10912 => x"00000000",
 10913 => x"00000000",
 10914 => x"00000000",
 10915 => x"00000000",
 10916 => x"00000000",
 10917 => x"00000000",
 10918 => x"00000000",
 10919 => x"00000000",
 10920 => x"00000000",
 10921 => x"00000000",
 10922 => x"00000000",
 10923 => x"00000001",
 10924 => x"330eabcd",
 10925 => x"1234e66d",
 10926 => x"deec0005",
 10927 => x"000b0000",
 10928 => x"00000000",
 10929 => x"00000000",
 10930 => x"00000000",
 10931 => x"00000000",
 10932 => x"00000000",
 10933 => x"00000000",
 10934 => x"00000000",
 10935 => x"00000000",
 10936 => x"00000000",
 10937 => x"00000000",
 10938 => x"00000000",
 10939 => x"00000000",
 10940 => x"00000000",
 10941 => x"00000000",
 10942 => x"00000000",
 10943 => x"00000000",
 10944 => x"00000000",
 10945 => x"00000000",
 10946 => x"00000000",
 10947 => x"00000000",
 10948 => x"00000000",
 10949 => x"00000000",
 10950 => x"00000000",
 10951 => x"00000000",
 10952 => x"00000000",
 10953 => x"00000000",
 10954 => x"00000000",
 10955 => x"00000000",
 10956 => x"00000000",
 10957 => x"00000000",
 10958 => x"00000000",
 10959 => x"00000000",
 10960 => x"00000000",
 10961 => x"00000000",
 10962 => x"00000000",
 10963 => x"00000000",
 10964 => x"00000000",
 10965 => x"00000000",
 10966 => x"00000000",
 10967 => x"00000000",
 10968 => x"00000000",
 10969 => x"00000000",
 10970 => x"00000000",
 10971 => x"00000000",
 10972 => x"00000000",
 10973 => x"00000000",
 10974 => x"00000000",
 10975 => x"00000000",
 10976 => x"00000000",
 10977 => x"00000000",
 10978 => x"00000000",
 10979 => x"00000000",
 10980 => x"00000000",
 10981 => x"00000000",
 10982 => x"00000000",
 10983 => x"00000000",
 10984 => x"00000000",
 10985 => x"00000000",
 10986 => x"00000000",
 10987 => x"00000000",
 10988 => x"00000000",
 10989 => x"00000000",
 10990 => x"00000000",
 10991 => x"00000000",
 10992 => x"00000000",
 10993 => x"00000000",
 10994 => x"00000000",
 10995 => x"00000000",
 10996 => x"00000000",
 10997 => x"00000000",
 10998 => x"00000000",
 10999 => x"00000000",
 11000 => x"00000000",
 11001 => x"00000000",
 11002 => x"00000000",
 11003 => x"00000000",
 11004 => x"00000000",
 11005 => x"00000000",
 11006 => x"00000000",
 11007 => x"00000000",
 11008 => x"00000000",
 11009 => x"00000000",
 11010 => x"00000000",
 11011 => x"00000000",
 11012 => x"00000000",
 11013 => x"00000000",
 11014 => x"00000000",
 11015 => x"00000000",
 11016 => x"00000000",
 11017 => x"00000000",
 11018 => x"00000000",
 11019 => x"00000000",
 11020 => x"00000000",
 11021 => x"00000000",
 11022 => x"00000000",
 11023 => x"00000000",
 11024 => x"00000000",
 11025 => x"00000000",
 11026 => x"00000000",
 11027 => x"00000000",
 11028 => x"00000000",
 11029 => x"00000000",
 11030 => x"00000000",
 11031 => x"00000000",
 11032 => x"00000000",
 11033 => x"00000000",
 11034 => x"00000000",
 11035 => x"00000000",
 11036 => x"00000000",
 11037 => x"00000000",
 11038 => x"00000000",
 11039 => x"00000000",
 11040 => x"00000000",
 11041 => x"00000000",
 11042 => x"00000000",
 11043 => x"00000000",
 11044 => x"00000000",
 11045 => x"00000000",
 11046 => x"00000000",
 11047 => x"00000000",
 11048 => x"00000000",
 11049 => x"00000000",
 11050 => x"00000000",
 11051 => x"00000000",
 11052 => x"00000000",
 11053 => x"00000000",
 11054 => x"00000000",
 11055 => x"00000000",
 11056 => x"00000000",
 11057 => x"00000000",
 11058 => x"00000000",
 11059 => x"00000000",
 11060 => x"00000000",
 11061 => x"00000000",
 11062 => x"00000000",
 11063 => x"00000000",
 11064 => x"00000000",
 11065 => x"00000000",
 11066 => x"00000000",
 11067 => x"00000000",
 11068 => x"00000000",
 11069 => x"00000000",
 11070 => x"00000000",
 11071 => x"00000000",
 11072 => x"00000000",
 11073 => x"00000000",
 11074 => x"00000000",
 11075 => x"00000000",
 11076 => x"00000000",
 11077 => x"00000000",
 11078 => x"00000000",
 11079 => x"00000000",
 11080 => x"00000000",
 11081 => x"00000000",
 11082 => x"00000000",
 11083 => x"00000000",
 11084 => x"00000000",
 11085 => x"00000000",
 11086 => x"00000000",
 11087 => x"00000000",
 11088 => x"00000000",
 11089 => x"00000000",
 11090 => x"00000000",
 11091 => x"00000000",
 11092 => x"00000000",
 11093 => x"00000000",
 11094 => x"00000000",
 11095 => x"00000000",
 11096 => x"00000000",
 11097 => x"00000000",
 11098 => x"00000000",
 11099 => x"00000000",
 11100 => x"00000000",
 11101 => x"00000000",
 11102 => x"00000000",
 11103 => x"00000000",
 11104 => x"43000000",
 11105 => x"00000000",
 11106 => x"00000000",
 11107 => x"00000000",
 11108 => x"00000000",
 11109 => x"00000000",
 11110 => x"00000001",
 11111 => x"0000a414",
 11112 => x"0000a574",
 11113 => x"ffffffff",
 11114 => x"00000000",
 11115 => x"ffffffff",
 11116 => x"00000000",
 11117 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
