-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0b97e00c",
     3 => x"3a0b0b0b",
     4 => x"94ec0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b95ac2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b97",
   162 => x"cc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b90",
   171 => x"f02d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b92",
   179 => x"a22d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0b97dc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f8e",
   257 => x"cc3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"53510497",
   280 => x"dc08802e",
   281 => x"a13897e0",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"9f900c82",
   286 => x"a0800b9f",
   287 => x"940c8290",
   288 => x"800b9f98",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0b9f",
   292 => x"900cf880",
   293 => x"8082800b",
   294 => x"9f940cf8",
   295 => x"80808480",
   296 => x"0b9f980c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0b9f90",
   300 => x"0c80c0a8",
   301 => x"80940b9f",
   302 => x"940c0b0b",
   303 => x"0b96fc0b",
   304 => x"9f980c04",
   305 => x"ff3d0d9f",
   306 => x"9c335170",
   307 => x"a33897e8",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"97e80c70",
   312 => x"2d97e808",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0b9f9c34",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0b9f",
   319 => x"8c08802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0b9f8c",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"fd3d0d97",
   330 => x"f00876b0",
   331 => x"ea299412",
   332 => x"0c54850b",
   333 => x"98150c98",
   334 => x"14087081",
   335 => x"06515372",
   336 => x"f638853d",
   337 => x"0d04ff3d",
   338 => x"0d97f008",
   339 => x"74101075",
   340 => x"10059412",
   341 => x"0c52850b",
   342 => x"98130c98",
   343 => x"12087081",
   344 => x"06515170",
   345 => x"f638833d",
   346 => x"0d04803d",
   347 => x"0d725180",
   348 => x"71278738",
   349 => x"ff115170",
   350 => x"fb38823d",
   351 => x"0d04803d",
   352 => x"0d97f008",
   353 => x"51870b84",
   354 => x"120c823d",
   355 => x"0d04803d",
   356 => x"0d97f408",
   357 => x"51b60b8c",
   358 => x"120c830b",
   359 => x"88120c82",
   360 => x"3d0d04ff",
   361 => x"3d0d97f4",
   362 => x"08528412",
   363 => x"08708106",
   364 => x"51517080",
   365 => x"2ef43871",
   366 => x"087081ff",
   367 => x"06800c51",
   368 => x"833d0d04",
   369 => x"fe3d0d02",
   370 => x"93053397",
   371 => x"f4085353",
   372 => x"84120870",
   373 => x"822a7081",
   374 => x"06515151",
   375 => x"70802ef0",
   376 => x"3872720c",
   377 => x"843d0d04",
   378 => x"fe3d0d02",
   379 => x"93053353",
   380 => x"728a2e9d",
   381 => x"3897f408",
   382 => x"52841208",
   383 => x"70822a70",
   384 => x"81065151",
   385 => x"5170802e",
   386 => x"f0387272",
   387 => x"0c843d0d",
   388 => x"0497f408",
   389 => x"52841208",
   390 => x"70822a70",
   391 => x"81065151",
   392 => x"5170802e",
   393 => x"f0388d72",
   394 => x"0c841208",
   395 => x"70822a70",
   396 => x"81065151",
   397 => x"5170802e",
   398 => x"c038cf39",
   399 => x"fd3d0d75",
   400 => x"70335254",
   401 => x"70802ea9",
   402 => x"387097f4",
   403 => x"08535381",
   404 => x"1454728a",
   405 => x"2e9f3884",
   406 => x"12087082",
   407 => x"2a708106",
   408 => x"51515170",
   409 => x"802ef038",
   410 => x"72720c73",
   411 => x"335372df",
   412 => x"38853d0d",
   413 => x"04841208",
   414 => x"70822a70",
   415 => x"81065151",
   416 => x"5170802e",
   417 => x"f0388d72",
   418 => x"0c841208",
   419 => x"70822a70",
   420 => x"81065151",
   421 => x"5170802e",
   422 => x"ffbd38cc",
   423 => x"39803d0d",
   424 => x"97ec0851",
   425 => x"81ff0b88",
   426 => x"120c823d",
   427 => x"0d04fb3d",
   428 => x"0d8880e0",
   429 => x"870b97ec",
   430 => x"0897f008",
   431 => x"7284130c",
   432 => x"565755af",
   433 => x"d7c20b94",
   434 => x"150c850b",
   435 => x"98150c98",
   436 => x"14087081",
   437 => x"06515372",
   438 => x"f638749f",
   439 => x"2a751007",
   440 => x"7084180c",
   441 => x"55afd7c2",
   442 => x"0b94150c",
   443 => x"850b9815",
   444 => x"0cdd39fe",
   445 => x"3d0d97f0",
   446 => x"085382fd",
   447 => x"bc900ba4",
   448 => x"140c97f4",
   449 => x"0852a813",
   450 => x"08708106",
   451 => x"515170f6",
   452 => x"38841208",
   453 => x"70822a70",
   454 => x"81065151",
   455 => x"5170802e",
   456 => x"f03880e1",
   457 => x"720c850b",
   458 => x"a8140ca8",
   459 => x"13087081",
   460 => x"06515170",
   461 => x"d138da39",
   462 => x"ff3d0d97",
   463 => x"ec085271",
   464 => x"08708f06",
   465 => x"7071842b",
   466 => x"0784150c",
   467 => x"51517108",
   468 => x"708f0670",
   469 => x"71842b07",
   470 => x"84150c51",
   471 => x"51e139fa",
   472 => x"3d0d97f0",
   473 => x"0854870b",
   474 => x"84150c97",
   475 => x"f40855b6",
   476 => x"0b8c160c",
   477 => x"830b8816",
   478 => x"0c97800b",
   479 => x"97803354",
   480 => x"5772802e",
   481 => x"a6387256",
   482 => x"81175775",
   483 => x"8a2e818e",
   484 => x"38841508",
   485 => x"70822a70",
   486 => x"81065151",
   487 => x"5372802e",
   488 => x"f0387575",
   489 => x"0c763356",
   490 => x"75de3897",
   491 => x"980b9798",
   492 => x"33545772",
   493 => x"802ea638",
   494 => x"72568117",
   495 => x"57758a2e",
   496 => x"81853884",
   497 => x"15087082",
   498 => x"2a708106",
   499 => x"51515372",
   500 => x"802ef038",
   501 => x"75750c76",
   502 => x"335675de",
   503 => x"3897ec08",
   504 => x"5681ff0b",
   505 => x"88170c88",
   506 => x"80e08770",
   507 => x"84180c55",
   508 => x"afd7c20b",
   509 => x"94150c85",
   510 => x"0b98150c",
   511 => x"98140881",
   512 => x"065776f8",
   513 => x"38749f2a",
   514 => x"75100770",
   515 => x"84180c55",
   516 => x"afd7c20b",
   517 => x"94150c85",
   518 => x"0b98150c",
   519 => x"df398415",
   520 => x"0870822a",
   521 => x"70810651",
   522 => x"51537280",
   523 => x"2ef0388d",
   524 => x"750c8415",
   525 => x"0870822a",
   526 => x"70810651",
   527 => x"51537280",
   528 => x"2efece38",
   529 => x"fedc3984",
   530 => x"15087082",
   531 => x"2a708106",
   532 => x"51515372",
   533 => x"802ef038",
   534 => x"8d750c84",
   535 => x"15087082",
   536 => x"2a708106",
   537 => x"51515372",
   538 => x"802efed7",
   539 => x"38fee539",
   540 => x"8c08028c",
   541 => x"0cf93d0d",
   542 => x"800b8c08",
   543 => x"fc050c8c",
   544 => x"08880508",
   545 => x"8025ab38",
   546 => x"8c088805",
   547 => x"08308c08",
   548 => x"88050c80",
   549 => x"0b8c08f4",
   550 => x"050c8c08",
   551 => x"fc050888",
   552 => x"38810b8c",
   553 => x"08f4050c",
   554 => x"8c08f405",
   555 => x"088c08fc",
   556 => x"050c8c08",
   557 => x"8c050880",
   558 => x"25ab388c",
   559 => x"088c0508",
   560 => x"308c088c",
   561 => x"050c800b",
   562 => x"8c08f005",
   563 => x"0c8c08fc",
   564 => x"05088838",
   565 => x"810b8c08",
   566 => x"f0050c8c",
   567 => x"08f00508",
   568 => x"8c08fc05",
   569 => x"0c80538c",
   570 => x"088c0508",
   571 => x"528c0888",
   572 => x"05085181",
   573 => x"a73f8008",
   574 => x"708c08f8",
   575 => x"050c548c",
   576 => x"08fc0508",
   577 => x"802e8c38",
   578 => x"8c08f805",
   579 => x"08308c08",
   580 => x"f8050c8c",
   581 => x"08f80508",
   582 => x"70800c54",
   583 => x"893d0d8c",
   584 => x"0c048c08",
   585 => x"028c0cfb",
   586 => x"3d0d800b",
   587 => x"8c08fc05",
   588 => x"0c8c0888",
   589 => x"05088025",
   590 => x"93388c08",
   591 => x"88050830",
   592 => x"8c088805",
   593 => x"0c810b8c",
   594 => x"08fc050c",
   595 => x"8c088c05",
   596 => x"0880258c",
   597 => x"388c088c",
   598 => x"0508308c",
   599 => x"088c050c",
   600 => x"81538c08",
   601 => x"8c050852",
   602 => x"8c088805",
   603 => x"0851ad3f",
   604 => x"8008708c",
   605 => x"08f8050c",
   606 => x"548c08fc",
   607 => x"0508802e",
   608 => x"8c388c08",
   609 => x"f8050830",
   610 => x"8c08f805",
   611 => x"0c8c08f8",
   612 => x"05087080",
   613 => x"0c54873d",
   614 => x"0d8c0c04",
   615 => x"8c08028c",
   616 => x"0cfd3d0d",
   617 => x"810b8c08",
   618 => x"fc050c80",
   619 => x"0b8c08f8",
   620 => x"050c8c08",
   621 => x"8c05088c",
   622 => x"08880508",
   623 => x"27ac388c",
   624 => x"08fc0508",
   625 => x"802ea338",
   626 => x"800b8c08",
   627 => x"8c050824",
   628 => x"99388c08",
   629 => x"8c050810",
   630 => x"8c088c05",
   631 => x"0c8c08fc",
   632 => x"0508108c",
   633 => x"08fc050c",
   634 => x"c9398c08",
   635 => x"fc050880",
   636 => x"2e80c938",
   637 => x"8c088c05",
   638 => x"088c0888",
   639 => x"050826a1",
   640 => x"388c0888",
   641 => x"05088c08",
   642 => x"8c050831",
   643 => x"8c088805",
   644 => x"0c8c08f8",
   645 => x"05088c08",
   646 => x"fc050807",
   647 => x"8c08f805",
   648 => x"0c8c08fc",
   649 => x"0508812a",
   650 => x"8c08fc05",
   651 => x"0c8c088c",
   652 => x"0508812a",
   653 => x"8c088c05",
   654 => x"0cffaf39",
   655 => x"8c089005",
   656 => x"08802e8f",
   657 => x"388c0888",
   658 => x"0508708c",
   659 => x"08f4050c",
   660 => x"518d398c",
   661 => x"08f80508",
   662 => x"708c08f4",
   663 => x"050c518c",
   664 => x"08f40508",
   665 => x"800c853d",
   666 => x"0d8c0c04",
   667 => x"fd3d0d80",
   668 => x"0b97e008",
   669 => x"54547281",
   670 => x"2e983873",
   671 => x"9fa00cf3",
   672 => x"de3ff2fc",
   673 => x"3f97f852",
   674 => x"8151f9d3",
   675 => x"3f800851",
   676 => x"9e3f729f",
   677 => x"a00cf3c7",
   678 => x"3ff2e53f",
   679 => x"97f85281",
   680 => x"51f9bc3f",
   681 => x"80085187",
   682 => x"3f00ff39",
   683 => x"00ff39f7",
   684 => x"3d0d7b97",
   685 => x"fc0882c8",
   686 => x"11085a54",
   687 => x"5a77802e",
   688 => x"80d93881",
   689 => x"88188419",
   690 => x"08ff0581",
   691 => x"712b5955",
   692 => x"59807424",
   693 => x"80e93880",
   694 => x"7424b538",
   695 => x"73822b78",
   696 => x"11880556",
   697 => x"56818019",
   698 => x"08770653",
   699 => x"72802eb5",
   700 => x"38781670",
   701 => x"08535379",
   702 => x"51740853",
   703 => x"722dff14",
   704 => x"fc17fc17",
   705 => x"79812c5a",
   706 => x"57575473",
   707 => x"8025d638",
   708 => x"77085877",
   709 => x"ffad3897",
   710 => x"fc0853bc",
   711 => x"1308a538",
   712 => x"7951ff85",
   713 => x"3f740853",
   714 => x"722dff14",
   715 => x"fc17fc17",
   716 => x"79812c5a",
   717 => x"57575473",
   718 => x"8025ffa9",
   719 => x"38d23980",
   720 => x"57ff9439",
   721 => x"7251bc13",
   722 => x"0853722d",
   723 => x"7951fed9",
   724 => x"3fff3d0d",
   725 => x"9f800bfc",
   726 => x"05700852",
   727 => x"5270ff2e",
   728 => x"9138702d",
   729 => x"fc127008",
   730 => x"525270ff",
   731 => x"2e098106",
   732 => x"f138833d",
   733 => x"0d0404f2",
   734 => x"cb3f0400",
   735 => x"00000040",
   736 => x"536f432c",
   737 => x"205a5055",
   738 => x"20746573",
   739 => x"74207072",
   740 => x"6f677261",
   741 => x"6d0a0000",
   742 => x"636f6d70",
   743 => x"696c6564",
   744 => x"3a204175",
   745 => x"67202034",
   746 => x"20323031",
   747 => x"30202020",
   748 => x"31373a34",
   749 => x"363a3138",
   750 => x"0a000000",
   751 => x"64756d6d",
   752 => x"792e6578",
   753 => x"65000000",
   754 => x"43000000",
   755 => x"00ffffff",
   756 => x"ff00ffff",
   757 => x"ffff00ff",
   758 => x"ffffff00",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000f88",
   763 => x"80000800",
   764 => x"80000200",
   765 => x"80000100",
   766 => x"00000bbc",
   767 => x"00000c00",
   768 => x"00000000",
   769 => x"00000e68",
   770 => x"00000ec4",
   771 => x"00000f20",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000bc8",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
   785 => x"00000000",
   786 => x"00000000",
   787 => x"00000000",
   788 => x"00000000",
   789 => x"00000000",
   790 => x"00000000",
   791 => x"00000000",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
   799 => x"00000000",
   800 => x"00000000",
   801 => x"00000000",
   802 => x"00000000",
   803 => x"00000000",
   804 => x"00000000",
   805 => x"00000000",
   806 => x"00000000",
   807 => x"00000000",
   808 => x"00000000",
   809 => x"00000000",
   810 => x"00000001",
   811 => x"330eabcd",
   812 => x"1234e66d",
   813 => x"deec0005",
   814 => x"000b0000",
   815 => x"00000000",
   816 => x"00000000",
   817 => x"00000000",
   818 => x"00000000",
   819 => x"00000000",
   820 => x"00000000",
   821 => x"00000000",
   822 => x"00000000",
   823 => x"00000000",
   824 => x"00000000",
   825 => x"00000000",
   826 => x"00000000",
   827 => x"00000000",
   828 => x"00000000",
   829 => x"00000000",
   830 => x"00000000",
   831 => x"00000000",
   832 => x"00000000",
   833 => x"00000000",
   834 => x"00000000",
   835 => x"00000000",
   836 => x"00000000",
   837 => x"00000000",
   838 => x"00000000",
   839 => x"00000000",
   840 => x"00000000",
   841 => x"00000000",
   842 => x"00000000",
   843 => x"00000000",
   844 => x"00000000",
   845 => x"00000000",
   846 => x"00000000",
   847 => x"00000000",
   848 => x"00000000",
   849 => x"00000000",
   850 => x"00000000",
   851 => x"00000000",
   852 => x"00000000",
   853 => x"00000000",
   854 => x"00000000",
   855 => x"00000000",
   856 => x"00000000",
   857 => x"00000000",
   858 => x"00000000",
   859 => x"00000000",
   860 => x"00000000",
   861 => x"00000000",
   862 => x"00000000",
   863 => x"00000000",
   864 => x"00000000",
   865 => x"00000000",
   866 => x"00000000",
   867 => x"00000000",
   868 => x"00000000",
   869 => x"00000000",
   870 => x"00000000",
   871 => x"00000000",
   872 => x"00000000",
   873 => x"00000000",
   874 => x"00000000",
   875 => x"00000000",
   876 => x"00000000",
   877 => x"00000000",
   878 => x"00000000",
   879 => x"00000000",
   880 => x"00000000",
   881 => x"00000000",
   882 => x"00000000",
   883 => x"00000000",
   884 => x"00000000",
   885 => x"00000000",
   886 => x"00000000",
   887 => x"00000000",
   888 => x"00000000",
   889 => x"00000000",
   890 => x"00000000",
   891 => x"00000000",
   892 => x"00000000",
   893 => x"00000000",
   894 => x"00000000",
   895 => x"00000000",
   896 => x"00000000",
   897 => x"00000000",
   898 => x"00000000",
   899 => x"00000000",
   900 => x"00000000",
   901 => x"00000000",
   902 => x"00000000",
   903 => x"00000000",
   904 => x"00000000",
   905 => x"00000000",
   906 => x"00000000",
   907 => x"00000000",
   908 => x"00000000",
   909 => x"00000000",
   910 => x"00000000",
   911 => x"00000000",
   912 => x"00000000",
   913 => x"00000000",
   914 => x"00000000",
   915 => x"00000000",
   916 => x"00000000",
   917 => x"00000000",
   918 => x"00000000",
   919 => x"00000000",
   920 => x"00000000",
   921 => x"00000000",
   922 => x"00000000",
   923 => x"00000000",
   924 => x"00000000",
   925 => x"00000000",
   926 => x"00000000",
   927 => x"00000000",
   928 => x"00000000",
   929 => x"00000000",
   930 => x"00000000",
   931 => x"00000000",
   932 => x"00000000",
   933 => x"00000000",
   934 => x"00000000",
   935 => x"00000000",
   936 => x"00000000",
   937 => x"00000000",
   938 => x"00000000",
   939 => x"00000000",
   940 => x"00000000",
   941 => x"00000000",
   942 => x"00000000",
   943 => x"00000000",
   944 => x"00000000",
   945 => x"00000000",
   946 => x"00000000",
   947 => x"00000000",
   948 => x"00000000",
   949 => x"00000000",
   950 => x"00000000",
   951 => x"00000000",
   952 => x"00000000",
   953 => x"00000000",
   954 => x"00000000",
   955 => x"00000000",
   956 => x"00000000",
   957 => x"00000000",
   958 => x"00000000",
   959 => x"00000000",
   960 => x"00000000",
   961 => x"00000000",
   962 => x"00000000",
   963 => x"00000000",
   964 => x"00000000",
   965 => x"00000000",
   966 => x"00000000",
   967 => x"00000000",
   968 => x"00000000",
   969 => x"00000000",
   970 => x"00000000",
   971 => x"00000000",
   972 => x"00000000",
   973 => x"00000000",
   974 => x"00000000",
   975 => x"00000000",
   976 => x"00000000",
   977 => x"00000000",
   978 => x"00000000",
   979 => x"00000000",
   980 => x"00000000",
   981 => x"00000000",
   982 => x"00000000",
   983 => x"00000000",
   984 => x"00000000",
   985 => x"00000000",
   986 => x"00000000",
   987 => x"00000000",
   988 => x"00000000",
   989 => x"00000000",
   990 => x"00000000",
   991 => x"ffffffff",
   992 => x"00000000",
   993 => x"ffffffff",
   994 => x"00000000",
   995 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
