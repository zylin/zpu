-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80ebe00c",
     3 => x"3a0b0b80",
     4 => x"dbfa0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80dcc32d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80eb",
   162 => x"cc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80d6",
   171 => x"e52d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80d8",
   179 => x"972d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80ebdc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"d5e43f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80ebdc08",
   281 => x"802ea438",
   282 => x"80ebe008",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80f3",
   286 => x"a00c82a0",
   287 => x"800b80f3",
   288 => x"a40c8290",
   289 => x"800b80f3",
   290 => x"a80c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"f3a00cf8",
   294 => x"80808280",
   295 => x"0b80f3a4",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"f3a80c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80f3a00c",
   302 => x"80c0a880",
   303 => x"940b80f3",
   304 => x"a40c0b0b",
   305 => x"80de980b",
   306 => x"80f3a80c",
   307 => x"04ff3d0d",
   308 => x"80f3ac33",
   309 => x"5170a738",
   310 => x"80ebe808",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"ebe80c70",
   315 => x"2d80ebe8",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80f3",
   319 => x"ac34833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80f39c08",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"f39c510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404f83d",
   333 => x"0d7a7c59",
   334 => x"53807356",
   335 => x"57767324",
   336 => x"80de3877",
   337 => x"17548a52",
   338 => x"745180cb",
   339 => x"f33f8008",
   340 => x"b0055372",
   341 => x"74348117",
   342 => x"578a5274",
   343 => x"5180cbbb",
   344 => x"3f800855",
   345 => x"8008dc38",
   346 => x"8008779f",
   347 => x"2a187081",
   348 => x"2c5b5656",
   349 => x"8079259e",
   350 => x"387717ff",
   351 => x"05557518",
   352 => x"70335553",
   353 => x"74337334",
   354 => x"73753481",
   355 => x"16ff1656",
   356 => x"56787624",
   357 => x"e9387618",
   358 => x"56807634",
   359 => x"8a3d0d04",
   360 => x"ad787081",
   361 => x"055a3472",
   362 => x"30781855",
   363 => x"558a5274",
   364 => x"5180cb8c",
   365 => x"3f8008b0",
   366 => x"05537274",
   367 => x"34811757",
   368 => x"8a527451",
   369 => x"80cad43f",
   370 => x"80085580",
   371 => x"08fef438",
   372 => x"ff9639f9",
   373 => x"3d0d7970",
   374 => x"71337081",
   375 => x"ff065455",
   376 => x"55557080",
   377 => x"2eb13880",
   378 => x"ec840852",
   379 => x"7281ff06",
   380 => x"81155553",
   381 => x"728a2e80",
   382 => x"f5388412",
   383 => x"0870822a",
   384 => x"81065257",
   385 => x"70802ef2",
   386 => x"3872720c",
   387 => x"73337081",
   388 => x"ff065953",
   389 => x"77d63874",
   390 => x"75335256",
   391 => x"70802e80",
   392 => x"c9387080",
   393 => x"ebfc0859",
   394 => x"53811680",
   395 => x"f3b43370",
   396 => x"81ff0670",
   397 => x"10101180",
   398 => x"f3b83370",
   399 => x"81ff0672",
   400 => x"90291170",
   401 => x"882b7a07",
   402 => x"7f0c5359",
   403 => x"59545458",
   404 => x"56728a2e",
   405 => x"be387380",
   406 => x"cf2eb838",
   407 => x"81155372",
   408 => x"80f3b834",
   409 => x"75335372",
   410 => x"c038893d",
   411 => x"0d048412",
   412 => x"0870822a",
   413 => x"81065758",
   414 => x"75802ef2",
   415 => x"388d720c",
   416 => x"84120870",
   417 => x"822a8106",
   418 => x"52577080",
   419 => x"2efeeb38",
   420 => x"fef73971",
   421 => x"a3269938",
   422 => x"81175271",
   423 => x"80f3b434",
   424 => x"800b80f3",
   425 => x"b8347533",
   426 => x"5372fefd",
   427 => x"38ffbb39",
   428 => x"800b80f3",
   429 => x"b434800b",
   430 => x"80f3b834",
   431 => x"e939fd3d",
   432 => x"0d80ebf8",
   433 => x"085480d5",
   434 => x"0b84150c",
   435 => x"80ec8408",
   436 => x"52841208",
   437 => x"81065170",
   438 => x"802ef638",
   439 => x"71087081",
   440 => x"ff06f611",
   441 => x"52545170",
   442 => x"ae268c38",
   443 => x"70101080",
   444 => x"e9cc0551",
   445 => x"70080484",
   446 => x"12087082",
   447 => x"2a708106",
   448 => x"51515170",
   449 => x"802ef038",
   450 => x"ab720c72",
   451 => x"8a2eaa38",
   452 => x"84120870",
   453 => x"822a7081",
   454 => x"06515151",
   455 => x"70802ef0",
   456 => x"3872720c",
   457 => x"84120870",
   458 => x"822a8106",
   459 => x"51537280",
   460 => x"2ef238ad",
   461 => x"720cff99",
   462 => x"39841208",
   463 => x"70822a70",
   464 => x"81065151",
   465 => x"5170802e",
   466 => x"f0388d72",
   467 => x"0c841208",
   468 => x"70822a70",
   469 => x"81065151",
   470 => x"5170802e",
   471 => x"ffb238c1",
   472 => x"3981ff0b",
   473 => x"84150cfe",
   474 => x"e83980ff",
   475 => x"0b84150c",
   476 => x"fedf39bf",
   477 => x"0b84150c",
   478 => x"fed7399f",
   479 => x"0b84150c",
   480 => x"fecf398f",
   481 => x"0b84150c",
   482 => x"fec73987",
   483 => x"0b84150c",
   484 => x"febf3983",
   485 => x"0b84150c",
   486 => x"feb73981",
   487 => x"0b84150c",
   488 => x"feaf3980",
   489 => x"0b84150c",
   490 => x"fea739e6",
   491 => x"3d0d80eb",
   492 => x"fc085580",
   493 => x"0b84160c",
   494 => x"fe800a0b",
   495 => x"88160c80",
   496 => x"0b80f3b4",
   497 => x"34800b80",
   498 => x"f3b83497",
   499 => x"3d705380",
   500 => x"ebf0088c",
   501 => x"11085355",
   502 => x"5bfad73f",
   503 => x"80e1b40b",
   504 => x"80e1b433",
   505 => x"555a7380",
   506 => x"2e80cc38",
   507 => x"80ebfc08",
   508 => x"74575c81",
   509 => x"1a80f3b4",
   510 => x"337081ff",
   511 => x"06701010",
   512 => x"1180f3b8",
   513 => x"337081ff",
   514 => x"06729029",
   515 => x"1170882b",
   516 => x"7d07630c",
   517 => x"445c5c42",
   518 => x"575a5a75",
   519 => x"8a2e87b3",
   520 => x"387680cf",
   521 => x"2e87ac38",
   522 => x"81185776",
   523 => x"80f3b834",
   524 => x"79335675",
   525 => x"ffbd387a",
   526 => x"7b33555a",
   527 => x"73802e80",
   528 => x"cc3880eb",
   529 => x"fc087457",
   530 => x"5b811a80",
   531 => x"f3b43370",
   532 => x"81ff0670",
   533 => x"10101180",
   534 => x"f3b83370",
   535 => x"81ff0672",
   536 => x"90291170",
   537 => x"882b7d07",
   538 => x"620c465c",
   539 => x"5c57575a",
   540 => x"5a758a2e",
   541 => x"86fb3876",
   542 => x"80cf2e86",
   543 => x"f4388118",
   544 => x"597880f3",
   545 => x"b8347933",
   546 => x"5675ffbd",
   547 => x"3880e1c4",
   548 => x"0b80e1c4",
   549 => x"33555a73",
   550 => x"802e80cc",
   551 => x"3880ebfc",
   552 => x"0874575b",
   553 => x"811a80f3",
   554 => x"b4337081",
   555 => x"ff067010",
   556 => x"101180f3",
   557 => x"b8337081",
   558 => x"ff067290",
   559 => x"29117088",
   560 => x"2b7d0762",
   561 => x"0c445c5c",
   562 => x"42575a5a",
   563 => x"758a2e85",
   564 => x"e4387680",
   565 => x"cf2e85dd",
   566 => x"38811856",
   567 => x"7580f3b8",
   568 => x"34793356",
   569 => x"75ffbd38",
   570 => x"80ebf008",
   571 => x"7008963d",
   572 => x"5b585a8b",
   573 => x"5380de9c",
   574 => x"52785180",
   575 => x"c8e33f82",
   576 => x"02840580",
   577 => x"cd055956",
   578 => x"768f0654",
   579 => x"73892685",
   580 => x"88387518",
   581 => x"b0155555",
   582 => x"73753476",
   583 => x"842aff17",
   584 => x"7081ff06",
   585 => x"585c5775",
   586 => x"df387879",
   587 => x"33555a73",
   588 => x"802e80cc",
   589 => x"3880ebfc",
   590 => x"0874575b",
   591 => x"811a80f3",
   592 => x"b4337081",
   593 => x"ff067010",
   594 => x"101180f3",
   595 => x"b8337081",
   596 => x"ff067290",
   597 => x"29117088",
   598 => x"2b7d0762",
   599 => x"0c465c5c",
   600 => x"57575a5a",
   601 => x"758a2e87",
   602 => x"e9387680",
   603 => x"cf2e87e2",
   604 => x"38811859",
   605 => x"7880f3b8",
   606 => x"34793356",
   607 => x"75ffbd38",
   608 => x"80e1d00b",
   609 => x"80e1d033",
   610 => x"555a7380",
   611 => x"2e80cc38",
   612 => x"80ebfc08",
   613 => x"74575b81",
   614 => x"1a80f3b4",
   615 => x"337081ff",
   616 => x"06701010",
   617 => x"1180f3b8",
   618 => x"337081ff",
   619 => x"06729029",
   620 => x"1170882b",
   621 => x"7d07620c",
   622 => x"445c5c42",
   623 => x"575a5a75",
   624 => x"8a2e87ac",
   625 => x"387680cf",
   626 => x"2e87a538",
   627 => x"81185574",
   628 => x"80f3b834",
   629 => x"79335675",
   630 => x"ffbd3889",
   631 => x"0a5c8070",
   632 => x"933d028c",
   633 => x"0580c105",
   634 => x"41425e5f",
   635 => x"7cbf0656",
   636 => x"7585d538",
   637 => x"80e1980b",
   638 => x"80e19833",
   639 => x"555a7380",
   640 => x"2e80cc38",
   641 => x"80ebfc08",
   642 => x"74575b81",
   643 => x"1a80f3b4",
   644 => x"337081ff",
   645 => x"06701010",
   646 => x"1180f3b8",
   647 => x"337081ff",
   648 => x"06729029",
   649 => x"1170882b",
   650 => x"7d07620c",
   651 => x"535c5c57",
   652 => x"575a5a75",
   653 => x"8a2e84c7",
   654 => x"387680cf",
   655 => x"2e84c038",
   656 => x"81185978",
   657 => x"80f3b834",
   658 => x"79335675",
   659 => x"ffbd387b",
   660 => x"568b5380",
   661 => x"de9c527f",
   662 => x"5180c685",
   663 => x"3f885775",
   664 => x"8f065473",
   665 => x"892683d2",
   666 => x"38761eb0",
   667 => x"15555573",
   668 => x"75347584",
   669 => x"2aff1870",
   670 => x"81ff0659",
   671 => x"5b5676df",
   672 => x"387f6033",
   673 => x"555a7380",
   674 => x"2e85bf38",
   675 => x"80ebfc08",
   676 => x"74575b81",
   677 => x"1a80f3b4",
   678 => x"337081ff",
   679 => x"06701010",
   680 => x"1180f3b8",
   681 => x"337081ff",
   682 => x"06729029",
   683 => x"1170882b",
   684 => x"7d07620c",
   685 => x"535c5c57",
   686 => x"575a5a75",
   687 => x"8a2e83a1",
   688 => x"387680cf",
   689 => x"2e839a38",
   690 => x"81185574",
   691 => x"80f3b834",
   692 => x"79335675",
   693 => x"ffbd3880",
   694 => x"e1d40b80",
   695 => x"e1d43355",
   696 => x"5a73802e",
   697 => x"80c73873",
   698 => x"56811a80",
   699 => x"f3b43370",
   700 => x"81ff0670",
   701 => x"10101180",
   702 => x"f3b83370",
   703 => x"81ff0672",
   704 => x"90291170",
   705 => x"882b7d07",
   706 => x"620c535c",
   707 => x"5c57575a",
   708 => x"5a758a2e",
   709 => x"82ad3876",
   710 => x"80cf2e82",
   711 => x"a6388118",
   712 => x"577680f3",
   713 => x"b8347933",
   714 => x"5675ffbd",
   715 => x"387b087c",
   716 => x"32703071",
   717 => x"07709f2a",
   718 => x"7081ff06",
   719 => x"b0117081",
   720 => x"ff0680f3",
   721 => x"b4337081",
   722 => x"ff067010",
   723 => x"101180f3",
   724 => x"b8337081",
   725 => x"ff067290",
   726 => x"29117088",
   727 => x"2b770767",
   728 => x"0c535a57",
   729 => x"5c5d525a",
   730 => x"5d525a5b",
   731 => x"57748a2e",
   732 => x"83a43876",
   733 => x"80cf2e83",
   734 => x"9d388118",
   735 => x"547380f3",
   736 => x"b834791f",
   737 => x"811d811f",
   738 => x"5f5d5f8f",
   739 => x"ff7d27fc",
   740 => x"db387e80",
   741 => x"0c9c3d0d",
   742 => x"047518b7",
   743 => x"15555573",
   744 => x"75347684",
   745 => x"2aff1770",
   746 => x"81ff0658",
   747 => x"5c5775fa",
   748 => x"d738faf6",
   749 => x"3974a326",
   750 => x"80f13881",
   751 => x"19557480",
   752 => x"f3b43480",
   753 => x"0b80f3b8",
   754 => x"34793356",
   755 => x"75f9d538",
   756 => x"fa963974",
   757 => x"a32680c4",
   758 => x"38811956",
   759 => x"7580f3b4",
   760 => x"34800b80",
   761 => x"f3b83479",
   762 => x"335675f8",
   763 => x"8638f8c7",
   764 => x"3974a326",
   765 => x"99388119",
   766 => x"587780f3",
   767 => x"b434800b",
   768 => x"80f3b834",
   769 => x"79335675",
   770 => x"f8bf38f9",
   771 => x"8039800b",
   772 => x"80f3b434",
   773 => x"800b80f3",
   774 => x"b834e939",
   775 => x"800b80f3",
   776 => x"b434800b",
   777 => x"80f3b834",
   778 => x"ffbd3980",
   779 => x"0b80f3b4",
   780 => x"34800b80",
   781 => x"f3b834ff",
   782 => x"9039761e",
   783 => x"b7155555",
   784 => x"fcad3974",
   785 => x"a32680f1",
   786 => x"38811956",
   787 => x"7580f3b4",
   788 => x"34800b80",
   789 => x"f3b83479",
   790 => x"335675fd",
   791 => x"8c38fdcd",
   792 => x"3974a326",
   793 => x"80c43881",
   794 => x"19587780",
   795 => x"f3b43480",
   796 => x"0b80f3b8",
   797 => x"34793356",
   798 => x"75fc9838",
   799 => x"fcd93974",
   800 => x"a3269938",
   801 => x"81195776",
   802 => x"80f3b434",
   803 => x"800b80f3",
   804 => x"b8347933",
   805 => x"5675faf3",
   806 => x"38fbb439",
   807 => x"800b80f3",
   808 => x"b434800b",
   809 => x"80f3b834",
   810 => x"e939800b",
   811 => x"80f3b434",
   812 => x"800b80f3",
   813 => x"b834ffbd",
   814 => x"39800b80",
   815 => x"f3b43480",
   816 => x"0b80f3b8",
   817 => x"34ff9039",
   818 => x"80ebfc08",
   819 => x"7c087d32",
   820 => x"70307107",
   821 => x"709f2a70",
   822 => x"81ff06b0",
   823 => x"117081ff",
   824 => x"0680f3b4",
   825 => x"337081ff",
   826 => x"06701010",
   827 => x"1180f3b8",
   828 => x"337081ff",
   829 => x"06729029",
   830 => x"1170882b",
   831 => x"77077d0c",
   832 => x"535a575d",
   833 => x"5e525b5e",
   834 => x"525b5c58",
   835 => x"5b748a2e",
   836 => x"098106fc",
   837 => x"de3875a3",
   838 => x"26a23881",
   839 => x"195b7a80",
   840 => x"f3b43480",
   841 => x"0b80f3b8",
   842 => x"34791f81",
   843 => x"1d811f5f",
   844 => x"5d5f8fff",
   845 => x"7d27f9b4",
   846 => x"38fcd739",
   847 => x"800b80f3",
   848 => x"b434800b",
   849 => x"80f3b834",
   850 => x"e03980eb",
   851 => x"fc085bfb",
   852 => x"863974a3",
   853 => x"2680c438",
   854 => x"81195776",
   855 => x"80f3b434",
   856 => x"800b80f3",
   857 => x"b8347933",
   858 => x"5675f7d0",
   859 => x"38f89139",
   860 => x"74a32699",
   861 => x"38811958",
   862 => x"7780f3b4",
   863 => x"34800b80",
   864 => x"f3b83479",
   865 => x"335675f8",
   866 => x"8e38f8cf",
   867 => x"39800b80",
   868 => x"f3b43480",
   869 => x"0b80f3b8",
   870 => x"34e93980",
   871 => x"0b80f3b4",
   872 => x"34800b80",
   873 => x"f3b834ff",
   874 => x"bd39dd3d",
   875 => x"0d80e1d8",
   876 => x"51f0a03f",
   877 => x"80ebec08",
   878 => x"700880e1",
   879 => x"e8535d55",
   880 => x"f0913fa0",
   881 => x"3d70537c",
   882 => x"81ffff06",
   883 => x"525deee2",
   884 => x"3f7c51ef",
   885 => x"fe3f80e1",
   886 => x"fc51eff7",
   887 => x"3f7b8f2a",
   888 => x"81069e3d",
   889 => x"5a568b53",
   890 => x"80de9c52",
   891 => x"7851bef1",
   892 => x"3f820284",
   893 => x"0580f105",
   894 => x"5957758f",
   895 => x"06547389",
   896 => x"2687fc38",
   897 => x"7618b015",
   898 => x"55557375",
   899 => x"3475842a",
   900 => x"ff187081",
   901 => x"ff06595b",
   902 => x"5676df38",
   903 => x"78793355",
   904 => x"5773802e",
   905 => x"a9387380",
   906 => x"ec840856",
   907 => x"56811757",
   908 => x"758a2e87",
   909 => x"e6388415",
   910 => x"0870822a",
   911 => x"81065b5b",
   912 => x"79802ef2",
   913 => x"3875750c",
   914 => x"76335675",
   915 => x"e0387879",
   916 => x"33555a73",
   917 => x"802e80cc",
   918 => x"387380eb",
   919 => x"fc085c56",
   920 => x"811a80f3",
   921 => x"b4337081",
   922 => x"ff067010",
   923 => x"101180f3",
   924 => x"b8337081",
   925 => x"ff067290",
   926 => x"29117088",
   927 => x"2b7d0762",
   928 => x"0c535c5c",
   929 => x"57575a5a",
   930 => x"758a2e87",
   931 => x"cf387680",
   932 => x"cf2e87c8",
   933 => x"38811857",
   934 => x"7680f3b8",
   935 => x"34793356",
   936 => x"75ffbd38",
   937 => x"80e29051",
   938 => x"eea93f7b",
   939 => x"902a8106",
   940 => x"9b3d5a56",
   941 => x"8b5380de",
   942 => x"9c527851",
   943 => x"bda33f82",
   944 => x"02840580",
   945 => x"e5055957",
   946 => x"758f0654",
   947 => x"73892686",
   948 => x"ef387618",
   949 => x"b0155555",
   950 => x"73753475",
   951 => x"842aff18",
   952 => x"7081ff06",
   953 => x"59565676",
   954 => x"df387879",
   955 => x"33555773",
   956 => x"802ea938",
   957 => x"80ec8408",
   958 => x"74575581",
   959 => x"1757758a",
   960 => x"2e878438",
   961 => x"84150870",
   962 => x"822a8106",
   963 => x"55587380",
   964 => x"2ef23875",
   965 => x"750c7633",
   966 => x"5675e038",
   967 => x"78793355",
   968 => x"5a73802e",
   969 => x"80cc3880",
   970 => x"ebfc0874",
   971 => x"575b811a",
   972 => x"80f3b433",
   973 => x"7081ff06",
   974 => x"70101011",
   975 => x"80f3b833",
   976 => x"7081ff06",
   977 => x"72902911",
   978 => x"70882b7d",
   979 => x"07620c53",
   980 => x"5c5c5757",
   981 => x"5a5a758a",
   982 => x"2e8fd738",
   983 => x"7680cf2e",
   984 => x"8fd03881",
   985 => x"18577680",
   986 => x"f3b83479",
   987 => x"335675ff",
   988 => x"bd3880e2",
   989 => x"a451ecdb",
   990 => x"3f7b952a",
   991 => x"83065473",
   992 => x"812e90bd",
   993 => x"38817426",
   994 => x"908f3873",
   995 => x"822e90cf",
   996 => x"3873832e",
   997 => x"8ce73880",
   998 => x"e2b851ec",
   999 => x"b63f7c52",
  1000 => x"7b972a87",
  1001 => x"06830581",
  1002 => x"712b525a",
  1003 => x"eb843f7c",
  1004 => x"51eca03f",
  1005 => x"80e2cc51",
  1006 => x"ec993f80",
  1007 => x"e2d451ec",
  1008 => x"923f7c52",
  1009 => x"7b9a2a81",
  1010 => x"06810551",
  1011 => x"eae43f7c",
  1012 => x"51ec803f",
  1013 => x"80e2e851",
  1014 => x"ebf93f7c",
  1015 => x"527b9b2a",
  1016 => x"87068305",
  1017 => x"51eacb3f",
  1018 => x"7c51ebe7",
  1019 => x"3f80e2fc",
  1020 => x"51ebe03f",
  1021 => x"7c527b9e",
  1022 => x"2a820751",
  1023 => x"eab43f7c",
  1024 => x"51ebd03f",
  1025 => x"80e39051",
  1026 => x"ebc93f7b",
  1027 => x"9f2a983d",
  1028 => x"5a568b53",
  1029 => x"80de9c52",
  1030 => x"7851bac5",
  1031 => x"3f820284",
  1032 => x"0580d905",
  1033 => x"5957758f",
  1034 => x"06547389",
  1035 => x"268ce738",
  1036 => x"7618b015",
  1037 => x"55557375",
  1038 => x"3475842a",
  1039 => x"ff187081",
  1040 => x"ff06595d",
  1041 => x"5676df38",
  1042 => x"78793355",
  1043 => x"5773802e",
  1044 => x"a93880ec",
  1045 => x"84087457",
  1046 => x"55811757",
  1047 => x"758a2e84",
  1048 => x"cb388415",
  1049 => x"0870822a",
  1050 => x"81065954",
  1051 => x"77802ef2",
  1052 => x"3875750c",
  1053 => x"76335675",
  1054 => x"e0387879",
  1055 => x"33555a73",
  1056 => x"802e80cc",
  1057 => x"3880ebfc",
  1058 => x"0874575b",
  1059 => x"811a80f3",
  1060 => x"b4337081",
  1061 => x"ff067010",
  1062 => x"101180f3",
  1063 => x"b8337081",
  1064 => x"ff067290",
  1065 => x"29117088",
  1066 => x"2b7d0762",
  1067 => x"0c5a5c5c",
  1068 => x"5f575a5a",
  1069 => x"758a2e8c",
  1070 => x"9f387680",
  1071 => x"cf2e8c98",
  1072 => x"38811857",
  1073 => x"7680f3b8",
  1074 => x"34793356",
  1075 => x"75ffbd38",
  1076 => x"80ebec08",
  1077 => x"84110880",
  1078 => x"e3a45356",
  1079 => x"58e9f43f",
  1080 => x"7c52749f",
  1081 => x"ff0651e8",
  1082 => x"c93f7c51",
  1083 => x"e9e53f80",
  1084 => x"e3b851e9",
  1085 => x"de3f7c52",
  1086 => x"748c2a87",
  1087 => x"06830581",
  1088 => x"712b525b",
  1089 => x"e8ac3f7c",
  1090 => x"51e9c83f",
  1091 => x"80e3cc51",
  1092 => x"e9c13f74",
  1093 => x"8f2a8106",
  1094 => x"953d5a56",
  1095 => x"8b5380de",
  1096 => x"9c527851",
  1097 => x"b8bb3f82",
  1098 => x"02840580",
  1099 => x"cd055957",
  1100 => x"758f0654",
  1101 => x"7389268a",
  1102 => x"f8387618",
  1103 => x"b0155555",
  1104 => x"73753475",
  1105 => x"842aff18",
  1106 => x"7081ff06",
  1107 => x"59555676",
  1108 => x"df387879",
  1109 => x"33555773",
  1110 => x"802ea938",
  1111 => x"80ec8408",
  1112 => x"74575581",
  1113 => x"1757758a",
  1114 => x"2e82e638",
  1115 => x"84150870",
  1116 => x"822a8106",
  1117 => x"595c7780",
  1118 => x"2ef23875",
  1119 => x"750c7633",
  1120 => x"5675e038",
  1121 => x"78793355",
  1122 => x"5a73802e",
  1123 => x"80cc3880",
  1124 => x"ebfc0874",
  1125 => x"575b811a",
  1126 => x"80f3b433",
  1127 => x"7081ff06",
  1128 => x"70101011",
  1129 => x"80f3b833",
  1130 => x"7081ff06",
  1131 => x"72902911",
  1132 => x"70882b7d",
  1133 => x"07620c42",
  1134 => x"5c5c5757",
  1135 => x"5a5a758a",
  1136 => x"2e89f738",
  1137 => x"7680cf2e",
  1138 => x"89f03881",
  1139 => x"18577680",
  1140 => x"f3b83479",
  1141 => x"335675ff",
  1142 => x"bd3880eb",
  1143 => x"ec088811",
  1144 => x"0880e3e0",
  1145 => x"535659e7",
  1146 => x"ea3f7487",
  1147 => x"06547386",
  1148 => x"26828338",
  1149 => x"73101080",
  1150 => x"eb88055b",
  1151 => x"7a080476",
  1152 => x"18b71555",
  1153 => x"55737534",
  1154 => x"75842aff",
  1155 => x"187081ff",
  1156 => x"06595b56",
  1157 => x"76f7e338",
  1158 => x"f8823984",
  1159 => x"15087082",
  1160 => x"2a810659",
  1161 => x"5477802e",
  1162 => x"f2388d75",
  1163 => x"0c841508",
  1164 => x"70822a81",
  1165 => x"065b5b79",
  1166 => x"802ef7fa",
  1167 => x"38f88639",
  1168 => x"7618b715",
  1169 => x"55557375",
  1170 => x"3475842a",
  1171 => x"ff187081",
  1172 => x"ff065956",
  1173 => x"5676f8f0",
  1174 => x"38f98f39",
  1175 => x"74a32699",
  1176 => x"38811956",
  1177 => x"7580f3b4",
  1178 => x"34800b80",
  1179 => x"f3b83479",
  1180 => x"335675f7",
  1181 => x"eb38f8ac",
  1182 => x"39800b80",
  1183 => x"f3b43480",
  1184 => x"0b80f3b8",
  1185 => x"34e93984",
  1186 => x"15087082",
  1187 => x"2a81065b",
  1188 => x"5b79802e",
  1189 => x"f2388d75",
  1190 => x"0c841508",
  1191 => x"70822a81",
  1192 => x"06555873",
  1193 => x"802ef8dc",
  1194 => x"38f8e839",
  1195 => x"84150870",
  1196 => x"822a8106",
  1197 => x"555a7380",
  1198 => x"2ef2388d",
  1199 => x"750c8415",
  1200 => x"0870822a",
  1201 => x"81065954",
  1202 => x"77802efb",
  1203 => x"9538fba1",
  1204 => x"39841508",
  1205 => x"70822a81",
  1206 => x"065d5a7b",
  1207 => x"802ef238",
  1208 => x"8d750c84",
  1209 => x"15087082",
  1210 => x"2a810659",
  1211 => x"5c77802e",
  1212 => x"fcfa38fd",
  1213 => x"863980e3",
  1214 => x"f451e5d7",
  1215 => x"3f80e3fc",
  1216 => x"51e5d03f",
  1217 => x"80e48451",
  1218 => x"e5c93f74",
  1219 => x"832a8306",
  1220 => x"5473812e",
  1221 => x"89a13881",
  1222 => x"74268991",
  1223 => x"3873822e",
  1224 => x"89a93873",
  1225 => x"832e85a7",
  1226 => x"3880e498",
  1227 => x"51e5a43f",
  1228 => x"80e49c51",
  1229 => x"e59d3f74",
  1230 => x"852a8706",
  1231 => x"5473812e",
  1232 => x"85b13881",
  1233 => x"742688db",
  1234 => x"3873822e",
  1235 => x"89873873",
  1236 => x"832e84f1",
  1237 => x"3880e4b0",
  1238 => x"51e4f83f",
  1239 => x"74902a87",
  1240 => x"06547385",
  1241 => x"268c3873",
  1242 => x"101080eb",
  1243 => x"a4055473",
  1244 => x"080480e3",
  1245 => x"f451e4db",
  1246 => x"3f80e4c4",
  1247 => x"51e4d43f",
  1248 => x"7c527493",
  1249 => x"2a830682",
  1250 => x"0751e3a6",
  1251 => x"3f7c51e4",
  1252 => x"c23f80e4",
  1253 => x"d851e4bb",
  1254 => x"3f7c5274",
  1255 => x"942a8f06",
  1256 => x"51e38f3f",
  1257 => x"7c51e4ab",
  1258 => x"3f80e4ec",
  1259 => x"51e4a43f",
  1260 => x"7c527498",
  1261 => x"2a810681",
  1262 => x"0551e2f6",
  1263 => x"3f7c51e4",
  1264 => x"923f80e5",
  1265 => x"8051e48b",
  1266 => x"3f7c5274",
  1267 => x"9e2a8207",
  1268 => x"51e2df3f",
  1269 => x"7c51e3fb",
  1270 => x"3f80e594",
  1271 => x"51e3f43f",
  1272 => x"749f2a92",
  1273 => x"3d5a568b",
  1274 => x"5380de9c",
  1275 => x"527851b2",
  1276 => x"f03f8202",
  1277 => x"840580c1",
  1278 => x"05595775",
  1279 => x"8f065473",
  1280 => x"892685a4",
  1281 => x"387618b0",
  1282 => x"15555573",
  1283 => x"75347584",
  1284 => x"2aff1870",
  1285 => x"81ff0659",
  1286 => x"5e5676df",
  1287 => x"38787933",
  1288 => x"55577380",
  1289 => x"2ea93880",
  1290 => x"ec840874",
  1291 => x"57558117",
  1292 => x"57758a2e",
  1293 => x"82c53884",
  1294 => x"15087082",
  1295 => x"2a81065d",
  1296 => x"5d7b802e",
  1297 => x"f2387575",
  1298 => x"0c763356",
  1299 => x"75e03878",
  1300 => x"7933555a",
  1301 => x"73802e80",
  1302 => x"cc3880eb",
  1303 => x"fc087457",
  1304 => x"5b811a80",
  1305 => x"f3b43370",
  1306 => x"81ff0670",
  1307 => x"10101180",
  1308 => x"f3b83370",
  1309 => x"81ff0672",
  1310 => x"90291170",
  1311 => x"882b7d07",
  1312 => x"620c5a5c",
  1313 => x"5c40575a",
  1314 => x"5a758a2e",
  1315 => x"85863876",
  1316 => x"80cf2e84",
  1317 => x"ff388118",
  1318 => x"567580f3",
  1319 => x"b8347933",
  1320 => x"5675ffbd",
  1321 => x"3880ebec",
  1322 => x"08901108",
  1323 => x"80e5a853",
  1324 => x"5859e29f",
  1325 => x"3f768f3d",
  1326 => x"5a568b53",
  1327 => x"80de9c52",
  1328 => x"7851b19d",
  1329 => x"3f880284",
  1330 => x"05b50559",
  1331 => x"57758f06",
  1332 => x"54738926",
  1333 => x"83c93876",
  1334 => x"18b01555",
  1335 => x"55737534",
  1336 => x"75842aff",
  1337 => x"187081ff",
  1338 => x"06595c56",
  1339 => x"76df3878",
  1340 => x"79335557",
  1341 => x"73802ea9",
  1342 => x"3880ec84",
  1343 => x"08745755",
  1344 => x"81175775",
  1345 => x"8a2e8198",
  1346 => x"38841508",
  1347 => x"70822a81",
  1348 => x"06555b73",
  1349 => x"802ef238",
  1350 => x"75750c76",
  1351 => x"335675e0",
  1352 => x"38787933",
  1353 => x"555a7380",
  1354 => x"2e80cc38",
  1355 => x"80ebfc08",
  1356 => x"74575b81",
  1357 => x"1a80f3b4",
  1358 => x"337081ff",
  1359 => x"06701010",
  1360 => x"1180f3b8",
  1361 => x"337081ff",
  1362 => x"06729029",
  1363 => x"1170882b",
  1364 => x"7d07620c",
  1365 => x"5a5c5c40",
  1366 => x"575a5a75",
  1367 => x"8a2e8396",
  1368 => x"387680cf",
  1369 => x"2e838f38",
  1370 => x"81185675",
  1371 => x"80f3b834",
  1372 => x"79335675",
  1373 => x"ffbd38a5",
  1374 => x"3d0d0484",
  1375 => x"15087082",
  1376 => x"2a81065c",
  1377 => x"587a802e",
  1378 => x"f2388d75",
  1379 => x"0c841508",
  1380 => x"70822a81",
  1381 => x"065d5d7b",
  1382 => x"802efd9b",
  1383 => x"38fda739",
  1384 => x"84150870",
  1385 => x"822a8106",
  1386 => x"5b5c7980",
  1387 => x"2ef2388d",
  1388 => x"750c8415",
  1389 => x"0870822a",
  1390 => x"8106555b",
  1391 => x"73802efe",
  1392 => x"c838fed4",
  1393 => x"3980e5bc",
  1394 => x"51e0883f",
  1395 => x"fb873980",
  1396 => x"e5c051df",
  1397 => x"fe3f80e4",
  1398 => x"9851dff7",
  1399 => x"3f80e49c",
  1400 => x"51dff03f",
  1401 => x"74852a87",
  1402 => x"06547381",
  1403 => x"2e098106",
  1404 => x"fad13880",
  1405 => x"e5c451df",
  1406 => x"da3ffad9",
  1407 => x"3980e5cc",
  1408 => x"51dfd03f",
  1409 => x"80e2b851",
  1410 => x"dfc93f7c",
  1411 => x"527b972a",
  1412 => x"87068305",
  1413 => x"81712b52",
  1414 => x"5ade973f",
  1415 => x"7c51dfb3",
  1416 => x"3f80e2cc",
  1417 => x"51dfac3f",
  1418 => x"80e2d451",
  1419 => x"dfa53f7c",
  1420 => x"527b9a2a",
  1421 => x"81068105",
  1422 => x"51ddf73f",
  1423 => x"7c51df93",
  1424 => x"3f80e2e8",
  1425 => x"51df8c3f",
  1426 => x"7c527b9b",
  1427 => x"2a870683",
  1428 => x"0551ddde",
  1429 => x"3f7c51de",
  1430 => x"fa3f80e2",
  1431 => x"fc51def3",
  1432 => x"3f7c527b",
  1433 => x"9e2a8207",
  1434 => x"51ddc73f",
  1435 => x"7c51dee3",
  1436 => x"3f80e390",
  1437 => x"51dedc3f",
  1438 => x"7b9f2a98",
  1439 => x"3d5a568b",
  1440 => x"5380de9c",
  1441 => x"527851ad",
  1442 => x"d83f8202",
  1443 => x"840580d9",
  1444 => x"055957f3",
  1445 => x"91397618",
  1446 => x"b7155555",
  1447 => x"f3983976",
  1448 => x"18b71555",
  1449 => x"55fcb639",
  1450 => x"7618b715",
  1451 => x"5555fadb",
  1452 => x"397618b7",
  1453 => x"155555f5",
  1454 => x"873974a3",
  1455 => x"2681cb38",
  1456 => x"81195675",
  1457 => x"80f3b434",
  1458 => x"800b80f3",
  1459 => x"b8347933",
  1460 => x"5675f5c2",
  1461 => x"38f68339",
  1462 => x"74a32681",
  1463 => x"9e388119",
  1464 => x"567580f3",
  1465 => x"b434800b",
  1466 => x"80f3b834",
  1467 => x"79335675",
  1468 => x"f39a38f3",
  1469 => x"db3974a3",
  1470 => x"2680f138",
  1471 => x"81195574",
  1472 => x"80f3b434",
  1473 => x"800b80f3",
  1474 => x"b8347933",
  1475 => x"5675fca3",
  1476 => x"38fce439",
  1477 => x"74a32680",
  1478 => x"c4388119",
  1479 => x"557480f3",
  1480 => x"b434800b",
  1481 => x"80f3b834",
  1482 => x"79335675",
  1483 => x"fab338fa",
  1484 => x"f43974a3",
  1485 => x"26993881",
  1486 => x"19567580",
  1487 => x"f3b43480",
  1488 => x"0b80f3b8",
  1489 => x"34793356",
  1490 => x"75efe338",
  1491 => x"f0a43980",
  1492 => x"0b80f3b4",
  1493 => x"34800b80",
  1494 => x"f3b834e9",
  1495 => x"39800b80",
  1496 => x"f3b43480",
  1497 => x"0b80f3b8",
  1498 => x"34ffbd39",
  1499 => x"800b80f3",
  1500 => x"b434800b",
  1501 => x"80f3b834",
  1502 => x"ff903980",
  1503 => x"0b80f3b4",
  1504 => x"34800b80",
  1505 => x"f3b834fe",
  1506 => x"e339800b",
  1507 => x"80f3b434",
  1508 => x"800b80f3",
  1509 => x"b834feb6",
  1510 => x"3980e5d4",
  1511 => x"51dcb43f",
  1512 => x"fce23980",
  1513 => x"e5dc51dc",
  1514 => x"aa3ff7a9",
  1515 => x"3980e5e4",
  1516 => x"51dca03f",
  1517 => x"fca03980",
  1518 => x"e5e851dc",
  1519 => x"963ffc96",
  1520 => x"3980e5ec",
  1521 => x"51dc8c3f",
  1522 => x"fcba3980",
  1523 => x"e5f451dc",
  1524 => x"823ffc82",
  1525 => x"3980e5f8",
  1526 => x"51dbf83f",
  1527 => x"f6f73980",
  1528 => x"e5fc51db",
  1529 => x"ee3ffc9c",
  1530 => x"3980e684",
  1531 => x"51f68b39",
  1532 => x"80e5f851",
  1533 => x"f6843980",
  1534 => x"e68851f5",
  1535 => x"fd3980e6",
  1536 => x"8c51f5f6",
  1537 => x"3980e690",
  1538 => x"51dbc83f",
  1539 => x"80e4c451",
  1540 => x"dbc13f7c",
  1541 => x"5274932a",
  1542 => x"83068207",
  1543 => x"51da933f",
  1544 => x"7c51dbaf",
  1545 => x"3f80e4d8",
  1546 => x"51dba83f",
  1547 => x"7c527494",
  1548 => x"2a8f0651",
  1549 => x"d9fc3f7c",
  1550 => x"51db983f",
  1551 => x"80e4ec51",
  1552 => x"db913f7c",
  1553 => x"5274982a",
  1554 => x"81068105",
  1555 => x"51d9e33f",
  1556 => x"7c51daff",
  1557 => x"3f80e580",
  1558 => x"51daf83f",
  1559 => x"7c52749e",
  1560 => x"2a820751",
  1561 => x"d9cc3f7c",
  1562 => x"51dae83f",
  1563 => x"80e59451",
  1564 => x"dae13f74",
  1565 => x"9f2a923d",
  1566 => x"5a568b53",
  1567 => x"80de9c52",
  1568 => x"7851a9dd",
  1569 => x"3f820284",
  1570 => x"0580c105",
  1571 => x"5957f6eb",
  1572 => x"3980e6a0",
  1573 => x"51dabc3f",
  1574 => x"80e4c451",
  1575 => x"dab53f7c",
  1576 => x"5274932a",
  1577 => x"83068207",
  1578 => x"51d9873f",
  1579 => x"7c51daa3",
  1580 => x"3f80e4d8",
  1581 => x"51da9c3f",
  1582 => x"7c527494",
  1583 => x"2a8f0651",
  1584 => x"d8f03f7c",
  1585 => x"51da8c3f",
  1586 => x"80e4ec51",
  1587 => x"da853f7c",
  1588 => x"5274982a",
  1589 => x"81068105",
  1590 => x"51d8d73f",
  1591 => x"7c51d9f3",
  1592 => x"3f80e580",
  1593 => x"51d9ec3f",
  1594 => x"7c52749e",
  1595 => x"2a820751",
  1596 => x"d8c03f7c",
  1597 => x"51d9dc3f",
  1598 => x"80e59451",
  1599 => x"d9d53f74",
  1600 => x"9f2a923d",
  1601 => x"5a568b53",
  1602 => x"80de9c52",
  1603 => x"7851a8d1",
  1604 => x"3f820284",
  1605 => x"0580c105",
  1606 => x"5957f5df",
  1607 => x"3980e6ac",
  1608 => x"51d9b03f",
  1609 => x"80e4c451",
  1610 => x"d9a93f7c",
  1611 => x"5274932a",
  1612 => x"83068207",
  1613 => x"51d7fb3f",
  1614 => x"7c51d997",
  1615 => x"3f80e4d8",
  1616 => x"51d9903f",
  1617 => x"7c527494",
  1618 => x"2a8f0651",
  1619 => x"d7e43f7c",
  1620 => x"51d9803f",
  1621 => x"80e4ec51",
  1622 => x"d8f93f7c",
  1623 => x"5274982a",
  1624 => x"81068105",
  1625 => x"51d7cb3f",
  1626 => x"7c51d8e7",
  1627 => x"3f80e580",
  1628 => x"51d8e03f",
  1629 => x"7c52749e",
  1630 => x"2a820751",
  1631 => x"d7b43f7c",
  1632 => x"51d8d03f",
  1633 => x"80e59451",
  1634 => x"d8c93f74",
  1635 => x"9f2a923d",
  1636 => x"5a568b53",
  1637 => x"80de9c52",
  1638 => x"7851a7c5",
  1639 => x"3f820284",
  1640 => x"0580c105",
  1641 => x"5957f4d3",
  1642 => x"3980e6bc",
  1643 => x"51d8a43f",
  1644 => x"80e4c451",
  1645 => x"d89d3f7c",
  1646 => x"5274932a",
  1647 => x"83068207",
  1648 => x"51d6ef3f",
  1649 => x"7c51d88b",
  1650 => x"3f80e4d8",
  1651 => x"51d8843f",
  1652 => x"7c527494",
  1653 => x"2a8f0651",
  1654 => x"d6d83f7c",
  1655 => x"51d7f43f",
  1656 => x"80e4ec51",
  1657 => x"d7ed3f7c",
  1658 => x"5274982a",
  1659 => x"81068105",
  1660 => x"51d6bf3f",
  1661 => x"7c51d7db",
  1662 => x"3f80e580",
  1663 => x"51d7d43f",
  1664 => x"7c52749e",
  1665 => x"2a820751",
  1666 => x"d6a83f7c",
  1667 => x"51d7c43f",
  1668 => x"80e59451",
  1669 => x"d7bd3f74",
  1670 => x"9f2a923d",
  1671 => x"5a568b53",
  1672 => x"80de9c52",
  1673 => x"7851a6b9",
  1674 => x"3f820284",
  1675 => x"0580c105",
  1676 => x"5957f3c7",
  1677 => x"3980e6c8",
  1678 => x"51d7983f",
  1679 => x"80e4c451",
  1680 => x"d7913f7c",
  1681 => x"5274932a",
  1682 => x"83068207",
  1683 => x"51d5e33f",
  1684 => x"7c51d6ff",
  1685 => x"3f80e4d8",
  1686 => x"51d6f83f",
  1687 => x"7c527494",
  1688 => x"2a8f0651",
  1689 => x"d5cc3f7c",
  1690 => x"51d6e83f",
  1691 => x"80e4ec51",
  1692 => x"d6e13f7c",
  1693 => x"5274982a",
  1694 => x"81068105",
  1695 => x"51d5b33f",
  1696 => x"7c51d6cf",
  1697 => x"3f80e580",
  1698 => x"51d6c83f",
  1699 => x"7c52749e",
  1700 => x"2a820751",
  1701 => x"d59c3f7c",
  1702 => x"51d6b83f",
  1703 => x"80e59451",
  1704 => x"d6b13f74",
  1705 => x"9f2a923d",
  1706 => x"5a568b53",
  1707 => x"80de9c52",
  1708 => x"7851a5ad",
  1709 => x"3f820284",
  1710 => x"0580c105",
  1711 => x"5957f2bb",
  1712 => x"39e53d0d",
  1713 => x"80ebec08",
  1714 => x"84110870",
  1715 => x"9fff0651",
  1716 => x"55558a55",
  1717 => x"bb742783",
  1718 => x"388f5573",
  1719 => x"5287e851",
  1720 => x"a0b93f80",
  1721 => x"08fd0575",
  1722 => x"297083ff",
  1723 => x"ff0680e6",
  1724 => x"e4534058",
  1725 => x"d5dd3fd9",
  1726 => x"b23f8008",
  1727 => x"83ffff06",
  1728 => x"80e78052",
  1729 => x"57d5cc3f",
  1730 => x"983d7053",
  1731 => x"80ebf008",
  1732 => x"8c110853",
  1733 => x"575dd49a",
  1734 => x"3f7c51d5",
  1735 => x"b63f80e1",
  1736 => x"d451d5af",
  1737 => x"3f76963d",
  1738 => x"5a568b53",
  1739 => x"80de9c52",
  1740 => x"7851a4ad",
  1741 => x"3f880284",
  1742 => x"0580d105",
  1743 => x"5957758f",
  1744 => x"06547389",
  1745 => x"2688aa38",
  1746 => x"7618b015",
  1747 => x"55557375",
  1748 => x"3475842a",
  1749 => x"ff187081",
  1750 => x"ff06595b",
  1751 => x"5676df38",
  1752 => x"78793355",
  1753 => x"5773802e",
  1754 => x"a9387380",
  1755 => x"ec840856",
  1756 => x"56811757",
  1757 => x"758a2e88",
  1758 => x"94388415",
  1759 => x"0870822a",
  1760 => x"81064142",
  1761 => x"7f802ef2",
  1762 => x"3875750c",
  1763 => x"76335675",
  1764 => x"e0387879",
  1765 => x"33555a73",
  1766 => x"802e80cc",
  1767 => x"387380eb",
  1768 => x"fc085c56",
  1769 => x"811a80f3",
  1770 => x"b4337081",
  1771 => x"ff067010",
  1772 => x"101180f3",
  1773 => x"b8337081",
  1774 => x"ff067290",
  1775 => x"29117088",
  1776 => x"2b7d0762",
  1777 => x"0c4a5c5c",
  1778 => x"57575a5a",
  1779 => x"758a2e87",
  1780 => x"e1387680",
  1781 => x"cf2e87da",
  1782 => x"38811859",
  1783 => x"7880f3b8",
  1784 => x"34793356",
  1785 => x"75ffbd38",
  1786 => x"90b43f80",
  1787 => x"e78c519d",
  1788 => x"8a3f80eb",
  1789 => x"f0087f30",
  1790 => x"57558c15",
  1791 => x"08577577",
  1792 => x"25963880",
  1793 => x"0b84160c",
  1794 => x"74085877",
  1795 => x"ed387408",
  1796 => x"5877802e",
  1797 => x"f338e339",
  1798 => x"800b8816",
  1799 => x"0c740856",
  1800 => x"75802ef9",
  1801 => x"3880750c",
  1802 => x"8ff43f80",
  1803 => x"e794519c",
  1804 => x"ca3f8252",
  1805 => x"805197da",
  1806 => x"3f7c5280",
  1807 => x"ebf0088c",
  1808 => x"1108525a",
  1809 => x"d1ec3f7c",
  1810 => x"519cb03f",
  1811 => x"a05196b0",
  1812 => x"3f82518d",
  1813 => x"ea3f83ff",
  1814 => x"ff0b80eb",
  1815 => x"f0088c11",
  1816 => x"08435640",
  1817 => x"805ed4cd",
  1818 => x"7e4542ab",
  1819 => x"b30b8c16",
  1820 => x"085c437a",
  1821 => x"7f2583ca",
  1822 => x"38800b88",
  1823 => x"160c7408",
  1824 => x"5c7b802e",
  1825 => x"f938d6a3",
  1826 => x"3f800883",
  1827 => x"ffff0680",
  1828 => x"e1980b80",
  1829 => x"e1983356",
  1830 => x"5b5c7380",
  1831 => x"2e80cc38",
  1832 => x"80ebfc08",
  1833 => x"74575b81",
  1834 => x"1a80f3b4",
  1835 => x"337081ff",
  1836 => x"06701010",
  1837 => x"1180f3b8",
  1838 => x"337081ff",
  1839 => x"06729029",
  1840 => x"1170882b",
  1841 => x"7d07620c",
  1842 => x"535c5c57",
  1843 => x"575a5a75",
  1844 => x"8a2e86f1",
  1845 => x"387680cf",
  1846 => x"2e86ea38",
  1847 => x"81185978",
  1848 => x"80f3b834",
  1849 => x"79335675",
  1850 => x"ffbd387b",
  1851 => x"60278c38",
  1852 => x"7b80ebf0",
  1853 => x"088c1108",
  1854 => x"4358407b",
  1855 => x"30708025",
  1856 => x"55587d97",
  1857 => x"38817075",
  1858 => x"06575575",
  1859 => x"802e8c38",
  1860 => x"7480ebf0",
  1861 => x"088c1108",
  1862 => x"445b5e7b",
  1863 => x"30708025",
  1864 => x"555b7d80",
  1865 => x"2e973881",
  1866 => x"70750655",
  1867 => x"5573802e",
  1868 => x"8c387480",
  1869 => x"ebf0088c",
  1870 => x"11084556",
  1871 => x"4480e198",
  1872 => x"51d1903f",
  1873 => x"82528051",
  1874 => x"95c83f7c",
  1875 => x"5280ebf0",
  1876 => x"088c1108",
  1877 => x"5259cfda",
  1878 => x"3f7c519a",
  1879 => x"9e3fa051",
  1880 => x"949e3f7c",
  1881 => x"7d335557",
  1882 => x"73802ea9",
  1883 => x"3880ec84",
  1884 => x"08745755",
  1885 => x"81175775",
  1886 => x"8a2e84e1",
  1887 => x"38841508",
  1888 => x"70822a81",
  1889 => x"06555873",
  1890 => x"802ef238",
  1891 => x"75750c76",
  1892 => x"335675e0",
  1893 => x"3880e7a0",
  1894 => x"0b80e7a0",
  1895 => x"33555773",
  1896 => x"802ea938",
  1897 => x"80ec8408",
  1898 => x"74575581",
  1899 => x"1757758a",
  1900 => x"2e84cf38",
  1901 => x"84150870",
  1902 => x"822a8106",
  1903 => x"5a5a7880",
  1904 => x"2ef23875",
  1905 => x"750c7633",
  1906 => x"5675e038",
  1907 => x"7c527b51",
  1908 => x"cee03f7c",
  1909 => x"51cffc3f",
  1910 => x"80e7a40b",
  1911 => x"80e7a433",
  1912 => x"555a7380",
  1913 => x"2e80cc38",
  1914 => x"80ebfc08",
  1915 => x"74575b81",
  1916 => x"1a80f3b4",
  1917 => x"337081ff",
  1918 => x"06701010",
  1919 => x"1180f3b8",
  1920 => x"337081ff",
  1921 => x"06729029",
  1922 => x"1170882b",
  1923 => x"7d07620c",
  1924 => x"5a5c5c5f",
  1925 => x"575a5a75",
  1926 => x"8a2e848b",
  1927 => x"387680cf",
  1928 => x"2e848438",
  1929 => x"81185675",
  1930 => x"80f3b834",
  1931 => x"79335675",
  1932 => x"ffbd3880",
  1933 => x"ebf0088c",
  1934 => x"11085c55",
  1935 => x"7e7b24fc",
  1936 => x"b8388bda",
  1937 => x"3f80e7ac",
  1938 => x"5198b03f",
  1939 => x"63802e84",
  1940 => x"ae387d80",
  1941 => x"2e84a838",
  1942 => x"62623170",
  1943 => x"9f2a1170",
  1944 => x"812c6571",
  1945 => x"3180ebf0",
  1946 => x"088c1108",
  1947 => x"70733153",
  1948 => x"40535941",
  1949 => x"56578076",
  1950 => x"259938ff",
  1951 => x"1656800b",
  1952 => x"84160c74",
  1953 => x"085978ee",
  1954 => x"38740859",
  1955 => x"78802ef3",
  1956 => x"38e43980",
  1957 => x"e19851ce",
  1958 => x"ba3f7d80",
  1959 => x"2e85b338",
  1960 => x"80e7b851",
  1961 => x"cead3f80",
  1962 => x"e19851ce",
  1963 => x"a63f6380",
  1964 => x"2e83e238",
  1965 => x"80e7c451",
  1966 => x"ce993f80",
  1967 => x"e7d051ce",
  1968 => x"923f7c52",
  1969 => x"6151ccea",
  1970 => x"3f7c51ce",
  1971 => x"863f80e7",
  1972 => x"e051cdff",
  1973 => x"3f7c5262",
  1974 => x"51ccd73f",
  1975 => x"7c51cdf3",
  1976 => x"3f80e198",
  1977 => x"51cdec3f",
  1978 => x"80e7f051",
  1979 => x"cde53f7c",
  1980 => x"527651cc",
  1981 => x"bd3f7c51",
  1982 => x"cdd93f80",
  1983 => x"e88051cd",
  1984 => x"d23f7c52",
  1985 => x"769f2a17",
  1986 => x"70812c52",
  1987 => x"42cca33f",
  1988 => x"7c51cdbf",
  1989 => x"3f80e198",
  1990 => x"51cdb83f",
  1991 => x"80e89051",
  1992 => x"cdb13f7c",
  1993 => x"527f51cc",
  1994 => x"893f7c51",
  1995 => x"cda53f80",
  1996 => x"e8a051cd",
  1997 => x"9e3f7c52",
  1998 => x"6051cbf6",
  1999 => x"3f7c51cd",
  2000 => x"923f80e1",
  2001 => x"9851cd8b",
  2002 => x"3f80e8b0",
  2003 => x"51cd843f",
  2004 => x"7c5280eb",
  2005 => x"f0088c11",
  2006 => x"08525ecb",
  2007 => x"d53f7c51",
  2008 => x"ccf13f89",
  2009 => x"b93f80e8",
  2010 => x"c051968f",
  2011 => x"3f9d3d0d",
  2012 => x"047618b7",
  2013 => x"15555573",
  2014 => x"75347584",
  2015 => x"2aff1870",
  2016 => x"81ff0659",
  2017 => x"5b5676f7",
  2018 => x"b538f7d4",
  2019 => x"39841508",
  2020 => x"70822a81",
  2021 => x"065c5e7a",
  2022 => x"802ef238",
  2023 => x"8d750c84",
  2024 => x"15087082",
  2025 => x"2a810641",
  2026 => x"427f802e",
  2027 => x"f7cc38f7",
  2028 => x"d83974a3",
  2029 => x"26993881",
  2030 => x"19557480",
  2031 => x"f3b43480",
  2032 => x"0b80f3b8",
  2033 => x"34793356",
  2034 => x"75f7d938",
  2035 => x"f89a3980",
  2036 => x"0b80f3b4",
  2037 => x"34800b80",
  2038 => x"f3b834e9",
  2039 => x"39841508",
  2040 => x"70822a81",
  2041 => x"06595b77",
  2042 => x"802ef238",
  2043 => x"8d750c84",
  2044 => x"15087082",
  2045 => x"2a810655",
  2046 => x"5873802e",
  2047 => x"faff38fb",
  2048 => x"8b398415",
  2049 => x"0870822a",
  2050 => x"81065b54",
  2051 => x"79802ef2",
  2052 => x"388d750c",
  2053 => x"84150870",
  2054 => x"822a8106",
  2055 => x"5a5a7880",
  2056 => x"2efb9138",
  2057 => x"fb9d3974",
  2058 => x"a32680c4",
  2059 => x"38811957",
  2060 => x"7680f3b4",
  2061 => x"34800b80",
  2062 => x"f3b83479",
  2063 => x"335675fb",
  2064 => x"ae38fbef",
  2065 => x"3974a326",
  2066 => x"99388119",
  2067 => x"557480f3",
  2068 => x"b434800b",
  2069 => x"80f3b834",
  2070 => x"79335675",
  2071 => x"f8c938f9",
  2072 => x"8a39800b",
  2073 => x"80f3b434",
  2074 => x"800b80f3",
  2075 => x"b834e939",
  2076 => x"800b80f3",
  2077 => x"b434800b",
  2078 => x"80f3b834",
  2079 => x"ffbd3960",
  2080 => x"63633180",
  2081 => x"ebf0088c",
  2082 => x"11087074",
  2083 => x"31545e57",
  2084 => x"5856fbe2",
  2085 => x"3980e8d4",
  2086 => x"51cab83f",
  2087 => x"80e7d051",
  2088 => x"cab13f7c",
  2089 => x"526151c9",
  2090 => x"893f7c51",
  2091 => x"caa53f80",
  2092 => x"e7e051ca",
  2093 => x"9e3f7c52",
  2094 => x"6251c8f6",
  2095 => x"3f7c51ca",
  2096 => x"923f80e1",
  2097 => x"9851ca8b",
  2098 => x"3f80e7f0",
  2099 => x"51ca843f",
  2100 => x"7c527651",
  2101 => x"c8dc3f7c",
  2102 => x"51c9f83f",
  2103 => x"80e88051",
  2104 => x"c9f13f7c",
  2105 => x"52769f2a",
  2106 => x"1770812c",
  2107 => x"5242c8c2",
  2108 => x"3f7c51c9",
  2109 => x"de3f80e1",
  2110 => x"9851c9d7",
  2111 => x"3f80e890",
  2112 => x"51c9d03f",
  2113 => x"7c527f51",
  2114 => x"c8a83f7c",
  2115 => x"51c9c43f",
  2116 => x"80e8a051",
  2117 => x"c9bd3f7c",
  2118 => x"526051c8",
  2119 => x"953f7c51",
  2120 => x"c9b13f80",
  2121 => x"e19851c9",
  2122 => x"aa3f80e8",
  2123 => x"b051c9a3",
  2124 => x"3f7c5280",
  2125 => x"ebf0088c",
  2126 => x"1108525e",
  2127 => x"c7f43f7c",
  2128 => x"51c9903f",
  2129 => x"85d83f80",
  2130 => x"e8c05192",
  2131 => x"ae3f9d3d",
  2132 => x"0d0480e8",
  2133 => x"e451facc",
  2134 => x"39f83d0d",
  2135 => x"80ebf808",
  2136 => x"7008810a",
  2137 => x"0680f3b0",
  2138 => x"0c5385a1",
  2139 => x"3f86bd3f",
  2140 => x"80ebfc08",
  2141 => x"52800b84",
  2142 => x"130cfe80",
  2143 => x"0a0b8813",
  2144 => x"0c800b80",
  2145 => x"f3b43480",
  2146 => x"0b80f3b8",
  2147 => x"3480ec84",
  2148 => x"0853b60b",
  2149 => x"8c140c83",
  2150 => x"0b88140c",
  2151 => x"80ebf808",
  2152 => x"88110881",
  2153 => x"ff078812",
  2154 => x"0c5380eb",
  2155 => x"f40853ff",
  2156 => x"0b84140c",
  2157 => x"fc94800b",
  2158 => x"88140c82",
  2159 => x"d0affdfb",
  2160 => x"0b8c140c",
  2161 => x"80c0730c",
  2162 => x"72087086",
  2163 => x"2a810651",
  2164 => x"5271f538",
  2165 => x"90130870",
  2166 => x"832a8106",
  2167 => x"515473f4",
  2168 => x"3881fc80",
  2169 => x"810b9014",
  2170 => x"0c901308",
  2171 => x"70832a81",
  2172 => x"06515271",
  2173 => x"f43880fd",
  2174 => x"c0810b90",
  2175 => x"140c849e",
  2176 => x"3f80e1a0",
  2177 => x"5190f43f",
  2178 => x"890a5283",
  2179 => x"ffff5371",
  2180 => x"720c8412",
  2181 => x"ff145452",
  2182 => x"728025f3",
  2183 => x"3880e8f4",
  2184 => x"5190d83f",
  2185 => x"80e0e851",
  2186 => x"c7a93f80",
  2187 => x"0b80ebfc",
  2188 => x"08555372",
  2189 => x"882b740c",
  2190 => x"81135397",
  2191 => x"907326f3",
  2192 => x"38800b80",
  2193 => x"f3b43480",
  2194 => x"0b80f3b8",
  2195 => x"3480e980",
  2196 => x"51c7803f",
  2197 => x"80f3b008",
  2198 => x"802e81b9",
  2199 => x"3880e988",
  2200 => x"51c6f03f",
  2201 => x"80e99851",
  2202 => x"c6e93fd6",
  2203 => x"bd3f8551",
  2204 => x"81cd3ff0",
  2205 => x"cc3f8a51",
  2206 => x"81c53f80",
  2207 => x"0b80ebfc",
  2208 => x"08555372",
  2209 => x"882b740c",
  2210 => x"81135397",
  2211 => x"907326f3",
  2212 => x"38800b80",
  2213 => x"f3b43480",
  2214 => x"0b80f3b8",
  2215 => x"34ca8c3f",
  2216 => x"80ebf808",
  2217 => x"70087087",
  2218 => x"2a810651",
  2219 => x"55537380",
  2220 => x"2e8b3880",
  2221 => x"ebf00852",
  2222 => x"800b8413",
  2223 => x"0c720870",
  2224 => x"842a8106",
  2225 => x"51547380",
  2226 => x"2e8b3880",
  2227 => x"ebf00852",
  2228 => x"800b8813",
  2229 => x"0c720870",
  2230 => x"852a8106",
  2231 => x"54527280",
  2232 => x"2effba38",
  2233 => x"82b83f80",
  2234 => x"e1a0518f",
  2235 => x"8e3f890a",
  2236 => x"5283ffff",
  2237 => x"5371720c",
  2238 => x"8412ff14",
  2239 => x"54528073",
  2240 => x"24ff9a38",
  2241 => x"71720c84",
  2242 => x"12ff1454",
  2243 => x"52728025",
  2244 => x"e438ff89",
  2245 => x"3980e9bc",
  2246 => x"51fec639",
  2247 => x"fd3d0d80",
  2248 => x"ec800876",
  2249 => x"b0ea2994",
  2250 => x"120c5485",
  2251 => x"0b98150c",
  2252 => x"98140870",
  2253 => x"81065153",
  2254 => x"72f63885",
  2255 => x"3d0d04fb",
  2256 => x"3d0d7756",
  2257 => x"80557476",
  2258 => x"27819938",
  2259 => x"80ec8008",
  2260 => x"54bfa9bc",
  2261 => x"0b94150c",
  2262 => x"850b9815",
  2263 => x"0c981408",
  2264 => x"70810651",
  2265 => x"5372f638",
  2266 => x"bfa9bc0b",
  2267 => x"94150c85",
  2268 => x"0b98150c",
  2269 => x"98140870",
  2270 => x"81065153",
  2271 => x"72f638bf",
  2272 => x"a9bc0b94",
  2273 => x"150c850b",
  2274 => x"98150c98",
  2275 => x"14087081",
  2276 => x"06515372",
  2277 => x"f638bfa9",
  2278 => x"bc0b9415",
  2279 => x"0c850b98",
  2280 => x"150c9814",
  2281 => x"08708106",
  2282 => x"515372f6",
  2283 => x"38bfa9bc",
  2284 => x"0b94150c",
  2285 => x"850b9815",
  2286 => x"0c981408",
  2287 => x"70810651",
  2288 => x"5372f638",
  2289 => x"bfa9bc0b",
  2290 => x"94150c85",
  2291 => x"0b98150c",
  2292 => x"98140870",
  2293 => x"81065153",
  2294 => x"72f63881",
  2295 => x"15557575",
  2296 => x"26feee38",
  2297 => x"873d0d04",
  2298 => x"ff3d0d80",
  2299 => x"ec800874",
  2300 => x"10107510",
  2301 => x"0594120c",
  2302 => x"52850b98",
  2303 => x"130c9812",
  2304 => x"08708106",
  2305 => x"515170f6",
  2306 => x"38833d0d",
  2307 => x"04803d0d",
  2308 => x"80ec8008",
  2309 => x"51870b84",
  2310 => x"120c823d",
  2311 => x"0d04fd3d",
  2312 => x"0d810b80",
  2313 => x"ebf80884",
  2314 => x"110870fe",
  2315 => x"ffff0684",
  2316 => x"130c5484",
  2317 => x"110870e1",
  2318 => x"ff068413",
  2319 => x"0c548411",
  2320 => x"0884120c",
  2321 => x"84110870",
  2322 => x"80c08007",
  2323 => x"84130c54",
  2324 => x"54705254",
  2325 => x"ff923f80",
  2326 => x"ebf80884",
  2327 => x"110870ff",
  2328 => x"bfff0684",
  2329 => x"130c5384",
  2330 => x"110870e1",
  2331 => x"ff068413",
  2332 => x"0c538411",
  2333 => x"08708280",
  2334 => x"0784130c",
  2335 => x"53841108",
  2336 => x"7080c080",
  2337 => x"0784130c",
  2338 => x"53537351",
  2339 => x"feda3f80",
  2340 => x"ebf80884",
  2341 => x"1108ffbf",
  2342 => x"ff068412",
  2343 => x"0c53aa51",
  2344 => x"fec63f82",
  2345 => x"51fcf53f",
  2346 => x"853d0d04",
  2347 => x"fd3d0d80",
  2348 => x"ebf80888",
  2349 => x"110883de",
  2350 => x"80078812",
  2351 => x"0c841108",
  2352 => x"fca1ff06",
  2353 => x"84120c53",
  2354 => x"8f51fcd0",
  2355 => x"3f80ebf8",
  2356 => x"08841108",
  2357 => x"e1ff0684",
  2358 => x"120c8411",
  2359 => x"08868007",
  2360 => x"84120c84",
  2361 => x"110880c0",
  2362 => x"80078412",
  2363 => x"0c538151",
  2364 => x"fdf63f80",
  2365 => x"ebf80884",
  2366 => x"1108ffbf",
  2367 => x"ff068412",
  2368 => x"0c538551",
  2369 => x"fc963f80",
  2370 => x"ebf80884",
  2371 => x"110880c0",
  2372 => x"80078412",
  2373 => x"0c538151",
  2374 => x"fdce3f80",
  2375 => x"ebf80884",
  2376 => x"1108ffbf",
  2377 => x"ff068412",
  2378 => x"0c538151",
  2379 => x"fbee3f80",
  2380 => x"ebf80884",
  2381 => x"110880c0",
  2382 => x"80078412",
  2383 => x"0c538151",
  2384 => x"fda63f80",
  2385 => x"ebf80884",
  2386 => x"1108ffbf",
  2387 => x"ff068412",
  2388 => x"0c538151",
  2389 => x"fbc63f80",
  2390 => x"ebf80884",
  2391 => x"1108e1ff",
  2392 => x"0684120c",
  2393 => x"5384800b",
  2394 => x"84140870",
  2395 => x"72078416",
  2396 => x"0c538414",
  2397 => x"087080c0",
  2398 => x"80078416",
  2399 => x"0c535481",
  2400 => x"51fce53f",
  2401 => x"80ebf808",
  2402 => x"84110870",
  2403 => x"ffbfff06",
  2404 => x"84130c53",
  2405 => x"538551fb",
  2406 => x"833f80eb",
  2407 => x"f8088411",
  2408 => x"0870feff",
  2409 => x"ff068413",
  2410 => x"0c538411",
  2411 => x"0870e1ff",
  2412 => x"0684130c",
  2413 => x"53841108",
  2414 => x"70760784",
  2415 => x"130c5384",
  2416 => x"110880c0",
  2417 => x"80078412",
  2418 => x"0c538151",
  2419 => x"fc9a3f80",
  2420 => x"ebf80884",
  2421 => x"1108ffbf",
  2422 => x"ff068412",
  2423 => x"0c841108",
  2424 => x"e1ff0684",
  2425 => x"120c8411",
  2426 => x"08908007",
  2427 => x"84120c84",
  2428 => x"110880c0",
  2429 => x"80078412",
  2430 => x"0c548151",
  2431 => x"fbea3f80",
  2432 => x"ebf80884",
  2433 => x"1108ffbf",
  2434 => x"ff068412",
  2435 => x"0c54aa51",
  2436 => x"fbd63f80",
  2437 => x"ebf80884",
  2438 => x"1108feff",
  2439 => x"ff068412",
  2440 => x"0c841108",
  2441 => x"e1ff0684",
  2442 => x"120c8411",
  2443 => x"0884120c",
  2444 => x"84110880",
  2445 => x"c0800784",
  2446 => x"120c5481",
  2447 => x"51fba93f",
  2448 => x"80ebf808",
  2449 => x"841108ff",
  2450 => x"bfff0684",
  2451 => x"120c8411",
  2452 => x"08e1ff06",
  2453 => x"84120c84",
  2454 => x"11089880",
  2455 => x"0784120c",
  2456 => x"84110880",
  2457 => x"c0800784",
  2458 => x"120c5481",
  2459 => x"51faf93f",
  2460 => x"80ebf808",
  2461 => x"841108ff",
  2462 => x"bfff0684",
  2463 => x"120c54aa",
  2464 => x"51fae53f",
  2465 => x"80ebf808",
  2466 => x"841108fe",
  2467 => x"ffff0684",
  2468 => x"120c8411",
  2469 => x"08e1ff06",
  2470 => x"84120c84",
  2471 => x"11088412",
  2472 => x"0c841108",
  2473 => x"80c08007",
  2474 => x"84120c54",
  2475 => x"8151fab8",
  2476 => x"3f80ebf8",
  2477 => x"08841108",
  2478 => x"ffbfff06",
  2479 => x"84120c84",
  2480 => x"1108e1ff",
  2481 => x"0684120c",
  2482 => x"8411088c",
  2483 => x"80078412",
  2484 => x"0c841108",
  2485 => x"80c08007",
  2486 => x"84120c54",
  2487 => x"8151fa88",
  2488 => x"3f80ebf8",
  2489 => x"08841108",
  2490 => x"ffbfff06",
  2491 => x"84120c54",
  2492 => x"aa51f9f4",
  2493 => x"3f810b80",
  2494 => x"ebf80884",
  2495 => x"110870fe",
  2496 => x"ffff0684",
  2497 => x"130c5484",
  2498 => x"110870e1",
  2499 => x"ff068413",
  2500 => x"0c548411",
  2501 => x"0884120c",
  2502 => x"84110870",
  2503 => x"80c08007",
  2504 => x"84130c54",
  2505 => x"54705254",
  2506 => x"f9be3f80",
  2507 => x"ebf80884",
  2508 => x"110870ff",
  2509 => x"bfff0684",
  2510 => x"130c5384",
  2511 => x"110870e1",
  2512 => x"ff068413",
  2513 => x"0c538411",
  2514 => x"08708280",
  2515 => x"0784130c",
  2516 => x"53841108",
  2517 => x"7080c080",
  2518 => x"0784130c",
  2519 => x"53537351",
  2520 => x"f9863f80",
  2521 => x"ebf80884",
  2522 => x"1108ffbf",
  2523 => x"ff068412",
  2524 => x"0c53aa51",
  2525 => x"f8f23f82",
  2526 => x"51f7a13f",
  2527 => x"853d0d04",
  2528 => x"fb3d0d02",
  2529 => x"9f053380",
  2530 => x"ebf80884",
  2531 => x"11088180",
  2532 => x"80078412",
  2533 => x"0c545581",
  2534 => x"f00b8414",
  2535 => x"08e1ff06",
  2536 => x"84150c70",
  2537 => x"7606842b",
  2538 => x"84150870",
  2539 => x"72078417",
  2540 => x"0c548415",
  2541 => x"0880c080",
  2542 => x"0784160c",
  2543 => x"55568151",
  2544 => x"f8a63f80",
  2545 => x"ebf80884",
  2546 => x"1108ffbf",
  2547 => x"ff068412",
  2548 => x"0c841108",
  2549 => x"e1ff0684",
  2550 => x"120c7588",
  2551 => x"2b77842b",
  2552 => x"06841208",
  2553 => x"71078413",
  2554 => x"0c841208",
  2555 => x"80c08007",
  2556 => x"84130c56",
  2557 => x"538151f7",
  2558 => x"ef3f80eb",
  2559 => x"f8088411",
  2560 => x"08ffbfff",
  2561 => x"0684120c",
  2562 => x"53ae51f7",
  2563 => x"db3f873d",
  2564 => x"0d04fc3d",
  2565 => x"0d029b05",
  2566 => x"33028405",
  2567 => x"9f053354",
  2568 => x"5272822e",
  2569 => x"81ad3882",
  2570 => x"73259138",
  2571 => x"72832e83",
  2572 => x"bc387284",
  2573 => x"2e82a938",
  2574 => x"863d0d04",
  2575 => x"72812e09",
  2576 => x"8106f538",
  2577 => x"ff801270",
  2578 => x"81ff0680",
  2579 => x"ebf80884",
  2580 => x"1108feff",
  2581 => x"ff068412",
  2582 => x"0c841108",
  2583 => x"e1ff0684",
  2584 => x"120c7184",
  2585 => x"2b9e8006",
  2586 => x"84120870",
  2587 => x"72078414",
  2588 => x"0c548412",
  2589 => x"0880c080",
  2590 => x"0784130c",
  2591 => x"57555652",
  2592 => x"8151f6e4",
  2593 => x"3f80ebf8",
  2594 => x"08841108",
  2595 => x"ffbfff06",
  2596 => x"84120c84",
  2597 => x"1108e1ff",
  2598 => x"0684120c",
  2599 => x"75882b9e",
  2600 => x"80068412",
  2601 => x"08710784",
  2602 => x"130c8412",
  2603 => x"0880c080",
  2604 => x"0784130c",
  2605 => x"55538151",
  2606 => x"f6ae3f80",
  2607 => x"ebf80884",
  2608 => x"1108ffbf",
  2609 => x"ff068412",
  2610 => x"0c53aa51",
  2611 => x"f69a3f86",
  2612 => x"3d0d04c0",
  2613 => x"127081ff",
  2614 => x"0680ebf8",
  2615 => x"08841108",
  2616 => x"feffff06",
  2617 => x"84120c84",
  2618 => x"1108e1ff",
  2619 => x"0684120c",
  2620 => x"71842b9e",
  2621 => x"80068412",
  2622 => x"08707207",
  2623 => x"84140c54",
  2624 => x"84120880",
  2625 => x"c0800784",
  2626 => x"130c5755",
  2627 => x"56528151",
  2628 => x"f5d63f80",
  2629 => x"ebf80884",
  2630 => x"1108ffbf",
  2631 => x"ff068412",
  2632 => x"0c841108",
  2633 => x"e1ff0684",
  2634 => x"120c7588",
  2635 => x"2b9e8006",
  2636 => x"84120871",
  2637 => x"0784130c",
  2638 => x"84120880",
  2639 => x"c0800784",
  2640 => x"130c5553",
  2641 => x"8151f5a0",
  2642 => x"3f80ebf8",
  2643 => x"08841108",
  2644 => x"ffbfff06",
  2645 => x"84120c53",
  2646 => x"aa51f58c",
  2647 => x"3ffef039",
  2648 => x"d0127081",
  2649 => x"ff0680eb",
  2650 => x"f8088411",
  2651 => x"08feffff",
  2652 => x"0684120c",
  2653 => x"841108e1",
  2654 => x"ff068412",
  2655 => x"0c71842b",
  2656 => x"9e800684",
  2657 => x"12087072",
  2658 => x"0784140c",
  2659 => x"54841208",
  2660 => x"80c08007",
  2661 => x"84130c57",
  2662 => x"55565281",
  2663 => x"51f4c93f",
  2664 => x"80ebf808",
  2665 => x"841108ff",
  2666 => x"bfff0684",
  2667 => x"120c8411",
  2668 => x"08e1ff06",
  2669 => x"84120c75",
  2670 => x"882b9e80",
  2671 => x"06841208",
  2672 => x"71078413",
  2673 => x"0c841208",
  2674 => x"80c08007",
  2675 => x"84130c55",
  2676 => x"538151f4",
  2677 => x"933f80eb",
  2678 => x"f8088411",
  2679 => x"08ffbfff",
  2680 => x"0684120c",
  2681 => x"53aa51f3",
  2682 => x"ff3ffde3",
  2683 => x"39ff9012",
  2684 => x"7081ff06",
  2685 => x"80ebf808",
  2686 => x"841108fe",
  2687 => x"ffff0684",
  2688 => x"120c8411",
  2689 => x"08e1ff06",
  2690 => x"84120c71",
  2691 => x"842b9e80",
  2692 => x"06841208",
  2693 => x"70720784",
  2694 => x"140c5484",
  2695 => x"120880c0",
  2696 => x"80078413",
  2697 => x"0c575556",
  2698 => x"528151f3",
  2699 => x"bb3f80eb",
  2700 => x"f8088411",
  2701 => x"08ffbfff",
  2702 => x"0684120c",
  2703 => x"841108e1",
  2704 => x"ff068412",
  2705 => x"0c75882b",
  2706 => x"9e800684",
  2707 => x"12087107",
  2708 => x"84130c84",
  2709 => x"120880c0",
  2710 => x"80078413",
  2711 => x"0c555381",
  2712 => x"51f3853f",
  2713 => x"80ebf808",
  2714 => x"841108ff",
  2715 => x"bfff0684",
  2716 => x"120c53aa",
  2717 => x"51f2f13f",
  2718 => x"fcd539fb",
  2719 => x"3d0d7770",
  2720 => x"33535671",
  2721 => x"802e818f",
  2722 => x"38715581",
  2723 => x"1680ebf8",
  2724 => x"08841108",
  2725 => x"81808007",
  2726 => x"84120c84",
  2727 => x"1108e1ff",
  2728 => x"0684120c",
  2729 => x"76842b9e",
  2730 => x"80068412",
  2731 => x"08707207",
  2732 => x"84140c55",
  2733 => x"84120880",
  2734 => x"c0800784",
  2735 => x"130c5654",
  2736 => x"568151f2",
  2737 => x"a33f80eb",
  2738 => x"f8088411",
  2739 => x"08ffbfff",
  2740 => x"0684120c",
  2741 => x"841108e1",
  2742 => x"ff068412",
  2743 => x"0c75882b",
  2744 => x"9e800684",
  2745 => x"12087107",
  2746 => x"84130c84",
  2747 => x"120880c0",
  2748 => x"80078413",
  2749 => x"0c555381",
  2750 => x"51f1ed3f",
  2751 => x"80ebf808",
  2752 => x"841108ff",
  2753 => x"bfff0684",
  2754 => x"120c53ae",
  2755 => x"51f1d93f",
  2756 => x"75335574",
  2757 => x"fef53887",
  2758 => x"3d0d048c",
  2759 => x"08028c0c",
  2760 => x"fd3d0d80",
  2761 => x"538c088c",
  2762 => x"0508528c",
  2763 => x"08880508",
  2764 => x"5182de3f",
  2765 => x"80087080",
  2766 => x"0c54853d",
  2767 => x"0d8c0c04",
  2768 => x"8c08028c",
  2769 => x"0cfd3d0d",
  2770 => x"81538c08",
  2771 => x"8c050852",
  2772 => x"8c088805",
  2773 => x"085182b9",
  2774 => x"3f800870",
  2775 => x"800c5485",
  2776 => x"3d0d8c0c",
  2777 => x"048c0802",
  2778 => x"8c0cf93d",
  2779 => x"0d800b8c",
  2780 => x"08fc050c",
  2781 => x"8c088805",
  2782 => x"088025ab",
  2783 => x"388c0888",
  2784 => x"0508308c",
  2785 => x"0888050c",
  2786 => x"800b8c08",
  2787 => x"f4050c8c",
  2788 => x"08fc0508",
  2789 => x"8838810b",
  2790 => x"8c08f405",
  2791 => x"0c8c08f4",
  2792 => x"05088c08",
  2793 => x"fc050c8c",
  2794 => x"088c0508",
  2795 => x"8025ab38",
  2796 => x"8c088c05",
  2797 => x"08308c08",
  2798 => x"8c050c80",
  2799 => x"0b8c08f0",
  2800 => x"050c8c08",
  2801 => x"fc050888",
  2802 => x"38810b8c",
  2803 => x"08f0050c",
  2804 => x"8c08f005",
  2805 => x"088c08fc",
  2806 => x"050c8053",
  2807 => x"8c088c05",
  2808 => x"08528c08",
  2809 => x"88050851",
  2810 => x"81a73f80",
  2811 => x"08708c08",
  2812 => x"f8050c54",
  2813 => x"8c08fc05",
  2814 => x"08802e8c",
  2815 => x"388c08f8",
  2816 => x"0508308c",
  2817 => x"08f8050c",
  2818 => x"8c08f805",
  2819 => x"0870800c",
  2820 => x"54893d0d",
  2821 => x"8c0c048c",
  2822 => x"08028c0c",
  2823 => x"fb3d0d80",
  2824 => x"0b8c08fc",
  2825 => x"050c8c08",
  2826 => x"88050880",
  2827 => x"2593388c",
  2828 => x"08880508",
  2829 => x"308c0888",
  2830 => x"050c810b",
  2831 => x"8c08fc05",
  2832 => x"0c8c088c",
  2833 => x"05088025",
  2834 => x"8c388c08",
  2835 => x"8c050830",
  2836 => x"8c088c05",
  2837 => x"0c81538c",
  2838 => x"088c0508",
  2839 => x"528c0888",
  2840 => x"050851ad",
  2841 => x"3f800870",
  2842 => x"8c08f805",
  2843 => x"0c548c08",
  2844 => x"fc050880",
  2845 => x"2e8c388c",
  2846 => x"08f80508",
  2847 => x"308c08f8",
  2848 => x"050c8c08",
  2849 => x"f8050870",
  2850 => x"800c5487",
  2851 => x"3d0d8c0c",
  2852 => x"048c0802",
  2853 => x"8c0cfd3d",
  2854 => x"0d810b8c",
  2855 => x"08fc050c",
  2856 => x"800b8c08",
  2857 => x"f8050c8c",
  2858 => x"088c0508",
  2859 => x"8c088805",
  2860 => x"0827ac38",
  2861 => x"8c08fc05",
  2862 => x"08802ea3",
  2863 => x"38800b8c",
  2864 => x"088c0508",
  2865 => x"2499388c",
  2866 => x"088c0508",
  2867 => x"108c088c",
  2868 => x"050c8c08",
  2869 => x"fc050810",
  2870 => x"8c08fc05",
  2871 => x"0cc9398c",
  2872 => x"08fc0508",
  2873 => x"802e80c9",
  2874 => x"388c088c",
  2875 => x"05088c08",
  2876 => x"88050826",
  2877 => x"a1388c08",
  2878 => x"8805088c",
  2879 => x"088c0508",
  2880 => x"318c0888",
  2881 => x"050c8c08",
  2882 => x"f805088c",
  2883 => x"08fc0508",
  2884 => x"078c08f8",
  2885 => x"050c8c08",
  2886 => x"fc050881",
  2887 => x"2a8c08fc",
  2888 => x"050c8c08",
  2889 => x"8c050881",
  2890 => x"2a8c088c",
  2891 => x"050cffaf",
  2892 => x"398c0890",
  2893 => x"0508802e",
  2894 => x"8f388c08",
  2895 => x"88050870",
  2896 => x"8c08f405",
  2897 => x"0c518d39",
  2898 => x"8c08f805",
  2899 => x"08708c08",
  2900 => x"f4050c51",
  2901 => x"8c08f405",
  2902 => x"08800c85",
  2903 => x"3d0d8c0c",
  2904 => x"04fc3d0d",
  2905 => x"7670797b",
  2906 => x"55555555",
  2907 => x"8f72278c",
  2908 => x"38727507",
  2909 => x"83065170",
  2910 => x"802ea738",
  2911 => x"ff125271",
  2912 => x"ff2e9838",
  2913 => x"72708105",
  2914 => x"54337470",
  2915 => x"81055634",
  2916 => x"ff125271",
  2917 => x"ff2e0981",
  2918 => x"06ea3874",
  2919 => x"800c863d",
  2920 => x"0d047451",
  2921 => x"72708405",
  2922 => x"54087170",
  2923 => x"8405530c",
  2924 => x"72708405",
  2925 => x"54087170",
  2926 => x"8405530c",
  2927 => x"72708405",
  2928 => x"54087170",
  2929 => x"8405530c",
  2930 => x"72708405",
  2931 => x"54087170",
  2932 => x"8405530c",
  2933 => x"f0125271",
  2934 => x"8f26c938",
  2935 => x"83722795",
  2936 => x"38727084",
  2937 => x"05540871",
  2938 => x"70840553",
  2939 => x"0cfc1252",
  2940 => x"718326ed",
  2941 => x"387054ff",
  2942 => x"8339fd3d",
  2943 => x"0d800b80",
  2944 => x"ebe00854",
  2945 => x"5472812e",
  2946 => x"9c387380",
  2947 => x"f3bc0cff",
  2948 => x"acce3fff",
  2949 => x"abea3f80",
  2950 => x"ec885281",
  2951 => x"51e6ba3f",
  2952 => x"800851a2",
  2953 => x"3f7280f3",
  2954 => x"bc0cffac",
  2955 => x"b33fffab",
  2956 => x"cf3f80ec",
  2957 => x"88528151",
  2958 => x"e69f3f80",
  2959 => x"0851873f",
  2960 => x"00ff3900",
  2961 => x"ff39f73d",
  2962 => x"0d7b80ec",
  2963 => x"8c0882c8",
  2964 => x"11085a54",
  2965 => x"5a77802e",
  2966 => x"80da3881",
  2967 => x"88188419",
  2968 => x"08ff0581",
  2969 => x"712b5955",
  2970 => x"59807424",
  2971 => x"80ea3880",
  2972 => x"7424b538",
  2973 => x"73822b78",
  2974 => x"11880556",
  2975 => x"56818019",
  2976 => x"08770653",
  2977 => x"72802eb6",
  2978 => x"38781670",
  2979 => x"08535379",
  2980 => x"51740853",
  2981 => x"722dff14",
  2982 => x"fc17fc17",
  2983 => x"79812c5a",
  2984 => x"57575473",
  2985 => x"8025d638",
  2986 => x"77085877",
  2987 => x"ffad3880",
  2988 => x"ec8c0853",
  2989 => x"bc1308a5",
  2990 => x"387951ff",
  2991 => x"833f7408",
  2992 => x"53722dff",
  2993 => x"14fc17fc",
  2994 => x"1779812c",
  2995 => x"5a575754",
  2996 => x"738025ff",
  2997 => x"a838d139",
  2998 => x"8057ff93",
  2999 => x"397251bc",
  3000 => x"13085372",
  3001 => x"2d7951fe",
  3002 => x"d73fff3d",
  3003 => x"0d80f390",
  3004 => x"0bfc0570",
  3005 => x"08525270",
  3006 => x"ff2e9138",
  3007 => x"702dfc12",
  3008 => x"70085252",
  3009 => x"70ff2e09",
  3010 => x"8106f138",
  3011 => x"833d0d04",
  3012 => x"04ffabb9",
  3013 => x"3f040000",
  3014 => x"00000040",
  3015 => x"30782020",
  3016 => x"20202020",
  3017 => x"20200000",
  3018 => x"0a677265",
  3019 => x"74682072",
  3020 => x"65676973",
  3021 => x"74657273",
  3022 => x"3a000000",
  3023 => x"0a636f6e",
  3024 => x"74726f6c",
  3025 => x"3a202020",
  3026 => x"20202000",
  3027 => x"0a737461",
  3028 => x"7475733a",
  3029 => x"20202020",
  3030 => x"20202000",
  3031 => x"0a6d6163",
  3032 => x"5f6d7362",
  3033 => x"3a202020",
  3034 => x"20202000",
  3035 => x"0a6d6163",
  3036 => x"5f6c7362",
  3037 => x"3a202020",
  3038 => x"20202000",
  3039 => x"0a6d6469",
  3040 => x"6f5f636f",
  3041 => x"6e74726f",
  3042 => x"6c3a2000",
  3043 => x"0a74785f",
  3044 => x"706f696e",
  3045 => x"7465723a",
  3046 => x"20202000",
  3047 => x"0a72785f",
  3048 => x"706f696e",
  3049 => x"7465723a",
  3050 => x"20202000",
  3051 => x"0a656463",
  3052 => x"6c5f6970",
  3053 => x"3a202020",
  3054 => x"20202000",
  3055 => x"0a686173",
  3056 => x"685f6d73",
  3057 => x"623a2020",
  3058 => x"20202000",
  3059 => x"0a686173",
  3060 => x"685f6c73",
  3061 => x"623a2020",
  3062 => x"20202000",
  3063 => x"0a6d6469",
  3064 => x"6f207068",
  3065 => x"79207265",
  3066 => x"67697374",
  3067 => x"65727300",
  3068 => x"0a206d64",
  3069 => x"696f2070",
  3070 => x"68793a20",
  3071 => x"00000000",
  3072 => x"0a202072",
  3073 => x"65673a20",
  3074 => x"00000000",
  3075 => x"2d3e2000",
  3076 => x"0a677265",
  3077 => x"74682d3e",
  3078 => x"636f6e74",
  3079 => x"726f6c20",
  3080 => x"3a000000",
  3081 => x"0a677265",
  3082 => x"74682d3e",
  3083 => x"73746174",
  3084 => x"75732020",
  3085 => x"3a000000",
  3086 => x"0a646573",
  3087 => x"63722d3e",
  3088 => x"636f6e74",
  3089 => x"726f6c20",
  3090 => x"3a000000",
  3091 => x"77726974",
  3092 => x"65206164",
  3093 => x"64726573",
  3094 => x"733a2000",
  3095 => x"20206c65",
  3096 => x"6e677468",
  3097 => x"3a200000",
  3098 => x"0a0a0000",
  3099 => x"72656164",
  3100 => x"20206164",
  3101 => x"64726573",
  3102 => x"733a2000",
  3103 => x"20206578",
  3104 => x"70656374",
  3105 => x"3a200000",
  3106 => x"2020676f",
  3107 => x"743a2000",
  3108 => x"20657272",
  3109 => x"6f720000",
  3110 => x"0a000000",
  3111 => x"206f6b00",
  3112 => x"6d656d6f",
  3113 => x"72792074",
  3114 => x"65737420",
  3115 => x"696e6974",
  3116 => x"00000000",
  3117 => x"70686173",
  3118 => x"65207368",
  3119 => x"6966743a",
  3120 => x"20000000",
  3121 => x"20207374",
  3122 => x"61747573",
  3123 => x"3a200000",
  3124 => x"20202020",
  3125 => x"20000000",
  3126 => x"44445220",
  3127 => x"6d656d6f",
  3128 => x"72792069",
  3129 => x"6e666f00",
  3130 => x"0a617574",
  3131 => x"6f20745f",
  3132 => x"52455245",
  3133 => x"5348203a",
  3134 => x"00000000",
  3135 => x"0a636c6f",
  3136 => x"636b2065",
  3137 => x"6e61626c",
  3138 => x"6520203a",
  3139 => x"00000000",
  3140 => x"0a696e69",
  3141 => x"74616c69",
  3142 => x"7a652020",
  3143 => x"2020203a",
  3144 => x"00000000",
  3145 => x"0a636f6c",
  3146 => x"756d6e20",
  3147 => x"73697a65",
  3148 => x"2020203a",
  3149 => x"00000000",
  3150 => x"0a62616e",
  3151 => x"6b73697a",
  3152 => x"65202020",
  3153 => x"2020203a",
  3154 => x"00000000",
  3155 => x"4d627974",
  3156 => x"65000000",
  3157 => x"0a745f52",
  3158 => x"43442020",
  3159 => x"20202020",
  3160 => x"2020203a",
  3161 => x"00000000",
  3162 => x"0a745f52",
  3163 => x"46432020",
  3164 => x"20202020",
  3165 => x"2020203a",
  3166 => x"00000000",
  3167 => x"0a745f52",
  3168 => x"50202020",
  3169 => x"20202020",
  3170 => x"2020203a",
  3171 => x"00000000",
  3172 => x"0a726566",
  3173 => x"72657368",
  3174 => x"20656e2e",
  3175 => x"2020203a",
  3176 => x"00000000",
  3177 => x"0a444452",
  3178 => x"20667265",
  3179 => x"7175656e",
  3180 => x"6379203a",
  3181 => x"00000000",
  3182 => x"0a444452",
  3183 => x"20646174",
  3184 => x"61207769",
  3185 => x"6474683a",
  3186 => x"00000000",
  3187 => x"0a6d6f62",
  3188 => x"696c6520",
  3189 => x"73757070",
  3190 => x"6f72743a",
  3191 => x"00000000",
  3192 => x"0a73656c",
  3193 => x"66207265",
  3194 => x"66726573",
  3195 => x"6820203a",
  3196 => x"00000000",
  3197 => x"756e6b6e",
  3198 => x"6f776e00",
  3199 => x"20617272",
  3200 => x"61790000",
  3201 => x"0a74656d",
  3202 => x"702d636f",
  3203 => x"6d702072",
  3204 => x"6566723a",
  3205 => x"00000000",
  3206 => x"c2b04300",
  3207 => x"0a647269",
  3208 => x"76652073",
  3209 => x"7472656e",
  3210 => x"6774683a",
  3211 => x"00000000",
  3212 => x"0a706f77",
  3213 => x"65722073",
  3214 => x"6176696e",
  3215 => x"6720203a",
  3216 => x"00000000",
  3217 => x"0a745f58",
  3218 => x"50202020",
  3219 => x"20202020",
  3220 => x"2020203a",
  3221 => x"00000000",
  3222 => x"0a745f58",
  3223 => x"53522020",
  3224 => x"20202020",
  3225 => x"2020203a",
  3226 => x"00000000",
  3227 => x"0a745f43",
  3228 => x"4b452020",
  3229 => x"20202020",
  3230 => x"2020203a",
  3231 => x"00000000",
  3232 => x"0a434153",
  3233 => x"206c6174",
  3234 => x"656e6379",
  3235 => x"2020203a",
  3236 => x"00000000",
  3237 => x"0a6d6f62",
  3238 => x"696c6520",
  3239 => x"656e6162",
  3240 => x"6c65643a",
  3241 => x"00000000",
  3242 => x"0a737461",
  3243 => x"74757320",
  3244 => x"72656164",
  3245 => x"2020203a",
  3246 => x"00000000",
  3247 => x"332f3400",
  3248 => x"38350000",
  3249 => x"68616c66",
  3250 => x"00000000",
  3251 => x"34303639",
  3252 => x"00000000",
  3253 => x"20353132",
  3254 => x"00000000",
  3255 => x"66756c6c",
  3256 => x"00000000",
  3257 => x"37300000",
  3258 => x"34350000",
  3259 => x"31303234",
  3260 => x"00000000",
  3261 => x"31350000",
  3262 => x"312f3400",
  3263 => x"32303438",
  3264 => x"00000000",
  3265 => x"312f3800",
  3266 => x"312f3200",
  3267 => x"312f3100",
  3268 => x"64656570",
  3269 => x"20706f77",
  3270 => x"65722064",
  3271 => x"6f776e00",
  3272 => x"636c6f63",
  3273 => x"6b207374",
  3274 => x"6f700000",
  3275 => x"73656c66",
  3276 => x"20726566",
  3277 => x"72657368",
  3278 => x"00000000",
  3279 => x"706f7765",
  3280 => x"7220646f",
  3281 => x"776e0000",
  3282 => x"6e6f6e65",
  3283 => x"00000000",
  3284 => x"61646472",
  3285 => x"6573733a",
  3286 => x"20000000",
  3287 => x"20646174",
  3288 => x"613a2000",
  3289 => x"0a0a4443",
  3290 => x"4d207068",
  3291 => x"61736520",
  3292 => x"73686966",
  3293 => x"74207465",
  3294 => x"7374696e",
  3295 => x"67000000",
  3296 => x"0a696e69",
  3297 => x"7469616c",
  3298 => x"3a200000",
  3299 => x"676f2064",
  3300 => x"6f776e00",
  3301 => x"7363616e",
  3302 => x"2072616e",
  3303 => x"67650000",
  3304 => x"09000000",
  3305 => x"20202020",
  3306 => x"00000000",
  3307 => x"676f2074",
  3308 => x"6f206579",
  3309 => x"65000000",
  3310 => x"6c6f7720",
  3311 => x"666f756e",
  3312 => x"64000000",
  3313 => x"68696768",
  3314 => x"20666f75",
  3315 => x"6e640000",
  3316 => x"0a6c6f77",
  3317 => x"3a202020",
  3318 => x"20202020",
  3319 => x"20200000",
  3320 => x"0a686967",
  3321 => x"683a2020",
  3322 => x"20202020",
  3323 => x"20200000",
  3324 => x"0a646966",
  3325 => x"663a2020",
  3326 => x"20202020",
  3327 => x"20200000",
  3328 => x"0a646966",
  3329 => x"662f323a",
  3330 => x"20202020",
  3331 => x"20200000",
  3332 => x"0a6d696e",
  3333 => x"5f657272",
  3334 => x"3a202020",
  3335 => x"20200000",
  3336 => x"0a6d696e",
  3337 => x"5f657272",
  3338 => x"5f706f73",
  3339 => x"3a200000",
  3340 => x"0a66696e",
  3341 => x"616c3a20",
  3342 => x"20202020",
  3343 => x"20200000",
  3344 => x"64636d5f",
  3345 => x"74657374",
  3346 => x"5f707320",
  3347 => x"646f6e65",
  3348 => x"00000000",
  3349 => x"68696768",
  3350 => x"204e4f54",
  3351 => x"20666f75",
  3352 => x"6e640000",
  3353 => x"6c6f7720",
  3354 => x"4e4f5420",
  3355 => x"666f756e",
  3356 => x"64000000",
  3357 => x"696e6974",
  3358 => x"20646f6e",
  3359 => x"652e0000",
  3360 => x"74657374",
  3361 => x"2e632000",
  3362 => x"286f6e20",
  3363 => x"73696d75",
  3364 => x"6c61746f",
  3365 => x"72290a00",
  3366 => x"636f6d70",
  3367 => x"696c6564",
  3368 => x"3a205365",
  3369 => x"70203330",
  3370 => x"20323031",
  3371 => x"30202031",
  3372 => x"363a3334",
  3373 => x"3a30330a",
  3374 => x"00000000",
  3375 => x"286f6e20",
  3376 => x"68617264",
  3377 => x"77617265",
  3378 => x"290a0000",
  3379 => x"000006d1",
  3380 => x"000006f7",
  3381 => x"000006f7",
  3382 => x"000006d1",
  3383 => x"000006f7",
  3384 => x"000006f7",
  3385 => x"000006f7",
  3386 => x"000006f7",
  3387 => x"000006f7",
  3388 => x"000006f7",
  3389 => x"000006f7",
  3390 => x"000006f7",
  3391 => x"000006f7",
  3392 => x"000006f7",
  3393 => x"000006f7",
  3394 => x"000006f7",
  3395 => x"000006f7",
  3396 => x"000006f7",
  3397 => x"000006f7",
  3398 => x"000006f7",
  3399 => x"000006f7",
  3400 => x"000006f7",
  3401 => x"000006f7",
  3402 => x"000006f7",
  3403 => x"000006f7",
  3404 => x"000006f7",
  3405 => x"000006f7",
  3406 => x"000006f7",
  3407 => x"000006f7",
  3408 => x"000006f7",
  3409 => x"000006f7",
  3410 => x"000006f7",
  3411 => x"000006f7",
  3412 => x"000006f7",
  3413 => x"000006f7",
  3414 => x"000006f7",
  3415 => x"000006f7",
  3416 => x"000006f7",
  3417 => x"000007a3",
  3418 => x"0000079b",
  3419 => x"00000793",
  3420 => x"0000078b",
  3421 => x"00000783",
  3422 => x"0000077b",
  3423 => x"00000773",
  3424 => x"0000076a",
  3425 => x"00000761",
  3426 => x"000017fe",
  3427 => x"000017f7",
  3428 => x"000017f0",
  3429 => x"000012f6",
  3430 => x"000012f6",
  3431 => x"000017e9",
  3432 => x"000017e9",
  3433 => x"00001a35",
  3434 => x"000019a9",
  3435 => x"0000191d",
  3436 => x"00001372",
  3437 => x"00001891",
  3438 => x"00001805",
  3439 => x"64756d6d",
  3440 => x"792e6578",
  3441 => x"65000000",
  3442 => x"43000000",
  3443 => x"00ffffff",
  3444 => x"ff00ffff",
  3445 => x"ffff00ff",
  3446 => x"ffffff00",
  3447 => x"00000000",
  3448 => x"00000000",
  3449 => x"00000000",
  3450 => x"00003998",
  3451 => x"fff00000",
  3452 => x"80000e00",
  3453 => x"80000c00",
  3454 => x"80000800",
  3455 => x"80000600",
  3456 => x"80000200",
  3457 => x"80000100",
  3458 => x"000035bc",
  3459 => x"00003610",
  3460 => x"00000000",
  3461 => x"00003878",
  3462 => x"000038d4",
  3463 => x"00003930",
  3464 => x"00000000",
  3465 => x"00000000",
  3466 => x"00000000",
  3467 => x"00000000",
  3468 => x"00000000",
  3469 => x"00000000",
  3470 => x"00000000",
  3471 => x"00000000",
  3472 => x"00000000",
  3473 => x"000035c8",
  3474 => x"00000000",
  3475 => x"00000000",
  3476 => x"00000000",
  3477 => x"00000000",
  3478 => x"00000000",
  3479 => x"00000000",
  3480 => x"00000000",
  3481 => x"00000000",
  3482 => x"00000000",
  3483 => x"00000000",
  3484 => x"00000000",
  3485 => x"00000000",
  3486 => x"00000000",
  3487 => x"00000000",
  3488 => x"00000000",
  3489 => x"00000000",
  3490 => x"00000000",
  3491 => x"00000000",
  3492 => x"00000000",
  3493 => x"00000000",
  3494 => x"00000000",
  3495 => x"00000000",
  3496 => x"00000000",
  3497 => x"00000000",
  3498 => x"00000000",
  3499 => x"00000000",
  3500 => x"00000000",
  3501 => x"00000000",
  3502 => x"00000001",
  3503 => x"330eabcd",
  3504 => x"1234e66d",
  3505 => x"deec0005",
  3506 => x"000b0000",
  3507 => x"00000000",
  3508 => x"00000000",
  3509 => x"00000000",
  3510 => x"00000000",
  3511 => x"00000000",
  3512 => x"00000000",
  3513 => x"00000000",
  3514 => x"00000000",
  3515 => x"00000000",
  3516 => x"00000000",
  3517 => x"00000000",
  3518 => x"00000000",
  3519 => x"00000000",
  3520 => x"00000000",
  3521 => x"00000000",
  3522 => x"00000000",
  3523 => x"00000000",
  3524 => x"00000000",
  3525 => x"00000000",
  3526 => x"00000000",
  3527 => x"00000000",
  3528 => x"00000000",
  3529 => x"00000000",
  3530 => x"00000000",
  3531 => x"00000000",
  3532 => x"00000000",
  3533 => x"00000000",
  3534 => x"00000000",
  3535 => x"00000000",
  3536 => x"00000000",
  3537 => x"00000000",
  3538 => x"00000000",
  3539 => x"00000000",
  3540 => x"00000000",
  3541 => x"00000000",
  3542 => x"00000000",
  3543 => x"00000000",
  3544 => x"00000000",
  3545 => x"00000000",
  3546 => x"00000000",
  3547 => x"00000000",
  3548 => x"00000000",
  3549 => x"00000000",
  3550 => x"00000000",
  3551 => x"00000000",
  3552 => x"00000000",
  3553 => x"00000000",
  3554 => x"00000000",
  3555 => x"00000000",
  3556 => x"00000000",
  3557 => x"00000000",
  3558 => x"00000000",
  3559 => x"00000000",
  3560 => x"00000000",
  3561 => x"00000000",
  3562 => x"00000000",
  3563 => x"00000000",
  3564 => x"00000000",
  3565 => x"00000000",
  3566 => x"00000000",
  3567 => x"00000000",
  3568 => x"00000000",
  3569 => x"00000000",
  3570 => x"00000000",
  3571 => x"00000000",
  3572 => x"00000000",
  3573 => x"00000000",
  3574 => x"00000000",
  3575 => x"00000000",
  3576 => x"00000000",
  3577 => x"00000000",
  3578 => x"00000000",
  3579 => x"00000000",
  3580 => x"00000000",
  3581 => x"00000000",
  3582 => x"00000000",
  3583 => x"00000000",
  3584 => x"00000000",
  3585 => x"00000000",
  3586 => x"00000000",
  3587 => x"00000000",
  3588 => x"00000000",
  3589 => x"00000000",
  3590 => x"00000000",
  3591 => x"00000000",
  3592 => x"00000000",
  3593 => x"00000000",
  3594 => x"00000000",
  3595 => x"00000000",
  3596 => x"00000000",
  3597 => x"00000000",
  3598 => x"00000000",
  3599 => x"00000000",
  3600 => x"00000000",
  3601 => x"00000000",
  3602 => x"00000000",
  3603 => x"00000000",
  3604 => x"00000000",
  3605 => x"00000000",
  3606 => x"00000000",
  3607 => x"00000000",
  3608 => x"00000000",
  3609 => x"00000000",
  3610 => x"00000000",
  3611 => x"00000000",
  3612 => x"00000000",
  3613 => x"00000000",
  3614 => x"00000000",
  3615 => x"00000000",
  3616 => x"00000000",
  3617 => x"00000000",
  3618 => x"00000000",
  3619 => x"00000000",
  3620 => x"00000000",
  3621 => x"00000000",
  3622 => x"00000000",
  3623 => x"00000000",
  3624 => x"00000000",
  3625 => x"00000000",
  3626 => x"00000000",
  3627 => x"00000000",
  3628 => x"00000000",
  3629 => x"00000000",
  3630 => x"00000000",
  3631 => x"00000000",
  3632 => x"00000000",
  3633 => x"00000000",
  3634 => x"00000000",
  3635 => x"00000000",
  3636 => x"00000000",
  3637 => x"00000000",
  3638 => x"00000000",
  3639 => x"00000000",
  3640 => x"00000000",
  3641 => x"00000000",
  3642 => x"00000000",
  3643 => x"00000000",
  3644 => x"00000000",
  3645 => x"00000000",
  3646 => x"00000000",
  3647 => x"00000000",
  3648 => x"00000000",
  3649 => x"00000000",
  3650 => x"00000000",
  3651 => x"00000000",
  3652 => x"00000000",
  3653 => x"00000000",
  3654 => x"00000000",
  3655 => x"00000000",
  3656 => x"00000000",
  3657 => x"00000000",
  3658 => x"00000000",
  3659 => x"00000000",
  3660 => x"00000000",
  3661 => x"00000000",
  3662 => x"00000000",
  3663 => x"00000000",
  3664 => x"00000000",
  3665 => x"00000000",
  3666 => x"00000000",
  3667 => x"00000000",
  3668 => x"00000000",
  3669 => x"00000000",
  3670 => x"00000000",
  3671 => x"00000000",
  3672 => x"00000000",
  3673 => x"00000000",
  3674 => x"00000000",
  3675 => x"00000000",
  3676 => x"00000000",
  3677 => x"00000000",
  3678 => x"00000000",
  3679 => x"00000000",
  3680 => x"00000000",
  3681 => x"00000000",
  3682 => x"00000000",
  3683 => x"ffffffff",
  3684 => x"00000000",
  3685 => x"ffffffff",
  3686 => x"00000000",
  3687 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
