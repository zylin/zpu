package version is

    constant version_time_c : string( 1 to 21) := "Feb 10 2012  14:45:31";

end package version;
