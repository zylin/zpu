-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80d6f40c",
     3 => x"3a0b0b80",
     4 => x"cfd60400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80d09f2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80d6",
   162 => x"e0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80ca",
   171 => x"c12d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80cb",
   179 => x"f32d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80d6f00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"c9c03f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80d6f008",
   281 => x"802ea438",
   282 => x"80d6f408",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80de",
   286 => x"ac0c82a0",
   287 => x"800b80de",
   288 => x"b00c8290",
   289 => x"800b80de",
   290 => x"b40c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"deac0cf8",
   294 => x"80808280",
   295 => x"0b80deb0",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"deb40c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80deac0c",
   302 => x"80c0a880",
   303 => x"940b80de",
   304 => x"b00c0b0b",
   305 => x"80d1f40b",
   306 => x"80deb40c",
   307 => x"04ff3d0d",
   308 => x"80deb833",
   309 => x"5170a738",
   310 => x"80d6fc08",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"d6fc0c70",
   315 => x"2d80d6fc",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80de",
   319 => x"b834833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80dea808",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"dea8510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404ff3d",
   333 => x"0d028f05",
   334 => x"33705252",
   335 => x"98e43f71",
   336 => x"5199da3f",
   337 => x"71800c83",
   338 => x"3d0d04f6",
   339 => x"3d0d7c57",
   340 => x"80707179",
   341 => x"08700870",
   342 => x"9b2a8106",
   343 => x"8c1d0c70",
   344 => x"9f2a7094",
   345 => x"1e0c5859",
   346 => x"5b5d5b59",
   347 => x"72792e09",
   348 => x"81069138",
   349 => x"80c0780c",
   350 => x"77087086",
   351 => x"2a810657",
   352 => x"5575f538",
   353 => x"90187008",
   354 => x"708b2a9f",
   355 => x"06901a0c",
   356 => x"5556850a",
   357 => x"0b98180c",
   358 => x"850a0b9c",
   359 => x"180c9418",
   360 => x"53850a73",
   361 => x"0c981854",
   362 => x"850a740c",
   363 => x"800ba018",
   364 => x"0c800ba4",
   365 => x"180c800b",
   366 => x"a8180c80",
   367 => x"0bac180c",
   368 => x"80765555",
   369 => x"94170875",
   370 => x"2e098106",
   371 => x"84de3890",
   372 => x"17085475",
   373 => x"0870832a",
   374 => x"81065153",
   375 => x"72f53873",
   376 => x"8b2bf880",
   377 => x"80808107",
   378 => x"760c7508",
   379 => x"70832a81",
   380 => x"06555573",
   381 => x"f5389018",
   382 => x"56901708",
   383 => x"54750870",
   384 => x"832a8106",
   385 => x"515372f5",
   386 => x"38738b2b",
   387 => x"8207760c",
   388 => x"75087083",
   389 => x"2a810654",
   390 => x"5472f538",
   391 => x"73842a81",
   392 => x"0653ff54",
   393 => x"72883875",
   394 => x"0870902a",
   395 => x"5553738f",
   396 => x"2a810653",
   397 => x"72c33872",
   398 => x"748c2a81",
   399 => x"06575575",
   400 => x"802e859a",
   401 => x"38901708",
   402 => x"90195754",
   403 => x"75087083",
   404 => x"2a810651",
   405 => x"5b7af538",
   406 => x"738b2b80",
   407 => x"c207760c",
   408 => x"75087083",
   409 => x"2a81065c",
   410 => x"547af538",
   411 => x"73842a81",
   412 => x"065bff54",
   413 => x"7a883875",
   414 => x"0870902a",
   415 => x"555b7385",
   416 => x"2c810654",
   417 => x"73963881",
   418 => x"15558386",
   419 => x"d07525ff",
   420 => x"b43880d1",
   421 => x"f8518f85",
   422 => x"3f760858",
   423 => x"800b9018",
   424 => x"08901a58",
   425 => x"555b7508",
   426 => x"70832a81",
   427 => x"06515574",
   428 => x"f538738b",
   429 => x"2b828207",
   430 => x"760c7508",
   431 => x"70832a81",
   432 => x"06565474",
   433 => x"f5387384",
   434 => x"2a810654",
   435 => x"ff557388",
   436 => x"38750870",
   437 => x"902a5653",
   438 => x"90170890",
   439 => x"19575475",
   440 => x"0870832a",
   441 => x"70810651",
   442 => x"515372f3",
   443 => x"38738b2b",
   444 => x"82c20776",
   445 => x"0c750870",
   446 => x"832a7081",
   447 => x"06515454",
   448 => x"72f33873",
   449 => x"842a7081",
   450 => x"065153ff",
   451 => x"54728838",
   452 => x"75087090",
   453 => x"2a555374",
   454 => x"882a8106",
   455 => x"5675802e",
   456 => x"90387388",
   457 => x"2a810656",
   458 => x"75802e85",
   459 => x"3881705b",
   460 => x"5974872a",
   461 => x"81065675",
   462 => x"802e9038",
   463 => x"73872a81",
   464 => x"06567580",
   465 => x"2e853881",
   466 => x"5a805974",
   467 => x"862a8106",
   468 => x"5574802e",
   469 => x"8e387386",
   470 => x"2a810654",
   471 => x"73802e83",
   472 => x"38815978",
   473 => x"842b7a87",
   474 => x"2b077b88",
   475 => x"2b07780c",
   476 => x"80d29451",
   477 => x"8da73f8c",
   478 => x"1708802e",
   479 => x"81c03880",
   480 => x"d29c518d",
   481 => x"983f80d2",
   482 => x"a8518d91",
   483 => x"3f760852",
   484 => x"a0518dac",
   485 => x"3f80d2c0",
   486 => x"518d823f",
   487 => x"79802e81",
   488 => x"be3880d2",
   489 => x"cc518cf5",
   490 => x"3f80d2d0",
   491 => x"518cee3f",
   492 => x"78802e81",
   493 => x"bc3880d2",
   494 => x"d8518ce1",
   495 => x"3f80d2e0",
   496 => x"518cda3f",
   497 => x"84175b81",
   498 => x"1b338518",
   499 => x"34821b33",
   500 => x"86183483",
   501 => x"1b338718",
   502 => x"34841b33",
   503 => x"88183485",
   504 => x"1b338918",
   505 => x"34760888",
   506 => x"117c3381",
   507 => x"1e337188",
   508 => x"2b07720c",
   509 => x"555b8c05",
   510 => x"821c3383",
   511 => x"1d337198",
   512 => x"2b71902b",
   513 => x"07841f33",
   514 => x"70882b72",
   515 => x"07608505",
   516 => x"33710776",
   517 => x"0c5e5c56",
   518 => x"59575a81",
   519 => x"0b800c8c",
   520 => x"3d0d0481",
   521 => x"15557482",
   522 => x"24fec538",
   523 => x"73087083",
   524 => x"2a810659",
   525 => x"5677802e",
   526 => x"ea388055",
   527 => x"ef3980d2",
   528 => x"ec518bd9",
   529 => x"3f80d2a8",
   530 => x"518bd23f",
   531 => x"760852a0",
   532 => x"518bed3f",
   533 => x"80d2c051",
   534 => x"8bc33f79",
   535 => x"fec43880",
   536 => x"d2f4518b",
   537 => x"b83f80d2",
   538 => x"d0518bb1",
   539 => x"3f78fec6",
   540 => x"3880d2f8",
   541 => x"518ba63f",
   542 => x"80d2e051",
   543 => x"8b9f3f84",
   544 => x"175b811b",
   545 => x"33851834",
   546 => x"821b3386",
   547 => x"1834831b",
   548 => x"33871834",
   549 => x"841b3388",
   550 => x"1834851b",
   551 => x"33891834",
   552 => x"76088811",
   553 => x"7c33811e",
   554 => x"3371882b",
   555 => x"07720c55",
   556 => x"5b8c0582",
   557 => x"1c33831d",
   558 => x"3371982b",
   559 => x"71902b07",
   560 => x"841f3370",
   561 => x"882b7207",
   562 => x"60850533",
   563 => x"7107760c",
   564 => x"5e5c5659",
   565 => x"575a810b",
   566 => x"800c8c3d",
   567 => x"0d049017",
   568 => x"08901957",
   569 => x"54750870",
   570 => x"832a8106",
   571 => x"5a5378f5",
   572 => x"38738b2b",
   573 => x"8207760c",
   574 => x"75087083",
   575 => x"2a810656",
   576 => x"5474f538",
   577 => x"73842a81",
   578 => x"0654ff55",
   579 => x"73883875",
   580 => x"0870902a",
   581 => x"5653748d",
   582 => x"2a548c17",
   583 => x"08802e92",
   584 => x"38738106",
   585 => x"56758b38",
   586 => x"74862a81",
   587 => x"06597880",
   588 => x"c9387381",
   589 => x"06567580",
   590 => x"2ea43874",
   591 => x"862a8106",
   592 => x"53729b38",
   593 => x"725b815a",
   594 => x"74882a81",
   595 => x"06597884",
   596 => x"2b7a872b",
   597 => x"077b882b",
   598 => x"07780cfc",
   599 => x"93397381",
   600 => x"065372e4",
   601 => x"3874862a",
   602 => x"81065372",
   603 => x"db387273",
   604 => x"76882a81",
   605 => x"065b5c5a",
   606 => x"d5398176",
   607 => x"76882a81",
   608 => x"065b5b5b",
   609 => x"c939ff3d",
   610 => x"0d739811",
   611 => x"085151bf",
   612 => x"5280710c",
   613 => x"ff128812",
   614 => x"52527180",
   615 => x"25f33883",
   616 => x"3d0d04fb",
   617 => x"3d0d777a",
   618 => x"981108a0",
   619 => x"12081010",
   620 => x"10117008",
   621 => x"708b2a81",
   622 => x"06515956",
   623 => x"54555680",
   624 => x"5174712e",
   625 => x"098106ad",
   626 => x"38788414",
   627 => x"0ca01408",
   628 => x"5170bf2e",
   629 => x"a7387010",
   630 => x"10101276",
   631 => x"90800771",
   632 => x"0c55a014",
   633 => x"088105a0",
   634 => x"150c7308",
   635 => x"70088107",
   636 => x"710c5681",
   637 => x"5170800c",
   638 => x"873d0d04",
   639 => x"83f81276",
   640 => x"b0800771",
   641 => x"0c5274a0",
   642 => x"150c7308",
   643 => x"70088107",
   644 => x"710c5681",
   645 => x"51df39fd",
   646 => x"3d0d75a8",
   647 => x"11087010",
   648 => x"10109813",
   649 => x"08057008",
   650 => x"708b2c70",
   651 => x"81065152",
   652 => x"57535353",
   653 => x"80547074",
   654 => x"2e098106",
   655 => x"8d3871bf",
   656 => x"2e8f3881",
   657 => x"12a8140c",
   658 => x"81547380",
   659 => x"0c853d0d",
   660 => x"0470a814",
   661 => x"0c8154f2",
   662 => x"39ee3d0d",
   663 => x"80d78408",
   664 => x"7008810a",
   665 => x"065c5781",
   666 => x"ff0b8818",
   667 => x"0c8f8a3f",
   668 => x"8de93f8e",
   669 => x"973f9bed",
   670 => x"567a8438",
   671 => x"8ab25675",
   672 => x"80deec0c",
   673 => x"80d38051",
   674 => x"87933f7a",
   675 => x"802e8589",
   676 => x"3880d38c",
   677 => x"5187863f",
   678 => x"f8808098",
   679 => x"800b80de",
   680 => x"bc0c800b",
   681 => x"fa808085",
   682 => x"80349b0b",
   683 => x"fa808085",
   684 => x"8134a10b",
   685 => x"fa808085",
   686 => x"823480e7",
   687 => x"0bfa8080",
   688 => x"858334ff",
   689 => x"b80bfa80",
   690 => x"80858434",
   691 => x"ffb80bfa",
   692 => x"80808585",
   693 => x"34de0bfa",
   694 => x"80808586",
   695 => x"34ffad0b",
   696 => x"fa808085",
   697 => x"8734ffbe",
   698 => x"0bfa8080",
   699 => x"858834ef",
   700 => x"0bfa8080",
   701 => x"85893480",
   702 => x"0bfa8080",
   703 => x"858a34a0",
   704 => x"0bfa8080",
   705 => x"858b3485",
   706 => x"0bfa8080",
   707 => x"858c34dc",
   708 => x"0bfa8080",
   709 => x"858d3480",
   710 => x"d7840858",
   711 => x"810b8419",
   712 => x"0c8653fa",
   713 => x"80808586",
   714 => x"5280dec0",
   715 => x"51b88e3f",
   716 => x"80d78408",
   717 => x"56820b84",
   718 => x"170c8059",
   719 => x"8e5a7aab",
   720 => x"38fa8080",
   721 => x"85801a5d",
   722 => x"797d3481",
   723 => x"1a7a7126",
   724 => x"7a057072",
   725 => x"5d5b5858",
   726 => x"7680268a",
   727 => x"3876e238",
   728 => x"8be97827",
   729 => x"dc3880d7",
   730 => x"84085683",
   731 => x"0b84170c",
   732 => x"80debc51",
   733 => x"f3d53f80",
   734 => x"debc51fc",
   735 => x"893f80d7",
   736 => x"84085984",
   737 => x"0b841a0c",
   738 => x"80d39851",
   739 => x"858f3f80",
   740 => x"59805afa",
   741 => x"80808580",
   742 => x"1a703353",
   743 => x"5e885185",
   744 => x"9f3f7886",
   745 => x"3879852e",
   746 => x"8638ba51",
   747 => x"84d53f81",
   748 => x"1a7a7126",
   749 => x"7a057072",
   750 => x"5d5b5858",
   751 => x"76802689",
   752 => x"3876d038",
   753 => x"857827cb",
   754 => x"388a5184",
   755 => x"b63f805d",
   756 => x"80c05e7a",
   757 => x"8738805d",
   758 => x"90800a5e",
   759 => x"a85184a3",
   760 => x"3f7d5185",
   761 => x"fd3f80d3",
   762 => x"b85184b1",
   763 => x"3f805b80",
   764 => x"0b80d784",
   765 => x"08585c85",
   766 => x"0b84180c",
   767 => x"8ab13f80",
   768 => x"085f7c80",
   769 => x"268b387c",
   770 => x"80d13880",
   771 => x"7e2780cb",
   772 => x"387a982b",
   773 => x"7c882a07",
   774 => x"81ff0680",
   775 => x"d784085b",
   776 => x"841b0c80",
   777 => x"debc53fa",
   778 => x"80808580",
   779 => x"528bea51",
   780 => x"faf13f80",
   781 => x"089f2c80",
   782 => x"081d7d71",
   783 => x"265a5b7b",
   784 => x"05780570",
   785 => x"7b5e5c59",
   786 => x"7c7926c5",
   787 => x"387c792e",
   788 => x"09810687",
   789 => x"387d7a26",
   790 => x"ffb73880",
   791 => x"5b805c7b",
   792 => x"81ff0680",
   793 => x"d784085b",
   794 => x"841b0c80",
   795 => x"debc51fb",
   796 => x"a63f8008",
   797 => x"9f2c8008",
   798 => x"1d7d7126",
   799 => x"595b7b05",
   800 => x"7705707b",
   801 => x"5e5c5978",
   802 => x"80268938",
   803 => x"78d138bf",
   804 => x"7a27cc38",
   805 => x"89993f80",
   806 => x"d7840857",
   807 => x"81ff0b84",
   808 => x"180c7e80",
   809 => x"083180d3",
   810 => x"c4525982",
   811 => x"f03f7851",
   812 => x"85ec3f80",
   813 => x"d3d05182",
   814 => x"e43f923d",
   815 => x"5a805c80",
   816 => x"dde07c55",
   817 => x"557c527d",
   818 => x"5379518b",
   819 => x"d33f805d",
   820 => x"87e87d55",
   821 => x"55616359",
   822 => x"52775379",
   823 => x"518bc13f",
   824 => x"80547855",
   825 => x"61635f52",
   826 => x"7d53943d",
   827 => x"f005518f",
   828 => x"8b3f6080",
   829 => x"d3d8525b",
   830 => x"82a33f7a",
   831 => x"56807b24",
   832 => x"81d23875",
   833 => x"8a2c5183",
   834 => x"d93f80d3",
   835 => x"e451828d",
   836 => x"3f800b80",
   837 => x"0c943d0d",
   838 => x"0480d3ec",
   839 => x"5181fe3f",
   840 => x"80d3fc51",
   841 => x"81f73ff8",
   842 => x"80809880",
   843 => x"0b80debc",
   844 => x"0c800bfa",
   845 => x"80808580",
   846 => x"349b0bfa",
   847 => x"80808581",
   848 => x"34a10bfa",
   849 => x"80808582",
   850 => x"3480e70b",
   851 => x"fa808085",
   852 => x"8334ffb8",
   853 => x"0bfa8080",
   854 => x"858434ff",
   855 => x"b80bfa80",
   856 => x"80858534",
   857 => x"de0bfa80",
   858 => x"80858634",
   859 => x"ffad0bfa",
   860 => x"80808587",
   861 => x"34ffbe0b",
   862 => x"fa808085",
   863 => x"8834ef0b",
   864 => x"fa808085",
   865 => x"8934800b",
   866 => x"fa808085",
   867 => x"8a34a00b",
   868 => x"fa808085",
   869 => x"8b34850b",
   870 => x"fa808085",
   871 => x"8c34dc0b",
   872 => x"fa808085",
   873 => x"8d3480d7",
   874 => x"84085881",
   875 => x"0b84190c",
   876 => x"8653fa80",
   877 => x"80858652",
   878 => x"80dec051",
   879 => x"b2ff3f80",
   880 => x"d7840856",
   881 => x"820b8417",
   882 => x"0c80598e",
   883 => x"5a7afb9b",
   884 => x"38faee39",
   885 => x"87ff1b70",
   886 => x"8a2c5256",
   887 => x"82843f80",
   888 => x"d3e451b9",
   889 => x"3f800b80",
   890 => x"0c943d0d",
   891 => x"04ff3d0d",
   892 => x"028f0533",
   893 => x"80d78008",
   894 => x"52710c80",
   895 => x"0b800c83",
   896 => x"3d0d04ff",
   897 => x"3d0d028f",
   898 => x"05335180",
   899 => x"deec0852",
   900 => x"712d8008",
   901 => x"81ff0680",
   902 => x"0c833d0d",
   903 => x"04fe3d0d",
   904 => x"74703353",
   905 => x"5371802e",
   906 => x"93388113",
   907 => x"725280de",
   908 => x"ec085353",
   909 => x"712d7233",
   910 => x"5271ef38",
   911 => x"843d0d04",
   912 => x"f43d0d7f",
   913 => x"028405bb",
   914 => x"05335557",
   915 => x"880b8c3d",
   916 => x"5a5a8953",
   917 => x"80d4c452",
   918 => x"7851b1e1",
   919 => x"3f737a2e",
   920 => x"80fa3879",
   921 => x"5673902e",
   922 => x"80e73802",
   923 => x"a7055876",
   924 => x"8f065473",
   925 => x"8926bf38",
   926 => x"7518b015",
   927 => x"55557375",
   928 => x"3476842a",
   929 => x"ff177081",
   930 => x"ff065855",
   931 => x"5775e038",
   932 => x"79195575",
   933 => x"75347870",
   934 => x"33555573",
   935 => x"802e9338",
   936 => x"81157452",
   937 => x"80deec08",
   938 => x"5755752d",
   939 => x"74335473",
   940 => x"ef388e3d",
   941 => x"0d047518",
   942 => x"b7155555",
   943 => x"73753476",
   944 => x"842aff17",
   945 => x"7081ff06",
   946 => x"58555775",
   947 => x"ffa138c0",
   948 => x"39847057",
   949 => x"5a02a705",
   950 => x"58ff9439",
   951 => x"8270575a",
   952 => x"f439f23d",
   953 => x"0d608c3d",
   954 => x"705b5b53",
   955 => x"80735657",
   956 => x"76732480",
   957 => x"f8387817",
   958 => x"548a5274",
   959 => x"51ac9d3f",
   960 => x"8008b005",
   961 => x"53727434",
   962 => x"8117578a",
   963 => x"527451ab",
   964 => x"e63f8008",
   965 => x"558008de",
   966 => x"38800877",
   967 => x"9f2a1870",
   968 => x"812c5a56",
   969 => x"56807825",
   970 => x"9e387817",
   971 => x"ff055575",
   972 => x"19703355",
   973 => x"53743373",
   974 => x"34737534",
   975 => x"8116ff16",
   976 => x"56567776",
   977 => x"24e93876",
   978 => x"19568076",
   979 => x"34797033",
   980 => x"54547280",
   981 => x"2e933881",
   982 => x"14735280",
   983 => x"deec0858",
   984 => x"54762d73",
   985 => x"335372ef",
   986 => x"38903d0d",
   987 => x"04ad7a34",
   988 => x"02a90573",
   989 => x"30711956",
   990 => x"56598a52",
   991 => x"7451ab9c",
   992 => x"3f8008b0",
   993 => x"05537274",
   994 => x"34811757",
   995 => x"8a527451",
   996 => x"aae53f80",
   997 => x"08558008",
   998 => x"fedc38fe",
   999 => x"fc39ec3d",
  1000 => x"0d665b87",
  1001 => x"e8527a51",
  1002 => x"aacd3f91",
  1003 => x"3d705a5a",
  1004 => x"800b8008",
  1005 => x"56577680",
  1006 => x"0824828e",
  1007 => x"38781754",
  1008 => x"8a527451",
  1009 => x"aad63f80",
  1010 => x"08b00553",
  1011 => x"72743481",
  1012 => x"17578a52",
  1013 => x"7451aa9f",
  1014 => x"3f800855",
  1015 => x"8008de38",
  1016 => x"8008779f",
  1017 => x"2a187081",
  1018 => x"2c5a5656",
  1019 => x"8078259e",
  1020 => x"387817ff",
  1021 => x"05557519",
  1022 => x"70335553",
  1023 => x"74337334",
  1024 => x"73753481",
  1025 => x"16ff1656",
  1026 => x"56777624",
  1027 => x"e9387619",
  1028 => x"56807634",
  1029 => x"79703354",
  1030 => x"5472802e",
  1031 => x"93388114",
  1032 => x"735280de",
  1033 => x"ec085854",
  1034 => x"762d7333",
  1035 => x"5372ef38",
  1036 => x"ae5180de",
  1037 => x"ec085877",
  1038 => x"2d87e852",
  1039 => x"7a51a9dc",
  1040 => x"3f8c3d70",
  1041 => x"5a5a800b",
  1042 => x"80085657",
  1043 => x"76800824",
  1044 => x"81ab3878",
  1045 => x"175b8a52",
  1046 => x"7451a9c0",
  1047 => x"3f8008b0",
  1048 => x"0554737b",
  1049 => x"34811757",
  1050 => x"8a527451",
  1051 => x"a9893f80",
  1052 => x"08558008",
  1053 => x"de388008",
  1054 => x"779f2a18",
  1055 => x"70812c5a",
  1056 => x"56568078",
  1057 => x"259e3878",
  1058 => x"17ff0555",
  1059 => x"75197033",
  1060 => x"5c537433",
  1061 => x"73347a75",
  1062 => x"348116ff",
  1063 => x"16565677",
  1064 => x"7624e938",
  1065 => x"76195680",
  1066 => x"76347970",
  1067 => x"33545472",
  1068 => x"802e9338",
  1069 => x"81147352",
  1070 => x"80deec08",
  1071 => x"5a54782d",
  1072 => x"73335372",
  1073 => x"ef38963d",
  1074 => x"0d04ad7a",
  1075 => x"340280c1",
  1076 => x"05800830",
  1077 => x"71195656",
  1078 => x"598a5274",
  1079 => x"51a8bd3f",
  1080 => x"8008b005",
  1081 => x"53727434",
  1082 => x"8117578a",
  1083 => x"527451a8",
  1084 => x"863f8008",
  1085 => x"558008fd",
  1086 => x"c438fde4",
  1087 => x"39ad7a34",
  1088 => x"02ad0580",
  1089 => x"08307119",
  1090 => x"5d56598a",
  1091 => x"527451a8",
  1092 => x"8b3f8008",
  1093 => x"b0055473",
  1094 => x"7b348117",
  1095 => x"578a5274",
  1096 => x"51a7d43f",
  1097 => x"80085580",
  1098 => x"08fea838",
  1099 => x"fec839fb",
  1100 => x"3d0d80d7",
  1101 => x"8c08a811",
  1102 => x"08fe06a8",
  1103 => x"120cb011",
  1104 => x"08a01208",
  1105 => x"a8130870",
  1106 => x"8107a815",
  1107 => x"0c567187",
  1108 => x"e8290580",
  1109 => x"0c575487",
  1110 => x"3d0d0480",
  1111 => x"3d0d80d7",
  1112 => x"8c085187",
  1113 => x"0b84120c",
  1114 => x"ff0bb412",
  1115 => x"0ca70bb8",
  1116 => x"120c87e8",
  1117 => x"0ba4120c",
  1118 => x"a70ba812",
  1119 => x"0cb0ea0b",
  1120 => x"94120c87",
  1121 => x"0b98120c",
  1122 => x"823d0d04",
  1123 => x"803d0d80",
  1124 => x"d7900851",
  1125 => x"b60b8c12",
  1126 => x"0c830b88",
  1127 => x"120c823d",
  1128 => x"0d04fe3d",
  1129 => x"0d029305",
  1130 => x"3353728a",
  1131 => x"2e9e3880",
  1132 => x"d7900852",
  1133 => x"84120870",
  1134 => x"822a7081",
  1135 => x"06515151",
  1136 => x"70802ef0",
  1137 => x"3872720c",
  1138 => x"843d0d04",
  1139 => x"80d79008",
  1140 => x"52841208",
  1141 => x"70822a70",
  1142 => x"81065151",
  1143 => x"5170802e",
  1144 => x"f0388d72",
  1145 => x"0c841208",
  1146 => x"70822a70",
  1147 => x"81065151",
  1148 => x"5170802e",
  1149 => x"ffbe38cd",
  1150 => x"39803d0d",
  1151 => x"80d78808",
  1152 => x"51800b84",
  1153 => x"120c83fe",
  1154 => x"800b8812",
  1155 => x"0c800b80",
  1156 => x"def03480",
  1157 => x"0b80def4",
  1158 => x"34823d0d",
  1159 => x"04fa3d0d",
  1160 => x"02a30533",
  1161 => x"80d78808",
  1162 => x"80def033",
  1163 => x"7081ff06",
  1164 => x"70101011",
  1165 => x"80def433",
  1166 => x"7081ff06",
  1167 => x"72902911",
  1168 => x"70882b78",
  1169 => x"07770c53",
  1170 => x"5b5b5555",
  1171 => x"59545473",
  1172 => x"8a2e9838",
  1173 => x"7480cf2e",
  1174 => x"9238738c",
  1175 => x"2ea43881",
  1176 => x"16537280",
  1177 => x"def43488",
  1178 => x"3d0d0471",
  1179 => x"a326a338",
  1180 => x"81175271",
  1181 => x"80def034",
  1182 => x"800b80de",
  1183 => x"f434883d",
  1184 => x"0d048052",
  1185 => x"71882b73",
  1186 => x"0c811252",
  1187 => x"97907226",
  1188 => x"f338800b",
  1189 => x"80def034",
  1190 => x"800b80de",
  1191 => x"f434df39",
  1192 => x"8c08028c",
  1193 => x"0ceb3d0d",
  1194 => x"800b8c08",
  1195 => x"f0050c80",
  1196 => x"0b8c08f4",
  1197 => x"050c8c08",
  1198 => x"8c05088c",
  1199 => x"08900508",
  1200 => x"5654738c",
  1201 => x"08f0050c",
  1202 => x"748c08f4",
  1203 => x"050c8c08",
  1204 => x"f8058c08",
  1205 => x"f0055656",
  1206 => x"88705475",
  1207 => x"53765254",
  1208 => x"a8db3f80",
  1209 => x"0b8c08e8",
  1210 => x"050c800b",
  1211 => x"8c08ec05",
  1212 => x"0c8c0894",
  1213 => x"05088c08",
  1214 => x"98050856",
  1215 => x"54738c08",
  1216 => x"e8050c74",
  1217 => x"8c08ec05",
  1218 => x"0c8c08f0",
  1219 => x"058c08e8",
  1220 => x"05565688",
  1221 => x"70547553",
  1222 => x"765254a8",
  1223 => x"a03f800b",
  1224 => x"8c08e805",
  1225 => x"0c800b8c",
  1226 => x"08ec050c",
  1227 => x"8c08fc05",
  1228 => x"0883ffff",
  1229 => x"068c08cc",
  1230 => x"050c8c08",
  1231 => x"fc050890",
  1232 => x"2a8c08c4",
  1233 => x"050c8c08",
  1234 => x"f4050883",
  1235 => x"ffff068c",
  1236 => x"08c8050c",
  1237 => x"8c08f405",
  1238 => x"08902a8c",
  1239 => x"08c0050c",
  1240 => x"8c08cc05",
  1241 => x"088c08c8",
  1242 => x"05082970",
  1243 => x"8c08dc05",
  1244 => x"0c8c08cc",
  1245 => x"05088c08",
  1246 => x"c0050829",
  1247 => x"708c08d8",
  1248 => x"050c8c08",
  1249 => x"c405088c",
  1250 => x"08c80508",
  1251 => x"29708c08",
  1252 => x"d4050c8c",
  1253 => x"08c40508",
  1254 => x"8c08c005",
  1255 => x"0829708c",
  1256 => x"08d0050c",
  1257 => x"8c08dc05",
  1258 => x"08902a8c",
  1259 => x"08d80508",
  1260 => x"118c08d8",
  1261 => x"050c8c08",
  1262 => x"d805088c",
  1263 => x"08d40508",
  1264 => x"058c08d8",
  1265 => x"050c5151",
  1266 => x"5151548c",
  1267 => x"08d80508",
  1268 => x"8c08d405",
  1269 => x"08278f38",
  1270 => x"8c08d005",
  1271 => x"08848080",
  1272 => x"058c08d0",
  1273 => x"050c8c08",
  1274 => x"d8050890",
  1275 => x"2a8c08d0",
  1276 => x"0508118c",
  1277 => x"08e0050c",
  1278 => x"8c08d805",
  1279 => x"0883ffff",
  1280 => x"0670902b",
  1281 => x"8c08dc05",
  1282 => x"0883ffff",
  1283 => x"0670128c",
  1284 => x"08e4050c",
  1285 => x"52575154",
  1286 => x"8c08e005",
  1287 => x"088c08e4",
  1288 => x"05085654",
  1289 => x"738c08e8",
  1290 => x"050c748c",
  1291 => x"08ec050c",
  1292 => x"8c08fc05",
  1293 => x"088c08f0",
  1294 => x"0508298c",
  1295 => x"08f80508",
  1296 => x"8c08f405",
  1297 => x"08297012",
  1298 => x"8c08e805",
  1299 => x"08118c08",
  1300 => x"e8050c51",
  1301 => x"55558c08",
  1302 => x"e805088c",
  1303 => x"08ec0508",
  1304 => x"8c088805",
  1305 => x"08585654",
  1306 => x"73760c74",
  1307 => x"84170c8c",
  1308 => x"08880508",
  1309 => x"800c973d",
  1310 => x"0d8c0c04",
  1311 => x"8c08028c",
  1312 => x"0cd43d0d",
  1313 => x"8c088c05",
  1314 => x"088c0890",
  1315 => x"05085553",
  1316 => x"728c08f8",
  1317 => x"050c738c",
  1318 => x"08fc050c",
  1319 => x"8c089405",
  1320 => x"088c0898",
  1321 => x"05085553",
  1322 => x"728c08f0",
  1323 => x"050c738c",
  1324 => x"08f4050c",
  1325 => x"800b8c08",
  1326 => x"ec050c80",
  1327 => x"0b8c08dc",
  1328 => x"050c800b",
  1329 => x"8c08e005",
  1330 => x"0c8c08f8",
  1331 => x"05088c08",
  1332 => x"fc050855",
  1333 => x"53728c08",
  1334 => x"dc050c73",
  1335 => x"8c08e005",
  1336 => x"0c800b8c",
  1337 => x"08d4050c",
  1338 => x"800b8c08",
  1339 => x"d8050c8c",
  1340 => x"08f00508",
  1341 => x"8c08f405",
  1342 => x"08555372",
  1343 => x"8c08d405",
  1344 => x"0c738c08",
  1345 => x"d8050c8c",
  1346 => x"08d80508",
  1347 => x"8c08c805",
  1348 => x"0c8c08d4",
  1349 => x"05088c08",
  1350 => x"c4050c8c",
  1351 => x"08e00508",
  1352 => x"8c08c005",
  1353 => x"0c8c08dc",
  1354 => x"05088c08",
  1355 => x"ffbc050c",
  1356 => x"8c08c405",
  1357 => x"0891a038",
  1358 => x"8c08ffbc",
  1359 => x"05088c08",
  1360 => x"c8050827",
  1361 => x"85fb388c",
  1362 => x"08c80508",
  1363 => x"8c08ffa4",
  1364 => x"050c8c08",
  1365 => x"ffa40508",
  1366 => x"83ffff26",
  1367 => x"a0388c08",
  1368 => x"ffa40508",
  1369 => x"81ff268b",
  1370 => x"38800b8c",
  1371 => x"08fef405",
  1372 => x"0ca93988",
  1373 => x"0b8c08fe",
  1374 => x"f4050c9f",
  1375 => x"398c08ff",
  1376 => x"a40508fe",
  1377 => x"800a268b",
  1378 => x"38900b8c",
  1379 => x"08fef405",
  1380 => x"0c893998",
  1381 => x"0b8c08fe",
  1382 => x"f4050c8c",
  1383 => x"08fef405",
  1384 => x"088c08ff",
  1385 => x"a0050c8c",
  1386 => x"08ffa405",
  1387 => x"088c08ff",
  1388 => x"a005082a",
  1389 => x"80d4d011",
  1390 => x"338c08ff",
  1391 => x"a0050811",
  1392 => x"a071318c",
  1393 => x"08ffa805",
  1394 => x"0c515153",
  1395 => x"8c08ffa8",
  1396 => x"0508802e",
  1397 => x"80cc388c",
  1398 => x"08c80508",
  1399 => x"8c08ffa8",
  1400 => x"05082b8c",
  1401 => x"08c8050c",
  1402 => x"8c08ffbc",
  1403 => x"05088c08",
  1404 => x"ffa80508",
  1405 => x"2ba00b8c",
  1406 => x"08ffa805",
  1407 => x"08318c08",
  1408 => x"c0050871",
  1409 => x"2a707307",
  1410 => x"8c08ffbc",
  1411 => x"050c8c08",
  1412 => x"c005088c",
  1413 => x"08ffa805",
  1414 => x"082b8c08",
  1415 => x"c0050c51",
  1416 => x"55538c08",
  1417 => x"c8050890",
  1418 => x"2a8c08ff",
  1419 => x"a0050c8c",
  1420 => x"08c80508",
  1421 => x"83ffff06",
  1422 => x"8c08ffa4",
  1423 => x"050c8c08",
  1424 => x"ffbc0508",
  1425 => x"8c08ffa0",
  1426 => x"05085370",
  1427 => x"52539dcc",
  1428 => x"3f800870",
  1429 => x"8c08ff94",
  1430 => x"050c8c08",
  1431 => x"ffa00508",
  1432 => x"538c08ff",
  1433 => x"bc050852",
  1434 => x"539d8c3f",
  1435 => x"8008708c",
  1436 => x"08ff9c05",
  1437 => x"0c8c08ff",
  1438 => x"9c05088c",
  1439 => x"08ffa405",
  1440 => x"0829708c",
  1441 => x"08ff8c05",
  1442 => x"0c8c08ff",
  1443 => x"94050870",
  1444 => x"902b8c08",
  1445 => x"c0050890",
  1446 => x"2a707207",
  1447 => x"8c08ff94",
  1448 => x"050c5257",
  1449 => x"5151538c",
  1450 => x"08ff9405",
  1451 => x"088c08ff",
  1452 => x"8c050827",
  1453 => x"80de388c",
  1454 => x"08ff9c05",
  1455 => x"08ff058c",
  1456 => x"08ff9c05",
  1457 => x"0c8c08ff",
  1458 => x"9405088c",
  1459 => x"08c80508",
  1460 => x"058c08ff",
  1461 => x"94050c8c",
  1462 => x"08c80508",
  1463 => x"8c08ff94",
  1464 => x"050826b0",
  1465 => x"388c08ff",
  1466 => x"9405088c",
  1467 => x"08ff8c05",
  1468 => x"0827a138",
  1469 => x"8c08ff9c",
  1470 => x"0508ff05",
  1471 => x"8c08ff9c",
  1472 => x"050c8c08",
  1473 => x"ff940508",
  1474 => x"8c08c805",
  1475 => x"08058c08",
  1476 => x"ff94050c",
  1477 => x"8c08ff94",
  1478 => x"05088c08",
  1479 => x"ff8c0508",
  1480 => x"318c08ff",
  1481 => x"94050c8c",
  1482 => x"08ff9405",
  1483 => x"088c08ff",
  1484 => x"a0050853",
  1485 => x"7052539b",
  1486 => x"e33f8008",
  1487 => x"708c08ff",
  1488 => x"90050c8c",
  1489 => x"08ffa005",
  1490 => x"08538c08",
  1491 => x"ff940508",
  1492 => x"52539ba3",
  1493 => x"3f800870",
  1494 => x"8c08ff98",
  1495 => x"050c8c08",
  1496 => x"ff980508",
  1497 => x"8c08ffa4",
  1498 => x"05082970",
  1499 => x"8c08ff8c",
  1500 => x"050c8c08",
  1501 => x"ff900508",
  1502 => x"70902b8c",
  1503 => x"08c00508",
  1504 => x"83ffff06",
  1505 => x"7072078c",
  1506 => x"08ff9005",
  1507 => x"0c525751",
  1508 => x"51538c08",
  1509 => x"ff900508",
  1510 => x"8c08ff8c",
  1511 => x"05082780",
  1512 => x"de388c08",
  1513 => x"ff980508",
  1514 => x"ff058c08",
  1515 => x"ff98050c",
  1516 => x"8c08ff90",
  1517 => x"05088c08",
  1518 => x"c8050805",
  1519 => x"8c08ff90",
  1520 => x"050c8c08",
  1521 => x"c805088c",
  1522 => x"08ff9005",
  1523 => x"0826b038",
  1524 => x"8c08ff90",
  1525 => x"05088c08",
  1526 => x"ff8c0508",
  1527 => x"27a1388c",
  1528 => x"08ff9805",
  1529 => x"08ff058c",
  1530 => x"08ff9805",
  1531 => x"0c8c08ff",
  1532 => x"9005088c",
  1533 => x"08c80508",
  1534 => x"058c08ff",
  1535 => x"90050c8c",
  1536 => x"08ff9005",
  1537 => x"088c08ff",
  1538 => x"8c050831",
  1539 => x"8c08ff90",
  1540 => x"050c8c08",
  1541 => x"ff9c0508",
  1542 => x"70902b70",
  1543 => x"8c08ff98",
  1544 => x"0508078c",
  1545 => x"08ffb405",
  1546 => x"0c8c08ff",
  1547 => x"9005088c",
  1548 => x"08c0050c",
  1549 => x"5153800b",
  1550 => x"8c08ffb0",
  1551 => x"050c8ad9",
  1552 => x"398c08c8",
  1553 => x"05089538",
  1554 => x"8c08c805",
  1555 => x"08528151",
  1556 => x"99a53f80",
  1557 => x"08708c08",
  1558 => x"c8050c53",
  1559 => x"8c08c805",
  1560 => x"088c08ff",
  1561 => x"8c050c8c",
  1562 => x"08ff8c05",
  1563 => x"0883ffff",
  1564 => x"26a0388c",
  1565 => x"08ff8c05",
  1566 => x"0881ff26",
  1567 => x"8b38800b",
  1568 => x"8c08fef0",
  1569 => x"050ca939",
  1570 => x"880b8c08",
  1571 => x"fef0050c",
  1572 => x"9f398c08",
  1573 => x"ff8c0508",
  1574 => x"fe800a26",
  1575 => x"8b38900b",
  1576 => x"8c08fef0",
  1577 => x"050c8939",
  1578 => x"980b8c08",
  1579 => x"fef0050c",
  1580 => x"8c08fef0",
  1581 => x"05088c08",
  1582 => x"ff90050c",
  1583 => x"8c08ff8c",
  1584 => x"05088c08",
  1585 => x"ff900508",
  1586 => x"2a80d4d0",
  1587 => x"11338c08",
  1588 => x"ff900508",
  1589 => x"11a07131",
  1590 => x"8c08ffa8",
  1591 => x"050c5151",
  1592 => x"538c08ff",
  1593 => x"a805089e",
  1594 => x"388c08ff",
  1595 => x"bc05088c",
  1596 => x"08c80508",
  1597 => x"318c08ff",
  1598 => x"bc050c81",
  1599 => x"0b8c08ff",
  1600 => x"b0050c85",
  1601 => x"8039a00b",
  1602 => x"8c08ffa8",
  1603 => x"0508318c",
  1604 => x"08ffac05",
  1605 => x"0c8c08c8",
  1606 => x"05088c08",
  1607 => x"ffa80508",
  1608 => x"2b8c08c8",
  1609 => x"050c8c08",
  1610 => x"ffbc0508",
  1611 => x"8c08ffac",
  1612 => x"05082a8c",
  1613 => x"08ffb805",
  1614 => x"0c8c08ff",
  1615 => x"bc05088c",
  1616 => x"08ffa805",
  1617 => x"082b8c08",
  1618 => x"c005088c",
  1619 => x"08ffac05",
  1620 => x"082a7072",
  1621 => x"078c08ff",
  1622 => x"bc050c8c",
  1623 => x"08c00508",
  1624 => x"8c08ffa8",
  1625 => x"05082b8c",
  1626 => x"08c0050c",
  1627 => x"8c08c805",
  1628 => x"08902a8c",
  1629 => x"08ff8c05",
  1630 => x"0c8c08c8",
  1631 => x"050883ff",
  1632 => x"ff068c08",
  1633 => x"ff90050c",
  1634 => x"8c08ffb8",
  1635 => x"05088c08",
  1636 => x"ff8c0508",
  1637 => x"55705451",
  1638 => x"54549780",
  1639 => x"3f800870",
  1640 => x"8c08ff9c",
  1641 => x"050c8c08",
  1642 => x"ff8c0508",
  1643 => x"538c08ff",
  1644 => x"b8050852",
  1645 => x"5396c03f",
  1646 => x"8008708c",
  1647 => x"08ff9405",
  1648 => x"0c8c08ff",
  1649 => x"9405088c",
  1650 => x"08ff9005",
  1651 => x"0829708c",
  1652 => x"08ffa405",
  1653 => x"0c8c08ff",
  1654 => x"9c050870",
  1655 => x"902b8c08",
  1656 => x"ffbc0508",
  1657 => x"902a7072",
  1658 => x"078c08ff",
  1659 => x"9c050c52",
  1660 => x"57515153",
  1661 => x"8c08ff9c",
  1662 => x"05088c08",
  1663 => x"ffa40508",
  1664 => x"2780de38",
  1665 => x"8c08ff94",
  1666 => x"0508ff05",
  1667 => x"8c08ff94",
  1668 => x"050c8c08",
  1669 => x"ff9c0508",
  1670 => x"8c08c805",
  1671 => x"08058c08",
  1672 => x"ff9c050c",
  1673 => x"8c08c805",
  1674 => x"088c08ff",
  1675 => x"9c050826",
  1676 => x"b0388c08",
  1677 => x"ff9c0508",
  1678 => x"8c08ffa4",
  1679 => x"050827a1",
  1680 => x"388c08ff",
  1681 => x"940508ff",
  1682 => x"058c08ff",
  1683 => x"94050c8c",
  1684 => x"08ff9c05",
  1685 => x"088c08c8",
  1686 => x"0508058c",
  1687 => x"08ff9c05",
  1688 => x"0c8c08ff",
  1689 => x"9c05088c",
  1690 => x"08ffa405",
  1691 => x"08318c08",
  1692 => x"ff9c050c",
  1693 => x"8c08ff9c",
  1694 => x"05088c08",
  1695 => x"ff8c0508",
  1696 => x"53705253",
  1697 => x"95963f80",
  1698 => x"08708c08",
  1699 => x"ffa0050c",
  1700 => x"8c08ff8c",
  1701 => x"0508538c",
  1702 => x"08ff9c05",
  1703 => x"08525394",
  1704 => x"d63f8008",
  1705 => x"708c08ff",
  1706 => x"98050c8c",
  1707 => x"08ff9805",
  1708 => x"088c08ff",
  1709 => x"90050829",
  1710 => x"708c08ff",
  1711 => x"a4050c8c",
  1712 => x"08ffa005",
  1713 => x"0870902b",
  1714 => x"8c08ffbc",
  1715 => x"050883ff",
  1716 => x"ff067072",
  1717 => x"078c08ff",
  1718 => x"a0050c52",
  1719 => x"57515153",
  1720 => x"8c08ffa0",
  1721 => x"05088c08",
  1722 => x"ffa40508",
  1723 => x"2780de38",
  1724 => x"8c08ff98",
  1725 => x"0508ff05",
  1726 => x"8c08ff98",
  1727 => x"050c8c08",
  1728 => x"ffa00508",
  1729 => x"8c08c805",
  1730 => x"08058c08",
  1731 => x"ffa0050c",
  1732 => x"8c08c805",
  1733 => x"088c08ff",
  1734 => x"a0050826",
  1735 => x"b0388c08",
  1736 => x"ffa00508",
  1737 => x"8c08ffa4",
  1738 => x"050827a1",
  1739 => x"388c08ff",
  1740 => x"980508ff",
  1741 => x"058c08ff",
  1742 => x"98050c8c",
  1743 => x"08ffa005",
  1744 => x"088c08c8",
  1745 => x"0508058c",
  1746 => x"08ffa005",
  1747 => x"0c8c08ff",
  1748 => x"a005088c",
  1749 => x"08ffa405",
  1750 => x"08318c08",
  1751 => x"ffa0050c",
  1752 => x"8c08ff94",
  1753 => x"05087090",
  1754 => x"2b708c08",
  1755 => x"ff980508",
  1756 => x"078c08ff",
  1757 => x"b0050c8c",
  1758 => x"08ffa005",
  1759 => x"088c08ff",
  1760 => x"bc050c51",
  1761 => x"538c08c8",
  1762 => x"0508902a",
  1763 => x"8c08ff8c",
  1764 => x"050c8c08",
  1765 => x"c8050883",
  1766 => x"ffff068c",
  1767 => x"08ff9005",
  1768 => x"0c8c08ff",
  1769 => x"bc05088c",
  1770 => x"08ff8c05",
  1771 => x"08537052",
  1772 => x"5392e93f",
  1773 => x"8008708c",
  1774 => x"08ff9c05",
  1775 => x"0c8c08ff",
  1776 => x"8c050853",
  1777 => x"8c08ffbc",
  1778 => x"05085253",
  1779 => x"92a93f80",
  1780 => x"08708c08",
  1781 => x"ff94050c",
  1782 => x"8c08ff94",
  1783 => x"05088c08",
  1784 => x"ff900508",
  1785 => x"29708c08",
  1786 => x"ffa4050c",
  1787 => x"8c08ff9c",
  1788 => x"05087090",
  1789 => x"2b8c08c0",
  1790 => x"0508902a",
  1791 => x"7072078c",
  1792 => x"08ff9c05",
  1793 => x"0c525751",
  1794 => x"51538c08",
  1795 => x"ff9c0508",
  1796 => x"8c08ffa4",
  1797 => x"05082780",
  1798 => x"de388c08",
  1799 => x"ff940508",
  1800 => x"ff058c08",
  1801 => x"ff94050c",
  1802 => x"8c08ff9c",
  1803 => x"05088c08",
  1804 => x"c8050805",
  1805 => x"8c08ff9c",
  1806 => x"050c8c08",
  1807 => x"c805088c",
  1808 => x"08ff9c05",
  1809 => x"0826b038",
  1810 => x"8c08ff9c",
  1811 => x"05088c08",
  1812 => x"ffa40508",
  1813 => x"27a1388c",
  1814 => x"08ff9405",
  1815 => x"08ff058c",
  1816 => x"08ff9405",
  1817 => x"0c8c08ff",
  1818 => x"9c05088c",
  1819 => x"08c80508",
  1820 => x"058c08ff",
  1821 => x"9c050c8c",
  1822 => x"08ff9c05",
  1823 => x"088c08ff",
  1824 => x"a4050831",
  1825 => x"8c08ff9c",
  1826 => x"050c8c08",
  1827 => x"ff9c0508",
  1828 => x"8c08ff8c",
  1829 => x"05085370",
  1830 => x"52539180",
  1831 => x"3f800870",
  1832 => x"8c08ffa0",
  1833 => x"050c8c08",
  1834 => x"ff8c0508",
  1835 => x"538c08ff",
  1836 => x"9c050852",
  1837 => x"5390c03f",
  1838 => x"8008708c",
  1839 => x"08ff9805",
  1840 => x"0c8c08ff",
  1841 => x"9805088c",
  1842 => x"08ff9005",
  1843 => x"0829708c",
  1844 => x"08ffa405",
  1845 => x"0c8c08ff",
  1846 => x"a0050870",
  1847 => x"902b8c08",
  1848 => x"c0050883",
  1849 => x"ffff0670",
  1850 => x"72078c08",
  1851 => x"ffa0050c",
  1852 => x"52575151",
  1853 => x"538c08ff",
  1854 => x"a005088c",
  1855 => x"08ffa405",
  1856 => x"082780de",
  1857 => x"388c08ff",
  1858 => x"980508ff",
  1859 => x"058c08ff",
  1860 => x"98050c8c",
  1861 => x"08ffa005",
  1862 => x"088c08c8",
  1863 => x"0508058c",
  1864 => x"08ffa005",
  1865 => x"0c8c08c8",
  1866 => x"05088c08",
  1867 => x"ffa00508",
  1868 => x"26b0388c",
  1869 => x"08ffa005",
  1870 => x"088c08ff",
  1871 => x"a4050827",
  1872 => x"a1388c08",
  1873 => x"ff980508",
  1874 => x"ff058c08",
  1875 => x"ff98050c",
  1876 => x"8c08ffa0",
  1877 => x"05088c08",
  1878 => x"c8050805",
  1879 => x"8c08ffa0",
  1880 => x"050c8c08",
  1881 => x"ffa00508",
  1882 => x"8c08ffa4",
  1883 => x"0508318c",
  1884 => x"08ffa005",
  1885 => x"0c8c08ff",
  1886 => x"94050870",
  1887 => x"902b708c",
  1888 => x"08ff9805",
  1889 => x"08078c08",
  1890 => x"ffb4050c",
  1891 => x"8c08ffa0",
  1892 => x"05088c08",
  1893 => x"c0050c51",
  1894 => x"538c08ec",
  1895 => x"0508802e",
  1896 => x"8ded388c",
  1897 => x"08c00508",
  1898 => x"8c08ffa8",
  1899 => x"05082a8c",
  1900 => x"08d0050c",
  1901 => x"800b8c08",
  1902 => x"cc050c8c",
  1903 => x"08ec0508",
  1904 => x"558c08cc",
  1905 => x"05088c08",
  1906 => x"d0050855",
  1907 => x"5372750c",
  1908 => x"7384160c",
  1909 => x"8db9398c",
  1910 => x"08ffbc05",
  1911 => x"088c08c4",
  1912 => x"05082780",
  1913 => x"cc38800b",
  1914 => x"8c08ffb4",
  1915 => x"050c800b",
  1916 => x"8c08ffb0",
  1917 => x"050c8c08",
  1918 => x"ec050880",
  1919 => x"2e8d9038",
  1920 => x"8c08c005",
  1921 => x"088c08d0",
  1922 => x"050c8c08",
  1923 => x"ffbc0508",
  1924 => x"8c08cc05",
  1925 => x"0c8c08ec",
  1926 => x"0508558c",
  1927 => x"08cc0508",
  1928 => x"8c08d005",
  1929 => x"08555372",
  1930 => x"750c7384",
  1931 => x"160c8cdf",
  1932 => x"398c08c4",
  1933 => x"05088c08",
  1934 => x"ff8c050c",
  1935 => x"8c08ff8c",
  1936 => x"050883ff",
  1937 => x"ff26a038",
  1938 => x"8c08ff8c",
  1939 => x"050881ff",
  1940 => x"268b3880",
  1941 => x"0b8c08fe",
  1942 => x"ec050ca9",
  1943 => x"39880b8c",
  1944 => x"08feec05",
  1945 => x"0c9f398c",
  1946 => x"08ff8c05",
  1947 => x"08fe800a",
  1948 => x"268b3890",
  1949 => x"0b8c08fe",
  1950 => x"ec050c89",
  1951 => x"39980b8c",
  1952 => x"08feec05",
  1953 => x"0c8c08fe",
  1954 => x"ec05088c",
  1955 => x"08ff9005",
  1956 => x"0c8c08ff",
  1957 => x"8c05088c",
  1958 => x"08ff9005",
  1959 => x"082a80d4",
  1960 => x"d011338c",
  1961 => x"08ff9005",
  1962 => x"0811a071",
  1963 => x"318c08ff",
  1964 => x"a8050c51",
  1965 => x"51538c08",
  1966 => x"ffa80508",
  1967 => x"81cc388c",
  1968 => x"08ffbc05",
  1969 => x"088c08c4",
  1970 => x"05082691",
  1971 => x"388c08c0",
  1972 => x"05088c08",
  1973 => x"c8050827",
  1974 => x"843880e3",
  1975 => x"39810b8c",
  1976 => x"08ffb405",
  1977 => x"0c8c08c0",
  1978 => x"05088c08",
  1979 => x"c8050831",
  1980 => x"8c08ff8c",
  1981 => x"050c8c08",
  1982 => x"ffbc0508",
  1983 => x"8c08c405",
  1984 => x"0831708c",
  1985 => x"08fee805",
  1986 => x"0c538c08",
  1987 => x"c005088c",
  1988 => x"08ff8c05",
  1989 => x"08278f38",
  1990 => x"8c08fee8",
  1991 => x"0508ff05",
  1992 => x"8c08fee8",
  1993 => x"050c8c08",
  1994 => x"fee80508",
  1995 => x"8c08ffbc",
  1996 => x"050c8c08",
  1997 => x"ff8c0508",
  1998 => x"8c08c005",
  1999 => x"0c893980",
  2000 => x"0b8c08ff",
  2001 => x"b4050c80",
  2002 => x"0b8c08ff",
  2003 => x"b0050c8c",
  2004 => x"08ec0508",
  2005 => x"802e8ab7",
  2006 => x"388c08c0",
  2007 => x"05088c08",
  2008 => x"d0050c8c",
  2009 => x"08ffbc05",
  2010 => x"088c08cc",
  2011 => x"050c8c08",
  2012 => x"ec050855",
  2013 => x"8c08cc05",
  2014 => x"088c08d0",
  2015 => x"05085553",
  2016 => x"72750c73",
  2017 => x"84160c8a",
  2018 => x"8639a00b",
  2019 => x"8c08ffa8",
  2020 => x"0508318c",
  2021 => x"08ffac05",
  2022 => x"0c8c08c4",
  2023 => x"05088c08",
  2024 => x"ffa80508",
  2025 => x"2b8c08c8",
  2026 => x"05088c08",
  2027 => x"ffac0508",
  2028 => x"2a707207",
  2029 => x"8c08c405",
  2030 => x"0c8c08c8",
  2031 => x"05088c08",
  2032 => x"ffa80508",
  2033 => x"2b8c08c8",
  2034 => x"050c8c08",
  2035 => x"ffbc0508",
  2036 => x"8c08ffac",
  2037 => x"05082a8c",
  2038 => x"08ffb805",
  2039 => x"0c8c08ff",
  2040 => x"bc05088c",
  2041 => x"08ffa805",
  2042 => x"082b8c08",
  2043 => x"c005088c",
  2044 => x"08ffac05",
  2045 => x"082a7072",
  2046 => x"078c08ff",
  2047 => x"bc050c8c",
  2048 => x"08c00508",
  2049 => x"8c08ffa8",
  2050 => x"05082b8c",
  2051 => x"08c0050c",
  2052 => x"8c08c405",
  2053 => x"08902a8c",
  2054 => x"08ff9405",
  2055 => x"0c8c08c4",
  2056 => x"050883ff",
  2057 => x"ff068c08",
  2058 => x"ff98050c",
  2059 => x"8c08ffb8",
  2060 => x"05088c08",
  2061 => x"ff940508",
  2062 => x"57705651",
  2063 => x"52525454",
  2064 => x"89da3f80",
  2065 => x"08708c08",
  2066 => x"ffa4050c",
  2067 => x"8c08ff94",
  2068 => x"0508538c",
  2069 => x"08ffb805",
  2070 => x"08525389",
  2071 => x"9a3f8008",
  2072 => x"708c08ff",
  2073 => x"9c050c8c",
  2074 => x"08ff9c05",
  2075 => x"088c08ff",
  2076 => x"98050829",
  2077 => x"708c08ff",
  2078 => x"84050c8c",
  2079 => x"08ffa405",
  2080 => x"0870902b",
  2081 => x"8c08ffbc",
  2082 => x"0508902a",
  2083 => x"7072078c",
  2084 => x"08ffa405",
  2085 => x"0c525751",
  2086 => x"51538c08",
  2087 => x"ffa40508",
  2088 => x"8c08ff84",
  2089 => x"05082780",
  2090 => x"de388c08",
  2091 => x"ff9c0508",
  2092 => x"ff058c08",
  2093 => x"ff9c050c",
  2094 => x"8c08ffa4",
  2095 => x"05088c08",
  2096 => x"c4050805",
  2097 => x"8c08ffa4",
  2098 => x"050c8c08",
  2099 => x"c405088c",
  2100 => x"08ffa405",
  2101 => x"0826b038",
  2102 => x"8c08ffa4",
  2103 => x"05088c08",
  2104 => x"ff840508",
  2105 => x"27a1388c",
  2106 => x"08ff9c05",
  2107 => x"08ff058c",
  2108 => x"08ff9c05",
  2109 => x"0c8c08ff",
  2110 => x"a405088c",
  2111 => x"08c40508",
  2112 => x"058c08ff",
  2113 => x"a4050c8c",
  2114 => x"08ffa405",
  2115 => x"088c08ff",
  2116 => x"84050831",
  2117 => x"8c08ffa4",
  2118 => x"050c8c08",
  2119 => x"ffa40508",
  2120 => x"8c08ff94",
  2121 => x"05085370",
  2122 => x"525387f0",
  2123 => x"3f800870",
  2124 => x"8c08ff88",
  2125 => x"050c8c08",
  2126 => x"ff940508",
  2127 => x"538c08ff",
  2128 => x"a4050852",
  2129 => x"5387b03f",
  2130 => x"8008708c",
  2131 => x"08ffa005",
  2132 => x"0c8c08ff",
  2133 => x"a005088c",
  2134 => x"08ff9805",
  2135 => x"0829708c",
  2136 => x"08ff8405",
  2137 => x"0c8c08ff",
  2138 => x"88050870",
  2139 => x"902b8c08",
  2140 => x"ffbc0508",
  2141 => x"83ffff06",
  2142 => x"7072078c",
  2143 => x"08ff8805",
  2144 => x"0c525751",
  2145 => x"51538c08",
  2146 => x"ff880508",
  2147 => x"8c08ff84",
  2148 => x"05082780",
  2149 => x"de388c08",
  2150 => x"ffa00508",
  2151 => x"ff058c08",
  2152 => x"ffa0050c",
  2153 => x"8c08ff88",
  2154 => x"05088c08",
  2155 => x"c4050805",
  2156 => x"8c08ff88",
  2157 => x"050c8c08",
  2158 => x"c405088c",
  2159 => x"08ff8805",
  2160 => x"0826b038",
  2161 => x"8c08ff88",
  2162 => x"05088c08",
  2163 => x"ff840508",
  2164 => x"27a1388c",
  2165 => x"08ffa005",
  2166 => x"08ff058c",
  2167 => x"08ffa005",
  2168 => x"0c8c08ff",
  2169 => x"8805088c",
  2170 => x"08c40508",
  2171 => x"058c08ff",
  2172 => x"88050c8c",
  2173 => x"08ff8805",
  2174 => x"088c08ff",
  2175 => x"84050831",
  2176 => x"8c08ff88",
  2177 => x"050c8c08",
  2178 => x"ff9c0508",
  2179 => x"70902b70",
  2180 => x"8c08ffa0",
  2181 => x"0508078c",
  2182 => x"08ffb405",
  2183 => x"0c8c08ff",
  2184 => x"8805088c",
  2185 => x"08ffbc05",
  2186 => x"0c8c08ff",
  2187 => x"b4050883",
  2188 => x"ffff068c",
  2189 => x"08ff9c05",
  2190 => x"0c8c08ff",
  2191 => x"b4050890",
  2192 => x"2a8c08ff",
  2193 => x"a4050c8c",
  2194 => x"08c80508",
  2195 => x"83ffff06",
  2196 => x"8c08ffa0",
  2197 => x"050c8c08",
  2198 => x"c8050890",
  2199 => x"2a8c08ff",
  2200 => x"80050c8c",
  2201 => x"08ff9c05",
  2202 => x"088c08ff",
  2203 => x"a0050829",
  2204 => x"708c08ff",
  2205 => x"84050c8c",
  2206 => x"08ff9c05",
  2207 => x"088c08ff",
  2208 => x"80050829",
  2209 => x"708c08ff",
  2210 => x"88050c8c",
  2211 => x"08ffa405",
  2212 => x"088c08ff",
  2213 => x"a0050829",
  2214 => x"708c08ff",
  2215 => x"94050c8c",
  2216 => x"08ffa405",
  2217 => x"088c08ff",
  2218 => x"80050829",
  2219 => x"708c08ff",
  2220 => x"98050c8c",
  2221 => x"08ff8405",
  2222 => x"08902a8c",
  2223 => x"08ff8805",
  2224 => x"08118c08",
  2225 => x"ff88050c",
  2226 => x"8c08ff88",
  2227 => x"05088c08",
  2228 => x"ff940508",
  2229 => x"058c08ff",
  2230 => x"88050c51",
  2231 => x"51515151",
  2232 => x"51538c08",
  2233 => x"ff880508",
  2234 => x"8c08ff94",
  2235 => x"05082791",
  2236 => x"388c08ff",
  2237 => x"98050884",
  2238 => x"8080058c",
  2239 => x"08ff9805",
  2240 => x"0c8c08ff",
  2241 => x"88050890",
  2242 => x"2a8c08ff",
  2243 => x"98050811",
  2244 => x"8c08ff8c",
  2245 => x"050c8c08",
  2246 => x"ff880508",
  2247 => x"83ffff06",
  2248 => x"70902b8c",
  2249 => x"08ff8405",
  2250 => x"0883ffff",
  2251 => x"0670128c",
  2252 => x"08ff9005",
  2253 => x"0c525651",
  2254 => x"538c08ff",
  2255 => x"8c05088c",
  2256 => x"08ffbc05",
  2257 => x"0826a538",
  2258 => x"8c08ff8c",
  2259 => x"05088c08",
  2260 => x"ffbc0508",
  2261 => x"2e098106",
  2262 => x"80fb388c",
  2263 => x"08ff9005",
  2264 => x"088c08c0",
  2265 => x"05082684",
  2266 => x"3880ea39",
  2267 => x"8c08ffb4",
  2268 => x"0508ff05",
  2269 => x"8c08ffb4",
  2270 => x"050c8c08",
  2271 => x"ff900508",
  2272 => x"8c08c805",
  2273 => x"08318c08",
  2274 => x"ff80050c",
  2275 => x"8c08ff8c",
  2276 => x"05088c08",
  2277 => x"c4050831",
  2278 => x"708c08fe",
  2279 => x"e4050c53",
  2280 => x"8c08ff90",
  2281 => x"05088c08",
  2282 => x"ff800508",
  2283 => x"278f388c",
  2284 => x"08fee405",
  2285 => x"08ff058c",
  2286 => x"08fee405",
  2287 => x"0c8c08fe",
  2288 => x"e405088c",
  2289 => x"08ff8c05",
  2290 => x"0c8c08ff",
  2291 => x"8005088c",
  2292 => x"08ff9005",
  2293 => x"0c800b8c",
  2294 => x"08ffb005",
  2295 => x"0c8c08ec",
  2296 => x"0508802e",
  2297 => x"81a9388c",
  2298 => x"08c00508",
  2299 => x"8c08ff90",
  2300 => x"0508318c",
  2301 => x"08ff8005",
  2302 => x"0c8c08ff",
  2303 => x"bc05088c",
  2304 => x"08ff8c05",
  2305 => x"0831708c",
  2306 => x"08fee005",
  2307 => x"0c538c08",
  2308 => x"c005088c",
  2309 => x"08ff8005",
  2310 => x"08278f38",
  2311 => x"8c08fee0",
  2312 => x"0508ff05",
  2313 => x"8c08fee0",
  2314 => x"050c8c08",
  2315 => x"fee00508",
  2316 => x"8c08ffbc",
  2317 => x"050c8c08",
  2318 => x"ff800508",
  2319 => x"8c08c005",
  2320 => x"0c8c08ff",
  2321 => x"bc05088c",
  2322 => x"08ffac05",
  2323 => x"082b8c08",
  2324 => x"c005088c",
  2325 => x"08ffa805",
  2326 => x"082a7072",
  2327 => x"078c08d0",
  2328 => x"050c8c08",
  2329 => x"ffbc0508",
  2330 => x"8c08ffa8",
  2331 => x"05082a8c",
  2332 => x"08cc050c",
  2333 => x"8c08ec05",
  2334 => x"08575454",
  2335 => x"8c08cc05",
  2336 => x"088c08d0",
  2337 => x"05085553",
  2338 => x"72750c73",
  2339 => x"84160c80",
  2340 => x"0b8c08fe",
  2341 => x"f8050c80",
  2342 => x"0b8c08fe",
  2343 => x"fc050c8c",
  2344 => x"08ffb005",
  2345 => x"088c08fe",
  2346 => x"f8050c8c",
  2347 => x"08ffb405",
  2348 => x"088c08fe",
  2349 => x"fc050c8c",
  2350 => x"08fef805",
  2351 => x"088c08fe",
  2352 => x"fc050855",
  2353 => x"53728c08",
  2354 => x"e4050c73",
  2355 => x"8c08e805",
  2356 => x"0c8c08e4",
  2357 => x"05088c08",
  2358 => x"e805088c",
  2359 => x"08880508",
  2360 => x"57555372",
  2361 => x"750c7384",
  2362 => x"160c8c08",
  2363 => x"88050880",
  2364 => x"0cae3d0d",
  2365 => x"8c0c048c",
  2366 => x"08028c0c",
  2367 => x"fd3d0d80",
  2368 => x"538c088c",
  2369 => x"0508528c",
  2370 => x"08880508",
  2371 => x"5182de3f",
  2372 => x"80087080",
  2373 => x"0c54853d",
  2374 => x"0d8c0c04",
  2375 => x"8c08028c",
  2376 => x"0cfd3d0d",
  2377 => x"81538c08",
  2378 => x"8c050852",
  2379 => x"8c088805",
  2380 => x"085182b9",
  2381 => x"3f800870",
  2382 => x"800c5485",
  2383 => x"3d0d8c0c",
  2384 => x"048c0802",
  2385 => x"8c0cf93d",
  2386 => x"0d800b8c",
  2387 => x"08fc050c",
  2388 => x"8c088805",
  2389 => x"088025ab",
  2390 => x"388c0888",
  2391 => x"0508308c",
  2392 => x"0888050c",
  2393 => x"800b8c08",
  2394 => x"f4050c8c",
  2395 => x"08fc0508",
  2396 => x"8838810b",
  2397 => x"8c08f405",
  2398 => x"0c8c08f4",
  2399 => x"05088c08",
  2400 => x"fc050c8c",
  2401 => x"088c0508",
  2402 => x"8025ab38",
  2403 => x"8c088c05",
  2404 => x"08308c08",
  2405 => x"8c050c80",
  2406 => x"0b8c08f0",
  2407 => x"050c8c08",
  2408 => x"fc050888",
  2409 => x"38810b8c",
  2410 => x"08f0050c",
  2411 => x"8c08f005",
  2412 => x"088c08fc",
  2413 => x"050c8053",
  2414 => x"8c088c05",
  2415 => x"08528c08",
  2416 => x"88050851",
  2417 => x"81a73f80",
  2418 => x"08708c08",
  2419 => x"f8050c54",
  2420 => x"8c08fc05",
  2421 => x"08802e8c",
  2422 => x"388c08f8",
  2423 => x"0508308c",
  2424 => x"08f8050c",
  2425 => x"8c08f805",
  2426 => x"0870800c",
  2427 => x"54893d0d",
  2428 => x"8c0c048c",
  2429 => x"08028c0c",
  2430 => x"fb3d0d80",
  2431 => x"0b8c08fc",
  2432 => x"050c8c08",
  2433 => x"88050880",
  2434 => x"2593388c",
  2435 => x"08880508",
  2436 => x"308c0888",
  2437 => x"050c810b",
  2438 => x"8c08fc05",
  2439 => x"0c8c088c",
  2440 => x"05088025",
  2441 => x"8c388c08",
  2442 => x"8c050830",
  2443 => x"8c088c05",
  2444 => x"0c81538c",
  2445 => x"088c0508",
  2446 => x"528c0888",
  2447 => x"050851ad",
  2448 => x"3f800870",
  2449 => x"8c08f805",
  2450 => x"0c548c08",
  2451 => x"fc050880",
  2452 => x"2e8c388c",
  2453 => x"08f80508",
  2454 => x"308c08f8",
  2455 => x"050c8c08",
  2456 => x"f8050870",
  2457 => x"800c5487",
  2458 => x"3d0d8c0c",
  2459 => x"048c0802",
  2460 => x"8c0cfd3d",
  2461 => x"0d810b8c",
  2462 => x"08fc050c",
  2463 => x"800b8c08",
  2464 => x"f8050c8c",
  2465 => x"088c0508",
  2466 => x"8c088805",
  2467 => x"0827ac38",
  2468 => x"8c08fc05",
  2469 => x"08802ea3",
  2470 => x"38800b8c",
  2471 => x"088c0508",
  2472 => x"2499388c",
  2473 => x"088c0508",
  2474 => x"108c088c",
  2475 => x"050c8c08",
  2476 => x"fc050810",
  2477 => x"8c08fc05",
  2478 => x"0cc9398c",
  2479 => x"08fc0508",
  2480 => x"802e80c9",
  2481 => x"388c088c",
  2482 => x"05088c08",
  2483 => x"88050826",
  2484 => x"a1388c08",
  2485 => x"8805088c",
  2486 => x"088c0508",
  2487 => x"318c0888",
  2488 => x"050c8c08",
  2489 => x"f805088c",
  2490 => x"08fc0508",
  2491 => x"078c08f8",
  2492 => x"050c8c08",
  2493 => x"fc050881",
  2494 => x"2a8c08fc",
  2495 => x"050c8c08",
  2496 => x"8c050881",
  2497 => x"2a8c088c",
  2498 => x"050cffaf",
  2499 => x"398c0890",
  2500 => x"0508802e",
  2501 => x"8f388c08",
  2502 => x"88050870",
  2503 => x"8c08f405",
  2504 => x"0c518d39",
  2505 => x"8c08f805",
  2506 => x"08708c08",
  2507 => x"f4050c51",
  2508 => x"8c08f405",
  2509 => x"08800c85",
  2510 => x"3d0d8c0c",
  2511 => x"04fc3d0d",
  2512 => x"7670797b",
  2513 => x"55555555",
  2514 => x"8f72278c",
  2515 => x"38727507",
  2516 => x"83065170",
  2517 => x"802ea738",
  2518 => x"ff125271",
  2519 => x"ff2e9838",
  2520 => x"72708105",
  2521 => x"54337470",
  2522 => x"81055634",
  2523 => x"ff125271",
  2524 => x"ff2e0981",
  2525 => x"06ea3874",
  2526 => x"800c863d",
  2527 => x"0d047451",
  2528 => x"72708405",
  2529 => x"54087170",
  2530 => x"8405530c",
  2531 => x"72708405",
  2532 => x"54087170",
  2533 => x"8405530c",
  2534 => x"72708405",
  2535 => x"54087170",
  2536 => x"8405530c",
  2537 => x"72708405",
  2538 => x"54087170",
  2539 => x"8405530c",
  2540 => x"f0125271",
  2541 => x"8f26c938",
  2542 => x"83722795",
  2543 => x"38727084",
  2544 => x"05540871",
  2545 => x"70840553",
  2546 => x"0cfc1252",
  2547 => x"718326ed",
  2548 => x"387054ff",
  2549 => x"8339fd3d",
  2550 => x"0d800b80",
  2551 => x"d6f40854",
  2552 => x"5472812e",
  2553 => x"9c387380",
  2554 => x"def80cff",
  2555 => x"b8f23fff",
  2556 => x"b88e3f80",
  2557 => x"d7945281",
  2558 => x"51c4de3f",
  2559 => x"800851a2",
  2560 => x"3f7280de",
  2561 => x"f80cffb8",
  2562 => x"d73fffb7",
  2563 => x"f33f80d7",
  2564 => x"94528151",
  2565 => x"c4c33f80",
  2566 => x"0851873f",
  2567 => x"00ff3900",
  2568 => x"ff39f73d",
  2569 => x"0d7b80d7",
  2570 => x"980882c8",
  2571 => x"11085a54",
  2572 => x"5a77802e",
  2573 => x"80da3881",
  2574 => x"88188419",
  2575 => x"08ff0581",
  2576 => x"712b5955",
  2577 => x"59807424",
  2578 => x"80ea3880",
  2579 => x"7424b538",
  2580 => x"73822b78",
  2581 => x"11880556",
  2582 => x"56818019",
  2583 => x"08770653",
  2584 => x"72802eb6",
  2585 => x"38781670",
  2586 => x"08535379",
  2587 => x"51740853",
  2588 => x"722dff14",
  2589 => x"fc17fc17",
  2590 => x"79812c5a",
  2591 => x"57575473",
  2592 => x"8025d638",
  2593 => x"77085877",
  2594 => x"ffad3880",
  2595 => x"d7980853",
  2596 => x"bc1308a5",
  2597 => x"387951ff",
  2598 => x"833f7408",
  2599 => x"53722dff",
  2600 => x"14fc17fc",
  2601 => x"1779812c",
  2602 => x"5a575754",
  2603 => x"738025ff",
  2604 => x"a838d139",
  2605 => x"8057ff93",
  2606 => x"397251bc",
  2607 => x"13085372",
  2608 => x"2d7951fe",
  2609 => x"d73fff3d",
  2610 => x"0d80de9c",
  2611 => x"0bfc0570",
  2612 => x"08525270",
  2613 => x"ff2e9138",
  2614 => x"702dfc12",
  2615 => x"70085252",
  2616 => x"70ff2e09",
  2617 => x"8106f138",
  2618 => x"833d0d04",
  2619 => x"04ffb7dd",
  2620 => x"3f040000",
  2621 => x"00000040",
  2622 => x"4175746f",
  2623 => x"2d6e6567",
  2624 => x"6f746961",
  2625 => x"74696f6e",
  2626 => x"20666169",
  2627 => x"6c65640a",
  2628 => x"00000000",
  2629 => x"47524554",
  2630 => x"48280000",
  2631 => x"31302f31",
  2632 => x"30302f31",
  2633 => x"30303000",
  2634 => x"29204574",
  2635 => x"6865726e",
  2636 => x"6574204d",
  2637 => x"41432061",
  2638 => x"74205b30",
  2639 => x"78000000",
  2640 => x"5d2e2052",
  2641 => x"756e6e69",
  2642 => x"6e672000",
  2643 => x"31303000",
  2644 => x"204d6270",
  2645 => x"73200000",
  2646 => x"66756c6c",
  2647 => x"00000000",
  2648 => x"20647570",
  2649 => x"6c65780a",
  2650 => x"00000000",
  2651 => x"31302f31",
  2652 => x"30300000",
  2653 => x"31300000",
  2654 => x"68616c66",
  2655 => x"00000000",
  2656 => x"0c677265",
  2657 => x"74682e63",
  2658 => x"00000000",
  2659 => x"20286f6e",
  2660 => x"2073696d",
  2661 => x"290a0000",
  2662 => x"0a53656e",
  2663 => x"64696e67",
  2664 => x"20313530",
  2665 => x"30204d62",
  2666 => x"79746520",
  2667 => x"6f662064",
  2668 => x"61746120",
  2669 => x"746f2000",
  2670 => x"20706163",
  2671 => x"6b657473",
  2672 => x"290a0a00",
  2673 => x"54696d65",
  2674 => x"20202020",
  2675 => x"3a200000",
  2676 => x"20736563",
  2677 => x"0a000000",
  2678 => x"42697472",
  2679 => x"61746520",
  2680 => x"3a200000",
  2681 => x"206b6270",
  2682 => x"730a0000",
  2683 => x"20286f6e",
  2684 => x"20686172",
  2685 => x"64776172",
  2686 => x"65290a00",
  2687 => x"636f6d70",
  2688 => x"696c6564",
  2689 => x"3a204a61",
  2690 => x"6e202037",
  2691 => x"20323031",
  2692 => x"31202031",
  2693 => x"343a3430",
  2694 => x"3a34360a",
  2695 => x"00000000",
  2696 => x"30622020",
  2697 => x"20202020",
  2698 => x"20202020",
  2699 => x"20202020",
  2700 => x"20202020",
  2701 => x"20202020",
  2702 => x"20202020",
  2703 => x"20202020",
  2704 => x"20200000",
  2705 => x"20202020",
  2706 => x"20202020",
  2707 => x"00000000",
  2708 => x"00010202",
  2709 => x"03030303",
  2710 => x"04040404",
  2711 => x"04040404",
  2712 => x"05050505",
  2713 => x"05050505",
  2714 => x"05050505",
  2715 => x"05050505",
  2716 => x"06060606",
  2717 => x"06060606",
  2718 => x"06060606",
  2719 => x"06060606",
  2720 => x"06060606",
  2721 => x"06060606",
  2722 => x"06060606",
  2723 => x"06060606",
  2724 => x"07070707",
  2725 => x"07070707",
  2726 => x"07070707",
  2727 => x"07070707",
  2728 => x"07070707",
  2729 => x"07070707",
  2730 => x"07070707",
  2731 => x"07070707",
  2732 => x"07070707",
  2733 => x"07070707",
  2734 => x"07070707",
  2735 => x"07070707",
  2736 => x"07070707",
  2737 => x"07070707",
  2738 => x"07070707",
  2739 => x"07070707",
  2740 => x"08080808",
  2741 => x"08080808",
  2742 => x"08080808",
  2743 => x"08080808",
  2744 => x"08080808",
  2745 => x"08080808",
  2746 => x"08080808",
  2747 => x"08080808",
  2748 => x"08080808",
  2749 => x"08080808",
  2750 => x"08080808",
  2751 => x"08080808",
  2752 => x"08080808",
  2753 => x"08080808",
  2754 => x"08080808",
  2755 => x"08080808",
  2756 => x"08080808",
  2757 => x"08080808",
  2758 => x"08080808",
  2759 => x"08080808",
  2760 => x"08080808",
  2761 => x"08080808",
  2762 => x"08080808",
  2763 => x"08080808",
  2764 => x"08080808",
  2765 => x"08080808",
  2766 => x"08080808",
  2767 => x"08080808",
  2768 => x"08080808",
  2769 => x"08080808",
  2770 => x"08080808",
  2771 => x"08080808",
  2772 => x"64756d6d",
  2773 => x"792e6578",
  2774 => x"65000000",
  2775 => x"43000000",
  2776 => x"00ffffff",
  2777 => x"ff00ffff",
  2778 => x"ffff00ff",
  2779 => x"ffffff00",
  2780 => x"00000000",
  2781 => x"00000000",
  2782 => x"00000000",
  2783 => x"00002f24",
  2784 => x"80000d00",
  2785 => x"80000800",
  2786 => x"80000600",
  2787 => x"80000200",
  2788 => x"80000100",
  2789 => x"00002b50",
  2790 => x"00002b9c",
  2791 => x"00000000",
  2792 => x"00002e04",
  2793 => x"00002e60",
  2794 => x"00002ebc",
  2795 => x"00000000",
  2796 => x"00000000",
  2797 => x"00000000",
  2798 => x"00000000",
  2799 => x"00000000",
  2800 => x"00000000",
  2801 => x"00000000",
  2802 => x"00000000",
  2803 => x"00000000",
  2804 => x"00002b5c",
  2805 => x"00000000",
  2806 => x"00000000",
  2807 => x"00000000",
  2808 => x"00000000",
  2809 => x"00000000",
  2810 => x"00000000",
  2811 => x"00000000",
  2812 => x"00000000",
  2813 => x"00000000",
  2814 => x"00000000",
  2815 => x"00000000",
  2816 => x"00000000",
  2817 => x"00000000",
  2818 => x"00000000",
  2819 => x"00000000",
  2820 => x"00000000",
  2821 => x"00000000",
  2822 => x"00000000",
  2823 => x"00000000",
  2824 => x"00000000",
  2825 => x"00000000",
  2826 => x"00000000",
  2827 => x"00000000",
  2828 => x"00000000",
  2829 => x"00000000",
  2830 => x"00000000",
  2831 => x"00000000",
  2832 => x"00000000",
  2833 => x"00000001",
  2834 => x"330eabcd",
  2835 => x"1234e66d",
  2836 => x"deec0005",
  2837 => x"000b0000",
  2838 => x"00000000",
  2839 => x"00000000",
  2840 => x"00000000",
  2841 => x"00000000",
  2842 => x"00000000",
  2843 => x"00000000",
  2844 => x"00000000",
  2845 => x"00000000",
  2846 => x"00000000",
  2847 => x"00000000",
  2848 => x"00000000",
  2849 => x"00000000",
  2850 => x"00000000",
  2851 => x"00000000",
  2852 => x"00000000",
  2853 => x"00000000",
  2854 => x"00000000",
  2855 => x"00000000",
  2856 => x"00000000",
  2857 => x"00000000",
  2858 => x"00000000",
  2859 => x"00000000",
  2860 => x"00000000",
  2861 => x"00000000",
  2862 => x"00000000",
  2863 => x"00000000",
  2864 => x"00000000",
  2865 => x"00000000",
  2866 => x"00000000",
  2867 => x"00000000",
  2868 => x"00000000",
  2869 => x"00000000",
  2870 => x"00000000",
  2871 => x"00000000",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000000",
  2884 => x"00000000",
  2885 => x"00000000",
  2886 => x"00000000",
  2887 => x"00000000",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000000",
  2895 => x"00000000",
  2896 => x"00000000",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000000",
  2900 => x"00000000",
  2901 => x"00000000",
  2902 => x"00000000",
  2903 => x"00000000",
  2904 => x"00000000",
  2905 => x"00000000",
  2906 => x"00000000",
  2907 => x"00000000",
  2908 => x"00000000",
  2909 => x"00000000",
  2910 => x"00000000",
  2911 => x"00000000",
  2912 => x"00000000",
  2913 => x"00000000",
  2914 => x"00000000",
  2915 => x"00000000",
  2916 => x"00000000",
  2917 => x"00000000",
  2918 => x"00000000",
  2919 => x"00000000",
  2920 => x"00000000",
  2921 => x"00000000",
  2922 => x"00000000",
  2923 => x"00000000",
  2924 => x"00000000",
  2925 => x"00000000",
  2926 => x"00000000",
  2927 => x"00000000",
  2928 => x"00000000",
  2929 => x"00000000",
  2930 => x"00000000",
  2931 => x"00000000",
  2932 => x"00000000",
  2933 => x"00000000",
  2934 => x"00000000",
  2935 => x"00000000",
  2936 => x"00000000",
  2937 => x"00000000",
  2938 => x"00000000",
  2939 => x"00000000",
  2940 => x"00000000",
  2941 => x"00000000",
  2942 => x"00000000",
  2943 => x"00000000",
  2944 => x"00000000",
  2945 => x"00000000",
  2946 => x"00000000",
  2947 => x"00000000",
  2948 => x"00000000",
  2949 => x"00000000",
  2950 => x"00000000",
  2951 => x"00000000",
  2952 => x"00000000",
  2953 => x"00000000",
  2954 => x"00000000",
  2955 => x"00000000",
  2956 => x"00000000",
  2957 => x"00000000",
  2958 => x"00000000",
  2959 => x"00000000",
  2960 => x"00000000",
  2961 => x"00000000",
  2962 => x"00000000",
  2963 => x"00000000",
  2964 => x"00000000",
  2965 => x"00000000",
  2966 => x"00000000",
  2967 => x"00000000",
  2968 => x"00000000",
  2969 => x"00000000",
  2970 => x"00000000",
  2971 => x"00000000",
  2972 => x"00000000",
  2973 => x"00000000",
  2974 => x"00000000",
  2975 => x"00000000",
  2976 => x"00000000",
  2977 => x"00000000",
  2978 => x"00000000",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00000000",
  2983 => x"00000000",
  2984 => x"00000000",
  2985 => x"00000000",
  2986 => x"00000000",
  2987 => x"00000000",
  2988 => x"00000000",
  2989 => x"00000000",
  2990 => x"00000000",
  2991 => x"00000000",
  2992 => x"00000000",
  2993 => x"00000000",
  2994 => x"00000000",
  2995 => x"00000000",
  2996 => x"00000000",
  2997 => x"00000000",
  2998 => x"00000000",
  2999 => x"00000000",
  3000 => x"00000000",
  3001 => x"00000000",
  3002 => x"00000000",
  3003 => x"00000000",
  3004 => x"00000000",
  3005 => x"00000000",
  3006 => x"00000000",
  3007 => x"00000000",
  3008 => x"00000000",
  3009 => x"00000000",
  3010 => x"00000000",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"ffffffff",
  3015 => x"00000000",
  3016 => x"ffffffff",
  3017 => x"00000000",
  3018 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
