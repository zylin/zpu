
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 15;
constant bytes : integer := 17892;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B0BBA";
    when 16#00001# => romdata <= X"C5040000";
    when 16#00002# => romdata <= X"00000000";
    when 16#00003# => romdata <= X"00000000";
    when 16#00004# => romdata <= X"00000000";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"0B0B0BBD";
    when 16#00009# => romdata <= X"AA040000";
    when 16#0000A# => romdata <= X"00000000";
    when 16#0000B# => romdata <= X"00000000";
    when 16#0000C# => romdata <= X"00000000";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B0BBC";
    when 16#00049# => romdata <= X"DE040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B0BBCC1";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B80FB";
    when 16#000A2# => romdata <= X"F0738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B0B";
    when 16#000A5# => romdata <= X"BCC40400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"0B0B0BBD";
    when 16#000A9# => romdata <= X"92040000";
    when 16#000AA# => romdata <= X"00000000";
    when 16#000AB# => romdata <= X"00000000";
    when 16#000AC# => romdata <= X"00000000";
    when 16#000AD# => romdata <= X"00000000";
    when 16#000AE# => romdata <= X"00000000";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"0B0B0BBC";
    when 16#000B1# => romdata <= X"FA040000";
    when 16#000B2# => romdata <= X"00000000";
    when 16#000B3# => romdata <= X"00000000";
    when 16#000B4# => romdata <= X"00000000";
    when 16#000B5# => romdata <= X"00000000";
    when 16#000B6# => romdata <= X"00000000";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"80FC800C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"FF3D0D02";
    when 16#00101# => romdata <= X"8F053351";
    when 16#00102# => romdata <= X"BADE3F71";
    when 16#00103# => romdata <= X"B00C833D";
    when 16#00104# => romdata <= X"0D04FD3D";
    when 16#00105# => romdata <= X"0D818BE4";
    when 16#00106# => romdata <= X"0852F881";
    when 16#00107# => romdata <= X"C08E800B";
    when 16#00108# => romdata <= X"80FC8C08";
    when 16#00109# => romdata <= X"55537180";
    when 16#0010A# => romdata <= X"2E80F738";
    when 16#0010B# => romdata <= X"7281FF06";
    when 16#0010C# => romdata <= X"84150C80";
    when 16#0010D# => romdata <= X"FBE03370";
    when 16#0010E# => romdata <= X"81FF0651";
    when 16#0010F# => romdata <= X"5271802E";
    when 16#00110# => romdata <= X"80C23872";
    when 16#00111# => romdata <= X"9F2A7310";
    when 16#00112# => romdata <= X"0753818B";
    when 16#00113# => romdata <= X"E8337081";
    when 16#00114# => romdata <= X"FF065152";
    when 16#00115# => romdata <= X"71802ED4";
    when 16#00116# => romdata <= X"38800B81";
    when 16#00117# => romdata <= X"8BE83493";
    when 16#00118# => romdata <= X"EE3F80FB";
    when 16#00119# => romdata <= X"DC335473";
    when 16#0011A# => romdata <= X"80E23880";
    when 16#0011B# => romdata <= X"FC8C0873";
    when 16#0011C# => romdata <= X"81FF0684";
    when 16#0011D# => romdata <= X"120C80FB";
    when 16#0011E# => romdata <= X"E0337081";
    when 16#0011F# => romdata <= X"FF065153";
    when 16#00120# => romdata <= X"5471C038";
    when 16#00121# => romdata <= X"72812A73";
    when 16#00122# => romdata <= X"9F2B0753";
    when 16#00123# => romdata <= X"FFBC3972";
    when 16#00124# => romdata <= X"812A739F";
    when 16#00125# => romdata <= X"2B075380";
    when 16#00126# => romdata <= X"FD51B8B5";
    when 16#00127# => romdata <= X"3F80FC8C";
    when 16#00128# => romdata <= X"08547281";
    when 16#00129# => romdata <= X"FF068415";
    when 16#0012A# => romdata <= X"0C80FBE0";
    when 16#0012B# => romdata <= X"337081FF";
    when 16#0012C# => romdata <= X"06535471";
    when 16#0012D# => romdata <= X"802ED838";
    when 16#0012E# => romdata <= X"729F2A73";
    when 16#0012F# => romdata <= X"10075380";
    when 16#00130# => romdata <= X"FD51B88D";
    when 16#00131# => romdata <= X"3F80FC8C";
    when 16#00132# => romdata <= X"0854D739";
    when 16#00133# => romdata <= X"800BB00C";
    when 16#00134# => romdata <= X"853D0D04";
    when 16#00135# => romdata <= X"FB3D0D8A";
    when 16#00136# => romdata <= X"51B3F53F";
    when 16#00137# => romdata <= X"8AD73FAC";
    when 16#00138# => romdata <= X"87530B0B";
    when 16#00139# => romdata <= X"80E5EC52";
    when 16#0013A# => romdata <= X"0B0B80E5";
    when 16#0013B# => romdata <= X"FC518AD8";
    when 16#0013C# => romdata <= X"3FAC9E53";
    when 16#0013D# => romdata <= X"0B0B80E6";
    when 16#0013E# => romdata <= X"84520B0B";
    when 16#0013F# => romdata <= X"80E6A051";
    when 16#00140# => romdata <= X"8AC63FB4";
    when 16#00141# => romdata <= X"AF530B0B";
    when 16#00142# => romdata <= X"80E6A852";
    when 16#00143# => romdata <= X"0B0B80F2";
    when 16#00144# => romdata <= X"84518AB4";
    when 16#00145# => romdata <= X"3FB69753";
    when 16#00146# => romdata <= X"0B0B80E6";
    when 16#00147# => romdata <= X"C0520B0B";
    when 16#00148# => romdata <= X"80E6B851";
    when 16#00149# => romdata <= X"8AA23FB8";
    when 16#0014A# => romdata <= X"B8530B0B";
    when 16#0014B# => romdata <= X"80E6CC52";
    when 16#0014C# => romdata <= X"0B0B80E6";
    when 16#0014D# => romdata <= X"EC518A90";
    when 16#0014E# => romdata <= X"3FB9A353";
    when 16#0014F# => romdata <= X"0B0B80E6";
    when 16#00150# => romdata <= X"F4520B0B";
    when 16#00151# => romdata <= X"80E79851";
    when 16#00152# => romdata <= X"89FE3FB9";
    when 16#00153# => romdata <= X"DC530B0B";
    when 16#00154# => romdata <= X"80E7A052";
    when 16#00155# => romdata <= X"0B0B80E7";
    when 16#00156# => romdata <= X"BC5189EC";
    when 16#00157# => romdata <= X"3FBA9253";
    when 16#00158# => romdata <= X"0B0B80E7";
    when 16#00159# => romdata <= X"C4520B0B";
    when 16#0015A# => romdata <= X"80E7E851";
    when 16#0015B# => romdata <= X"89DA3FB8";
    when 16#0015C# => romdata <= X"F8530B0B";
    when 16#0015D# => romdata <= X"80E7F052";
    when 16#0015E# => romdata <= X"0B0B80E8";
    when 16#0015F# => romdata <= X"885189C8";
    when 16#00160# => romdata <= X"3FB99153";
    when 16#00161# => romdata <= X"0B0B80E8";
    when 16#00162# => romdata <= X"90520B0B";
    when 16#00163# => romdata <= X"80E8AC51";
    when 16#00164# => romdata <= X"89B63FB7";
    when 16#00165# => romdata <= X"8D530B0B";
    when 16#00166# => romdata <= X"80E8B452";
    when 16#00167# => romdata <= X"0B0B80E8";
    when 16#00168# => romdata <= X"CC5189A4";
    when 16#00169# => romdata <= X"3FB7E353";
    when 16#0016A# => romdata <= X"0B0B80E8";
    when 16#0016B# => romdata <= X"D4520B0B";
    when 16#0016C# => romdata <= X"80E8F051";
    when 16#0016D# => romdata <= X"89923F91";
    when 16#0016E# => romdata <= X"A2530B0B";
    when 16#0016F# => romdata <= X"80E8F852";
    when 16#00170# => romdata <= X"0B0B80E9";
    when 16#00171# => romdata <= X"8C518980";
    when 16#00172# => romdata <= X"3F90E253";
    when 16#00173# => romdata <= X"0B0B80E9";
    when 16#00174# => romdata <= X"94520B0B";
    when 16#00175# => romdata <= X"80E9BC51";
    when 16#00176# => romdata <= X"88EE3FB3";
    when 16#00177# => romdata <= X"90530B0B";
    when 16#00178# => romdata <= X"80E9C452";
    when 16#00179# => romdata <= X"0B0B80E9";
    when 16#0017A# => romdata <= X"D85188DC";
    when 16#0017B# => romdata <= X"3F889253";
    when 16#0017C# => romdata <= X"0B0B80E9";
    when 16#0017D# => romdata <= X"E0520B0B";
    when 16#0017E# => romdata <= X"80E9F051";
    when 16#0017F# => romdata <= X"88CA3FA6";
    when 16#00180# => romdata <= X"C0530B0B";
    when 16#00181# => romdata <= X"80E9F452";
    when 16#00182# => romdata <= X"0B0B80EA";
    when 16#00183# => romdata <= X"885188B8";
    when 16#00184# => romdata <= X"3FA9C853";
    when 16#00185# => romdata <= X"0B0B80EA";
    when 16#00186# => romdata <= X"8C520B0B";
    when 16#00187# => romdata <= X"80EAB451";
    when 16#00188# => romdata <= X"88A63FB4";
    when 16#00189# => romdata <= X"83530B0B";
    when 16#0018A# => romdata <= X"80EABC52";
    when 16#0018B# => romdata <= X"0B0B80EA";
    when 16#0018C# => romdata <= X"CC518894";
    when 16#0018D# => romdata <= X"3F929C53";
    when 16#0018E# => romdata <= X"0B0B80EA";
    when 16#0018F# => romdata <= X"D0520B0B";
    when 16#00190# => romdata <= X"80EAE851";
    when 16#00191# => romdata <= X"88823FAA";
    when 16#00192# => romdata <= X"82530B0B";
    when 16#00193# => romdata <= X"80EAF052";
    when 16#00194# => romdata <= X"0B0B80EA";
    when 16#00195# => romdata <= X"FC5187F0";
    when 16#00196# => romdata <= X"3FABB153";
    when 16#00197# => romdata <= X"0B0B80EB";
    when 16#00198# => romdata <= X"80520B0B";
    when 16#00199# => romdata <= X"80EBA851";
    when 16#0019A# => romdata <= X"87DE3FAA";
    when 16#0019B# => romdata <= X"82530B0B";
    when 16#0019C# => romdata <= X"80EBB052";
    when 16#0019D# => romdata <= X"0B0B80EB";
    when 16#0019E# => romdata <= X"D05187CC";
    when 16#0019F# => romdata <= X"3FABF753";
    when 16#001A0# => romdata <= X"0B0B80EB";
    when 16#001A1# => romdata <= X"D4520B0B";
    when 16#001A2# => romdata <= X"80EBE451";
    when 16#001A3# => romdata <= X"87BA3F90";
    when 16#001A4# => romdata <= X"AE530B0B";
    when 16#001A5# => romdata <= X"80F5FC52";
    when 16#001A6# => romdata <= X"0B0B80E5";
    when 16#001A7# => romdata <= X"E45187A8";
    when 16#001A8# => romdata <= X"3F8E8C3F";
    when 16#001A9# => romdata <= X"87FF3F81";
    when 16#001AA# => romdata <= X"0B81A3D8";
    when 16#001AB# => romdata <= X"34818BE8";
    when 16#001AC# => romdata <= X"337081FF";
    when 16#001AD# => romdata <= X"06555573";
    when 16#001AE# => romdata <= X"81EA38B4";
    when 16#001AF# => romdata <= X"F63FB008";
    when 16#001B0# => romdata <= X"81D33887";
    when 16#001B1# => romdata <= X"EE3F80FC";
    when 16#001B2# => romdata <= X"8C087008";
    when 16#001B3# => romdata <= X"70842A81";
    when 16#001B4# => romdata <= X"06515556";
    when 16#001B5# => romdata <= X"73802E80";
    when 16#001B6# => romdata <= X"F238F881";
    when 16#001B7# => romdata <= X"C08E8055";
    when 16#001B8# => romdata <= X"818BE408";
    when 16#001B9# => romdata <= X"802E8183";
    when 16#001BA# => romdata <= X"387481FF";
    when 16#001BB# => romdata <= X"0684170C";
    when 16#001BC# => romdata <= X"80FBE033";
    when 16#001BD# => romdata <= X"7081FF06";
    when 16#001BE# => romdata <= X"51547380";
    when 16#001BF# => romdata <= X"2E80C138";
    when 16#001C0# => romdata <= X"749F2A75";
    when 16#001C1# => romdata <= X"10075581";
    when 16#001C2# => romdata <= X"8BE83370";
    when 16#001C3# => romdata <= X"81FF0651";
    when 16#001C4# => romdata <= X"5473802E";
    when 16#001C5# => romdata <= X"D438800B";
    when 16#001C6# => romdata <= X"818BE834";
    when 16#001C7# => romdata <= X"8EB13F80";
    when 16#001C8# => romdata <= X"FBDC3356";
    when 16#001C9# => romdata <= X"75A53880";
    when 16#001CA# => romdata <= X"FC8C0875";
    when 16#001CB# => romdata <= X"81FF0684";
    when 16#001CC# => romdata <= X"120C80FB";
    when 16#001CD# => romdata <= X"E0337081";
    when 16#001CE# => romdata <= X"FF065155";
    when 16#001CF# => romdata <= X"5673C138";
    when 16#001D0# => romdata <= X"74812A75";
    when 16#001D1# => romdata <= X"9F2B0755";
    when 16#001D2# => romdata <= X"FFBD3981";
    when 16#001D3# => romdata <= X"A3D83355";
    when 16#001D4# => romdata <= X"74FEDA38";
    when 16#001D5# => romdata <= X"873D0D04";
    when 16#001D6# => romdata <= X"74812A75";
    when 16#001D7# => romdata <= X"9F2B0755";
    when 16#001D8# => romdata <= X"80FD51B2";
    when 16#001D9# => romdata <= X"EC3F80FC";
    when 16#001DA# => romdata <= X"8C085674";
    when 16#001DB# => romdata <= X"81FF0684";
    when 16#001DC# => romdata <= X"170C80FB";
    when 16#001DD# => romdata <= X"E0337081";
    when 16#001DE# => romdata <= X"FF065754";
    when 16#001DF# => romdata <= X"75802ED8";
    when 16#001E0# => romdata <= X"38749F2A";
    when 16#001E1# => romdata <= X"75100755";
    when 16#001E2# => romdata <= X"80FD51B2";
    when 16#001E3# => romdata <= X"C43F80FC";
    when 16#001E4# => romdata <= X"8C0856D7";
    when 16#001E5# => romdata <= X"39B3AF3F";
    when 16#001E6# => romdata <= X"B00881FF";
    when 16#001E7# => romdata <= X"06518781";
    when 16#001E8# => romdata <= X"3FFEA039";
    when 16#001E9# => romdata <= X"800B818B";
    when 16#001EA# => romdata <= X"E8348DA3";
    when 16#001EB# => romdata <= X"3FB3843F";
    when 16#001EC# => romdata <= X"B008802E";
    when 16#001ED# => romdata <= X"FE8D38DD";
    when 16#001EE# => romdata <= X"39803D0D";
    when 16#001EF# => romdata <= X"0B0B80EB";
    when 16#001F0# => romdata <= X"EC51AEA6";
    when 16#001F1# => romdata <= X"3F8C51AE";
    when 16#001F2# => romdata <= X"873F0B0B";
    when 16#001F3# => romdata <= X"80EBF051";
    when 16#001F4# => romdata <= X"AE983F81";
    when 16#001F5# => romdata <= X"8BE40880";
    when 16#001F6# => romdata <= X"2E8E380B";
    when 16#001F7# => romdata <= X"0B80EC88";
    when 16#001F8# => romdata <= X"51AE873F";
    when 16#001F9# => romdata <= X"823D0D04";
    when 16#001FA# => romdata <= X"0B0B80EC";
    when 16#001FB# => romdata <= X"9451ADFA";
    when 16#001FC# => romdata <= X"3F810A51";
    when 16#001FD# => romdata <= X"ADF43F0B";
    when 16#001FE# => romdata <= X"0B80ECA8";
    when 16#001FF# => romdata <= X"51ADEB3F";
    when 16#00200# => romdata <= X"0B0B80EC";
    when 16#00201# => romdata <= X"D051ADE2";
    when 16#00202# => romdata <= X"3F80E451";
    when 16#00203# => romdata <= X"AFA63F0B";
    when 16#00204# => romdata <= X"0B80ECE4";
    when 16#00205# => romdata <= X"51ADD33F";
    when 16#00206# => romdata <= X"0B0B80EC";
    when 16#00207# => romdata <= X"EC51ADCA";
    when 16#00208# => romdata <= X"3F0B0B80";
    when 16#00209# => romdata <= X"ECF851AD";
    when 16#0020A# => romdata <= X"C13F823D";
    when 16#0020B# => romdata <= X"0D04FF89";
    when 16#0020C# => romdata <= X"3F8AFC3F";
    when 16#0020D# => romdata <= X"800BB00C";
    when 16#0020E# => romdata <= X"04FE3D0D";
    when 16#0020F# => romdata <= X"80FC9008";
    when 16#00210# => romdata <= X"98110870";
    when 16#00211# => romdata <= X"842A7081";
    when 16#00212# => romdata <= X"06515353";
    when 16#00213# => romdata <= X"5370802E";
    when 16#00214# => romdata <= X"8D3871EF";
    when 16#00215# => romdata <= X"0698140C";
    when 16#00216# => romdata <= X"810B818B";
    when 16#00217# => romdata <= X"E834843D";
    when 16#00218# => romdata <= X"0D04F93D";
    when 16#00219# => romdata <= X"0D815189";
    when 16#0021A# => romdata <= X"943FB008";
    when 16#0021B# => romdata <= X"55825189";
    when 16#0021C# => romdata <= X"8C3F74B0";
    when 16#0021D# => romdata <= X"08075399";
    when 16#0021E# => romdata <= X"CC57FCE2";
    when 16#0021F# => romdata <= X"97F68058";
    when 16#00220# => romdata <= X"72802E90";
    when 16#00221# => romdata <= X"38747554";
    when 16#00222# => romdata <= X"57805480";
    when 16#00223# => romdata <= X"770774B0";
    when 16#00224# => romdata <= X"08075957";
    when 16#00225# => romdata <= X"76517752";
    when 16#00226# => romdata <= X"9BFA3F72";
    when 16#00227# => romdata <= X"B00C893D";
    when 16#00228# => romdata <= X"0D04FB3D";
    when 16#00229# => romdata <= X"0D815187";
    when 16#0022A# => romdata <= X"A23FB008";
    when 16#0022B# => romdata <= X"56815382";
    when 16#0022C# => romdata <= X"528051A5";
    when 16#0022D# => romdata <= X"A83F80FB";
    when 16#0022E# => romdata <= X"EC085589";
    when 16#0022F# => romdata <= X"750C80FC";
    when 16#00230# => romdata <= X"8C088411";
    when 16#00231# => romdata <= X"0870810A";
    when 16#00232# => romdata <= X"0784130C";
    when 16#00233# => romdata <= X"55557551";
    when 16#00234# => romdata <= X"AFD93F80";
    when 16#00235# => romdata <= X"FC8C0884";
    when 16#00236# => romdata <= X"110870FE";
    when 16#00237# => romdata <= X"0A068413";
    when 16#00238# => romdata <= X"0C555581";
    when 16#00239# => romdata <= X"53825280";
    when 16#0023A# => romdata <= X"51A4F23F";
    when 16#0023B# => romdata <= X"80FBEC08";
    when 16#0023C# => romdata <= X"5589750C";
    when 16#0023D# => romdata <= X"80FC8C08";
    when 16#0023E# => romdata <= X"84110870";
    when 16#0023F# => romdata <= X"810A0784";
    when 16#00240# => romdata <= X"130C5555";
    when 16#00241# => romdata <= X"7551AFA3";
    when 16#00242# => romdata <= X"3F80FC8C";
    when 16#00243# => romdata <= X"08841108";
    when 16#00244# => romdata <= X"70FE0A06";
    when 16#00245# => romdata <= X"84130C55";
    when 16#00246# => romdata <= X"55FF9239";
    when 16#00247# => romdata <= X"FE3D0D81";
    when 16#00248# => romdata <= X"5186A83F";
    when 16#00249# => romdata <= X"80FC8C08";
    when 16#0024A# => romdata <= X"84110870";
    when 16#0024B# => romdata <= X"810A0784";
    when 16#0024C# => romdata <= X"130C5353";
    when 16#0024D# => romdata <= X"B00851AE";
    when 16#0024E# => romdata <= X"F23F80FC";
    when 16#0024F# => romdata <= X"8C088411";
    when 16#00250# => romdata <= X"0870FE0A";
    when 16#00251# => romdata <= X"06708414";
    when 16#00252# => romdata <= X"0CB00C53";
    when 16#00253# => romdata <= X"53843D0D";
    when 16#00254# => romdata <= X"04FC3D0D";
    when 16#00255# => romdata <= X"80FC8C08";
    when 16#00256# => romdata <= X"7008810A";
    when 16#00257# => romdata <= X"06818BE4";
    when 16#00258# => romdata <= X"0C54AF91";
    when 16#00259# => romdata <= X"3FAFB53F";
    when 16#0025A# => romdata <= X"8AC53F93";
    when 16#0025B# => romdata <= X"8C3F80FC";
    when 16#0025C# => romdata <= X"90089811";
    when 16#0025D# => romdata <= X"08708807";
    when 16#0025E# => romdata <= X"98130C55";
    when 16#0025F# => romdata <= X"55818BE4";
    when 16#00260# => romdata <= X"0880D538";
    when 16#00261# => romdata <= X"88800B81";
    when 16#00262# => romdata <= X"A4B40CFC";
    when 16#00263# => romdata <= X"AC3F818B";
    when 16#00264# => romdata <= X"E408802E";
    when 16#00265# => romdata <= X"80D33881";
    when 16#00266# => romdata <= X"53825280";
    when 16#00267# => romdata <= X"51A3BE3F";
    when 16#00268# => romdata <= X"80FBEC08";
    when 16#00269# => romdata <= X"5589750C";
    when 16#0026A# => romdata <= X"80FC8C08";
    when 16#0026B# => romdata <= X"84110870";
    when 16#0026C# => romdata <= X"810A0784";
    when 16#0026D# => romdata <= X"130C5555";
    when 16#0026E# => romdata <= X"8051ADEF";
    when 16#0026F# => romdata <= X"3F80FC8C";
    when 16#00270# => romdata <= X"08841108";
    when 16#00271# => romdata <= X"70FE0A06";
    when 16#00272# => romdata <= X"84130C55";
    when 16#00273# => romdata <= X"5580FBEC";
    when 16#00274# => romdata <= X"08558075";
    when 16#00275# => romdata <= X"0CB0AB3F";
    when 16#00276# => romdata <= X"BDBA0B81";
    when 16#00277# => romdata <= X"A4B40CFB";
    when 16#00278# => romdata <= X"D83F818B";
    when 16#00279# => romdata <= X"E408FFAF";
    when 16#0027A# => romdata <= X"3880C2E8";
    when 16#0027B# => romdata <= X"0B81A4B4";
    when 16#0027C# => romdata <= X"0CF5E13F";
    when 16#0027D# => romdata <= X"81538252";
    when 16#0027E# => romdata <= X"8051A2E1";
    when 16#0027F# => romdata <= X"3F80FBEC";
    when 16#00280# => romdata <= X"08558975";
    when 16#00281# => romdata <= X"0C80FC8C";
    when 16#00282# => romdata <= X"08841108";
    when 16#00283# => romdata <= X"70810A07";
    when 16#00284# => romdata <= X"84130C55";
    when 16#00285# => romdata <= X"558051AD";
    when 16#00286# => romdata <= X"923F80FC";
    when 16#00287# => romdata <= X"8C088411";
    when 16#00288# => romdata <= X"0870FE0A";
    when 16#00289# => romdata <= X"0684130C";
    when 16#0028A# => romdata <= X"555580FB";
    when 16#0028B# => romdata <= X"EC085580";
    when 16#0028C# => romdata <= X"750CAFCE";
    when 16#0028D# => romdata <= X"3F800B81";
    when 16#0028E# => romdata <= X"A3D03480";
    when 16#0028F# => romdata <= X"0B81A3CC";
    when 16#00290# => romdata <= X"34800B81";
    when 16#00291# => romdata <= X"A3D40C04";
    when 16#00292# => romdata <= X"FC3D0D81";
    when 16#00293# => romdata <= X"A3CC3353";
    when 16#00294# => romdata <= X"72A72680";
    when 16#00295# => romdata <= X"C5387652";
    when 16#00296# => romdata <= X"72101010";
    when 16#00297# => romdata <= X"73100581";
    when 16#00298# => romdata <= X"8BEC0551";
    when 16#00299# => romdata <= X"B4B73F77";
    when 16#0029A# => romdata <= X"5281A3CC";
    when 16#0029B# => romdata <= X"33709029";
    when 16#0029C# => romdata <= X"71317010";
    when 16#0029D# => romdata <= X"10818EFC";
    when 16#0029E# => romdata <= X"05535654";
    when 16#0029F# => romdata <= X"B49F3F81";
    when 16#002A0# => romdata <= X"A3CC3370";
    when 16#002A1# => romdata <= X"101081A1";
    when 16#002A2# => romdata <= X"DC057A71";
    when 16#002A3# => romdata <= X"0C548105";
    when 16#002A4# => romdata <= X"537281A3";
    when 16#002A5# => romdata <= X"CC34863D";
    when 16#002A6# => romdata <= X"0D0480ED";
    when 16#002A7# => romdata <= X"8051A8CA";
    when 16#002A8# => romdata <= X"3F863D0D";
    when 16#002A9# => romdata <= X"04803D0D";
    when 16#002AA# => romdata <= X"80ED9C51";
    when 16#002AB# => romdata <= X"A8BC3F82";
    when 16#002AC# => romdata <= X"3D0D04FE";
    when 16#002AD# => romdata <= X"3D0D81A3";
    when 16#002AE# => romdata <= X"D4085372";
    when 16#002AF# => romdata <= X"8538843D";
    when 16#002B0# => romdata <= X"0D04722D";
    when 16#002B1# => romdata <= X"B0085380";
    when 16#002B2# => romdata <= X"0B81A3D4";
    when 16#002B3# => romdata <= X"0CB0088C";
    when 16#002B4# => romdata <= X"3880ED9C";
    when 16#002B5# => romdata <= X"51A8933F";
    when 16#002B6# => romdata <= X"843D0D04";
    when 16#002B7# => romdata <= X"80F8CC51";
    when 16#002B8# => romdata <= X"A8883F72";
    when 16#002B9# => romdata <= X"83FFFF26";
    when 16#002BA# => romdata <= X"AA3881FF";
    when 16#002BB# => romdata <= X"73279638";
    when 16#002BC# => romdata <= X"72529051";
    when 16#002BD# => romdata <= X"A8973F8A";
    when 16#002BE# => romdata <= X"51A7D53F";
    when 16#002BF# => romdata <= X"80ED9C51";
    when 16#002C0# => romdata <= X"A7E83FD4";
    when 16#002C1# => romdata <= X"39725288";
    when 16#002C2# => romdata <= X"51A8823F";
    when 16#002C3# => romdata <= X"8A51A7C0";
    when 16#002C4# => romdata <= X"3FEA3972";
    when 16#002C5# => romdata <= X"52A051A7";
    when 16#002C6# => romdata <= X"F43F8A51";
    when 16#002C7# => romdata <= X"A7B23FDC";
    when 16#002C8# => romdata <= X"39FA3D0D";
    when 16#002C9# => romdata <= X"02A30533";
    when 16#002CA# => romdata <= X"56758D2E";
    when 16#002CB# => romdata <= X"80F43875";
    when 16#002CC# => romdata <= X"88327030";
    when 16#002CD# => romdata <= X"7780FF32";
    when 16#002CE# => romdata <= X"70307280";
    when 16#002CF# => romdata <= X"25718025";
    when 16#002D0# => romdata <= X"07545156";
    when 16#002D1# => romdata <= X"58557495";
    when 16#002D2# => romdata <= X"389F7627";
    when 16#002D3# => romdata <= X"8C3881A3";
    when 16#002D4# => romdata <= X"D0335580";
    when 16#002D5# => romdata <= X"CE7527AE";
    when 16#002D6# => romdata <= X"38883D0D";
    when 16#002D7# => romdata <= X"0481A3D0";
    when 16#002D8# => romdata <= X"33567580";
    when 16#002D9# => romdata <= X"2EF33888";
    when 16#002DA# => romdata <= X"51A6E53F";
    when 16#002DB# => romdata <= X"A051A6E0";
    when 16#002DC# => romdata <= X"3F8851A6";
    when 16#002DD# => romdata <= X"DB3F81A3";
    when 16#002DE# => romdata <= X"D033FF05";
    when 16#002DF# => romdata <= X"577681A3";
    when 16#002E0# => romdata <= X"D034883D";
    when 16#002E1# => romdata <= X"0D047551";
    when 16#002E2# => romdata <= X"A6C63F81";
    when 16#002E3# => romdata <= X"A3D03381";
    when 16#002E4# => romdata <= X"11555773";
    when 16#002E5# => romdata <= X"81A3D034";
    when 16#002E6# => romdata <= X"7581A2FC";
    when 16#002E7# => romdata <= X"1834883D";
    when 16#002E8# => romdata <= X"0D048A51";
    when 16#002E9# => romdata <= X"A6AA3F81";
    when 16#002EA# => romdata <= X"A3D03381";
    when 16#002EB# => romdata <= X"11565474";
    when 16#002EC# => romdata <= X"81A3D034";
    when 16#002ED# => romdata <= X"800B81A2";
    when 16#002EE# => romdata <= X"FC153480";
    when 16#002EF# => romdata <= X"56800B81";
    when 16#002F0# => romdata <= X"A2FC1733";
    when 16#002F1# => romdata <= X"565474A0";
    when 16#002F2# => romdata <= X"2E833881";
    when 16#002F3# => romdata <= X"5474802E";
    when 16#002F4# => romdata <= X"90387380";
    when 16#002F5# => romdata <= X"2E8B3881";
    when 16#002F6# => romdata <= X"167081FF";
    when 16#002F7# => romdata <= X"065757DD";
    when 16#002F8# => romdata <= X"3975802E";
    when 16#002F9# => romdata <= X"BF38800B";
    when 16#002FA# => romdata <= X"81A3CC33";
    when 16#002FB# => romdata <= X"55557474";
    when 16#002FC# => romdata <= X"27AB3873";
    when 16#002FD# => romdata <= X"57741010";
    when 16#002FE# => romdata <= X"10751005";
    when 16#002FF# => romdata <= X"765481A2";
    when 16#00300# => romdata <= X"FC53818B";
    when 16#00301# => romdata <= X"EC0551B2";
    when 16#00302# => romdata <= X"E03FB008";
    when 16#00303# => romdata <= X"802EA638";
    when 16#00304# => romdata <= X"81157081";
    when 16#00305# => romdata <= X"FF065654";
    when 16#00306# => romdata <= X"767526D9";
    when 16#00307# => romdata <= X"3880EDA0";
    when 16#00308# => romdata <= X"51A5C73F";
    when 16#00309# => romdata <= X"80ED9C51";
    when 16#0030A# => romdata <= X"A5C03F80";
    when 16#0030B# => romdata <= X"0B81A3D0";
    when 16#0030C# => romdata <= X"34883D0D";
    when 16#0030D# => romdata <= X"04741010";
    when 16#0030E# => romdata <= X"81A1DC05";
    when 16#0030F# => romdata <= X"700881A3";
    when 16#00310# => romdata <= X"D40C5680";
    when 16#00311# => romdata <= X"0B81A3D0";
    when 16#00312# => romdata <= X"34E739F7";
    when 16#00313# => romdata <= X"3D0D02AF";
    when 16#00314# => romdata <= X"05335980";
    when 16#00315# => romdata <= X"0B81A2FC";
    when 16#00316# => romdata <= X"3381A2FC";
    when 16#00317# => romdata <= X"59555673";
    when 16#00318# => romdata <= X"A02E0981";
    when 16#00319# => romdata <= X"06963881";
    when 16#0031A# => romdata <= X"167081FF";
    when 16#0031B# => romdata <= X"0681A2FC";
    when 16#0031C# => romdata <= X"11703353";
    when 16#0031D# => romdata <= X"59575473";
    when 16#0031E# => romdata <= X"A02EEC38";
    when 16#0031F# => romdata <= X"80587779";
    when 16#00320# => romdata <= X"2780EA38";
    when 16#00321# => romdata <= X"80773356";
    when 16#00322# => romdata <= X"5474742E";
    when 16#00323# => romdata <= X"83388154";
    when 16#00324# => romdata <= X"74A02E9A";
    when 16#00325# => romdata <= X"387380C5";
    when 16#00326# => romdata <= X"3874A02E";
    when 16#00327# => romdata <= X"91388118";
    when 16#00328# => romdata <= X"7081FF06";
    when 16#00329# => romdata <= X"59557878";
    when 16#0032A# => romdata <= X"26DA3880";
    when 16#0032B# => romdata <= X"C0398116";
    when 16#0032C# => romdata <= X"7081FF06";
    when 16#0032D# => romdata <= X"81A2FC11";
    when 16#0032E# => romdata <= X"70335752";
    when 16#0032F# => romdata <= X"575773A0";
    when 16#00330# => romdata <= X"2E098106";
    when 16#00331# => romdata <= X"D9388116";
    when 16#00332# => romdata <= X"7081FF06";
    when 16#00333# => romdata <= X"81A2FC11";
    when 16#00334# => romdata <= X"70335752";
    when 16#00335# => romdata <= X"575773A0";
    when 16#00336# => romdata <= X"2ED438C2";
    when 16#00337# => romdata <= X"39811670";
    when 16#00338# => romdata <= X"81FF0681";
    when 16#00339# => romdata <= X"A2FC1159";
    when 16#0033A# => romdata <= X"5755FF98";
    when 16#0033B# => romdata <= X"3980538B";
    when 16#0033C# => romdata <= X"3DFC0552";
    when 16#0033D# => romdata <= X"7651B5B6";
    when 16#0033E# => romdata <= X"3F8B3D0D";
    when 16#0033F# => romdata <= X"04F73D0D";
    when 16#00340# => romdata <= X"02AF0533";
    when 16#00341# => romdata <= X"59800B81";
    when 16#00342# => romdata <= X"A2FC3381";
    when 16#00343# => romdata <= X"A2FC5955";
    when 16#00344# => romdata <= X"5673A02E";
    when 16#00345# => romdata <= X"09810696";
    when 16#00346# => romdata <= X"38811670";
    when 16#00347# => romdata <= X"81FF0681";
    when 16#00348# => romdata <= X"A2FC1170";
    when 16#00349# => romdata <= X"33535957";
    when 16#0034A# => romdata <= X"5473A02E";
    when 16#0034B# => romdata <= X"EC388058";
    when 16#0034C# => romdata <= X"77792780";
    when 16#0034D# => romdata <= X"EA388077";
    when 16#0034E# => romdata <= X"33565474";
    when 16#0034F# => romdata <= X"742E8338";
    when 16#00350# => romdata <= X"815474A0";
    when 16#00351# => romdata <= X"2E9A3873";
    when 16#00352# => romdata <= X"80C53874";
    when 16#00353# => romdata <= X"A02E9138";
    when 16#00354# => romdata <= X"81187081";
    when 16#00355# => romdata <= X"FF065955";
    when 16#00356# => romdata <= X"787826DA";
    when 16#00357# => romdata <= X"3880C039";
    when 16#00358# => romdata <= X"81167081";
    when 16#00359# => romdata <= X"FF0681A2";
    when 16#0035A# => romdata <= X"FC117033";
    when 16#0035B# => romdata <= X"57525757";
    when 16#0035C# => romdata <= X"73A02E09";
    when 16#0035D# => romdata <= X"8106D938";
    when 16#0035E# => romdata <= X"81167081";
    when 16#0035F# => romdata <= X"FF0681A2";
    when 16#00360# => romdata <= X"FC117033";
    when 16#00361# => romdata <= X"57525757";
    when 16#00362# => romdata <= X"73A02ED4";
    when 16#00363# => romdata <= X"38C23981";
    when 16#00364# => romdata <= X"167081FF";
    when 16#00365# => romdata <= X"0681A2FC";
    when 16#00366# => romdata <= X"11595755";
    when 16#00367# => romdata <= X"FF983990";
    when 16#00368# => romdata <= X"538B3DFC";
    when 16#00369# => romdata <= X"05527651";
    when 16#0036A# => romdata <= X"B7A13F8B";
    when 16#0036B# => romdata <= X"3D0D04FC";
    when 16#0036C# => romdata <= X"3D0D8A51";
    when 16#0036D# => romdata <= X"A29A3F80";
    when 16#0036E# => romdata <= X"EDB451A2";
    when 16#0036F# => romdata <= X"AD3F800B";
    when 16#00370# => romdata <= X"81A3CC33";
    when 16#00371# => romdata <= X"53537272";
    when 16#00372# => romdata <= X"2780F538";
    when 16#00373# => romdata <= X"72101010";
    when 16#00374# => romdata <= X"73100581";
    when 16#00375# => romdata <= X"8BEC0570";
    when 16#00376# => romdata <= X"5254A28E";
    when 16#00377# => romdata <= X"3F72842B";
    when 16#00378# => romdata <= X"70743182";
    when 16#00379# => romdata <= X"2B818EFC";
    when 16#0037A# => romdata <= X"11335153";
    when 16#0037B# => romdata <= X"5571802E";
    when 16#0037C# => romdata <= X"B7387351";
    when 16#0037D# => romdata <= X"AE943FB0";
    when 16#0037E# => romdata <= X"0881FF06";
    when 16#0037F# => romdata <= X"52718926";
    when 16#00380# => romdata <= X"9338A051";
    when 16#00381# => romdata <= X"A1CA3F81";
    when 16#00382# => romdata <= X"127081FF";
    when 16#00383# => romdata <= X"06535489";
    when 16#00384# => romdata <= X"7227EF38";
    when 16#00385# => romdata <= X"80EDCC51";
    when 16#00386# => romdata <= X"A1D03F74";
    when 16#00387# => romdata <= X"7331822B";
    when 16#00388# => romdata <= X"818EFC05";
    when 16#00389# => romdata <= X"51A1C33F";
    when 16#0038A# => romdata <= X"8A51A1A4";
    when 16#0038B# => romdata <= X"3F811370";
    when 16#0038C# => romdata <= X"81FF0681";
    when 16#0038D# => romdata <= X"A3CC3354";
    when 16#0038E# => romdata <= X"54557173";
    when 16#0038F# => romdata <= X"26FF8D38";
    when 16#00390# => romdata <= X"8A51A18C";
    when 16#00391# => romdata <= X"3F81A3CC";
    when 16#00392# => romdata <= X"33B00C86";
    when 16#00393# => romdata <= X"3D0D04FE";
    when 16#00394# => romdata <= X"3D0D81A4";
    when 16#00395# => romdata <= X"AC22FF05";
    when 16#00396# => romdata <= X"517081A4";
    when 16#00397# => romdata <= X"AC237083";
    when 16#00398# => romdata <= X"FFFF0651";
    when 16#00399# => romdata <= X"7080C438";
    when 16#0039A# => romdata <= X"81A4B033";
    when 16#0039B# => romdata <= X"517081FF";
    when 16#0039C# => romdata <= X"2EB93870";
    when 16#0039D# => romdata <= X"10101081";
    when 16#0039E# => romdata <= X"A3DC0552";
    when 16#0039F# => romdata <= X"713381A4";
    when 16#003A0# => romdata <= X"B034FE72";
    when 16#003A1# => romdata <= X"3481A4B0";
    when 16#003A2# => romdata <= X"33701010";
    when 16#003A3# => romdata <= X"1081A3DC";
    when 16#003A4# => romdata <= X"05525382";
    when 16#003A5# => romdata <= X"112281A4";
    when 16#003A6# => romdata <= X"AC238412";
    when 16#003A7# => romdata <= X"0853722D";
    when 16#003A8# => romdata <= X"81A4AC22";
    when 16#003A9# => romdata <= X"5170802E";
    when 16#003AA# => romdata <= X"FFBE3884";
    when 16#003AB# => romdata <= X"3D0D04FF";
    when 16#003AC# => romdata <= X"3D0D8A52";
    when 16#003AD# => romdata <= X"71101010";
    when 16#003AE# => romdata <= X"81A3D405";
    when 16#003AF# => romdata <= X"51FE7134";
    when 16#003B0# => romdata <= X"FF127081";
    when 16#003B1# => romdata <= X"FF065351";
    when 16#003B2# => romdata <= X"71EA38FF";
    when 16#003B3# => romdata <= X"0B81A4B0";
    when 16#003B4# => romdata <= X"34833D0D";
    when 16#003B5# => romdata <= X"04FE3D0D";
    when 16#003B6# => romdata <= X"02930533";
    when 16#003B7# => romdata <= X"02840597";
    when 16#003B8# => romdata <= X"05335452";
    when 16#003B9# => romdata <= X"71842E80";
    when 16#003BA# => romdata <= X"D1387184";
    when 16#003BB# => romdata <= X"24913871";
    when 16#003BC# => romdata <= X"812EAC38";
    when 16#003BD# => romdata <= X"80EDD051";
    when 16#003BE# => romdata <= X"9FF03F84";
    when 16#003BF# => romdata <= X"3D0D0471";
    when 16#003C0# => romdata <= X"80D52E09";
    when 16#003C1# => romdata <= X"8106ED38";
    when 16#003C2# => romdata <= X"80EDDC51";
    when 16#003C3# => romdata <= X"9FDC3F72";
    when 16#003C4# => romdata <= X"8C26B338";
    when 16#003C5# => romdata <= X"72101080";
    when 16#003C6# => romdata <= X"F2D00552";
    when 16#003C7# => romdata <= X"71080480";
    when 16#003C8# => romdata <= X"EDE8519F";
    when 16#003C9# => romdata <= X"C53FFA13";
    when 16#003CA# => romdata <= X"527180DB";
    when 16#003CB# => romdata <= X"26983871";
    when 16#003CC# => romdata <= X"101080F3";
    when 16#003CD# => romdata <= X"84055271";
    when 16#003CE# => romdata <= X"080480ED";
    when 16#003CF# => romdata <= X"F4519FAA";
    when 16#003D0# => romdata <= X"3F728F2E";
    when 16#003D1# => romdata <= X"8C3880EE";
    when 16#003D2# => romdata <= X"80519F9E";
    when 16#003D3# => romdata <= X"3F843D0D";
    when 16#003D4# => romdata <= X"0480EE90";
    when 16#003D5# => romdata <= X"519F933F";
    when 16#003D6# => romdata <= X"843D0D04";
    when 16#003D7# => romdata <= X"80EEA851";
    when 16#003D8# => romdata <= X"9F883F84";
    when 16#003D9# => romdata <= X"3D0D0480";
    when 16#003DA# => romdata <= X"EEB8519E";
    when 16#003DB# => romdata <= X"FD3F843D";
    when 16#003DC# => romdata <= X"0D0480EE";
    when 16#003DD# => romdata <= X"D0519EF2";
    when 16#003DE# => romdata <= X"3F843D0D";
    when 16#003DF# => romdata <= X"0480EEE0";
    when 16#003E0# => romdata <= X"519EE73F";
    when 16#003E1# => romdata <= X"843D0D04";
    when 16#003E2# => romdata <= X"80EF8051";
    when 16#003E3# => romdata <= X"9EDC3F84";
    when 16#003E4# => romdata <= X"3D0D0480";
    when 16#003E5# => romdata <= X"EF9C519E";
    when 16#003E6# => romdata <= X"D13F843D";
    when 16#003E7# => romdata <= X"0D0480EF";
    when 16#003E8# => romdata <= X"B8519EC6";
    when 16#003E9# => romdata <= X"3F843D0D";
    when 16#003EA# => romdata <= X"0480EFCC";
    when 16#003EB# => romdata <= X"519EBB3F";
    when 16#003EC# => romdata <= X"843D0D04";
    when 16#003ED# => romdata <= X"80EFE851";
    when 16#003EE# => romdata <= X"9EB03F84";
    when 16#003EF# => romdata <= X"3D0D0480";
    when 16#003F0# => romdata <= X"EFF8519E";
    when 16#003F1# => romdata <= X"A53F843D";
    when 16#003F2# => romdata <= X"0D0480F0";
    when 16#003F3# => romdata <= X"88519E9A";
    when 16#003F4# => romdata <= X"3F843D0D";
    when 16#003F5# => romdata <= X"0480F0A8";
    when 16#003F6# => romdata <= X"519E8F3F";
    when 16#003F7# => romdata <= X"843D0D04";
    when 16#003F8# => romdata <= X"80F0BC51";
    when 16#003F9# => romdata <= X"9E843F84";
    when 16#003FA# => romdata <= X"3D0D0480";
    when 16#003FB# => romdata <= X"F0D8519D";
    when 16#003FC# => romdata <= X"F93F843D";
    when 16#003FD# => romdata <= X"0D0480F0";
    when 16#003FE# => romdata <= X"F0519DEE";
    when 16#003FF# => romdata <= X"3F843D0D";
    when 16#00400# => romdata <= X"0480F184";
    when 16#00401# => romdata <= X"519DE33F";
    when 16#00402# => romdata <= X"843D0D04";
    when 16#00403# => romdata <= X"80F19451";
    when 16#00404# => romdata <= X"9DD83F84";
    when 16#00405# => romdata <= X"3D0D0480";
    when 16#00406# => romdata <= X"F1A8519D";
    when 16#00407# => romdata <= X"CD3F843D";
    when 16#00408# => romdata <= X"0D0480F1";
    when 16#00409# => romdata <= X"B8519DC2";
    when 16#0040A# => romdata <= X"3F843D0D";
    when 16#0040B# => romdata <= X"0480F1D0";
    when 16#0040C# => romdata <= X"519DB73F";
    when 16#0040D# => romdata <= X"843D0D04";
    when 16#0040E# => romdata <= X"80F1E451";
    when 16#0040F# => romdata <= X"9DAC3F84";
    when 16#00410# => romdata <= X"3D0D0480";
    when 16#00411# => romdata <= X"F1F4519D";
    when 16#00412# => romdata <= X"A13F843D";
    when 16#00413# => romdata <= X"0D04F73D";
    when 16#00414# => romdata <= X"0D02B305";
    when 16#00415# => romdata <= X"337C7008";
    when 16#00416# => romdata <= X"C0808006";
    when 16#00417# => romdata <= X"59545A80";
    when 16#00418# => romdata <= X"5675832B";
    when 16#00419# => romdata <= X"7707BFE0";
    when 16#0041A# => romdata <= X"80077070";
    when 16#0041B# => romdata <= X"84055208";
    when 16#0041C# => romdata <= X"71088C2A";
    when 16#0041D# => romdata <= X"BFFE8006";
    when 16#0041E# => romdata <= X"79077198";
    when 16#0041F# => romdata <= X"2A728C2A";
    when 16#00420# => romdata <= X"9FFF0673";
    when 16#00421# => romdata <= X"852A708F";
    when 16#00422# => romdata <= X"06759F06";
    when 16#00423# => romdata <= X"5651585D";
    when 16#00424# => romdata <= X"58525558";
    when 16#00425# => romdata <= X"748D3881";
    when 16#00426# => romdata <= X"16568F76";
    when 16#00427# => romdata <= X"27C3388B";
    when 16#00428# => romdata <= X"3D0D0480";
    when 16#00429# => romdata <= X"F28C519C";
    when 16#0042A# => romdata <= X"C13F7551";
    when 16#0042B# => romdata <= X"9E863F84";
    when 16#0042C# => romdata <= X"52B00851";
    when 16#0042D# => romdata <= X"9FC73F80";
    when 16#0042E# => romdata <= X"F298519C";
    when 16#0042F# => romdata <= X"AD3F7452";
    when 16#00430# => romdata <= X"88519CC9";
    when 16#00431# => romdata <= X"3F8452B0";
    when 16#00432# => romdata <= X"08519FB1";
    when 16#00433# => romdata <= X"3F80F2A0";
    when 16#00434# => romdata <= X"519C973F";
    when 16#00435# => romdata <= X"78529051";
    when 16#00436# => romdata <= X"9CB33F86";
    when 16#00437# => romdata <= X"52B00851";
    when 16#00438# => romdata <= X"9F9B3F80";
    when 16#00439# => romdata <= X"F2A8519C";
    when 16#0043A# => romdata <= X"813F7251";
    when 16#0043B# => romdata <= X"9DC63F84";
    when 16#0043C# => romdata <= X"52B00851";
    when 16#0043D# => romdata <= X"9F873F80";
    when 16#0043E# => romdata <= X"F2B0519B";
    when 16#0043F# => romdata <= X"ED3F7351";
    when 16#00440# => romdata <= X"9DB23F84";
    when 16#00441# => romdata <= X"52B00851";
    when 16#00442# => romdata <= X"9EF33F80";
    when 16#00443# => romdata <= X"F2B8519B";
    when 16#00444# => romdata <= X"D93F7752";
    when 16#00445# => romdata <= X"A0519BF5";
    when 16#00446# => romdata <= X"3F8A52B0";
    when 16#00447# => romdata <= X"08519EDD";
    when 16#00448# => romdata <= X"3F799238";
    when 16#00449# => romdata <= X"8A519BA8";
    when 16#0044A# => romdata <= X"3F811656";
    when 16#0044B# => romdata <= X"8F7627FE";
    when 16#0044C# => romdata <= X"B038FEEB";
    when 16#0044D# => romdata <= X"397881FF";
    when 16#0044E# => romdata <= X"06527451";
    when 16#0044F# => romdata <= X"FB973F8A";
    when 16#00450# => romdata <= X"519B8D3F";
    when 16#00451# => romdata <= X"E439F83D";
    when 16#00452# => romdata <= X"0D02AB05";
    when 16#00453# => romdata <= X"33598056";
    when 16#00454# => romdata <= X"75852BE0";
    when 16#00455# => romdata <= X"9011E080";
    when 16#00456# => romdata <= X"12087098";
    when 16#00457# => romdata <= X"2A718C2A";
    when 16#00458# => romdata <= X"9FFF0672";
    when 16#00459# => romdata <= X"852A708F";
    when 16#0045A# => romdata <= X"06749F06";
    when 16#0045B# => romdata <= X"5551585B";
    when 16#0045C# => romdata <= X"53565955";
    when 16#0045D# => romdata <= X"74802E81";
    when 16#0045E# => romdata <= X"A13875BF";
    when 16#0045F# => romdata <= X"2681A938";
    when 16#00460# => romdata <= X"80F2C051";
    when 16#00461# => romdata <= X"9AE43F75";
    when 16#00462# => romdata <= X"519CA93F";
    when 16#00463# => romdata <= X"8652B008";
    when 16#00464# => romdata <= X"519DEA3F";
    when 16#00465# => romdata <= X"80F29851";
    when 16#00466# => romdata <= X"9AD03F74";
    when 16#00467# => romdata <= X"5288519A";
    when 16#00468# => romdata <= X"EC3F8452";
    when 16#00469# => romdata <= X"B008519D";
    when 16#0046A# => romdata <= X"D43F80F2";
    when 16#0046B# => romdata <= X"A0519ABA";
    when 16#0046C# => romdata <= X"3F765290";
    when 16#0046D# => romdata <= X"519AD63F";
    when 16#0046E# => romdata <= X"8652B008";
    when 16#0046F# => romdata <= X"519DBE3F";
    when 16#00470# => romdata <= X"80F2A851";
    when 16#00471# => romdata <= X"9AA43F72";
    when 16#00472# => romdata <= X"519BE93F";
    when 16#00473# => romdata <= X"8452B008";
    when 16#00474# => romdata <= X"519DAA3F";
    when 16#00475# => romdata <= X"80F2B051";
    when 16#00476# => romdata <= X"9A903F73";
    when 16#00477# => romdata <= X"519BD53F";
    when 16#00478# => romdata <= X"8452B008";
    when 16#00479# => romdata <= X"519D963F";
    when 16#0047A# => romdata <= X"80F2B851";
    when 16#0047B# => romdata <= X"99FC3F77";
    when 16#0047C# => romdata <= X"08C08080";
    when 16#0047D# => romdata <= X"0652A051";
    when 16#0047E# => romdata <= X"9A933F8A";
    when 16#0047F# => romdata <= X"52B00851";
    when 16#00480# => romdata <= X"9CFB3F78";
    when 16#00481# => romdata <= X"81AC388A";
    when 16#00482# => romdata <= X"5199C53F";
    when 16#00483# => romdata <= X"80537481";
    when 16#00484# => romdata <= X"2E81D938";
    when 16#00485# => romdata <= X"76862E81";
    when 16#00486# => romdata <= X"B5388116";
    when 16#00487# => romdata <= X"5680FF76";
    when 16#00488# => romdata <= X"27FEAD38";
    when 16#00489# => romdata <= X"8A3D0D04";
    when 16#0048A# => romdata <= X"80F2C851";
    when 16#0048B# => romdata <= X"99BC3FC0";
    when 16#0048C# => romdata <= X"16519B80";
    when 16#0048D# => romdata <= X"3F8652B0";
    when 16#0048E# => romdata <= X"08519CC1";
    when 16#0048F# => romdata <= X"3F80F298";
    when 16#00490# => romdata <= X"5199A73F";
    when 16#00491# => romdata <= X"74528851";
    when 16#00492# => romdata <= X"99C33F84";
    when 16#00493# => romdata <= X"52B00851";
    when 16#00494# => romdata <= X"9CAB3F80";
    when 16#00495# => romdata <= X"F2A05199";
    when 16#00496# => romdata <= X"913F7652";
    when 16#00497# => romdata <= X"905199AD";
    when 16#00498# => romdata <= X"3F8652B0";
    when 16#00499# => romdata <= X"08519C95";
    when 16#0049A# => romdata <= X"3F80F2A8";
    when 16#0049B# => romdata <= X"5198FB3F";
    when 16#0049C# => romdata <= X"72519AC0";
    when 16#0049D# => romdata <= X"3F8452B0";
    when 16#0049E# => romdata <= X"08519C81";
    when 16#0049F# => romdata <= X"3F80F2B0";
    when 16#004A0# => romdata <= X"5198E73F";
    when 16#004A1# => romdata <= X"73519AAC";
    when 16#004A2# => romdata <= X"3F8452B0";
    when 16#004A3# => romdata <= X"08519BED";
    when 16#004A4# => romdata <= X"3F80F2B8";
    when 16#004A5# => romdata <= X"5198D33F";
    when 16#004A6# => romdata <= X"7708C080";
    when 16#004A7# => romdata <= X"800652A0";
    when 16#004A8# => romdata <= X"5198EA3F";
    when 16#004A9# => romdata <= X"8A52B008";
    when 16#004AA# => romdata <= X"519BD23F";
    when 16#004AB# => romdata <= X"78802EFE";
    when 16#004AC# => romdata <= X"D6387681";
    when 16#004AD# => romdata <= X"FF065274";
    when 16#004AE# => romdata <= X"51F89A3F";
    when 16#004AF# => romdata <= X"8A519890";
    when 16#004B0# => romdata <= X"3F805374";
    when 16#004B1# => romdata <= X"812E0981";
    when 16#004B2# => romdata <= X"06FEC938";
    when 16#004B3# => romdata <= X"9F397281";
    when 16#004B4# => romdata <= X"06577680";
    when 16#004B5# => romdata <= X"2EFEC338";
    when 16#004B6# => romdata <= X"78527751";
    when 16#004B7# => romdata <= X"FAF03F81";
    when 16#004B8# => romdata <= X"165680FF";
    when 16#004B9# => romdata <= X"7627FCE8";
    when 16#004BA# => romdata <= X"38FEB939";
    when 16#004BB# => romdata <= X"74537686";
    when 16#004BC# => romdata <= X"2E098106";
    when 16#004BD# => romdata <= X"FEA438D6";
    when 16#004BE# => romdata <= X"39803D0D";
    when 16#004BF# => romdata <= X"80FC8808";
    when 16#004C0# => romdata <= X"51B1710C";
    when 16#004C1# => romdata <= X"81800B84";
    when 16#004C2# => romdata <= X"120C823D";
    when 16#004C3# => romdata <= X"0D04FE3D";
    when 16#004C4# => romdata <= X"0D740284";
    when 16#004C5# => romdata <= X"05970533";
    when 16#004C6# => romdata <= X"0288059B";
    when 16#004C7# => romdata <= X"05338813";
    when 16#004C8# => romdata <= X"0C8C120C";
    when 16#004C9# => romdata <= X"538C1308";
    when 16#004CA# => romdata <= X"70812A81";
    when 16#004CB# => romdata <= X"06515271";
    when 16#004CC# => romdata <= X"F4388C13";
    when 16#004CD# => romdata <= X"087081FF";
    when 16#004CE# => romdata <= X"06B00C51";
    when 16#004CF# => romdata <= X"843D0D04";
    when 16#004D0# => romdata <= X"FB3D0D80";
    when 16#004D1# => romdata <= X"0B80F5F4";
    when 16#004D2# => romdata <= X"5256979E";
    when 16#004D3# => romdata <= X"3F755574";
    when 16#004D4# => romdata <= X"105381D0";
    when 16#004D5# => romdata <= X"5280FC88";
    when 16#004D6# => romdata <= X"0851FFB2";
    when 16#004D7# => romdata <= X"3FB00887";
    when 16#004D8# => romdata <= X"2A708106";
    when 16#004D9# => romdata <= X"51547380";
    when 16#004DA# => romdata <= X"2E993881";
    when 16#004DB# => romdata <= X"157081FF";
    when 16#004DC# => romdata <= X"0670982B";
    when 16#004DD# => romdata <= X"52565473";
    when 16#004DE# => romdata <= X"8025D438";
    when 16#004DF# => romdata <= X"75B00C87";
    when 16#004E0# => romdata <= X"3D0D0480";
    when 16#004E1# => romdata <= X"F6805196";
    when 16#004E2# => romdata <= X"E13F7452";
    when 16#004E3# => romdata <= X"885196FD";
    when 16#004E4# => romdata <= X"3F80F68C";
    when 16#004E5# => romdata <= X"5196D33F";
    when 16#004E6# => romdata <= X"81167083";
    when 16#004E7# => romdata <= X"FFFF0681";
    when 16#004E8# => romdata <= X"177081FF";
    when 16#004E9# => romdata <= X"0670982B";
    when 16#004EA# => romdata <= X"52585257";
    when 16#004EB# => romdata <= X"54738025";
    when 16#004EC# => romdata <= X"FF9D38C8";
    when 16#004ED# => romdata <= X"39F33D0D";
    when 16#004EE# => romdata <= X"7F028405";
    when 16#004EF# => romdata <= X"80C30533";
    when 16#004F0# => romdata <= X"02880580";
    when 16#004F1# => romdata <= X"C6052280";
    when 16#004F2# => romdata <= X"F69C545B";
    when 16#004F3# => romdata <= X"5558969A";
    when 16#004F4# => romdata <= X"3F785197";
    when 16#004F5# => romdata <= X"DF3F80F6";
    when 16#004F6# => romdata <= X"A851968E";
    when 16#004F7# => romdata <= X"3F735288";
    when 16#004F8# => romdata <= X"5196AA3F";
    when 16#004F9# => romdata <= X"80EBEC51";
    when 16#004FA# => romdata <= X"96803F80";
    when 16#004FB# => romdata <= X"57767927";
    when 16#004FC# => romdata <= X"81913873";
    when 16#004FD# => romdata <= X"108E3D5C";
    when 16#004FE# => romdata <= X"5A795381";
    when 16#004FF# => romdata <= X"90527751";
    when 16#00500# => romdata <= X"FE8C3F76";
    when 16#00501# => romdata <= X"882A5390";
    when 16#00502# => romdata <= X"527751FE";
    when 16#00503# => romdata <= X"813F7681";
    when 16#00504# => romdata <= X"FF065390";
    when 16#00505# => romdata <= X"527751FD";
    when 16#00506# => romdata <= X"F53F811A";
    when 16#00507# => romdata <= X"53819052";
    when 16#00508# => romdata <= X"7751FDEA";
    when 16#00509# => romdata <= X"3F805380";
    when 16#0050A# => romdata <= X"E0527751";
    when 16#0050B# => romdata <= X"FDE03FB0";
    when 16#0050C# => romdata <= X"08872A81";
    when 16#0050D# => romdata <= X"0654738A";
    when 16#0050E# => romdata <= X"38881808";
    when 16#0050F# => romdata <= X"7081FF06";
    when 16#00510# => romdata <= X"5D567B81";
    when 16#00511# => romdata <= X"FF0680F8";
    when 16#00512# => romdata <= X"CC525695";
    when 16#00513# => romdata <= X"9D3F7552";
    when 16#00514# => romdata <= X"885195B9";
    when 16#00515# => romdata <= X"3F80EDFC";
    when 16#00516# => romdata <= X"51958F3F";
    when 16#00517# => romdata <= X"E0165480";
    when 16#00518# => romdata <= X"DF7427B6";
    when 16#00519# => romdata <= X"38768706";
    when 16#0051A# => romdata <= X"701C5755";
    when 16#0051B# => romdata <= X"A0763474";
    when 16#0051C# => romdata <= X"872EB938";
    when 16#0051D# => romdata <= X"81177083";
    when 16#0051E# => romdata <= X"FFFF0658";
    when 16#0051F# => romdata <= X"55787726";
    when 16#00520# => romdata <= X"FEF73880";
    when 16#00521# => romdata <= X"E00B8C19";
    when 16#00522# => romdata <= X"0C8C1808";
    when 16#00523# => romdata <= X"70812A81";
    when 16#00524# => romdata <= X"06585A76";
    when 16#00525# => romdata <= X"F4388F3D";
    when 16#00526# => romdata <= X"0D047687";
    when 16#00527# => romdata <= X"06701C55";
    when 16#00528# => romdata <= X"55757434";
    when 16#00529# => romdata <= X"74872E09";
    when 16#0052A# => romdata <= X"8106C938";
    when 16#0052B# => romdata <= X"7A5194BA";
    when 16#0052C# => romdata <= X"3F8A5194";
    when 16#0052D# => romdata <= X"9B3F8117";
    when 16#0052E# => romdata <= X"7083FFFF";
    when 16#0052F# => romdata <= X"06585578";
    when 16#00530# => romdata <= X"7726FEB5";
    when 16#00531# => romdata <= X"38FFBC39";
    when 16#00532# => romdata <= X"FB3D0D81";
    when 16#00533# => romdata <= X"51EEFC3F";
    when 16#00534# => romdata <= X"8251F0A9";
    when 16#00535# => romdata <= X"3FB00881";
    when 16#00536# => romdata <= X"FF065683";
    when 16#00537# => romdata <= X"51EEEC3F";
    when 16#00538# => romdata <= X"B00883FF";
    when 16#00539# => romdata <= X"FF0680FC";
    when 16#0053A# => romdata <= X"88085654";
    when 16#0053B# => romdata <= X"73843881";
    when 16#0053C# => romdata <= X"80547353";
    when 16#0053D# => romdata <= X"75527451";
    when 16#0053E# => romdata <= X"FDBB3F73";
    when 16#0053F# => romdata <= X"B00C873D";
    when 16#00540# => romdata <= X"0D04FB3D";
    when 16#00541# => romdata <= X"0D8151EF";
    when 16#00542# => romdata <= X"F43FB008";
    when 16#00543# => romdata <= X"538251EF";
    when 16#00544# => romdata <= X"EC3FB008";
    when 16#00545# => romdata <= X"56B00883";
    when 16#00546# => romdata <= X"38905672";
    when 16#00547# => romdata <= X"FC065575";
    when 16#00548# => romdata <= X"812E80F1";
    when 16#00549# => romdata <= X"38805473";
    when 16#0054A# => romdata <= X"7627AA38";
    when 16#0054B# => romdata <= X"73830653";
    when 16#0054C# => romdata <= X"72802EAE";
    when 16#0054D# => romdata <= X"3880F8CC";
    when 16#0054E# => romdata <= X"5193AF3F";
    when 16#0054F# => romdata <= X"74708405";
    when 16#00550# => romdata <= X"560852A0";
    when 16#00551# => romdata <= X"5193C63F";
    when 16#00552# => romdata <= X"A0519384";
    when 16#00553# => romdata <= X"3F811454";
    when 16#00554# => romdata <= X"757426D8";
    when 16#00555# => romdata <= X"388A5192";
    when 16#00556# => romdata <= X"F73F800B";
    when 16#00557# => romdata <= X"B00C873D";
    when 16#00558# => romdata <= X"0D0480F6";
    when 16#00559# => romdata <= X"C4519382";
    when 16#0055A# => romdata <= X"3F7452A0";
    when 16#0055B# => romdata <= X"51939E3F";
    when 16#0055C# => romdata <= X"80F88C51";
    when 16#0055D# => romdata <= X"92F43F80";
    when 16#0055E# => romdata <= X"F8CC5192";
    when 16#0055F# => romdata <= X"ED3F7470";
    when 16#00560# => romdata <= X"84055608";
    when 16#00561# => romdata <= X"52A05193";
    when 16#00562# => romdata <= X"843FA051";
    when 16#00563# => romdata <= X"92C23F81";
    when 16#00564# => romdata <= X"1454FFBC";
    when 16#00565# => romdata <= X"3980F8CC";
    when 16#00566# => romdata <= X"5192CF3F";
    when 16#00567# => romdata <= X"740852A0";
    when 16#00568# => romdata <= X"5192EA3F";
    when 16#00569# => romdata <= X"8A5192A8";
    when 16#0056A# => romdata <= X"3F800BB0";
    when 16#0056B# => romdata <= X"0C873D0D";
    when 16#0056C# => romdata <= X"04FC3D0D";
    when 16#0056D# => romdata <= X"8151EEC5";
    when 16#0056E# => romdata <= X"3FB00852";
    when 16#0056F# => romdata <= X"8251ED8B";
    when 16#00570# => romdata <= X"3FB00881";
    when 16#00571# => romdata <= X"FF067256";
    when 16#00572# => romdata <= X"53835472";
    when 16#00573# => romdata <= X"802EA138";
    when 16#00574# => romdata <= X"7351EEA9";
    when 16#00575# => romdata <= X"3F811470";
    when 16#00576# => romdata <= X"81FF06FF";
    when 16#00577# => romdata <= X"157081FF";
    when 16#00578# => romdata <= X"06B00879";
    when 16#00579# => romdata <= X"7084055B";
    when 16#0057A# => romdata <= X"0C565255";
    when 16#0057B# => romdata <= X"5272E138";
    when 16#0057C# => romdata <= X"72B00C86";
    when 16#0057D# => romdata <= X"3D0D0480";
    when 16#0057E# => romdata <= X"3D0D8C51";
    when 16#0057F# => romdata <= X"91D23F80";
    when 16#00580# => romdata <= X"0BB00C82";
    when 16#00581# => romdata <= X"3D0D0480";
    when 16#00582# => romdata <= X"3D0D80FC";
    when 16#00583# => romdata <= X"980851F8";
    when 16#00584# => romdata <= X"BB9586A1";
    when 16#00585# => romdata <= X"710C810B";
    when 16#00586# => romdata <= X"B00C823D";
    when 16#00587# => romdata <= X"0D04803D";
    when 16#00588# => romdata <= X"0D8151EC";
    when 16#00589# => romdata <= X"A63FB008";
    when 16#0058A# => romdata <= X"81FF0651";
    when 16#0058B# => romdata <= X"F6983F80";
    when 16#0058C# => romdata <= X"0BB00C82";
    when 16#0058D# => romdata <= X"3D0D04FF";
    when 16#0058E# => romdata <= X"3D0D80FB";
    when 16#0058F# => romdata <= X"E408A011";
    when 16#00590# => romdata <= X"087080FF";
    when 16#00591# => romdata <= X"0A06A013";
    when 16#00592# => romdata <= X"0C5252BB";
    when 16#00593# => romdata <= X"C880800B";
    when 16#00594# => romdata <= X"A0130C83";
    when 16#00595# => romdata <= X"3D0D04FF";
    when 16#00596# => romdata <= X"3D0D028F";
    when 16#00597# => romdata <= X"05337098";
    when 16#00598# => romdata <= X"2B80FBE4";
    when 16#00599# => romdata <= X"0852B012";
    when 16#0059A# => romdata <= X"0C51833D";
    when 16#0059B# => romdata <= X"0D04FF3D";
    when 16#0059C# => romdata <= X"0D80FBE4";
    when 16#0059D# => romdata <= X"0852A412";
    when 16#0059E# => romdata <= X"0870892A";
    when 16#0059F# => romdata <= X"70810651";
    when 16#005A0# => romdata <= X"51517080";
    when 16#005A1# => romdata <= X"2EF038B4";
    when 16#005A2# => romdata <= X"12087090";
    when 16#005A3# => romdata <= X"2AB00C51";
    when 16#005A4# => romdata <= X"833D0D04";
    when 16#005A5# => romdata <= X"F83D0D7A";
    when 16#005A6# => romdata <= X"7C5755FF";
    when 16#005A7# => romdata <= X"9A3F80FC";
    when 16#005A8# => romdata <= X"8C088411";
    when 16#005A9# => romdata <= X"08828080";
    when 16#005AA# => romdata <= X"0784120C";
    when 16#005AB# => romdata <= X"841108FD";
    when 16#005AC# => romdata <= X"FFFF0684";
    when 16#005AD# => romdata <= X"120C8411";
    when 16#005AE# => romdata <= X"08818080";
    when 16#005AF# => romdata <= X"0784120C";
    when 16#005B0# => romdata <= X"841108FE";
    when 16#005B1# => romdata <= X"FFFF0684";
    when 16#005B2# => romdata <= X"120C5390";
    when 16#005B3# => romdata <= X"0B893D34";
    when 16#005B4# => romdata <= X"94028405";
    when 16#005B5# => romdata <= X"9D053480";
    when 16#005B6# => romdata <= X"0284059E";
    when 16#005B7# => romdata <= X"053480E1";
    when 16#005B8# => romdata <= X"0284059F";
    when 16#005B9# => romdata <= X"0534883D";
    when 16#005BA# => romdata <= X"80FBE408";
    when 16#005BB# => romdata <= X"5457A413";
    when 16#005BC# => romdata <= X"0870882A";
    when 16#005BD# => romdata <= X"81065152";
    when 16#005BE# => romdata <= X"71802EF2";
    when 16#005BF# => romdata <= X"388751FE";
    when 16#005C0# => romdata <= X"D63F800B";
    when 16#005C1# => romdata <= X"80F6CF33";
    when 16#005C2# => romdata <= X"53537272";
    when 16#005C3# => romdata <= X"27993871";
    when 16#005C4# => romdata <= X"54761370";
    when 16#005C5# => romdata <= X"335252FE";
    when 16#005C6# => romdata <= X"BE3F8113";
    when 16#005C7# => romdata <= X"7081FF06";
    when 16#005C8# => romdata <= X"54527373";
    when 16#005C9# => romdata <= X"26EB38FE";
    when 16#005CA# => romdata <= X"C53F800B";
    when 16#005CB# => romdata <= X"80F6CF33";
    when 16#005CC# => romdata <= X"53537272";
    when 16#005CD# => romdata <= X"27933871";
    when 16#005CE# => romdata <= X"54FEB33F";
    when 16#005CF# => romdata <= X"81137081";
    when 16#005D0# => romdata <= X"FF065452";
    when 16#005D1# => romdata <= X"737326F1";
    when 16#005D2# => romdata <= X"3874882A";
    when 16#005D3# => romdata <= X"5473893D";
    when 16#005D4# => romdata <= X"34740284";
    when 16#005D5# => romdata <= X"059D0534";
    when 16#005D6# => romdata <= X"74882B76";
    when 16#005D7# => romdata <= X"982A0752";
    when 16#005D8# => romdata <= X"71028405";
    when 16#005D9# => romdata <= X"9E053474";
    when 16#005DA# => romdata <= X"902B7690";
    when 16#005DB# => romdata <= X"2A075473";
    when 16#005DC# => romdata <= X"0284059F";
    when 16#005DD# => romdata <= X"05347498";
    when 16#005DE# => romdata <= X"2B76882A";
    when 16#005DF# => romdata <= X"0753728A";
    when 16#005E0# => romdata <= X"3D347502";
    when 16#005E1# => romdata <= X"8405A105";
    when 16#005E2# => romdata <= X"3480FBE4";
    when 16#005E3# => romdata <= X"0853A413";
    when 16#005E4# => romdata <= X"0870882A";
    when 16#005E5# => romdata <= X"81065652";
    when 16#005E6# => romdata <= X"74802EF2";
    when 16#005E7# => romdata <= X"388251FD";
    when 16#005E8# => romdata <= X"B63F800B";
    when 16#005E9# => romdata <= X"80F6CA33";
    when 16#005EA# => romdata <= X"53537272";
    when 16#005EB# => romdata <= X"27993871";
    when 16#005EC# => romdata <= X"54761370";
    when 16#005ED# => romdata <= X"335256FD";
    when 16#005EE# => romdata <= X"9E3F8113";
    when 16#005EF# => romdata <= X"7081FF06";
    when 16#005F0# => romdata <= X"54557373";
    when 16#005F1# => romdata <= X"26EB38FD";
    when 16#005F2# => romdata <= X"A53F800B";
    when 16#005F3# => romdata <= X"80F6CA33";
    when 16#005F4# => romdata <= X"53537272";
    when 16#005F5# => romdata <= X"27933871";
    when 16#005F6# => romdata <= X"54FD933F";
    when 16#005F7# => romdata <= X"81137081";
    when 16#005F8# => romdata <= X"FF065452";
    when 16#005F9# => romdata <= X"737326F1";
    when 16#005FA# => romdata <= X"388A0B89";
    when 16#005FB# => romdata <= X"3D34FF8C";
    when 16#005FC# => romdata <= X"0284059D";
    when 16#005FD# => romdata <= X"053480FB";
    when 16#005FE# => romdata <= X"E40853A4";
    when 16#005FF# => romdata <= X"13087088";
    when 16#00600# => romdata <= X"2A810655";
    when 16#00601# => romdata <= X"5673802E";
    when 16#00602# => romdata <= X"F2388851";
    when 16#00603# => romdata <= X"FCC93F80";
    when 16#00604# => romdata <= X"0B80F6D0";
    when 16#00605# => romdata <= X"33535372";
    when 16#00606# => romdata <= X"72279938";
    when 16#00607# => romdata <= X"71547613";
    when 16#00608# => romdata <= X"70335255";
    when 16#00609# => romdata <= X"FCB13F81";
    when 16#0060A# => romdata <= X"137081FF";
    when 16#0060B# => romdata <= X"06545273";
    when 16#0060C# => romdata <= X"7326EB38";
    when 16#0060D# => romdata <= X"FCB83F80";
    when 16#0060E# => romdata <= X"0B80F6D0";
    when 16#0060F# => romdata <= X"33535372";
    when 16#00610# => romdata <= X"72279338";
    when 16#00611# => romdata <= X"7154FCA6";
    when 16#00612# => romdata <= X"3F811370";
    when 16#00613# => romdata <= X"81FF0654";
    when 16#00614# => romdata <= X"56737326";
    when 16#00615# => romdata <= X"F1388A0B";
    when 16#00616# => romdata <= X"893D34FF";
    when 16#00617# => romdata <= X"8C028405";
    when 16#00618# => romdata <= X"9D053480";
    when 16#00619# => romdata <= X"FBE40853";
    when 16#0061A# => romdata <= X"A4130870";
    when 16#0061B# => romdata <= X"882A8106";
    when 16#0061C# => romdata <= X"55557380";
    when 16#0061D# => romdata <= X"2EF23889";
    when 16#0061E# => romdata <= X"51FBDC3F";
    when 16#0061F# => romdata <= X"800B80F6";
    when 16#00620# => romdata <= X"D1335353";
    when 16#00621# => romdata <= X"72722799";
    when 16#00622# => romdata <= X"38715476";
    when 16#00623# => romdata <= X"13703352";
    when 16#00624# => romdata <= X"52FBC43F";
    when 16#00625# => romdata <= X"81137081";
    when 16#00626# => romdata <= X"FF065456";
    when 16#00627# => romdata <= X"737326EB";
    when 16#00628# => romdata <= X"38FBCB3F";
    when 16#00629# => romdata <= X"800B80F6";
    when 16#0062A# => romdata <= X"D1335353";
    when 16#0062B# => romdata <= X"72722793";
    when 16#0062C# => romdata <= X"387154FB";
    when 16#0062D# => romdata <= X"B93F8113";
    when 16#0062E# => romdata <= X"7081FF06";
    when 16#0062F# => romdata <= X"54577373";
    when 16#00630# => romdata <= X"26F13880";
    when 16#00631# => romdata <= X"FC8C0884";
    when 16#00632# => romdata <= X"110880C0";
    when 16#00633# => romdata <= X"80078412";
    when 16#00634# => romdata <= X"0C841108";
    when 16#00635# => romdata <= X"FFBFFF06";
    when 16#00636# => romdata <= X"84120C54";
    when 16#00637# => romdata <= X"800BB00C";
    when 16#00638# => romdata <= X"8A3D0D04";
    when 16#00639# => romdata <= X"F83D0D02";
    when 16#0063A# => romdata <= X"AB053389";
    when 16#0063B# => romdata <= X"3D80FBE4";
    when 16#0063C# => romdata <= X"08565856";
    when 16#0063D# => romdata <= X"A4140870";
    when 16#0063E# => romdata <= X"882A8106";
    when 16#0063F# => romdata <= X"51537280";
    when 16#00640# => romdata <= X"2EF23875";
    when 16#00641# => romdata <= X"81800751";
    when 16#00642# => romdata <= X"FACD3F80";
    when 16#00643# => romdata <= X"0B80F6C8";
    when 16#00644# => romdata <= X"17335454";
    when 16#00645# => romdata <= X"73732795";
    when 16#00646# => romdata <= X"38725580";
    when 16#00647# => romdata <= X"51FAB83F";
    when 16#00648# => romdata <= X"81147081";
    when 16#00649# => romdata <= X"FF065553";
    when 16#0064A# => romdata <= X"747426EF";
    when 16#0064B# => romdata <= X"38FABF3F";
    when 16#0064C# => romdata <= X"800B80F6";
    when 16#0064D# => romdata <= X"C8173370";
    when 16#0064E# => romdata <= X"81FF0655";
    when 16#0064F# => romdata <= X"57547373";
    when 16#00650# => romdata <= X"279A3872";
    when 16#00651# => romdata <= X"55761453";
    when 16#00652# => romdata <= X"FAA43FB0";
    when 16#00653# => romdata <= X"08733481";
    when 16#00654# => romdata <= X"147081FF";
    when 16#00655# => romdata <= X"06555374";
    when 16#00656# => romdata <= X"7426EA38";
    when 16#00657# => romdata <= X"7581FF06";
    when 16#00658# => romdata <= X"80F8CC52";
    when 16#00659# => romdata <= X"558B833F";
    when 16#0065A# => romdata <= X"80547375";
    when 16#0065B# => romdata <= X"27993873";
    when 16#0065C# => romdata <= X"17703353";
    when 16#0065D# => romdata <= X"5388518B";
    when 16#0065E# => romdata <= X"943F8114";
    when 16#0065F# => romdata <= X"7081FF06";
    when 16#00660# => romdata <= X"55567474";
    when 16#00661# => romdata <= X"26E9388A";
    when 16#00662# => romdata <= X"518AC53F";
    when 16#00663# => romdata <= X"8A3D0D04";
    when 16#00664# => romdata <= X"FE3D0D80";
    when 16#00665# => romdata <= X"FC8C0884";
    when 16#00666# => romdata <= X"11087081";
    when 16#00667# => romdata <= X"80800784";
    when 16#00668# => romdata <= X"130C5484";
    when 16#00669# => romdata <= X"110870FE";
    when 16#0066A# => romdata <= X"FFFF0684";
    when 16#0066B# => romdata <= X"130C5452";
    when 16#0066C# => romdata <= X"F9853F80";
    when 16#0066D# => romdata <= X"F6D4518A";
    when 16#0066E# => romdata <= X"B13F8751";
    when 16#0066F# => romdata <= X"FEA63F80";
    when 16#00670# => romdata <= X"F6E4518A";
    when 16#00671# => romdata <= X"A53F8251";
    when 16#00672# => romdata <= X"FE9A3F80";
    when 16#00673# => romdata <= X"F6F4518A";
    when 16#00674# => romdata <= X"993F8551";
    when 16#00675# => romdata <= X"FE8E3F80";
    when 16#00676# => romdata <= X"F784518A";
    when 16#00677# => romdata <= X"8D3F8651";
    when 16#00678# => romdata <= X"FE823F80";
    when 16#00679# => romdata <= X"F794518A";
    when 16#0067A# => romdata <= X"813F8851";
    when 16#0067B# => romdata <= X"FDF63F80";
    when 16#0067C# => romdata <= X"F7A45189";
    when 16#0067D# => romdata <= X"F53F8951";
    when 16#0067E# => romdata <= X"FDEA3F80";
    when 16#0067F# => romdata <= X"0BB00C84";
    when 16#00680# => romdata <= X"3D0D04FE";
    when 16#00681# => romdata <= X"3D0D80FC";
    when 16#00682# => romdata <= X"8C088411";
    when 16#00683# => romdata <= X"08820A07";
    when 16#00684# => romdata <= X"84120C70";
    when 16#00685# => romdata <= X"0870902A";
    when 16#00686# => romdata <= X"84130870";
    when 16#00687# => romdata <= X"FD0A0684";
    when 16#00688# => romdata <= X"150C5481";
    when 16#00689# => romdata <= X"FFFF06B0";
    when 16#0068A# => romdata <= X"0C535384";
    when 16#0068B# => romdata <= X"3D0D04FF";
    when 16#0068C# => romdata <= X"3D0D80FB";
    when 16#0068D# => romdata <= X"EC087008";
    when 16#0068E# => romdata <= X"7081FF06";
    when 16#0068F# => romdata <= X"51515271";
    when 16#00690# => romdata <= X"89268C38";
    when 16#00691# => romdata <= X"71101080";
    when 16#00692# => romdata <= X"F8F40552";
    when 16#00693# => romdata <= X"71080480";
    when 16#00694# => romdata <= X"F7B45189";
    when 16#00695# => romdata <= X"953F8A51";
    when 16#00696# => romdata <= X"88F63F80";
    when 16#00697# => romdata <= X"0BB00C83";
    when 16#00698# => romdata <= X"3D0D0480";
    when 16#00699# => romdata <= X"E7E85189";
    when 16#0069A# => romdata <= X"813F8A51";
    when 16#0069B# => romdata <= X"88E23F80";
    when 16#0069C# => romdata <= X"0BB00C83";
    when 16#0069D# => romdata <= X"3D0D0480";
    when 16#0069E# => romdata <= X"F7BC5188";
    when 16#0069F# => romdata <= X"ED3F8A51";
    when 16#006A0# => romdata <= X"88CE3F80";
    when 16#006A1# => romdata <= X"0BB00C83";
    when 16#006A2# => romdata <= X"3D0D0480";
    when 16#006A3# => romdata <= X"F7C45188";
    when 16#006A4# => romdata <= X"D93F8A51";
    when 16#006A5# => romdata <= X"88BA3F80";
    when 16#006A6# => romdata <= X"0BB00C83";
    when 16#006A7# => romdata <= X"3D0D0480";
    when 16#006A8# => romdata <= X"F7D05188";
    when 16#006A9# => romdata <= X"C53F8A51";
    when 16#006AA# => romdata <= X"88A63F80";
    when 16#006AB# => romdata <= X"0BB00C83";
    when 16#006AC# => romdata <= X"3D0D0480";
    when 16#006AD# => romdata <= X"F7D85188";
    when 16#006AE# => romdata <= X"B13F8A51";
    when 16#006AF# => romdata <= X"88923F80";
    when 16#006B0# => romdata <= X"0BB00C83";
    when 16#006B1# => romdata <= X"3D0D0480";
    when 16#006B2# => romdata <= X"F7E05188";
    when 16#006B3# => romdata <= X"9D3F8A51";
    when 16#006B4# => romdata <= X"87FE3F80";
    when 16#006B5# => romdata <= X"0BB00C83";
    when 16#006B6# => romdata <= X"3D0D0480";
    when 16#006B7# => romdata <= X"F7E85188";
    when 16#006B8# => romdata <= X"893F8A51";
    when 16#006B9# => romdata <= X"87EA3F80";
    when 16#006BA# => romdata <= X"0BB00C83";
    when 16#006BB# => romdata <= X"3D0D0480";
    when 16#006BC# => romdata <= X"F7F05187";
    when 16#006BD# => romdata <= X"F53F8A51";
    when 16#006BE# => romdata <= X"87D63F80";
    when 16#006BF# => romdata <= X"0BB00C83";
    when 16#006C0# => romdata <= X"3D0D0480";
    when 16#006C1# => romdata <= X"F7F85187";
    when 16#006C2# => romdata <= X"E13F8A51";
    when 16#006C3# => romdata <= X"87C23F80";
    when 16#006C4# => romdata <= X"0BB00C83";
    when 16#006C5# => romdata <= X"3D0D04FE";
    when 16#006C6# => romdata <= X"3D0D80FB";
    when 16#006C7# => romdata <= X"EC088411";
    when 16#006C8# => romdata <= X"0880F880";
    when 16#006C9# => romdata <= X"53545287";
    when 16#006CA# => romdata <= X"C13F7282";
    when 16#006CB# => romdata <= X"2A810651";
    when 16#006CC# => romdata <= X"89823F80";
    when 16#006CD# => romdata <= X"F8905187";
    when 16#006CE# => romdata <= X"B13F7281";
    when 16#006CF# => romdata <= X"2A810651";
    when 16#006D0# => romdata <= X"88F23F80";
    when 16#006D1# => romdata <= X"F8A45187";
    when 16#006D2# => romdata <= X"A13F7281";
    when 16#006D3# => romdata <= X"065188E4";
    when 16#006D4# => romdata <= X"3F8A5186";
    when 16#006D5# => romdata <= X"FB3F72B0";
    when 16#006D6# => romdata <= X"0C843D0D";
    when 16#006D7# => romdata <= X"04FE3D0D";
    when 16#006D8# => romdata <= X"02930533";
    when 16#006D9# => romdata <= X"02840597";
    when 16#006DA# => romdata <= X"053380FB";
    when 16#006DB# => romdata <= X"EC085553";
    when 16#006DC# => romdata <= X"5180730C";
    when 16#006DD# => romdata <= X"7688140C";
    when 16#006DE# => romdata <= X"70832B72";
    when 16#006DF# => romdata <= X"078C140C";
    when 16#006E0# => romdata <= X"72085170";
    when 16#006E1# => romdata <= X"FB3870B0";
    when 16#006E2# => romdata <= X"0C843D0D";
    when 16#006E3# => romdata <= X"04FE3D0D";
    when 16#006E4# => romdata <= X"80F8B851";
    when 16#006E5# => romdata <= X"86D43F80";
    when 16#006E6# => romdata <= X"FBEC08A0";
    when 16#006E7# => romdata <= X"11085353";
    when 16#006E8# => romdata <= X"A05186E9";
    when 16#006E9# => romdata <= X"3F80FBEC";
    when 16#006EA# => romdata <= X"08A41108";
    when 16#006EB# => romdata <= X"5353A051";
    when 16#006EC# => romdata <= X"86DB3F80";
    when 16#006ED# => romdata <= X"F8D05186";
    when 16#006EE# => romdata <= X"B13F80FB";
    when 16#006EF# => romdata <= X"EC08A811";
    when 16#006F0# => romdata <= X"085353A0";
    when 16#006F1# => romdata <= X"5186C63F";
    when 16#006F2# => romdata <= X"80FBEC08";
    when 16#006F3# => romdata <= X"AC110853";
    when 16#006F4# => romdata <= X"53A05186";
    when 16#006F5# => romdata <= X"B83F8A51";
    when 16#006F6# => romdata <= X"85F63F80";
    when 16#006F7# => romdata <= X"0BB00C84";
    when 16#006F8# => romdata <= X"3D0D04FC";
    when 16#006F9# => romdata <= X"3D0D80FB";
    when 16#006FA# => romdata <= X"EC089C11";
    when 16#006FB# => romdata <= X"087081FF";
    when 16#006FC# => romdata <= X"0680F8E8";
    when 16#006FD# => romdata <= X"54575353";
    when 16#006FE# => romdata <= X"85F03F74";
    when 16#006FF# => romdata <= X"5187B53F";
    when 16#00700# => romdata <= X"8A5185CC";
    when 16#00701# => romdata <= X"3F800BFF";
    when 16#00702# => romdata <= X"16555372";
    when 16#00703# => romdata <= X"7425A238";
    when 16#00704# => romdata <= X"72101080";
    when 16#00705# => romdata <= X"FBE80805";
    when 16#00706# => romdata <= X"70085252";
    when 16#00707# => romdata <= X"87963F8A";
    when 16#00708# => romdata <= X"5185AD3F";
    when 16#00709# => romdata <= X"81137081";
    when 16#0070A# => romdata <= X"FF065452";
    when 16#0070B# => romdata <= X"737324E0";
    when 16#0070C# => romdata <= X"3874B00C";
    when 16#0070D# => romdata <= X"863D0D04";
    when 16#0070E# => romdata <= X"FD3D0D81";
    when 16#0070F# => romdata <= X"51E08C3F";
    when 16#00710# => romdata <= X"B00881FF";
    when 16#00711# => romdata <= X"06528251";
    when 16#00712# => romdata <= X"E1B33FB0";
    when 16#00713# => romdata <= X"0881FF06";
    when 16#00714# => romdata <= X"538351E1";
    when 16#00715# => romdata <= X"A83F80FB";
    when 16#00716# => romdata <= X"EC085480";
    when 16#00717# => romdata <= X"740CB008";
    when 16#00718# => romdata <= X"88150C71";
    when 16#00719# => romdata <= X"832B7307";
    when 16#0071A# => romdata <= X"8C150C73";
    when 16#0071B# => romdata <= X"085271FB";
    when 16#0071C# => romdata <= X"3871B00C";
    when 16#0071D# => romdata <= X"853D0D04";
    when 16#0071E# => romdata <= X"FF3D0D81";
    when 16#0071F# => romdata <= X"51DFCC3F";
    when 16#00720# => romdata <= X"80FBEC08";
    when 16#00721# => romdata <= X"B0089012";
    when 16#00722# => romdata <= X"0C528272";
    when 16#00723# => romdata <= X"0C833D0D";
    when 16#00724# => romdata <= X"04803D0D";
    when 16#00725# => romdata <= X"80FBEC08";
    when 16#00726# => romdata <= X"5180710C";
    when 16#00727# => romdata <= X"70B00C82";
    when 16#00728# => romdata <= X"3D0D04FD";
    when 16#00729# => romdata <= X"3D0D800B";
    when 16#0072A# => romdata <= X"80FBEC08";
    when 16#0072B# => romdata <= X"54548073";
    when 16#0072C# => romdata <= X"0CFECAC0";
    when 16#0072D# => romdata <= X"90860B88";
    when 16#0072E# => romdata <= X"140C7383";
    when 16#0072F# => romdata <= X"2B82078C";
    when 16#00730# => romdata <= X"140C7208";
    when 16#00731# => romdata <= X"5271FB38";
    when 16#00732# => romdata <= X"81147081";
    when 16#00733# => romdata <= X"FF065551";
    when 16#00734# => romdata <= X"A27427DA";
    when 16#00735# => romdata <= X"3871B00C";
    when 16#00736# => romdata <= X"853D0D04";
    when 16#00737# => romdata <= X"FD3D0D80";
    when 16#00738# => romdata <= X"0B80FBEC";
    when 16#00739# => romdata <= X"08545480";
    when 16#0073A# => romdata <= X"730C880A";
    when 16#0073B# => romdata <= X"0B88140C";
    when 16#0073C# => romdata <= X"73832B81";
    when 16#0073D# => romdata <= X"078C140C";
    when 16#0073E# => romdata <= X"72085271";
    when 16#0073F# => romdata <= X"FB388114";
    when 16#00740# => romdata <= X"7081FF06";
    when 16#00741# => romdata <= X"5551A274";
    when 16#00742# => romdata <= X"27DD3871";
    when 16#00743# => romdata <= X"B00C853D";
    when 16#00744# => romdata <= X"0D04FE3D";
    when 16#00745# => romdata <= X"0D8151DE";
    when 16#00746# => romdata <= X"B23F80FB";
    when 16#00747# => romdata <= X"EC085380";
    when 16#00748# => romdata <= X"730C810B";
    when 16#00749# => romdata <= X"88140CB0";
    when 16#0074A# => romdata <= X"08832B8F";
    when 16#0074B# => romdata <= X"F8067082";
    when 16#0074C# => romdata <= X"078C150C";
    when 16#0074D# => romdata <= X"52720852";
    when 16#0074E# => romdata <= X"71FB3889";
    when 16#0074F# => romdata <= X"730C71B0";
    when 16#00750# => romdata <= X"0C843D0D";
    when 16#00751# => romdata <= X"04D88A3F";
    when 16#00752# => romdata <= X"04FB3D0D";
    when 16#00753# => romdata <= X"77795555";
    when 16#00754# => romdata <= X"80567575";
    when 16#00755# => romdata <= X"24AB3880";
    when 16#00756# => romdata <= X"74249D38";
    when 16#00757# => romdata <= X"80537352";
    when 16#00758# => romdata <= X"745180E1";
    when 16#00759# => romdata <= X"3FB00854";
    when 16#0075A# => romdata <= X"75802E85";
    when 16#0075B# => romdata <= X"38B00830";
    when 16#0075C# => romdata <= X"5473B00C";
    when 16#0075D# => romdata <= X"873D0D04";
    when 16#0075E# => romdata <= X"73307681";
    when 16#0075F# => romdata <= X"325754DC";
    when 16#00760# => romdata <= X"39743055";
    when 16#00761# => romdata <= X"81567380";
    when 16#00762# => romdata <= X"25D238EC";
    when 16#00763# => romdata <= X"39FA3D0D";
    when 16#00764# => romdata <= X"787A5755";
    when 16#00765# => romdata <= X"80577675";
    when 16#00766# => romdata <= X"24A43875";
    when 16#00767# => romdata <= X"9F2C5481";
    when 16#00768# => romdata <= X"53757432";
    when 16#00769# => romdata <= X"74315274";
    when 16#0076A# => romdata <= X"519B3FB0";
    when 16#0076B# => romdata <= X"08547680";
    when 16#0076C# => romdata <= X"2E8538B0";
    when 16#0076D# => romdata <= X"08305473";
    when 16#0076E# => romdata <= X"B00C883D";
    when 16#0076F# => romdata <= X"0D047430";
    when 16#00770# => romdata <= X"558157D7";
    when 16#00771# => romdata <= X"39FC3D0D";
    when 16#00772# => romdata <= X"76785354";
    when 16#00773# => romdata <= X"81538074";
    when 16#00774# => romdata <= X"73265255";
    when 16#00775# => romdata <= X"72802E98";
    when 16#00776# => romdata <= X"3870802E";
    when 16#00777# => romdata <= X"A9388072";
    when 16#00778# => romdata <= X"24A43871";
    when 16#00779# => romdata <= X"10731075";
    when 16#0077A# => romdata <= X"72265354";
    when 16#0077B# => romdata <= X"5272EA38";
    when 16#0077C# => romdata <= X"73517883";
    when 16#0077D# => romdata <= X"38745170";
    when 16#0077E# => romdata <= X"B00C863D";
    when 16#0077F# => romdata <= X"0D047281";
    when 16#00780# => romdata <= X"2A72812A";
    when 16#00781# => romdata <= X"53537280";
    when 16#00782# => romdata <= X"2EE63871";
    when 16#00783# => romdata <= X"7426EF38";
    when 16#00784# => romdata <= X"73723175";
    when 16#00785# => romdata <= X"74077481";
    when 16#00786# => romdata <= X"2A74812A";
    when 16#00787# => romdata <= X"55555654";
    when 16#00788# => romdata <= X"E5391010";
    when 16#00789# => romdata <= X"10101010";
    when 16#0078A# => romdata <= X"10101010";
    when 16#0078B# => romdata <= X"10101010";
    when 16#0078C# => romdata <= X"10101010";
    when 16#0078D# => romdata <= X"10101010";
    when 16#0078E# => romdata <= X"10101010";
    when 16#0078F# => romdata <= X"10101010";
    when 16#00790# => romdata <= X"10535104";
    when 16#00791# => romdata <= X"7381FF06";
    when 16#00792# => romdata <= X"73830609";
    when 16#00793# => romdata <= X"81058305";
    when 16#00794# => romdata <= X"1010102B";
    when 16#00795# => romdata <= X"0772FC06";
    when 16#00796# => romdata <= X"0C515104";
    when 16#00797# => romdata <= X"3C047272";
    when 16#00798# => romdata <= X"80728106";
    when 16#00799# => romdata <= X"FF050972";
    when 16#0079A# => romdata <= X"06057110";
    when 16#0079B# => romdata <= X"52720A10";
    when 16#0079C# => romdata <= X"0A5372ED";
    when 16#0079D# => romdata <= X"38515153";
    when 16#0079E# => romdata <= X"5104B008";
    when 16#0079F# => romdata <= X"B408B808";
    when 16#007A0# => romdata <= X"7575BB8D";
    when 16#007A1# => romdata <= X"2D5050B0";
    when 16#007A2# => romdata <= X"0856B80C";
    when 16#007A3# => romdata <= X"B40CB00C";
    when 16#007A4# => romdata <= X"5104B008";
    when 16#007A5# => romdata <= X"B408B808";
    when 16#007A6# => romdata <= X"7575BAC9";
    when 16#007A7# => romdata <= X"2D5050B0";
    when 16#007A8# => romdata <= X"0856B80C";
    when 16#007A9# => romdata <= X"B40CB00C";
    when 16#007AA# => romdata <= X"5104B008";
    when 16#007AB# => romdata <= X"B408B808";
    when 16#007AC# => romdata <= X"90B92DB8";
    when 16#007AD# => romdata <= X"0CB40CB0";
    when 16#007AE# => romdata <= X"0C04FF3D";
    when 16#007AF# => romdata <= X"0D028F05";
    when 16#007B0# => romdata <= X"3380FC9C";
    when 16#007B1# => romdata <= X"0852710C";
    when 16#007B2# => romdata <= X"800BB00C";
    when 16#007B3# => romdata <= X"833D0D04";
    when 16#007B4# => romdata <= X"FF3D0D02";
    when 16#007B5# => romdata <= X"8F053351";
    when 16#007B6# => romdata <= X"81A4B408";
    when 16#007B7# => romdata <= X"52712DB0";
    when 16#007B8# => romdata <= X"0881FF06";
    when 16#007B9# => romdata <= X"B00C833D";
    when 16#007BA# => romdata <= X"0D04FE3D";
    when 16#007BB# => romdata <= X"0D747033";
    when 16#007BC# => romdata <= X"53537180";
    when 16#007BD# => romdata <= X"2E933881";
    when 16#007BE# => romdata <= X"13725281";
    when 16#007BF# => romdata <= X"A4B40853";
    when 16#007C0# => romdata <= X"53712D72";
    when 16#007C1# => romdata <= X"335271EF";
    when 16#007C2# => romdata <= X"38843D0D";
    when 16#007C3# => romdata <= X"04F43D0D";
    when 16#007C4# => romdata <= X"7F028405";
    when 16#007C5# => romdata <= X"BB053355";
    when 16#007C6# => romdata <= X"57880B8C";
    when 16#007C7# => romdata <= X"3D5B5989";
    when 16#007C8# => romdata <= X"5380F9C0";
    when 16#007C9# => romdata <= X"52795185";
    when 16#007CA# => romdata <= X"E63F7379";
    when 16#007CB# => romdata <= X"2E80FF38";
    when 16#007CC# => romdata <= X"78567390";
    when 16#007CD# => romdata <= X"2E80EC38";
    when 16#007CE# => romdata <= X"02A70558";
    when 16#007CF# => romdata <= X"768F0654";
    when 16#007D0# => romdata <= X"73892680";
    when 16#007D1# => romdata <= X"C2387518";
    when 16#007D2# => romdata <= X"B0155555";
    when 16#007D3# => romdata <= X"73753476";
    when 16#007D4# => romdata <= X"842AFF17";
    when 16#007D5# => romdata <= X"7081FF06";
    when 16#007D6# => romdata <= X"58555775";
    when 16#007D7# => romdata <= X"DF38781A";
    when 16#007D8# => romdata <= X"55757534";
    when 16#007D9# => romdata <= X"79703355";
    when 16#007DA# => romdata <= X"5573802E";
    when 16#007DB# => romdata <= X"93388115";
    when 16#007DC# => romdata <= X"745281A4";
    when 16#007DD# => romdata <= X"B4085755";
    when 16#007DE# => romdata <= X"752D7433";
    when 16#007DF# => romdata <= X"5473EF38";
    when 16#007E0# => romdata <= X"78B00C8E";
    when 16#007E1# => romdata <= X"3D0D0475";
    when 16#007E2# => romdata <= X"18B71555";
    when 16#007E3# => romdata <= X"55737534";
    when 16#007E4# => romdata <= X"76842AFF";
    when 16#007E5# => romdata <= X"177081FF";
    when 16#007E6# => romdata <= X"06585557";
    when 16#007E7# => romdata <= X"75FF9D38";
    when 16#007E8# => romdata <= X"FFBC3984";
    when 16#007E9# => romdata <= X"70575902";
    when 16#007EA# => romdata <= X"A70558FF";
    when 16#007EB# => romdata <= X"8F398270";
    when 16#007EC# => romdata <= X"5759F439";
    when 16#007ED# => romdata <= X"F13D0D61";
    when 16#007EE# => romdata <= X"8D3D705B";
    when 16#007EF# => romdata <= X"5C5A807A";
    when 16#007F0# => romdata <= X"5657767A";
    when 16#007F1# => romdata <= X"24818538";
    when 16#007F2# => romdata <= X"7817548A";
    when 16#007F3# => romdata <= X"52745184";
    when 16#007F4# => romdata <= X"8C3FB008";
    when 16#007F5# => romdata <= X"B0055372";
    when 16#007F6# => romdata <= X"74348117";
    when 16#007F7# => romdata <= X"578A5274";
    when 16#007F8# => romdata <= X"5183D53F";
    when 16#007F9# => romdata <= X"B00855B0";
    when 16#007FA# => romdata <= X"08DE38B0";
    when 16#007FB# => romdata <= X"08779F2A";
    when 16#007FC# => romdata <= X"1870812C";
    when 16#007FD# => romdata <= X"5A565680";
    when 16#007FE# => romdata <= X"78259E38";
    when 16#007FF# => romdata <= X"7817FF05";
    when 16#00800# => romdata <= X"55751970";
    when 16#00801# => romdata <= X"33555374";
    when 16#00802# => romdata <= X"33733473";
    when 16#00803# => romdata <= X"75348116";
    when 16#00804# => romdata <= X"FF165656";
    when 16#00805# => romdata <= X"777624E9";
    when 16#00806# => romdata <= X"38761958";
    when 16#00807# => romdata <= X"80783480";
    when 16#00808# => romdata <= X"7A241770";
    when 16#00809# => romdata <= X"81FF067C";
    when 16#0080A# => romdata <= X"70335657";
    when 16#0080B# => romdata <= X"55567280";
    when 16#0080C# => romdata <= X"2E933881";
    when 16#0080D# => romdata <= X"15735281";
    when 16#0080E# => romdata <= X"A4B40858";
    when 16#0080F# => romdata <= X"55762D74";
    when 16#00810# => romdata <= X"335372EF";
    when 16#00811# => romdata <= X"3873B00C";
    when 16#00812# => romdata <= X"913D0D04";
    when 16#00813# => romdata <= X"AD7B3402";
    when 16#00814# => romdata <= X"AD057A30";
    when 16#00815# => romdata <= X"71195656";
    when 16#00816# => romdata <= X"598A5274";
    when 16#00817# => romdata <= X"5182FE3F";
    when 16#00818# => romdata <= X"B008B005";
    when 16#00819# => romdata <= X"53727434";
    when 16#0081A# => romdata <= X"8117578A";
    when 16#0081B# => romdata <= X"52745182";
    when 16#0081C# => romdata <= X"C73FB008";
    when 16#0081D# => romdata <= X"55B008FE";
    when 16#0081E# => romdata <= X"CF38FEEF";
    when 16#0081F# => romdata <= X"39FD3D0D";
    when 16#00820# => romdata <= X"02970533";
    when 16#00821# => romdata <= X"0284059B";
    when 16#00822# => romdata <= X"05335553";
    when 16#00823# => romdata <= X"72742797";
    when 16#00824# => romdata <= X"38A05181";
    when 16#00825# => romdata <= X"A4B40852";
    when 16#00826# => romdata <= X"712D8113";
    when 16#00827# => romdata <= X"7081FF06";
    when 16#00828# => romdata <= X"54527373";
    when 16#00829# => romdata <= X"26EB3885";
    when 16#0082A# => romdata <= X"3D0D04FF";
    when 16#0082B# => romdata <= X"3D0D80FC";
    when 16#0082C# => romdata <= X"90087410";
    when 16#0082D# => romdata <= X"1570822B";
    when 16#0082E# => romdata <= X"94130C52";
    when 16#0082F# => romdata <= X"52850B98";
    when 16#00830# => romdata <= X"130C9812";
    when 16#00831# => romdata <= X"08708106";
    when 16#00832# => romdata <= X"515170F6";
    when 16#00833# => romdata <= X"38833D0D";
    when 16#00834# => romdata <= X"04FD3D0D";
    when 16#00835# => romdata <= X"80FC9008";
    when 16#00836# => romdata <= X"7680E1D4";
    when 16#00837# => romdata <= X"2994120C";
    when 16#00838# => romdata <= X"54850B98";
    when 16#00839# => romdata <= X"150C9814";
    when 16#0083A# => romdata <= X"08708106";
    when 16#0083B# => romdata <= X"515372F6";
    when 16#0083C# => romdata <= X"38853D0D";
    when 16#0083D# => romdata <= X"04803D0D";
    when 16#0083E# => romdata <= X"80FC9008";
    when 16#0083F# => romdata <= X"51870B84";
    when 16#00840# => romdata <= X"120CFF0B";
    when 16#00841# => romdata <= X"A4120CA7";
    when 16#00842# => romdata <= X"0BA8120C";
    when 16#00843# => romdata <= X"80E1D40B";
    when 16#00844# => romdata <= X"94120C87";
    when 16#00845# => romdata <= X"0B98120C";
    when 16#00846# => romdata <= X"823D0D04";
    when 16#00847# => romdata <= X"803D0D80";
    when 16#00848# => romdata <= X"FC940851";
    when 16#00849# => romdata <= X"80EC0B8C";
    when 16#0084A# => romdata <= X"120C830B";
    when 16#0084B# => romdata <= X"88120C82";
    when 16#0084C# => romdata <= X"3D0D0480";
    when 16#0084D# => romdata <= X"3D0D80FC";
    when 16#0084E# => romdata <= X"94088411";
    when 16#0084F# => romdata <= X"088106B0";
    when 16#00850# => romdata <= X"0C51823D";
    when 16#00851# => romdata <= X"0D04FF3D";
    when 16#00852# => romdata <= X"0D80FC94";
    when 16#00853# => romdata <= X"08528412";
    when 16#00854# => romdata <= X"08708106";
    when 16#00855# => romdata <= X"51517080";
    when 16#00856# => romdata <= X"2EF43871";
    when 16#00857# => romdata <= X"087081FF";
    when 16#00858# => romdata <= X"06B00C51";
    when 16#00859# => romdata <= X"833D0D04";
    when 16#0085A# => romdata <= X"FE3D0D02";
    when 16#0085B# => romdata <= X"93053353";
    when 16#0085C# => romdata <= X"728A2E9C";
    when 16#0085D# => romdata <= X"3880FC94";
    when 16#0085E# => romdata <= X"08528412";
    when 16#0085F# => romdata <= X"0870892A";
    when 16#00860# => romdata <= X"70810651";
    when 16#00861# => romdata <= X"515170F2";
    when 16#00862# => romdata <= X"3872720C";
    when 16#00863# => romdata <= X"843D0D04";
    when 16#00864# => romdata <= X"80FC9408";
    when 16#00865# => romdata <= X"52841208";
    when 16#00866# => romdata <= X"70892A70";
    when 16#00867# => romdata <= X"81065151";
    when 16#00868# => romdata <= X"5170F238";
    when 16#00869# => romdata <= X"8D720C84";
    when 16#0086A# => romdata <= X"12087089";
    when 16#0086B# => romdata <= X"2A708106";
    when 16#0086C# => romdata <= X"51515170";
    when 16#0086D# => romdata <= X"C538D239";
    when 16#0086E# => romdata <= X"BC0802BC";
    when 16#0086F# => romdata <= X"0CFD3D0D";
    when 16#00870# => romdata <= X"8053BC08";
    when 16#00871# => romdata <= X"8C050852";
    when 16#00872# => romdata <= X"BC088805";
    when 16#00873# => romdata <= X"0851F7F5";
    when 16#00874# => romdata <= X"3FB00870";
    when 16#00875# => romdata <= X"B00C5485";
    when 16#00876# => romdata <= X"3D0DBC0C";
    when 16#00877# => romdata <= X"04BC0802";
    when 16#00878# => romdata <= X"BC0CFD3D";
    when 16#00879# => romdata <= X"0D8153BC";
    when 16#0087A# => romdata <= X"088C0508";
    when 16#0087B# => romdata <= X"52BC0888";
    when 16#0087C# => romdata <= X"050851F7";
    when 16#0087D# => romdata <= X"D03FB008";
    when 16#0087E# => romdata <= X"70B00C54";
    when 16#0087F# => romdata <= X"853D0DBC";
    when 16#00880# => romdata <= X"0C04803D";
    when 16#00881# => romdata <= X"0D865184";
    when 16#00882# => romdata <= X"963F8151";
    when 16#00883# => romdata <= X"A1D33FFC";
    when 16#00884# => romdata <= X"3D0D7670";
    when 16#00885# => romdata <= X"797B5555";
    when 16#00886# => romdata <= X"55558F72";
    when 16#00887# => romdata <= X"278C3872";
    when 16#00888# => romdata <= X"75078306";
    when 16#00889# => romdata <= X"5170802E";
    when 16#0088A# => romdata <= X"A738FF12";
    when 16#0088B# => romdata <= X"5271FF2E";
    when 16#0088C# => romdata <= X"98387270";
    when 16#0088D# => romdata <= X"81055433";
    when 16#0088E# => romdata <= X"74708105";
    when 16#0088F# => romdata <= X"5634FF12";
    when 16#00890# => romdata <= X"5271FF2E";
    when 16#00891# => romdata <= X"098106EA";
    when 16#00892# => romdata <= X"3874B00C";
    when 16#00893# => romdata <= X"863D0D04";
    when 16#00894# => romdata <= X"74517270";
    when 16#00895# => romdata <= X"84055408";
    when 16#00896# => romdata <= X"71708405";
    when 16#00897# => romdata <= X"530C7270";
    when 16#00898# => romdata <= X"84055408";
    when 16#00899# => romdata <= X"71708405";
    when 16#0089A# => romdata <= X"530C7270";
    when 16#0089B# => romdata <= X"84055408";
    when 16#0089C# => romdata <= X"71708405";
    when 16#0089D# => romdata <= X"530C7270";
    when 16#0089E# => romdata <= X"84055408";
    when 16#0089F# => romdata <= X"71708405";
    when 16#008A0# => romdata <= X"530CF012";
    when 16#008A1# => romdata <= X"52718F26";
    when 16#008A2# => romdata <= X"C9388372";
    when 16#008A3# => romdata <= X"27953872";
    when 16#008A4# => romdata <= X"70840554";
    when 16#008A5# => romdata <= X"08717084";
    when 16#008A6# => romdata <= X"05530CFC";
    when 16#008A7# => romdata <= X"12527183";
    when 16#008A8# => romdata <= X"26ED3870";
    when 16#008A9# => romdata <= X"54FF8339";
    when 16#008AA# => romdata <= X"FD3D0D75";
    when 16#008AB# => romdata <= X"5384D813";
    when 16#008AC# => romdata <= X"08802E8A";
    when 16#008AD# => romdata <= X"38805372";
    when 16#008AE# => romdata <= X"B00C853D";
    when 16#008AF# => romdata <= X"0D048180";
    when 16#008B0# => romdata <= X"5272518D";
    when 16#008B1# => romdata <= X"9B3FB008";
    when 16#008B2# => romdata <= X"84D8140C";
    when 16#008B3# => romdata <= X"FF53B008";
    when 16#008B4# => romdata <= X"802EE438";
    when 16#008B5# => romdata <= X"B008549F";
    when 16#008B6# => romdata <= X"53807470";
    when 16#008B7# => romdata <= X"8405560C";
    when 16#008B8# => romdata <= X"FF135380";
    when 16#008B9# => romdata <= X"7324CE38";
    when 16#008BA# => romdata <= X"80747084";
    when 16#008BB# => romdata <= X"05560CFF";
    when 16#008BC# => romdata <= X"13537280";
    when 16#008BD# => romdata <= X"25E338FF";
    when 16#008BE# => romdata <= X"BC39FD3D";
    when 16#008BF# => romdata <= X"0D757755";
    when 16#008C0# => romdata <= X"539F7427";
    when 16#008C1# => romdata <= X"8D389673";
    when 16#008C2# => romdata <= X"0CFF5271";
    when 16#008C3# => romdata <= X"B00C853D";
    when 16#008C4# => romdata <= X"0D0484D8";
    when 16#008C5# => romdata <= X"13085271";
    when 16#008C6# => romdata <= X"802E9338";
    when 16#008C7# => romdata <= X"73101012";
    when 16#008C8# => romdata <= X"70087972";
    when 16#008C9# => romdata <= X"0C515271";
    when 16#008CA# => romdata <= X"B00C853D";
    when 16#008CB# => romdata <= X"0D047251";
    when 16#008CC# => romdata <= X"FEF63FFF";
    when 16#008CD# => romdata <= X"52B008D3";
    when 16#008CE# => romdata <= X"3884D813";
    when 16#008CF# => romdata <= X"08741010";
    when 16#008D0# => romdata <= X"1170087A";
    when 16#008D1# => romdata <= X"720C5151";
    when 16#008D2# => romdata <= X"52DD39F9";
    when 16#008D3# => romdata <= X"3D0D797B";
    when 16#008D4# => romdata <= X"5856769F";
    when 16#008D5# => romdata <= X"2680E838";
    when 16#008D6# => romdata <= X"84D81608";
    when 16#008D7# => romdata <= X"5473802E";
    when 16#008D8# => romdata <= X"AA387610";
    when 16#008D9# => romdata <= X"10147008";
    when 16#008DA# => romdata <= X"55557380";
    when 16#008DB# => romdata <= X"2EBA3880";
    when 16#008DC# => romdata <= X"5873812E";
    when 16#008DD# => romdata <= X"8F3873FF";
    when 16#008DE# => romdata <= X"2EA33880";
    when 16#008DF# => romdata <= X"750C7651";
    when 16#008E0# => romdata <= X"732D8058";
    when 16#008E1# => romdata <= X"77B00C89";
    when 16#008E2# => romdata <= X"3D0D0475";
    when 16#008E3# => romdata <= X"51FE993F";
    when 16#008E4# => romdata <= X"FF58B008";
    when 16#008E5# => romdata <= X"EF3884D8";
    when 16#008E6# => romdata <= X"160854C6";
    when 16#008E7# => romdata <= X"3996760C";
    when 16#008E8# => romdata <= X"810BB00C";
    when 16#008E9# => romdata <= X"893D0D04";
    when 16#008EA# => romdata <= X"755181ED";
    when 16#008EB# => romdata <= X"3F7653B0";
    when 16#008EC# => romdata <= X"08527551";
    when 16#008ED# => romdata <= X"81AD3FB0";
    when 16#008EE# => romdata <= X"08B00C89";
    when 16#008EF# => romdata <= X"3D0D0496";
    when 16#008F0# => romdata <= X"760CFF0B";
    when 16#008F1# => romdata <= X"B00C893D";
    when 16#008F2# => romdata <= X"0D04FC3D";
    when 16#008F3# => romdata <= X"0D767856";
    when 16#008F4# => romdata <= X"53FF5474";
    when 16#008F5# => romdata <= X"9F26B138";
    when 16#008F6# => romdata <= X"84D81308";
    when 16#008F7# => romdata <= X"5271802E";
    when 16#008F8# => romdata <= X"AE387410";
    when 16#008F9# => romdata <= X"10127008";
    when 16#008FA# => romdata <= X"53538154";
    when 16#008FB# => romdata <= X"71802E98";
    when 16#008FC# => romdata <= X"38825471";
    when 16#008FD# => romdata <= X"FF2E9138";
    when 16#008FE# => romdata <= X"83547181";
    when 16#008FF# => romdata <= X"2E8A3880";
    when 16#00900# => romdata <= X"730C7451";
    when 16#00901# => romdata <= X"712D8054";
    when 16#00902# => romdata <= X"73B00C86";
    when 16#00903# => romdata <= X"3D0D0472";
    when 16#00904# => romdata <= X"51FD953F";
    when 16#00905# => romdata <= X"B008F138";
    when 16#00906# => romdata <= X"84D81308";
    when 16#00907# => romdata <= X"52C439FF";
    when 16#00908# => romdata <= X"3D0D7352";
    when 16#00909# => romdata <= X"80FCA008";
    when 16#0090A# => romdata <= X"51FEA03F";
    when 16#0090B# => romdata <= X"833D0D04";
    when 16#0090C# => romdata <= X"FE3D0D75";
    when 16#0090D# => romdata <= X"53745280";
    when 16#0090E# => romdata <= X"FCA00851";
    when 16#0090F# => romdata <= X"FDBC3F84";
    when 16#00910# => romdata <= X"3D0D0480";
    when 16#00911# => romdata <= X"3D0D80FC";
    when 16#00912# => romdata <= X"A00851FC";
    when 16#00913# => romdata <= X"DB3F823D";
    when 16#00914# => romdata <= X"0D04FF3D";
    when 16#00915# => romdata <= X"0D735280";
    when 16#00916# => romdata <= X"FCA00851";
    when 16#00917# => romdata <= X"FEEC3F83";
    when 16#00918# => romdata <= X"3D0D04FC";
    when 16#00919# => romdata <= X"3D0D800B";
    when 16#0091A# => romdata <= X"81A4BC0C";
    when 16#0091B# => romdata <= X"78527751";
    when 16#0091C# => romdata <= X"9CAA3FB0";
    when 16#0091D# => romdata <= X"0854B008";
    when 16#0091E# => romdata <= X"FF2E8838";
    when 16#0091F# => romdata <= X"73B00C86";
    when 16#00920# => romdata <= X"3D0D0481";
    when 16#00921# => romdata <= X"A4BC0855";
    when 16#00922# => romdata <= X"74802EF0";
    when 16#00923# => romdata <= X"38767571";
    when 16#00924# => romdata <= X"0C5373B0";
    when 16#00925# => romdata <= X"0C863D0D";
    when 16#00926# => romdata <= X"049BFC3F";
    when 16#00927# => romdata <= X"04FC3D0D";
    when 16#00928# => romdata <= X"76707970";
    when 16#00929# => romdata <= X"73078306";
    when 16#0092A# => romdata <= X"54545455";
    when 16#0092B# => romdata <= X"7080C338";
    when 16#0092C# => romdata <= X"71700870";
    when 16#0092D# => romdata <= X"0970F7FB";
    when 16#0092E# => romdata <= X"FDFF1306";
    when 16#0092F# => romdata <= X"70F88482";
    when 16#00930# => romdata <= X"81800651";
    when 16#00931# => romdata <= X"51535354";
    when 16#00932# => romdata <= X"70A63884";
    when 16#00933# => romdata <= X"14727470";
    when 16#00934# => romdata <= X"8405560C";
    when 16#00935# => romdata <= X"70087009";
    when 16#00936# => romdata <= X"70F7FBFD";
    when 16#00937# => romdata <= X"FF130670";
    when 16#00938# => romdata <= X"F8848281";
    when 16#00939# => romdata <= X"80065151";
    when 16#0093A# => romdata <= X"53535470";
    when 16#0093B# => romdata <= X"802EDC38";
    when 16#0093C# => romdata <= X"73527170";
    when 16#0093D# => romdata <= X"81055333";
    when 16#0093E# => romdata <= X"51707370";
    when 16#0093F# => romdata <= X"81055534";
    when 16#00940# => romdata <= X"70F03874";
    when 16#00941# => romdata <= X"B00C863D";
    when 16#00942# => romdata <= X"0D04FD3D";
    when 16#00943# => romdata <= X"0D757071";
    when 16#00944# => romdata <= X"83065355";
    when 16#00945# => romdata <= X"5270B838";
    when 16#00946# => romdata <= X"71700870";
    when 16#00947# => romdata <= X"09F7FBFD";
    when 16#00948# => romdata <= X"FF120670";
    when 16#00949# => romdata <= X"F8848281";
    when 16#0094A# => romdata <= X"80065151";
    when 16#0094B# => romdata <= X"5253709D";
    when 16#0094C# => romdata <= X"38841370";
    when 16#0094D# => romdata <= X"087009F7";
    when 16#0094E# => romdata <= X"FBFDFF12";
    when 16#0094F# => romdata <= X"0670F884";
    when 16#00950# => romdata <= X"82818006";
    when 16#00951# => romdata <= X"51515253";
    when 16#00952# => romdata <= X"70802EE5";
    when 16#00953# => romdata <= X"38725271";
    when 16#00954# => romdata <= X"33517080";
    when 16#00955# => romdata <= X"2E8A3881";
    when 16#00956# => romdata <= X"12703352";
    when 16#00957# => romdata <= X"5270F838";
    when 16#00958# => romdata <= X"717431B0";
    when 16#00959# => romdata <= X"0C853D0D";
    when 16#0095A# => romdata <= X"04FA3D0D";
    when 16#0095B# => romdata <= X"787A7C70";
    when 16#0095C# => romdata <= X"54555552";
    when 16#0095D# => romdata <= X"72802E80";
    when 16#0095E# => romdata <= X"D9387174";
    when 16#0095F# => romdata <= X"07830651";
    when 16#00960# => romdata <= X"70802E80";
    when 16#00961# => romdata <= X"D438FF13";
    when 16#00962# => romdata <= X"5372FF2E";
    when 16#00963# => romdata <= X"B1387133";
    when 16#00964# => romdata <= X"74335651";
    when 16#00965# => romdata <= X"74712E09";
    when 16#00966# => romdata <= X"8106A938";
    when 16#00967# => romdata <= X"72802E81";
    when 16#00968# => romdata <= X"87387081";
    when 16#00969# => romdata <= X"FF065170";
    when 16#0096A# => romdata <= X"802E80FC";
    when 16#0096B# => romdata <= X"38811281";
    when 16#0096C# => romdata <= X"15FF1555";
    when 16#0096D# => romdata <= X"555272FF";
    when 16#0096E# => romdata <= X"2E098106";
    when 16#0096F# => romdata <= X"D1387133";
    when 16#00970# => romdata <= X"74335651";
    when 16#00971# => romdata <= X"7081FF06";
    when 16#00972# => romdata <= X"7581FF06";
    when 16#00973# => romdata <= X"71713151";
    when 16#00974# => romdata <= X"525270B0";
    when 16#00975# => romdata <= X"0C883D0D";
    when 16#00976# => romdata <= X"04717457";
    when 16#00977# => romdata <= X"55837327";
    when 16#00978# => romdata <= X"88387108";
    when 16#00979# => romdata <= X"74082E88";
    when 16#0097A# => romdata <= X"38747655";
    when 16#0097B# => romdata <= X"52FF9739";
    when 16#0097C# => romdata <= X"FC135372";
    when 16#0097D# => romdata <= X"802EB138";
    when 16#0097E# => romdata <= X"74087009";
    when 16#0097F# => romdata <= X"F7FBFDFF";
    when 16#00980# => romdata <= X"120670F8";
    when 16#00981# => romdata <= X"84828180";
    when 16#00982# => romdata <= X"06515151";
    when 16#00983# => romdata <= X"709A3884";
    when 16#00984# => romdata <= X"15841757";
    when 16#00985# => romdata <= X"55837327";
    when 16#00986# => romdata <= X"D0387408";
    when 16#00987# => romdata <= X"76082ED0";
    when 16#00988# => romdata <= X"38747655";
    when 16#00989# => romdata <= X"52FEDF39";
    when 16#0098A# => romdata <= X"800BB00C";
    when 16#0098B# => romdata <= X"883D0D04";
    when 16#0098C# => romdata <= X"F33D0D60";
    when 16#0098D# => romdata <= X"6264725A";
    when 16#0098E# => romdata <= X"5A5E5E80";
    when 16#0098F# => romdata <= X"5C767081";
    when 16#00990# => romdata <= X"05583380";
    when 16#00991# => romdata <= X"F9D51133";
    when 16#00992# => romdata <= X"70832A70";
    when 16#00993# => romdata <= X"81065155";
    when 16#00994# => romdata <= X"555672E9";
    when 16#00995# => romdata <= X"3875AD2E";
    when 16#00996# => romdata <= X"82883875";
    when 16#00997# => romdata <= X"AB2E8284";
    when 16#00998# => romdata <= X"38773070";
    when 16#00999# => romdata <= X"79078025";
    when 16#0099A# => romdata <= X"79903270";
    when 16#0099B# => romdata <= X"30707207";
    when 16#0099C# => romdata <= X"80257307";
    when 16#0099D# => romdata <= X"53575751";
    when 16#0099E# => romdata <= X"5372802E";
    when 16#0099F# => romdata <= X"873875B0";
    when 16#009A0# => romdata <= X"2E81EB38";
    when 16#009A1# => romdata <= X"778A3888";
    when 16#009A2# => romdata <= X"5875B02E";
    when 16#009A3# => romdata <= X"83388A58";
    when 16#009A4# => romdata <= X"810A5A7B";
    when 16#009A5# => romdata <= X"8438FE0A";
    when 16#009A6# => romdata <= X"5A775279";
    when 16#009A7# => romdata <= X"51F6BE3F";
    when 16#009A8# => romdata <= X"B0087853";
    when 16#009A9# => romdata <= X"7A525BF6";
    when 16#009AA# => romdata <= X"8F3FB008";
    when 16#009AB# => romdata <= X"5A807080";
    when 16#009AC# => romdata <= X"F9D51833";
    when 16#009AD# => romdata <= X"70822A70";
    when 16#009AE# => romdata <= X"81065156";
    when 16#009AF# => romdata <= X"565A5572";
    when 16#009B0# => romdata <= X"802E80C1";
    when 16#009B1# => romdata <= X"38D01656";
    when 16#009B2# => romdata <= X"75782580";
    when 16#009B3# => romdata <= X"D7388079";
    when 16#009B4# => romdata <= X"24757B26";
    when 16#009B5# => romdata <= X"07537293";
    when 16#009B6# => romdata <= X"38747A2E";
    when 16#009B7# => romdata <= X"80EB387A";
    when 16#009B8# => romdata <= X"762580ED";
    when 16#009B9# => romdata <= X"3872802E";
    when 16#009BA# => romdata <= X"80E738FF";
    when 16#009BB# => romdata <= X"77708105";
    when 16#009BC# => romdata <= X"59335759";
    when 16#009BD# => romdata <= X"80F9D516";
    when 16#009BE# => romdata <= X"3370822A";
    when 16#009BF# => romdata <= X"70810651";
    when 16#009C0# => romdata <= X"545472C1";
    when 16#009C1# => romdata <= X"38738306";
    when 16#009C2# => romdata <= X"5372802E";
    when 16#009C3# => romdata <= X"97387381";
    when 16#009C4# => romdata <= X"06C91755";
    when 16#009C5# => romdata <= X"53728538";
    when 16#009C6# => romdata <= X"FFA91654";
    when 16#009C7# => romdata <= X"73567776";
    when 16#009C8# => romdata <= X"24FFAB38";
    when 16#009C9# => romdata <= X"80792480";
    when 16#009CA# => romdata <= X"F0387B80";
    when 16#009CB# => romdata <= X"2E843874";
    when 16#009CC# => romdata <= X"30557C80";
    when 16#009CD# => romdata <= X"2E8C38FF";
    when 16#009CE# => romdata <= X"17537883";
    when 16#009CF# => romdata <= X"387D5372";
    when 16#009D0# => romdata <= X"7D0C74B0";
    when 16#009D1# => romdata <= X"0C8F3D0D";
    when 16#009D2# => romdata <= X"04815375";
    when 16#009D3# => romdata <= X"7B24FF95";
    when 16#009D4# => romdata <= X"38817579";
    when 16#009D5# => romdata <= X"29177870";
    when 16#009D6# => romdata <= X"81055A33";
    when 16#009D7# => romdata <= X"585659FF";
    when 16#009D8# => romdata <= X"9339815C";
    when 16#009D9# => romdata <= X"76708105";
    when 16#009DA# => romdata <= X"583356FD";
    when 16#009DB# => romdata <= X"F4398077";
    when 16#009DC# => romdata <= X"33545472";
    when 16#009DD# => romdata <= X"80F82EB2";
    when 16#009DE# => romdata <= X"387280D8";
    when 16#009DF# => romdata <= X"32703070";
    when 16#009E0# => romdata <= X"80257607";
    when 16#009E1# => romdata <= X"51515372";
    when 16#009E2# => romdata <= X"802EFDF8";
    when 16#009E3# => romdata <= X"38811733";
    when 16#009E4# => romdata <= X"82185856";
    when 16#009E5# => romdata <= X"9058FDF8";
    when 16#009E6# => romdata <= X"39810A55";
    when 16#009E7# => romdata <= X"7B8438FE";
    when 16#009E8# => romdata <= X"0A557F53";
    when 16#009E9# => romdata <= X"A2730CFF";
    when 16#009EA# => romdata <= X"89398154";
    when 16#009EB# => romdata <= X"CC39FD3D";
    when 16#009EC# => romdata <= X"0D775476";
    when 16#009ED# => romdata <= X"53755280";
    when 16#009EE# => romdata <= X"FCA00851";
    when 16#009EF# => romdata <= X"FCF23F85";
    when 16#009F0# => romdata <= X"3D0D04F3";
    when 16#009F1# => romdata <= X"3D0D6062";
    when 16#009F2# => romdata <= X"64725A5A";
    when 16#009F3# => romdata <= X"5D5D805E";
    when 16#009F4# => romdata <= X"76708105";
    when 16#009F5# => romdata <= X"583380F9";
    when 16#009F6# => romdata <= X"D5113370";
    when 16#009F7# => romdata <= X"832A7081";
    when 16#009F8# => romdata <= X"06515555";
    when 16#009F9# => romdata <= X"5672E938";
    when 16#009FA# => romdata <= X"75AD2E81";
    when 16#009FB# => romdata <= X"FF3875AB";
    when 16#009FC# => romdata <= X"2E81FB38";
    when 16#009FD# => romdata <= X"77307079";
    when 16#009FE# => romdata <= X"07802579";
    when 16#009FF# => romdata <= X"90327030";
    when 16#00A00# => romdata <= X"70720780";
    when 16#00A01# => romdata <= X"25730753";
    when 16#00A02# => romdata <= X"57575153";
    when 16#00A03# => romdata <= X"72802E87";
    when 16#00A04# => romdata <= X"3875B02E";
    when 16#00A05# => romdata <= X"81E23877";
    when 16#00A06# => romdata <= X"8A388858";
    when 16#00A07# => romdata <= X"75B02E83";
    when 16#00A08# => romdata <= X"388A5877";
    when 16#00A09# => romdata <= X"52FF51F3";
    when 16#00A0A# => romdata <= X"8F3FB008";
    when 16#00A0B# => romdata <= X"78535AFF";
    when 16#00A0C# => romdata <= X"51F3AA3F";
    when 16#00A0D# => romdata <= X"B0085B80";
    when 16#00A0E# => romdata <= X"705A5580";
    when 16#00A0F# => romdata <= X"F9D51633";
    when 16#00A10# => romdata <= X"70822A70";
    when 16#00A11# => romdata <= X"81065154";
    when 16#00A12# => romdata <= X"5472802E";
    when 16#00A13# => romdata <= X"80C138D0";
    when 16#00A14# => romdata <= X"16567578";
    when 16#00A15# => romdata <= X"2580D738";
    when 16#00A16# => romdata <= X"80792475";
    when 16#00A17# => romdata <= X"7B260753";
    when 16#00A18# => romdata <= X"72933874";
    when 16#00A19# => romdata <= X"7A2E80EB";
    when 16#00A1A# => romdata <= X"387A7625";
    when 16#00A1B# => romdata <= X"80ED3872";
    when 16#00A1C# => romdata <= X"802E80E7";
    when 16#00A1D# => romdata <= X"38FF7770";
    when 16#00A1E# => romdata <= X"81055933";
    when 16#00A1F# => romdata <= X"575980F9";
    when 16#00A20# => romdata <= X"D5163370";
    when 16#00A21# => romdata <= X"822A7081";
    when 16#00A22# => romdata <= X"06515454";
    when 16#00A23# => romdata <= X"72C13873";
    when 16#00A24# => romdata <= X"83065372";
    when 16#00A25# => romdata <= X"802E9738";
    when 16#00A26# => romdata <= X"738106C9";
    when 16#00A27# => romdata <= X"17555372";
    when 16#00A28# => romdata <= X"8538FFA9";
    when 16#00A29# => romdata <= X"16547356";
    when 16#00A2A# => romdata <= X"777624FF";
    when 16#00A2B# => romdata <= X"AB388079";
    when 16#00A2C# => romdata <= X"24818938";
    when 16#00A2D# => romdata <= X"7D802E84";
    when 16#00A2E# => romdata <= X"38743055";
    when 16#00A2F# => romdata <= X"7B802E8C";
    when 16#00A30# => romdata <= X"38FF1753";
    when 16#00A31# => romdata <= X"7883387C";
    when 16#00A32# => romdata <= X"53727C0C";
    when 16#00A33# => romdata <= X"74B00C8F";
    when 16#00A34# => romdata <= X"3D0D0481";
    when 16#00A35# => romdata <= X"53757B24";
    when 16#00A36# => romdata <= X"FF953881";
    when 16#00A37# => romdata <= X"75792917";
    when 16#00A38# => romdata <= X"78708105";
    when 16#00A39# => romdata <= X"5A335856";
    when 16#00A3A# => romdata <= X"59FF9339";
    when 16#00A3B# => romdata <= X"815E7670";
    when 16#00A3C# => romdata <= X"81055833";
    when 16#00A3D# => romdata <= X"56FDFD39";
    when 16#00A3E# => romdata <= X"80773354";
    when 16#00A3F# => romdata <= X"547280F8";
    when 16#00A40# => romdata <= X"2E80C338";
    when 16#00A41# => romdata <= X"7280D832";
    when 16#00A42# => romdata <= X"70307080";
    when 16#00A43# => romdata <= X"25760751";
    when 16#00A44# => romdata <= X"51537280";
    when 16#00A45# => romdata <= X"2EFE8038";
    when 16#00A46# => romdata <= X"81173382";
    when 16#00A47# => romdata <= X"18585690";
    when 16#00A48# => romdata <= X"705358FF";
    when 16#00A49# => romdata <= X"51F1913F";
    when 16#00A4A# => romdata <= X"B0087853";
    when 16#00A4B# => romdata <= X"5AFF51F1";
    when 16#00A4C# => romdata <= X"AC3FB008";
    when 16#00A4D# => romdata <= X"5B80705A";
    when 16#00A4E# => romdata <= X"55FE8039";
    when 16#00A4F# => romdata <= X"FF605455";
    when 16#00A50# => romdata <= X"A2730CFE";
    when 16#00A51# => romdata <= X"F7398154";
    when 16#00A52# => romdata <= X"FFBA39FD";
    when 16#00A53# => romdata <= X"3D0D7754";
    when 16#00A54# => romdata <= X"76537552";
    when 16#00A55# => romdata <= X"80FCA008";
    when 16#00A56# => romdata <= X"51FCE83F";
    when 16#00A57# => romdata <= X"853D0D04";
    when 16#00A58# => romdata <= X"F33D0D7F";
    when 16#00A59# => romdata <= X"618B1170";
    when 16#00A5A# => romdata <= X"F8065C55";
    when 16#00A5B# => romdata <= X"555E7296";
    when 16#00A5C# => romdata <= X"26833890";
    when 16#00A5D# => romdata <= X"59807924";
    when 16#00A5E# => romdata <= X"747A2607";
    when 16#00A5F# => romdata <= X"53805472";
    when 16#00A60# => romdata <= X"742E0981";
    when 16#00A61# => romdata <= X"0680CB38";
    when 16#00A62# => romdata <= X"7D518BCA";
    when 16#00A63# => romdata <= X"3F7883F7";
    when 16#00A64# => romdata <= X"2680C638";
    when 16#00A65# => romdata <= X"78832A70";
    when 16#00A66# => romdata <= X"10101081";
    when 16#00A67# => romdata <= X"83DC058C";
    when 16#00A68# => romdata <= X"11085959";
    when 16#00A69# => romdata <= X"5A76782E";
    when 16#00A6A# => romdata <= X"83B03884";
    when 16#00A6B# => romdata <= X"1708FC06";
    when 16#00A6C# => romdata <= X"568C1708";
    when 16#00A6D# => romdata <= X"88180871";
    when 16#00A6E# => romdata <= X"8C120C88";
    when 16#00A6F# => romdata <= X"120C5875";
    when 16#00A70# => romdata <= X"17841108";
    when 16#00A71# => romdata <= X"81078412";
    when 16#00A72# => romdata <= X"0C537D51";
    when 16#00A73# => romdata <= X"8B893F88";
    when 16#00A74# => romdata <= X"175473B0";
    when 16#00A75# => romdata <= X"0C8F3D0D";
    when 16#00A76# => romdata <= X"0478892A";
    when 16#00A77# => romdata <= X"79832A5B";
    when 16#00A78# => romdata <= X"5372802E";
    when 16#00A79# => romdata <= X"BF387886";
    when 16#00A7A# => romdata <= X"2AB8055A";
    when 16#00A7B# => romdata <= X"847327B4";
    when 16#00A7C# => romdata <= X"3880DB13";
    when 16#00A7D# => romdata <= X"5A947327";
    when 16#00A7E# => romdata <= X"AB38788C";
    when 16#00A7F# => romdata <= X"2A80EE05";
    when 16#00A80# => romdata <= X"5A80D473";
    when 16#00A81# => romdata <= X"279E3878";
    when 16#00A82# => romdata <= X"8F2A80F7";
    when 16#00A83# => romdata <= X"055A82D4";
    when 16#00A84# => romdata <= X"73279138";
    when 16#00A85# => romdata <= X"78922A80";
    when 16#00A86# => romdata <= X"FC055A8A";
    when 16#00A87# => romdata <= X"D4732784";
    when 16#00A88# => romdata <= X"3880FE5A";
    when 16#00A89# => romdata <= X"79101010";
    when 16#00A8A# => romdata <= X"8183DC05";
    when 16#00A8B# => romdata <= X"8C110858";
    when 16#00A8C# => romdata <= X"5576752E";
    when 16#00A8D# => romdata <= X"A3388417";
    when 16#00A8E# => romdata <= X"08FC0670";
    when 16#00A8F# => romdata <= X"7A315556";
    when 16#00A90# => romdata <= X"738F2488";
    when 16#00A91# => romdata <= X"D5387380";
    when 16#00A92# => romdata <= X"25FEE638";
    when 16#00A93# => romdata <= X"8C170857";
    when 16#00A94# => romdata <= X"76752E09";
    when 16#00A95# => romdata <= X"8106DF38";
    when 16#00A96# => romdata <= X"811A5A81";
    when 16#00A97# => romdata <= X"83EC0857";
    when 16#00A98# => romdata <= X"768183E4";
    when 16#00A99# => romdata <= X"2E82C038";
    when 16#00A9A# => romdata <= X"841708FC";
    when 16#00A9B# => romdata <= X"06707A31";
    when 16#00A9C# => romdata <= X"5556738F";
    when 16#00A9D# => romdata <= X"2481F938";
    when 16#00A9E# => romdata <= X"8183E40B";
    when 16#00A9F# => romdata <= X"8183F00C";
    when 16#00AA0# => romdata <= X"8183E40B";
    when 16#00AA1# => romdata <= X"8183EC0C";
    when 16#00AA2# => romdata <= X"738025FE";
    when 16#00AA3# => romdata <= X"B23883FF";
    when 16#00AA4# => romdata <= X"762783DF";
    when 16#00AA5# => romdata <= X"3875892A";
    when 16#00AA6# => romdata <= X"76832A55";
    when 16#00AA7# => romdata <= X"5372802E";
    when 16#00AA8# => romdata <= X"BF387586";
    when 16#00AA9# => romdata <= X"2AB80554";
    when 16#00AAA# => romdata <= X"847327B4";
    when 16#00AAB# => romdata <= X"3880DB13";
    when 16#00AAC# => romdata <= X"54947327";
    when 16#00AAD# => romdata <= X"AB38758C";
    when 16#00AAE# => romdata <= X"2A80EE05";
    when 16#00AAF# => romdata <= X"5480D473";
    when 16#00AB0# => romdata <= X"279E3875";
    when 16#00AB1# => romdata <= X"8F2A80F7";
    when 16#00AB2# => romdata <= X"055482D4";
    when 16#00AB3# => romdata <= X"73279138";
    when 16#00AB4# => romdata <= X"75922A80";
    when 16#00AB5# => romdata <= X"FC05548A";
    when 16#00AB6# => romdata <= X"D4732784";
    when 16#00AB7# => romdata <= X"3880FE54";
    when 16#00AB8# => romdata <= X"73101010";
    when 16#00AB9# => romdata <= X"8183DC05";
    when 16#00ABA# => romdata <= X"88110856";
    when 16#00ABB# => romdata <= X"5874782E";
    when 16#00ABC# => romdata <= X"86CF3884";
    when 16#00ABD# => romdata <= X"1508FC06";
    when 16#00ABE# => romdata <= X"53757327";
    when 16#00ABF# => romdata <= X"8D388815";
    when 16#00AC0# => romdata <= X"08557478";
    when 16#00AC1# => romdata <= X"2E098106";
    when 16#00AC2# => romdata <= X"EA388C15";
    when 16#00AC3# => romdata <= X"088183DC";
    when 16#00AC4# => romdata <= X"0B840508";
    when 16#00AC5# => romdata <= X"718C1A0C";
    when 16#00AC6# => romdata <= X"76881A0C";
    when 16#00AC7# => romdata <= X"7888130C";
    when 16#00AC8# => romdata <= X"788C180C";
    when 16#00AC9# => romdata <= X"5D587953";
    when 16#00ACA# => romdata <= X"807A2483";
    when 16#00ACB# => romdata <= X"E6387282";
    when 16#00ACC# => romdata <= X"2C81712B";
    when 16#00ACD# => romdata <= X"5C537A7C";
    when 16#00ACE# => romdata <= X"26819838";
    when 16#00ACF# => romdata <= X"7B7B0653";
    when 16#00AD0# => romdata <= X"7282F138";
    when 16#00AD1# => romdata <= X"79FC0684";
    when 16#00AD2# => romdata <= X"055A7A10";
    when 16#00AD3# => romdata <= X"707D0654";
    when 16#00AD4# => romdata <= X"5B7282E0";
    when 16#00AD5# => romdata <= X"38841A5A";
    when 16#00AD6# => romdata <= X"F1398817";
    when 16#00AD7# => romdata <= X"8C110858";
    when 16#00AD8# => romdata <= X"5876782E";
    when 16#00AD9# => romdata <= X"098106FC";
    when 16#00ADA# => romdata <= X"C238821A";
    when 16#00ADB# => romdata <= X"5AFDEC39";
    when 16#00ADC# => romdata <= X"78177981";
    when 16#00ADD# => romdata <= X"0784190C";
    when 16#00ADE# => romdata <= X"708183F0";
    when 16#00ADF# => romdata <= X"0C708183";
    when 16#00AE0# => romdata <= X"EC0C8183";
    when 16#00AE1# => romdata <= X"E40B8C12";
    when 16#00AE2# => romdata <= X"0C8C1108";
    when 16#00AE3# => romdata <= X"88120C74";
    when 16#00AE4# => romdata <= X"81078412";
    when 16#00AE5# => romdata <= X"0C741175";
    when 16#00AE6# => romdata <= X"710C5153";
    when 16#00AE7# => romdata <= X"7D5187B7";
    when 16#00AE8# => romdata <= X"3F881754";
    when 16#00AE9# => romdata <= X"FCAC3981";
    when 16#00AEA# => romdata <= X"83DC0B84";
    when 16#00AEB# => romdata <= X"05087A54";
    when 16#00AEC# => romdata <= X"5C798025";
    when 16#00AED# => romdata <= X"FEF83882";
    when 16#00AEE# => romdata <= X"DA397A09";
    when 16#00AEF# => romdata <= X"7C067081";
    when 16#00AF0# => romdata <= X"83DC0B84";
    when 16#00AF1# => romdata <= X"050C5C7A";
    when 16#00AF2# => romdata <= X"105B7A7C";
    when 16#00AF3# => romdata <= X"2685387A";
    when 16#00AF4# => romdata <= X"85B83881";
    when 16#00AF5# => romdata <= X"83DC0B88";
    when 16#00AF6# => romdata <= X"05087084";
    when 16#00AF7# => romdata <= X"1208FC06";
    when 16#00AF8# => romdata <= X"707C317C";
    when 16#00AF9# => romdata <= X"72268F72";
    when 16#00AFA# => romdata <= X"25075757";
    when 16#00AFB# => romdata <= X"5C5D5572";
    when 16#00AFC# => romdata <= X"802E80DB";
    when 16#00AFD# => romdata <= X"38797A16";
    when 16#00AFE# => romdata <= X"8183D408";
    when 16#00AFF# => romdata <= X"1B90115A";
    when 16#00B00# => romdata <= X"55575B81";
    when 16#00B01# => romdata <= X"83D008FF";
    when 16#00B02# => romdata <= X"2E8838A0";
    when 16#00B03# => romdata <= X"8F13E080";
    when 16#00B04# => romdata <= X"06577652";
    when 16#00B05# => romdata <= X"7D5186C0";
    when 16#00B06# => romdata <= X"3FB00854";
    when 16#00B07# => romdata <= X"B008FF2E";
    when 16#00B08# => romdata <= X"9038B008";
    when 16#00B09# => romdata <= X"76278299";
    when 16#00B0A# => romdata <= X"38748183";
    when 16#00B0B# => romdata <= X"DC2E8291";
    when 16#00B0C# => romdata <= X"388183DC";
    when 16#00B0D# => romdata <= X"0B880508";
    when 16#00B0E# => romdata <= X"55841508";
    when 16#00B0F# => romdata <= X"FC06707A";
    when 16#00B10# => romdata <= X"317A7226";
    when 16#00B11# => romdata <= X"8F722507";
    when 16#00B12# => romdata <= X"52555372";
    when 16#00B13# => romdata <= X"83E63874";
    when 16#00B14# => romdata <= X"79810784";
    when 16#00B15# => romdata <= X"170C7916";
    when 16#00B16# => romdata <= X"708183DC";
    when 16#00B17# => romdata <= X"0B88050C";
    when 16#00B18# => romdata <= X"75810784";
    when 16#00B19# => romdata <= X"120C547E";
    when 16#00B1A# => romdata <= X"525785EB";
    when 16#00B1B# => romdata <= X"3F881754";
    when 16#00B1C# => romdata <= X"FAE03975";
    when 16#00B1D# => romdata <= X"832A7054";
    when 16#00B1E# => romdata <= X"54807424";
    when 16#00B1F# => romdata <= X"819B3872";
    when 16#00B20# => romdata <= X"822C8171";
    when 16#00B21# => romdata <= X"2B8183E0";
    when 16#00B22# => romdata <= X"08077081";
    when 16#00B23# => romdata <= X"83DC0B84";
    when 16#00B24# => romdata <= X"050C7510";
    when 16#00B25# => romdata <= X"10108183";
    when 16#00B26# => romdata <= X"DC058811";
    when 16#00B27# => romdata <= X"08585A5D";
    when 16#00B28# => romdata <= X"53778C18";
    when 16#00B29# => romdata <= X"0C748818";
    when 16#00B2A# => romdata <= X"0C768819";
    when 16#00B2B# => romdata <= X"0C768C16";
    when 16#00B2C# => romdata <= X"0CFCF339";
    when 16#00B2D# => romdata <= X"797A1010";
    when 16#00B2E# => romdata <= X"108183DC";
    when 16#00B2F# => romdata <= X"05705759";
    when 16#00B30# => romdata <= X"5D8C1508";
    when 16#00B31# => romdata <= X"5776752E";
    when 16#00B32# => romdata <= X"A3388417";
    when 16#00B33# => romdata <= X"08FC0670";
    when 16#00B34# => romdata <= X"7A315556";
    when 16#00B35# => romdata <= X"738F2483";
    when 16#00B36# => romdata <= X"CA387380";
    when 16#00B37# => romdata <= X"25848138";
    when 16#00B38# => romdata <= X"8C170857";
    when 16#00B39# => romdata <= X"76752E09";
    when 16#00B3A# => romdata <= X"8106DF38";
    when 16#00B3B# => romdata <= X"8815811B";
    when 16#00B3C# => romdata <= X"70830655";
    when 16#00B3D# => romdata <= X"5B5572C9";
    when 16#00B3E# => romdata <= X"387C8306";
    when 16#00B3F# => romdata <= X"5372802E";
    when 16#00B40# => romdata <= X"FDB838FF";
    when 16#00B41# => romdata <= X"1DF81959";
    when 16#00B42# => romdata <= X"5D881808";
    when 16#00B43# => romdata <= X"782EEA38";
    when 16#00B44# => romdata <= X"FDB53983";
    when 16#00B45# => romdata <= X"1A53FC96";
    when 16#00B46# => romdata <= X"39831470";
    when 16#00B47# => romdata <= X"822C8171";
    when 16#00B48# => romdata <= X"2B8183E0";
    when 16#00B49# => romdata <= X"08077081";
    when 16#00B4A# => romdata <= X"83DC0B84";
    when 16#00B4B# => romdata <= X"050C7610";
    when 16#00B4C# => romdata <= X"10108183";
    when 16#00B4D# => romdata <= X"DC058811";
    when 16#00B4E# => romdata <= X"08595B5E";
    when 16#00B4F# => romdata <= X"5153FEE1";
    when 16#00B50# => romdata <= X"398183A0";
    when 16#00B51# => romdata <= X"081758B0";
    when 16#00B52# => romdata <= X"08762E81";
    when 16#00B53# => romdata <= X"8D388183";
    when 16#00B54# => romdata <= X"D008FF2E";
    when 16#00B55# => romdata <= X"83EC3873";
    when 16#00B56# => romdata <= X"76311881";
    when 16#00B57# => romdata <= X"83A00C73";
    when 16#00B58# => romdata <= X"87067057";
    when 16#00B59# => romdata <= X"5372802E";
    when 16#00B5A# => romdata <= X"88388873";
    when 16#00B5B# => romdata <= X"31701555";
    when 16#00B5C# => romdata <= X"5676149F";
    when 16#00B5D# => romdata <= X"FF06A080";
    when 16#00B5E# => romdata <= X"71311770";
    when 16#00B5F# => romdata <= X"547F5357";
    when 16#00B60# => romdata <= X"5383D53F";
    when 16#00B61# => romdata <= X"B00853B0";
    when 16#00B62# => romdata <= X"08FF2E81";
    when 16#00B63# => romdata <= X"A0388183";
    when 16#00B64# => romdata <= X"A0081670";
    when 16#00B65# => romdata <= X"8183A00C";
    when 16#00B66# => romdata <= X"74758183";
    when 16#00B67# => romdata <= X"DC0B8805";
    when 16#00B68# => romdata <= X"0C747631";
    when 16#00B69# => romdata <= X"18708107";
    when 16#00B6A# => romdata <= X"51555658";
    when 16#00B6B# => romdata <= X"7B8183DC";
    when 16#00B6C# => romdata <= X"2E839C38";
    when 16#00B6D# => romdata <= X"798F2682";
    when 16#00B6E# => romdata <= X"CB38810B";
    when 16#00B6F# => romdata <= X"84150C84";
    when 16#00B70# => romdata <= X"1508FC06";
    when 16#00B71# => romdata <= X"707A317A";
    when 16#00B72# => romdata <= X"72268F72";
    when 16#00B73# => romdata <= X"25075255";
    when 16#00B74# => romdata <= X"5372802E";
    when 16#00B75# => romdata <= X"FCF93880";
    when 16#00B76# => romdata <= X"DB39B008";
    when 16#00B77# => romdata <= X"9FFF0653";
    when 16#00B78# => romdata <= X"72FEEB38";
    when 16#00B79# => romdata <= X"778183A0";
    when 16#00B7A# => romdata <= X"0C8183DC";
    when 16#00B7B# => romdata <= X"0B880508";
    when 16#00B7C# => romdata <= X"7B188107";
    when 16#00B7D# => romdata <= X"84120C55";
    when 16#00B7E# => romdata <= X"8183CC08";
    when 16#00B7F# => romdata <= X"78278638";
    when 16#00B80# => romdata <= X"778183CC";
    when 16#00B81# => romdata <= X"0C8183C8";
    when 16#00B82# => romdata <= X"087827FC";
    when 16#00B83# => romdata <= X"AC387781";
    when 16#00B84# => romdata <= X"83C80C84";
    when 16#00B85# => romdata <= X"1508FC06";
    when 16#00B86# => romdata <= X"707A317A";
    when 16#00B87# => romdata <= X"72268F72";
    when 16#00B88# => romdata <= X"25075255";
    when 16#00B89# => romdata <= X"5372802E";
    when 16#00B8A# => romdata <= X"FCA53888";
    when 16#00B8B# => romdata <= X"39807454";
    when 16#00B8C# => romdata <= X"56FEDB39";
    when 16#00B8D# => romdata <= X"7D51829F";
    when 16#00B8E# => romdata <= X"3F800BB0";
    when 16#00B8F# => romdata <= X"0C8F3D0D";
    when 16#00B90# => romdata <= X"04735380";
    when 16#00B91# => romdata <= X"7424A938";
    when 16#00B92# => romdata <= X"72822C81";
    when 16#00B93# => romdata <= X"712B8183";
    when 16#00B94# => romdata <= X"E0080770";
    when 16#00B95# => romdata <= X"8183DC0B";
    when 16#00B96# => romdata <= X"84050C5D";
    when 16#00B97# => romdata <= X"53778C18";
    when 16#00B98# => romdata <= X"0C748818";
    when 16#00B99# => romdata <= X"0C768819";
    when 16#00B9A# => romdata <= X"0C768C16";
    when 16#00B9B# => romdata <= X"0CF9B739";
    when 16#00B9C# => romdata <= X"83147082";
    when 16#00B9D# => romdata <= X"2C81712B";
    when 16#00B9E# => romdata <= X"8183E008";
    when 16#00B9F# => romdata <= X"07708183";
    when 16#00BA0# => romdata <= X"DC0B8405";
    when 16#00BA1# => romdata <= X"0C5E5153";
    when 16#00BA2# => romdata <= X"D4397B7B";
    when 16#00BA3# => romdata <= X"065372FC";
    when 16#00BA4# => romdata <= X"A338841A";
    when 16#00BA5# => romdata <= X"7B105C5A";
    when 16#00BA6# => romdata <= X"F139FF1A";
    when 16#00BA7# => romdata <= X"8111515A";
    when 16#00BA8# => romdata <= X"F7B93978";
    when 16#00BA9# => romdata <= X"17798107";
    when 16#00BAA# => romdata <= X"84190C8C";
    when 16#00BAB# => romdata <= X"18088819";
    when 16#00BAC# => romdata <= X"08718C12";
    when 16#00BAD# => romdata <= X"0C88120C";
    when 16#00BAE# => romdata <= X"59708183";
    when 16#00BAF# => romdata <= X"F00C7081";
    when 16#00BB0# => romdata <= X"83EC0C81";
    when 16#00BB1# => romdata <= X"83E40B8C";
    when 16#00BB2# => romdata <= X"120C8C11";
    when 16#00BB3# => romdata <= X"0888120C";
    when 16#00BB4# => romdata <= X"74810784";
    when 16#00BB5# => romdata <= X"120C7411";
    when 16#00BB6# => romdata <= X"75710C51";
    when 16#00BB7# => romdata <= X"53F9BD39";
    when 16#00BB8# => romdata <= X"75178411";
    when 16#00BB9# => romdata <= X"08810784";
    when 16#00BBA# => romdata <= X"120C538C";
    when 16#00BBB# => romdata <= X"17088818";
    when 16#00BBC# => romdata <= X"08718C12";
    when 16#00BBD# => romdata <= X"0C88120C";
    when 16#00BBE# => romdata <= X"587D5180";
    when 16#00BBF# => romdata <= X"DA3F8817";
    when 16#00BC0# => romdata <= X"54F5CF39";
    when 16#00BC1# => romdata <= X"7284150C";
    when 16#00BC2# => romdata <= X"F41AF806";
    when 16#00BC3# => romdata <= X"70841E08";
    when 16#00BC4# => romdata <= X"81060784";
    when 16#00BC5# => romdata <= X"1E0C701D";
    when 16#00BC6# => romdata <= X"545B850B";
    when 16#00BC7# => romdata <= X"84140C85";
    when 16#00BC8# => romdata <= X"0B88140C";
    when 16#00BC9# => romdata <= X"8F7B27FD";
    when 16#00BCA# => romdata <= X"CF38881C";
    when 16#00BCB# => romdata <= X"527D5182";
    when 16#00BCC# => romdata <= X"903F8183";
    when 16#00BCD# => romdata <= X"DC0B8805";
    when 16#00BCE# => romdata <= X"088183A0";
    when 16#00BCF# => romdata <= X"085955FD";
    when 16#00BD0# => romdata <= X"B7397781";
    when 16#00BD1# => romdata <= X"83A00C73";
    when 16#00BD2# => romdata <= X"8183D00C";
    when 16#00BD3# => romdata <= X"FC913972";
    when 16#00BD4# => romdata <= X"84150CFD";
    when 16#00BD5# => romdata <= X"A3390404";
    when 16#00BD6# => romdata <= X"FD3D0D80";
    when 16#00BD7# => romdata <= X"0B81A4BC";
    when 16#00BD8# => romdata <= X"0C765186";
    when 16#00BD9# => romdata <= X"CB3FB008";
    when 16#00BDA# => romdata <= X"53B008FF";
    when 16#00BDB# => romdata <= X"2E883872";
    when 16#00BDC# => romdata <= X"B00C853D";
    when 16#00BDD# => romdata <= X"0D0481A4";
    when 16#00BDE# => romdata <= X"BC085473";
    when 16#00BDF# => romdata <= X"802EF038";
    when 16#00BE0# => romdata <= X"7574710C";
    when 16#00BE1# => romdata <= X"5272B00C";
    when 16#00BE2# => romdata <= X"853D0D04";
    when 16#00BE3# => romdata <= X"FB3D0D77";
    when 16#00BE4# => romdata <= X"705256C2";
    when 16#00BE5# => romdata <= X"3F8183DC";
    when 16#00BE6# => romdata <= X"0B880508";
    when 16#00BE7# => romdata <= X"841108FC";
    when 16#00BE8# => romdata <= X"06707B31";
    when 16#00BE9# => romdata <= X"9FEF05E0";
    when 16#00BEA# => romdata <= X"8006E080";
    when 16#00BEB# => romdata <= X"05565653";
    when 16#00BEC# => romdata <= X"A0807424";
    when 16#00BED# => romdata <= X"94388052";
    when 16#00BEE# => romdata <= X"7551FF9C";
    when 16#00BEF# => romdata <= X"3F8183E4";
    when 16#00BF0# => romdata <= X"08155372";
    when 16#00BF1# => romdata <= X"B0082E8F";
    when 16#00BF2# => romdata <= X"387551FF";
    when 16#00BF3# => romdata <= X"8A3F8053";
    when 16#00BF4# => romdata <= X"72B00C87";
    when 16#00BF5# => romdata <= X"3D0D0473";
    when 16#00BF6# => romdata <= X"30527551";
    when 16#00BF7# => romdata <= X"FEFA3FB0";
    when 16#00BF8# => romdata <= X"08FF2EA8";
    when 16#00BF9# => romdata <= X"388183DC";
    when 16#00BFA# => romdata <= X"0B880508";
    when 16#00BFB# => romdata <= X"75753181";
    when 16#00BFC# => romdata <= X"0784120C";
    when 16#00BFD# => romdata <= X"538183A0";
    when 16#00BFE# => romdata <= X"08743181";
    when 16#00BFF# => romdata <= X"83A00C75";
    when 16#00C00# => romdata <= X"51FED43F";
    when 16#00C01# => romdata <= X"810BB00C";
    when 16#00C02# => romdata <= X"873D0D04";
    when 16#00C03# => romdata <= X"80527551";
    when 16#00C04# => romdata <= X"FEC63F81";
    when 16#00C05# => romdata <= X"83DC0B88";
    when 16#00C06# => romdata <= X"0508B008";
    when 16#00C07# => romdata <= X"71315653";
    when 16#00C08# => romdata <= X"8F7525FF";
    when 16#00C09# => romdata <= X"A438B008";
    when 16#00C0A# => romdata <= X"8183D008";
    when 16#00C0B# => romdata <= X"318183A0";
    when 16#00C0C# => romdata <= X"0C748107";
    when 16#00C0D# => romdata <= X"84140C75";
    when 16#00C0E# => romdata <= X"51FE9C3F";
    when 16#00C0F# => romdata <= X"8053FF90";
    when 16#00C10# => romdata <= X"39F63D0D";
    when 16#00C11# => romdata <= X"7C7E545B";
    when 16#00C12# => romdata <= X"72802E82";
    when 16#00C13# => romdata <= X"83387A51";
    when 16#00C14# => romdata <= X"FE843FF8";
    when 16#00C15# => romdata <= X"13841108";
    when 16#00C16# => romdata <= X"70FE0670";
    when 16#00C17# => romdata <= X"13841108";
    when 16#00C18# => romdata <= X"FC065D58";
    when 16#00C19# => romdata <= X"59545881";
    when 16#00C1A# => romdata <= X"83E40875";
    when 16#00C1B# => romdata <= X"2E82DE38";
    when 16#00C1C# => romdata <= X"7884160C";
    when 16#00C1D# => romdata <= X"80738106";
    when 16#00C1E# => romdata <= X"545A727A";
    when 16#00C1F# => romdata <= X"2E81D538";
    when 16#00C20# => romdata <= X"78158411";
    when 16#00C21# => romdata <= X"08810651";
    when 16#00C22# => romdata <= X"5372A038";
    when 16#00C23# => romdata <= X"78175779";
    when 16#00C24# => romdata <= X"81E63888";
    when 16#00C25# => romdata <= X"15085372";
    when 16#00C26# => romdata <= X"8183E42E";
    when 16#00C27# => romdata <= X"82F9388C";
    when 16#00C28# => romdata <= X"1508708C";
    when 16#00C29# => romdata <= X"150C7388";
    when 16#00C2A# => romdata <= X"120C5676";
    when 16#00C2B# => romdata <= X"81078419";
    when 16#00C2C# => romdata <= X"0C761877";
    when 16#00C2D# => romdata <= X"710C5379";
    when 16#00C2E# => romdata <= X"81913883";
    when 16#00C2F# => romdata <= X"FF772781";
    when 16#00C30# => romdata <= X"C8387689";
    when 16#00C31# => romdata <= X"2A77832A";
    when 16#00C32# => romdata <= X"56537280";
    when 16#00C33# => romdata <= X"2EBF3876";
    when 16#00C34# => romdata <= X"862AB805";
    when 16#00C35# => romdata <= X"55847327";
    when 16#00C36# => romdata <= X"B43880DB";
    when 16#00C37# => romdata <= X"13559473";
    when 16#00C38# => romdata <= X"27AB3876";
    when 16#00C39# => romdata <= X"8C2A80EE";
    when 16#00C3A# => romdata <= X"055580D4";
    when 16#00C3B# => romdata <= X"73279E38";
    when 16#00C3C# => romdata <= X"768F2A80";
    when 16#00C3D# => romdata <= X"F7055582";
    when 16#00C3E# => romdata <= X"D4732791";
    when 16#00C3F# => romdata <= X"3876922A";
    when 16#00C40# => romdata <= X"80FC0555";
    when 16#00C41# => romdata <= X"8AD47327";
    when 16#00C42# => romdata <= X"843880FE";
    when 16#00C43# => romdata <= X"55741010";
    when 16#00C44# => romdata <= X"108183DC";
    when 16#00C45# => romdata <= X"05881108";
    when 16#00C46# => romdata <= X"55567376";
    when 16#00C47# => romdata <= X"2E82B338";
    when 16#00C48# => romdata <= X"841408FC";
    when 16#00C49# => romdata <= X"06537673";
    when 16#00C4A# => romdata <= X"278D3888";
    when 16#00C4B# => romdata <= X"14085473";
    when 16#00C4C# => romdata <= X"762E0981";
    when 16#00C4D# => romdata <= X"06EA388C";
    when 16#00C4E# => romdata <= X"1408708C";
    when 16#00C4F# => romdata <= X"1A0C7488";
    when 16#00C50# => romdata <= X"1A0C7888";
    when 16#00C51# => romdata <= X"120C5677";
    when 16#00C52# => romdata <= X"8C150C7A";
    when 16#00C53# => romdata <= X"51FC883F";
    when 16#00C54# => romdata <= X"8C3D0D04";
    when 16#00C55# => romdata <= X"77087871";
    when 16#00C56# => romdata <= X"31597705";
    when 16#00C57# => romdata <= X"88190854";
    when 16#00C58# => romdata <= X"57728183";
    when 16#00C59# => romdata <= X"E42E80E0";
    when 16#00C5A# => romdata <= X"388C1808";
    when 16#00C5B# => romdata <= X"708C150C";
    when 16#00C5C# => romdata <= X"7388120C";
    when 16#00C5D# => romdata <= X"56FE8939";
    when 16#00C5E# => romdata <= X"8815088C";
    when 16#00C5F# => romdata <= X"1608708C";
    when 16#00C60# => romdata <= X"130C5788";
    when 16#00C61# => romdata <= X"170CFEA3";
    when 16#00C62# => romdata <= X"3976832A";
    when 16#00C63# => romdata <= X"70545580";
    when 16#00C64# => romdata <= X"75248198";
    when 16#00C65# => romdata <= X"3872822C";
    when 16#00C66# => romdata <= X"81712B81";
    when 16#00C67# => romdata <= X"83E00807";
    when 16#00C68# => romdata <= X"8183DC0B";
    when 16#00C69# => romdata <= X"84050C53";
    when 16#00C6A# => romdata <= X"74101010";
    when 16#00C6B# => romdata <= X"8183DC05";
    when 16#00C6C# => romdata <= X"88110855";
    when 16#00C6D# => romdata <= X"56758C19";
    when 16#00C6E# => romdata <= X"0C738819";
    when 16#00C6F# => romdata <= X"0C778817";
    when 16#00C70# => romdata <= X"0C778C15";
    when 16#00C71# => romdata <= X"0CFF8439";
    when 16#00C72# => romdata <= X"815AFDB4";
    when 16#00C73# => romdata <= X"39781773";
    when 16#00C74# => romdata <= X"81065457";
    when 16#00C75# => romdata <= X"72983877";
    when 16#00C76# => romdata <= X"08787131";
    when 16#00C77# => romdata <= X"5977058C";
    when 16#00C78# => romdata <= X"1908881A";
    when 16#00C79# => romdata <= X"08718C12";
    when 16#00C7A# => romdata <= X"0C88120C";
    when 16#00C7B# => romdata <= X"57577681";
    when 16#00C7C# => romdata <= X"0784190C";
    when 16#00C7D# => romdata <= X"778183DC";
    when 16#00C7E# => romdata <= X"0B88050C";
    when 16#00C7F# => romdata <= X"8183D808";
    when 16#00C80# => romdata <= X"7726FEC7";
    when 16#00C81# => romdata <= X"388183D4";
    when 16#00C82# => romdata <= X"08527A51";
    when 16#00C83# => romdata <= X"FAFE3F7A";
    when 16#00C84# => romdata <= X"51FAC43F";
    when 16#00C85# => romdata <= X"FEBA3981";
    when 16#00C86# => romdata <= X"788C150C";
    when 16#00C87# => romdata <= X"7888150C";
    when 16#00C88# => romdata <= X"738C1A0C";
    when 16#00C89# => romdata <= X"73881A0C";
    when 16#00C8A# => romdata <= X"5AFD8039";
    when 16#00C8B# => romdata <= X"83157082";
    when 16#00C8C# => romdata <= X"2C81712B";
    when 16#00C8D# => romdata <= X"8183E008";
    when 16#00C8E# => romdata <= X"078183DC";
    when 16#00C8F# => romdata <= X"0B84050C";
    when 16#00C90# => romdata <= X"51537410";
    when 16#00C91# => romdata <= X"10108183";
    when 16#00C92# => romdata <= X"DC058811";
    when 16#00C93# => romdata <= X"085556FE";
    when 16#00C94# => romdata <= X"E4397453";
    when 16#00C95# => romdata <= X"807524A7";
    when 16#00C96# => romdata <= X"3872822C";
    when 16#00C97# => romdata <= X"81712B81";
    when 16#00C98# => romdata <= X"83E00807";
    when 16#00C99# => romdata <= X"8183DC0B";
    when 16#00C9A# => romdata <= X"84050C53";
    when 16#00C9B# => romdata <= X"758C190C";
    when 16#00C9C# => romdata <= X"7388190C";
    when 16#00C9D# => romdata <= X"7788170C";
    when 16#00C9E# => romdata <= X"778C150C";
    when 16#00C9F# => romdata <= X"FDCD3983";
    when 16#00CA0# => romdata <= X"1570822C";
    when 16#00CA1# => romdata <= X"81712B81";
    when 16#00CA2# => romdata <= X"83E00807";
    when 16#00CA3# => romdata <= X"8183DC0B";
    when 16#00CA4# => romdata <= X"84050C51";
    when 16#00CA5# => romdata <= X"53D63981";
    when 16#00CA6# => romdata <= X"0BB00C04";
    when 16#00CA7# => romdata <= X"803D0D72";
    when 16#00CA8# => romdata <= X"812E8938";
    when 16#00CA9# => romdata <= X"800BB00C";
    when 16#00CAA# => romdata <= X"823D0D04";
    when 16#00CAB# => romdata <= X"7351B23F";
    when 16#00CAC# => romdata <= X"FE3D0D81";
    when 16#00CAD# => romdata <= X"A4B80851";
    when 16#00CAE# => romdata <= X"708A3881";
    when 16#00CAF# => romdata <= X"A4C07081";
    when 16#00CB0# => romdata <= X"A4B80C51";
    when 16#00CB1# => romdata <= X"70751252";
    when 16#00CB2# => romdata <= X"52FF5370";
    when 16#00CB3# => romdata <= X"87FB8080";
    when 16#00CB4# => romdata <= X"26883870";
    when 16#00CB5# => romdata <= X"81A4B80C";
    when 16#00CB6# => romdata <= X"715372B0";
    when 16#00CB7# => romdata <= X"0C843D0D";
    when 16#00CB8# => romdata <= X"0400FF39";
    when 16#00CB9# => romdata <= X"68656C70";
    when 16#00CBA# => romdata <= X"00000000";
    when 16#00CBB# => romdata <= X"73797374";
    when 16#00CBC# => romdata <= X"656D2072";
    when 16#00CBD# => romdata <= X"65736574";
    when 16#00CBE# => romdata <= X"00000000";
    when 16#00CBF# => romdata <= X"72657365";
    when 16#00CC0# => romdata <= X"74000000";
    when 16#00CC1# => romdata <= X"73686F77";
    when 16#00CC2# => romdata <= X"20737973";
    when 16#00CC3# => romdata <= X"74656D20";
    when 16#00CC4# => romdata <= X"696E666F";
    when 16#00CC5# => romdata <= X"203C7665";
    when 16#00CC6# => romdata <= X"72626F73";
    when 16#00CC7# => romdata <= X"653E0000";
    when 16#00CC8# => romdata <= X"73797369";
    when 16#00CC9# => romdata <= X"6E666F00";
    when 16#00CCA# => romdata <= X"72656E61";
    when 16#00CCB# => romdata <= X"20636F6E";
    when 16#00CCC# => romdata <= X"74726F6C";
    when 16#00CCD# => romdata <= X"6C657220";
    when 16#00CCE# => romdata <= X"73746174";
    when 16#00CCF# => romdata <= X"75730000";
    when 16#00CD0# => romdata <= X"72656E61";
    when 16#00CD1# => romdata <= X"20737461";
    when 16#00CD2# => romdata <= X"74757300";
    when 16#00CD3# => romdata <= X"3C636861";
    when 16#00CD4# => romdata <= X"6E6E656C";
    when 16#00CD5# => romdata <= X"3E203C68";
    when 16#00CD6# => romdata <= X"6967683E";
    when 16#00CD7# => romdata <= X"203C6C6F";
    when 16#00CD8# => romdata <= X"775F636F";
    when 16#00CD9# => romdata <= X"6E666967";
    when 16#00CDA# => romdata <= X"3E000000";
    when 16#00CDB# => romdata <= X"636F6E66";
    when 16#00CDC# => romdata <= X"69670000";
    when 16#00CDD# => romdata <= X"646F2063";
    when 16#00CDE# => romdata <= X"6F6D706C";
    when 16#00CDF# => romdata <= X"65746520";
    when 16#00CE0# => romdata <= X"64656D6F";
    when 16#00CE1# => romdata <= X"20636F6E";
    when 16#00CE2# => romdata <= X"66696720";
    when 16#00CE3# => romdata <= X"666F7220";
    when 16#00CE4# => romdata <= X"52454E41";
    when 16#00CE5# => romdata <= X"00000000";
    when 16#00CE6# => romdata <= X"64656D6F";
    when 16#00CE7# => romdata <= X"00000000";
    when 16#00CE8# => romdata <= X"73657420";
    when 16#00CE9# => romdata <= X"52454E41";
    when 16#00CEA# => romdata <= X"20746F20";
    when 16#00CEB# => romdata <= X"706F7765";
    when 16#00CEC# => romdata <= X"7220646F";
    when 16#00CED# => romdata <= X"776E206D";
    when 16#00CEE# => romdata <= X"6F646500";
    when 16#00CEF# => romdata <= X"706F6666";
    when 16#00CF0# => romdata <= X"00000000";
    when 16#00CF1# => romdata <= X"73657420";
    when 16#00CF2# => romdata <= X"72656E61";
    when 16#00CF3# => romdata <= X"20636861";
    when 16#00CF4# => romdata <= X"6E6E656C";
    when 16#00CF5# => romdata <= X"20302074";
    when 16#00CF6# => romdata <= X"6F20666F";
    when 16#00CF7# => romdata <= X"6C6C6F77";
    when 16#00CF8# => romdata <= X"6572206D";
    when 16#00CF9# => romdata <= X"6F646500";
    when 16#00CFA# => romdata <= X"666F6C6C";
    when 16#00CFB# => romdata <= X"6F770000";
    when 16#00CFC# => romdata <= X"3C74696D";
    when 16#00CFD# => romdata <= X"653E2061";
    when 16#00CFE# => romdata <= X"63746976";
    when 16#00CFF# => romdata <= X"61746520";
    when 16#00D00# => romdata <= X"52454E41";
    when 16#00D01# => romdata <= X"00000000";
    when 16#00D02# => romdata <= X"61637175";
    when 16#00D03# => romdata <= X"69726500";
    when 16#00D04# => romdata <= X"73657420";
    when 16#00D05# => romdata <= X"52454E41";
    when 16#00D06# => romdata <= X"20636F6E";
    when 16#00D07# => romdata <= X"74726F6C";
    when 16#00D08# => romdata <= X"6C657220";
    when 16#00D09# => romdata <= X"746F2049";
    when 16#00D0A# => romdata <= X"444C4500";
    when 16#00D0B# => romdata <= X"73746F70";
    when 16#00D0C# => romdata <= X"00000000";
    when 16#00D0D# => romdata <= X"7072696E";
    when 16#00D0E# => romdata <= X"74207472";
    when 16#00D0F# => romdata <= X"69676765";
    when 16#00D10# => romdata <= X"72206368";
    when 16#00D11# => romdata <= X"61696E73";
    when 16#00D12# => romdata <= X"00000000";
    when 16#00D13# => romdata <= X"63686169";
    when 16#00D14# => romdata <= X"6E730000";
    when 16#00D15# => romdata <= X"7072696E";
    when 16#00D16# => romdata <= X"74207361";
    when 16#00D17# => romdata <= X"6D706C65";
    when 16#00D18# => romdata <= X"64205245";
    when 16#00D19# => romdata <= X"4E412074";
    when 16#00D1A# => romdata <= X"6F6B656E";
    when 16#00D1B# => romdata <= X"73000000";
    when 16#00D1C# => romdata <= X"746F6B65";
    when 16#00D1D# => romdata <= X"6E000000";
    when 16#00D1E# => romdata <= X"74726F75";
    when 16#00D1F# => romdata <= X"626C6573";
    when 16#00D20# => romdata <= X"65617263";
    when 16#00D21# => romdata <= X"68205245";
    when 16#00D22# => romdata <= X"4E410000";
    when 16#00D23# => romdata <= X"74726F75";
    when 16#00D24# => romdata <= X"626C6500";
    when 16#00D25# => romdata <= X"696E6974";
    when 16#00D26# => romdata <= X"616C697A";
    when 16#00D27# => romdata <= X"65204444";
    when 16#00D28# => romdata <= X"53206368";
    when 16#00D29# => romdata <= X"6970203C";
    when 16#00D2A# => romdata <= X"66726571";
    when 16#00D2B# => romdata <= X"2074756E";
    when 16#00D2C# => romdata <= X"696E6720";
    when 16#00D2D# => romdata <= X"776F7264";
    when 16#00D2E# => romdata <= X"3E000000";
    when 16#00D2F# => romdata <= X"64647369";
    when 16#00D30# => romdata <= X"6E697400";
    when 16#00D31# => romdata <= X"72656164";
    when 16#00D32# => romdata <= X"20646473";
    when 16#00D33# => romdata <= X"20726567";
    when 16#00D34# => romdata <= X"69737465";
    when 16#00D35# => romdata <= X"72730000";
    when 16#00D36# => romdata <= X"64647369";
    when 16#00D37# => romdata <= X"6E666F00";
    when 16#00D38# => romdata <= X"72756E6E";
    when 16#00D39# => romdata <= X"696E6720";
    when 16#00D3A# => romdata <= X"6C696768";
    when 16#00D3B# => romdata <= X"74000000";
    when 16#00D3C# => romdata <= X"72756E00";
    when 16#00D3D# => romdata <= X"63686563";
    when 16#00D3E# => romdata <= X"6B204932";
    when 16#00D3F# => romdata <= X"43206164";
    when 16#00D40# => romdata <= X"64726573";
    when 16#00D41# => romdata <= X"73000000";
    when 16#00D42# => romdata <= X"69326300";
    when 16#00D43# => romdata <= X"72656164";
    when 16#00D44# => romdata <= X"20454550";
    when 16#00D45# => romdata <= X"524F4D20";
    when 16#00D46# => romdata <= X"3C627573";
    when 16#00D47# => romdata <= X"3E203C69";
    when 16#00D48# => romdata <= X"32635F61";
    when 16#00D49# => romdata <= X"6464723E";
    when 16#00D4A# => romdata <= X"203C6C65";
    when 16#00D4B# => romdata <= X"6E677468";
    when 16#00D4C# => romdata <= X"3E000000";
    when 16#00D4D# => romdata <= X"65657072";
    when 16#00D4E# => romdata <= X"6F6D0000";
    when 16#00D4F# => romdata <= X"72656164";
    when 16#00D50# => romdata <= X"20616463";
    when 16#00D51# => romdata <= X"2076616C";
    when 16#00D52# => romdata <= X"75650000";
    when 16#00D53# => romdata <= X"61646300";
    when 16#00D54# => romdata <= X"67656E65";
    when 16#00D55# => romdata <= X"72617465";
    when 16#00D56# => romdata <= X"20746573";
    when 16#00D57# => romdata <= X"7420696D";
    when 16#00D58# => romdata <= X"70756C73";
    when 16#00D59# => romdata <= X"65000000";
    when 16#00D5A# => romdata <= X"74657374";
    when 16#00D5B# => romdata <= X"67656E00";
    when 16#00D5C# => romdata <= X"616C6961";
    when 16#00D5D# => romdata <= X"7320666F";
    when 16#00D5E# => romdata <= X"72207800";
    when 16#00D5F# => romdata <= X"6D656D00";
    when 16#00D60# => romdata <= X"77726974";
    when 16#00D61# => romdata <= X"6520776F";
    when 16#00D62# => romdata <= X"7264203C";
    when 16#00D63# => romdata <= X"61646472";
    when 16#00D64# => romdata <= X"3E203C6C";
    when 16#00D65# => romdata <= X"656E6774";
    when 16#00D66# => romdata <= X"683E203C";
    when 16#00D67# => romdata <= X"76616C75";
    when 16#00D68# => romdata <= X"65287329";
    when 16#00D69# => romdata <= X"3E000000";
    when 16#00D6A# => romdata <= X"776D656D";
    when 16#00D6B# => romdata <= X"00000000";
    when 16#00D6C# => romdata <= X"6558616D";
    when 16#00D6D# => romdata <= X"696E6520";
    when 16#00D6E# => romdata <= X"6D656D6F";
    when 16#00D6F# => romdata <= X"7279203C";
    when 16#00D70# => romdata <= X"61646472";
    when 16#00D71# => romdata <= X"3E203C6C";
    when 16#00D72# => romdata <= X"656E6774";
    when 16#00D73# => romdata <= X"683E0000";
    when 16#00D74# => romdata <= X"78000000";
    when 16#00D75# => romdata <= X"636C6561";
    when 16#00D76# => romdata <= X"72207363";
    when 16#00D77# => romdata <= X"7265656E";
    when 16#00D78# => romdata <= X"00000000";
    when 16#00D79# => romdata <= X"636C6561";
    when 16#00D7A# => romdata <= X"72000000";
    when 16#00D7B# => romdata <= X"0A0A0000";
    when 16#00D7C# => romdata <= X"72656E61";
    when 16#00D7D# => romdata <= X"3320636F";
    when 16#00D7E# => romdata <= X"6E74726F";
    when 16#00D7F# => romdata <= X"6C6C6572";
    when 16#00D80# => romdata <= X"20626F61";
    when 16#00D81# => romdata <= X"72640000";
    when 16#00D82# => romdata <= X"20286F6E";
    when 16#00D83# => romdata <= X"2073696D";
    when 16#00D84# => romdata <= X"290A0000";
    when 16#00D85# => romdata <= X"0A485720";
    when 16#00D86# => romdata <= X"73796E74";
    when 16#00D87# => romdata <= X"68657369";
    when 16#00D88# => romdata <= X"7A65643A";
    when 16#00D89# => romdata <= X"20000000";
    when 16#00D8A# => romdata <= X"0A535720";
    when 16#00D8B# => romdata <= X"636F6D70";
    when 16#00D8C# => romdata <= X"696C6564";
    when 16#00D8D# => romdata <= X"2020203A";
    when 16#00D8E# => romdata <= X"20446563";
    when 16#00D8F# => romdata <= X"20323120";
    when 16#00D90# => romdata <= X"32303131";
    when 16#00D91# => romdata <= X"20203135";
    when 16#00D92# => romdata <= X"3A30303A";
    when 16#00D93# => romdata <= X"35390000";
    when 16#00D94# => romdata <= X"0A737973";
    when 16#00D95# => romdata <= X"74656D20";
    when 16#00D96# => romdata <= X"636C6F63";
    when 16#00D97# => romdata <= X"6B20203A";
    when 16#00D98# => romdata <= X"20000000";
    when 16#00D99# => romdata <= X"204D487A";
    when 16#00D9A# => romdata <= X"0A000000";
    when 16#00D9B# => romdata <= X"44454255";
    when 16#00D9C# => romdata <= X"47204D4F";
    when 16#00D9D# => romdata <= X"44450000";
    when 16#00D9E# => romdata <= X"204F4E0A";
    when 16#00D9F# => romdata <= X"00000000";
    when 16#00DA0# => romdata <= X"4552524F";
    when 16#00DA1# => romdata <= X"523A2074";
    when 16#00DA2# => romdata <= X"6F6F206D";
    when 16#00DA3# => romdata <= X"75636820";
    when 16#00DA4# => romdata <= X"636F6D6D";
    when 16#00DA5# => romdata <= X"616E6473";
    when 16#00DA6# => romdata <= X"2E0A0000";
    when 16#00DA7# => romdata <= X"3E200000";
    when 16#00DA8# => romdata <= X"636F6D6D";
    when 16#00DA9# => romdata <= X"616E6420";
    when 16#00DAA# => romdata <= X"6E6F7420";
    when 16#00DAB# => romdata <= X"666F756E";
    when 16#00DAC# => romdata <= X"642E0A00";
    when 16#00DAD# => romdata <= X"73757070";
    when 16#00DAE# => romdata <= X"6F727465";
    when 16#00DAF# => romdata <= X"6420636F";
    when 16#00DB0# => romdata <= X"6D6D616E";
    when 16#00DB1# => romdata <= X"64733A0A";
    when 16#00DB2# => romdata <= X"0A000000";
    when 16#00DB3# => romdata <= X"202D2000";
    when 16#00DB4# => romdata <= X"76656E64";
    when 16#00DB5# => romdata <= X"6F723F20";
    when 16#00DB6# => romdata <= X"20000000";
    when 16#00DB7# => romdata <= X"485A4452";
    when 16#00DB8# => romdata <= X"20202020";
    when 16#00DB9# => romdata <= X"20000000";
    when 16#00DBA# => romdata <= X"67616973";
    when 16#00DBB# => romdata <= X"6C657220";
    when 16#00DBC# => romdata <= X"20000000";
    when 16#00DBD# => romdata <= X"45534120";
    when 16#00DBE# => romdata <= X"20202020";
    when 16#00DBF# => romdata <= X"20000000";
    when 16#00DC0# => romdata <= X"756E6B6E";
    when 16#00DC1# => romdata <= X"6F776E20";
    when 16#00DC2# => romdata <= X"64657669";
    when 16#00DC3# => romdata <= X"63650000";
    when 16#00DC4# => romdata <= X"4C656F6E";
    when 16#00DC5# => romdata <= X"32204D65";
    when 16#00DC6# => romdata <= X"6D6F7279";
    when 16#00DC7# => romdata <= X"20436F6E";
    when 16#00DC8# => romdata <= X"74726F6C";
    when 16#00DC9# => romdata <= X"6C657200";
    when 16#00DCA# => romdata <= X"56474120";
    when 16#00DCB# => romdata <= X"636F6E74";
    when 16#00DCC# => romdata <= X"726F6C6C";
    when 16#00DCD# => romdata <= X"65720000";
    when 16#00DCE# => romdata <= X"53504920";
    when 16#00DCF# => romdata <= X"4D656D6F";
    when 16#00DD0# => romdata <= X"72792043";
    when 16#00DD1# => romdata <= X"6F6E7472";
    when 16#00DD2# => romdata <= X"6F6C6C65";
    when 16#00DD3# => romdata <= X"72000000";
    when 16#00DD4# => romdata <= X"53504920";
    when 16#00DD5# => romdata <= X"436F6E74";
    when 16#00DD6# => romdata <= X"726F6C6C";
    when 16#00DD7# => romdata <= X"65720000";
    when 16#00DD8# => romdata <= X"414D4241";
    when 16#00DD9# => romdata <= X"20577261";
    when 16#00DDA# => romdata <= X"70706572";
    when 16#00DDB# => romdata <= X"20666F72";
    when 16#00DDC# => romdata <= X"204F4320";
    when 16#00DDD# => romdata <= X"4932432D";
    when 16#00DDE# => romdata <= X"6D617374";
    when 16#00DDF# => romdata <= X"65720000";
    when 16#00DE0# => romdata <= X"47522031";
    when 16#00DE1# => romdata <= X"302F3130";
    when 16#00DE2# => romdata <= X"30204D62";
    when 16#00DE3# => romdata <= X"69742045";
    when 16#00DE4# => romdata <= X"74686572";
    when 16#00DE5# => romdata <= X"6E657420";
    when 16#00DE6# => romdata <= X"4D414300";
    when 16#00DE7# => romdata <= X"47656E65";
    when 16#00DE8# => romdata <= X"72616C20";
    when 16#00DE9# => romdata <= X"50757270";
    when 16#00DEA# => romdata <= X"6F736520";
    when 16#00DEB# => romdata <= X"492F4F20";
    when 16#00DEC# => romdata <= X"706F7274";
    when 16#00DED# => romdata <= X"00000000";
    when 16#00DEE# => romdata <= X"4D6F6475";
    when 16#00DEF# => romdata <= X"6C617220";
    when 16#00DF0# => romdata <= X"54696D65";
    when 16#00DF1# => romdata <= X"7220556E";
    when 16#00DF2# => romdata <= X"69740000";
    when 16#00DF3# => romdata <= X"4475616C";
    when 16#00DF4# => romdata <= X"2D706F72";
    when 16#00DF5# => romdata <= X"74204148";
    when 16#00DF6# => romdata <= X"42205352";
    when 16#00DF7# => romdata <= X"414D206D";
    when 16#00DF8# => romdata <= X"6F64756C";
    when 16#00DF9# => romdata <= X"65000000";
    when 16#00DFA# => romdata <= X"47656E65";
    when 16#00DFB# => romdata <= X"72696320";
    when 16#00DFC# => romdata <= X"55415254";
    when 16#00DFD# => romdata <= X"00000000";
    when 16#00DFE# => romdata <= X"4148422F";
    when 16#00DFF# => romdata <= X"41504220";
    when 16#00E00# => romdata <= X"42726964";
    when 16#00E01# => romdata <= X"67650000";
    when 16#00E02# => romdata <= X"64696666";
    when 16#00E03# => romdata <= X"6572656E";
    when 16#00E04# => romdata <= X"7469616C";
    when 16#00E05# => romdata <= X"20637572";
    when 16#00E06# => romdata <= X"72656E74";
    when 16#00E07# => romdata <= X"206D6F6E";
    when 16#00E08# => romdata <= X"69746F72";
    when 16#00E09# => romdata <= X"00000000";
    when 16#00E0A# => romdata <= X"64656275";
    when 16#00E0B# => romdata <= X"67207472";
    when 16#00E0C# => romdata <= X"61636572";
    when 16#00E0D# => romdata <= X"206D656D";
    when 16#00E0E# => romdata <= X"6F727900";
    when 16#00E0F# => romdata <= X"4541444F";
    when 16#00E10# => romdata <= X"47533130";
    when 16#00E11# => romdata <= X"32206469";
    when 16#00E12# => romdata <= X"73706C61";
    when 16#00E13# => romdata <= X"79206472";
    when 16#00E14# => romdata <= X"69766572";
    when 16#00E15# => romdata <= X"00000000";
    when 16#00E16# => romdata <= X"64656275";
    when 16#00E17# => romdata <= X"67206275";
    when 16#00E18# => romdata <= X"66666572";
    when 16#00E19# => romdata <= X"20636F6E";
    when 16#00E1A# => romdata <= X"74726F6C";
    when 16#00E1B# => romdata <= X"00000000";
    when 16#00E1C# => romdata <= X"52454E41";
    when 16#00E1D# => romdata <= X"3320636F";
    when 16#00E1E# => romdata <= X"6E74726F";
    when 16#00E1F# => romdata <= X"6C6C6572";
    when 16#00E20# => romdata <= X"00000000";
    when 16#00E21# => romdata <= X"53465020";
    when 16#00E22# => romdata <= X"636F6E74";
    when 16#00E23# => romdata <= X"726F6C6C";
    when 16#00E24# => romdata <= X"65720000";
    when 16#00E25# => romdata <= X"5A505520";
    when 16#00E26# => romdata <= X"4D656D6F";
    when 16#00E27# => romdata <= X"72792077";
    when 16#00E28# => romdata <= X"72617070";
    when 16#00E29# => romdata <= X"65720000";
    when 16#00E2A# => romdata <= X"5A505520";
    when 16#00E2B# => romdata <= X"41484220";
    when 16#00E2C# => romdata <= X"57726170";
    when 16#00E2D# => romdata <= X"70657200";
    when 16#00E2E# => romdata <= X"6265616D";
    when 16#00E2F# => romdata <= X"20706F73";
    when 16#00E30# => romdata <= X"6974696F";
    when 16#00E31# => romdata <= X"6E206D6F";
    when 16#00E32# => romdata <= X"6E69746F";
    when 16#00E33# => romdata <= X"72000000";
    when 16#00E34# => romdata <= X"74726967";
    when 16#00E35# => romdata <= X"67657220";
    when 16#00E36# => romdata <= X"67656E65";
    when 16#00E37# => romdata <= X"7261746F";
    when 16#00E38# => romdata <= X"72000000";
    when 16#00E39# => romdata <= X"64656275";
    when 16#00E3A# => romdata <= X"6720636F";
    when 16#00E3B# => romdata <= X"6E736F6C";
    when 16#00E3C# => romdata <= X"65000000";
    when 16#00E3D# => romdata <= X"44434D20";
    when 16#00E3E# => romdata <= X"70686173";
    when 16#00E3F# => romdata <= X"65207368";
    when 16#00E40# => romdata <= X"69667420";
    when 16#00E41# => romdata <= X"636F6E74";
    when 16#00E42# => romdata <= X"726F6C00";
    when 16#00E43# => romdata <= X"20206170";
    when 16#00E44# => romdata <= X"62736C76";
    when 16#00E45# => romdata <= X"00000000";
    when 16#00E46# => romdata <= X"76656E64";
    when 16#00E47# => romdata <= X"20307800";
    when 16#00E48# => romdata <= X"64657620";
    when 16#00E49# => romdata <= X"30780000";
    when 16#00E4A# => romdata <= X"76657220";
    when 16#00E4B# => romdata <= X"00000000";
    when 16#00E4C# => romdata <= X"69727120";
    when 16#00E4D# => romdata <= X"00000000";
    when 16#00E4E# => romdata <= X"61646472";
    when 16#00E4F# => romdata <= X"20307800";
    when 16#00E50# => romdata <= X"6168626D";
    when 16#00E51# => romdata <= X"73740000";
    when 16#00E52# => romdata <= X"61686273";
    when 16#00E53# => romdata <= X"6C760000";
    when 16#00E54# => romdata <= X"00000F46";
    when 16#00E55# => romdata <= X"00001017";
    when 16#00E56# => romdata <= X"0000100C";
    when 16#00E57# => romdata <= X"00001043";
    when 16#00E58# => romdata <= X"00001038";
    when 16#00E59# => romdata <= X"0000102D";
    when 16#00E5A# => romdata <= X"00001022";
    when 16#00E5B# => romdata <= X"00000FEB";
    when 16#00E5C# => romdata <= X"00000FE0";
    when 16#00E5D# => romdata <= X"00000FD5";
    when 16#00E5E# => romdata <= X"00000FCA";
    when 16#00E5F# => romdata <= X"00001001";
    when 16#00E60# => romdata <= X"00000FF6";
    when 16#00E61# => romdata <= X"00000FBF";
    when 16#00E62# => romdata <= X"00000F46";
    when 16#00E63# => romdata <= X"00000F46";
    when 16#00E64# => romdata <= X"00000F46";
    when 16#00E65# => romdata <= X"00000F46";
    when 16#00E66# => romdata <= X"00000F46";
    when 16#00E67# => romdata <= X"00000FB4";
    when 16#00E68# => romdata <= X"00000F46";
    when 16#00E69# => romdata <= X"00000F46";
    when 16#00E6A# => romdata <= X"00000FA9";
    when 16#00E6B# => romdata <= X"00000F46";
    when 16#00E6C# => romdata <= X"00000F9E";
    when 16#00E6D# => romdata <= X"00000F46";
    when 16#00E6E# => romdata <= X"00000F46";
    when 16#00E6F# => romdata <= X"00000F46";
    when 16#00E70# => romdata <= X"00000F46";
    when 16#00E71# => romdata <= X"00000F46";
    when 16#00E72# => romdata <= X"00000F46";
    when 16#00E73# => romdata <= X"00000F46";
    when 16#00E74# => romdata <= X"00000F46";
    when 16#00E75# => romdata <= X"00000F93";
    when 16#00E76# => romdata <= X"00000F46";
    when 16#00E77# => romdata <= X"00000F46";
    when 16#00E78# => romdata <= X"00000F88";
    when 16#00E79# => romdata <= X"00000F46";
    when 16#00E7A# => romdata <= X"00000F46";
    when 16#00E7B# => romdata <= X"00000F46";
    when 16#00E7C# => romdata <= X"00000F46";
    when 16#00E7D# => romdata <= X"00000F46";
    when 16#00E7E# => romdata <= X"00000F46";
    when 16#00E7F# => romdata <= X"00000F46";
    when 16#00E80# => romdata <= X"00000F46";
    when 16#00E81# => romdata <= X"00000F46";
    when 16#00E82# => romdata <= X"00000F46";
    when 16#00E83# => romdata <= X"00000F7D";
    when 16#00E84# => romdata <= X"00000F46";
    when 16#00E85# => romdata <= X"00000F46";
    when 16#00E86# => romdata <= X"00000F46";
    when 16#00E87# => romdata <= X"00000F46";
    when 16#00E88# => romdata <= X"00000F72";
    when 16#00E89# => romdata <= X"00000F46";
    when 16#00E8A# => romdata <= X"00000F46";
    when 16#00E8B# => romdata <= X"00000F46";
    when 16#00E8C# => romdata <= X"00000F46";
    when 16#00E8D# => romdata <= X"00000F46";
    when 16#00E8E# => romdata <= X"00000F46";
    when 16#00E8F# => romdata <= X"00000F46";
    when 16#00E90# => romdata <= X"00000F46";
    when 16#00E91# => romdata <= X"00000F46";
    when 16#00E92# => romdata <= X"00000F46";
    when 16#00E93# => romdata <= X"00000F46";
    when 16#00E94# => romdata <= X"00000F46";
    when 16#00E95# => romdata <= X"00000F46";
    when 16#00E96# => romdata <= X"00000F46";
    when 16#00E97# => romdata <= X"00000F46";
    when 16#00E98# => romdata <= X"00000F46";
    when 16#00E99# => romdata <= X"00000F46";
    when 16#00E9A# => romdata <= X"00000F46";
    when 16#00E9B# => romdata <= X"00000F46";
    when 16#00E9C# => romdata <= X"00000F46";
    when 16#00E9D# => romdata <= X"00000F46";
    when 16#00E9E# => romdata <= X"00000F46";
    when 16#00E9F# => romdata <= X"00000F46";
    when 16#00EA0# => romdata <= X"00000F67";
    when 16#00EA1# => romdata <= X"00000F46";
    when 16#00EA2# => romdata <= X"00000F46";
    when 16#00EA3# => romdata <= X"00000F46";
    when 16#00EA4# => romdata <= X"00000F46";
    when 16#00EA5# => romdata <= X"00000F46";
    when 16#00EA6# => romdata <= X"00000F46";
    when 16#00EA7# => romdata <= X"00000F46";
    when 16#00EA8# => romdata <= X"00000F46";
    when 16#00EA9# => romdata <= X"00000F46";
    when 16#00EAA# => romdata <= X"00000F46";
    when 16#00EAB# => romdata <= X"00000F46";
    when 16#00EAC# => romdata <= X"00000F46";
    when 16#00EAD# => romdata <= X"00000F46";
    when 16#00EAE# => romdata <= X"00000F46";
    when 16#00EAF# => romdata <= X"00000F46";
    when 16#00EB0# => romdata <= X"00000F46";
    when 16#00EB1# => romdata <= X"00000F46";
    when 16#00EB2# => romdata <= X"00000F46";
    when 16#00EB3# => romdata <= X"00000F46";
    when 16#00EB4# => romdata <= X"00000F46";
    when 16#00EB5# => romdata <= X"00000F46";
    when 16#00EB6# => romdata <= X"00000F46";
    when 16#00EB7# => romdata <= X"00000F46";
    when 16#00EB8# => romdata <= X"00000F46";
    when 16#00EB9# => romdata <= X"00000F46";
    when 16#00EBA# => romdata <= X"00000F46";
    when 16#00EBB# => romdata <= X"00000F46";
    when 16#00EBC# => romdata <= X"00000F5C";
    when 16#00EBD# => romdata <= X"69326320";
    when 16#00EBE# => romdata <= X"464D430A";
    when 16#00EBF# => romdata <= X"00000000";
    when 16#00EC0# => romdata <= X"61646472";
    when 16#00EC1# => romdata <= X"6573733A";
    when 16#00EC2# => romdata <= X"20307800";
    when 16#00EC3# => romdata <= X"2020202D";
    when 16#00EC4# => romdata <= X"2D3E2020";
    when 16#00EC5# => romdata <= X"2041434B";
    when 16#00EC6# => romdata <= X"0A000000";
    when 16#00EC7# => romdata <= X"72656164";
    when 16#00EC8# => romdata <= X"20646174";
    when 16#00EC9# => romdata <= X"61202800";
    when 16#00ECA# => romdata <= X"20627974";
    when 16#00ECB# => romdata <= X"65732920";
    when 16#00ECC# => romdata <= X"66726F6D";
    when 16#00ECD# => romdata <= X"20493243";
    when 16#00ECE# => romdata <= X"2D616464";
    when 16#00ECF# => romdata <= X"72657373";
    when 16#00ED0# => romdata <= X"20307800";
    when 16#00ED1# => romdata <= X"0A307800";
    when 16#00ED2# => romdata <= X"02020606";
    when 16#00ED3# => romdata <= X"06040304";
    when 16#00ED4# => romdata <= X"02020102";
    when 16#00ED5# => romdata <= X"636F6E74";
    when 16#00ED6# => romdata <= X"726F6C20";
    when 16#00ED7# => romdata <= X"2020203A";
    when 16#00ED8# => romdata <= X"20000000";
    when 16#00ED9# => romdata <= X"66726571";
    when 16#00EDA# => romdata <= X"75656E63";
    when 16#00EDB# => romdata <= X"7920203A";
    when 16#00EDC# => romdata <= X"20000000";
    when 16#00EDD# => romdata <= X"75706461";
    when 16#00EDE# => romdata <= X"74652063";
    when 16#00EDF# => romdata <= X"6C6B203A";
    when 16#00EE0# => romdata <= X"20000000";
    when 16#00EE1# => romdata <= X"72616D70";
    when 16#00EE2# => romdata <= X"20726174";
    when 16#00EE3# => romdata <= X"6520203A";
    when 16#00EE4# => romdata <= X"20000000";
    when 16#00EE5# => romdata <= X"49206D75";
    when 16#00EE6# => romdata <= X"6C742072";
    when 16#00EE7# => romdata <= X"6567203A";
    when 16#00EE8# => romdata <= X"20000000";
    when 16#00EE9# => romdata <= X"51206D75";
    when 16#00EEA# => romdata <= X"6C742072";
    when 16#00EEB# => romdata <= X"6567203A";
    when 16#00EEC# => romdata <= X"20000000";
    when 16#00EED# => romdata <= X"554E4B4E";
    when 16#00EEE# => romdata <= X"4F574E00";
    when 16#00EEF# => romdata <= X"69646C65";
    when 16#00EF0# => romdata <= X"00000000";
    when 16#00EF1# => romdata <= X"636F6E66";
    when 16#00EF2# => romdata <= X"69677572";
    when 16#00EF3# => romdata <= X"65000000";
    when 16#00EF4# => romdata <= X"64657465";
    when 16#00EF5# => romdata <= X"63740000";
    when 16#00EF6# => romdata <= X"61717569";
    when 16#00EF7# => romdata <= X"72650000";
    when 16#00EF8# => romdata <= X"616E616C";
    when 16#00EF9# => romdata <= X"797A6500";
    when 16#00EFA# => romdata <= X"64657369";
    when 16#00EFB# => romdata <= X"72650000";
    when 16#00EFC# => romdata <= X"72656164";
    when 16#00EFD# => romdata <= X"6F757400";
    when 16#00EFE# => romdata <= X"72656164";
    when 16#00EFF# => romdata <= X"6C616700";
    when 16#00F00# => romdata <= X"66617374";
    when 16#00F01# => romdata <= X"20747269";
    when 16#00F02# => romdata <= X"67676572";
    when 16#00F03# => romdata <= X"203A2000";
    when 16#00F04# => romdata <= X"0A736C6F";
    when 16#00F05# => romdata <= X"77207472";
    when 16#00F06# => romdata <= X"69676765";
    when 16#00F07# => romdata <= X"72203A20";
    when 16#00F08# => romdata <= X"00000000";
    when 16#00F09# => romdata <= X"0A6F7665";
    when 16#00F0A# => romdata <= X"72666C6F";
    when 16#00F0B# => romdata <= X"77202020";
    when 16#00F0C# => romdata <= X"20203A20";
    when 16#00F0D# => romdata <= X"00000000";
    when 16#00F0E# => romdata <= X"66617374";
    when 16#00F0F# => romdata <= X"20747269";
    when 16#00F10# => romdata <= X"67676572";
    when 16#00F11# => romdata <= X"20636861";
    when 16#00F12# => romdata <= X"696E3A20";
    when 16#00F13# => romdata <= X"30780000";
    when 16#00F14# => romdata <= X"0A736C6F";
    when 16#00F15# => romdata <= X"77207472";
    when 16#00F16# => romdata <= X"69676765";
    when 16#00F17# => romdata <= X"72206368";
    when 16#00F18# => romdata <= X"61696E3A";
    when 16#00F19# => romdata <= X"20307800";
    when 16#00F1A# => romdata <= X"746F6B65";
    when 16#00F1B# => romdata <= X"6E733A20";
    when 16#00F1C# => romdata <= X"00000000";
    when 16#00F1D# => romdata <= X"00001A77";
    when 16#00F1E# => romdata <= X"00001A8B";
    when 16#00F1F# => romdata <= X"00001A4F";
    when 16#00F20# => romdata <= X"00001A9F";
    when 16#00F21# => romdata <= X"00001AB3";
    when 16#00F22# => romdata <= X"00001AC7";
    when 16#00F23# => romdata <= X"00001ADB";
    when 16#00F24# => romdata <= X"00001AEF";
    when 16#00F25# => romdata <= X"00001B03";
    when 16#00F26# => romdata <= X"00001A63";
    when 16#00F27# => romdata <= X"30622020";
    when 16#00F28# => romdata <= X"20202020";
    when 16#00F29# => romdata <= X"20202020";
    when 16#00F2A# => romdata <= X"20202020";
    when 16#00F2B# => romdata <= X"20202020";
    when 16#00F2C# => romdata <= X"20202020";
    when 16#00F2D# => romdata <= X"20202020";
    when 16#00F2E# => romdata <= X"20202020";
    when 16#00F2F# => romdata <= X"20200000";
    when 16#00F30# => romdata <= X"20202020";
    when 16#00F31# => romdata <= X"20202020";
    when 16#00F32# => romdata <= X"00000000";
    when 16#00F33# => romdata <= X"79657300";
    when 16#00F34# => romdata <= X"6E6F0000";
    when 16#00F35# => romdata <= X"00202020";
    when 16#00F36# => romdata <= X"20202020";
    when 16#00F37# => romdata <= X"20202828";
    when 16#00F38# => romdata <= X"28282820";
    when 16#00F39# => romdata <= X"20202020";
    when 16#00F3A# => romdata <= X"20202020";
    when 16#00F3B# => romdata <= X"20202020";
    when 16#00F3C# => romdata <= X"20202020";
    when 16#00F3D# => romdata <= X"20881010";
    when 16#00F3E# => romdata <= X"10101010";
    when 16#00F3F# => romdata <= X"10101010";
    when 16#00F40# => romdata <= X"10101010";
    when 16#00F41# => romdata <= X"10040404";
    when 16#00F42# => romdata <= X"04040404";
    when 16#00F43# => romdata <= X"04040410";
    when 16#00F44# => romdata <= X"10101010";
    when 16#00F45# => romdata <= X"10104141";
    when 16#00F46# => romdata <= X"41414141";
    when 16#00F47# => romdata <= X"01010101";
    when 16#00F48# => romdata <= X"01010101";
    when 16#00F49# => romdata <= X"01010101";
    when 16#00F4A# => romdata <= X"01010101";
    when 16#00F4B# => romdata <= X"01010101";
    when 16#00F4C# => romdata <= X"10101010";
    when 16#00F4D# => romdata <= X"10104242";
    when 16#00F4E# => romdata <= X"42424242";
    when 16#00F4F# => romdata <= X"02020202";
    when 16#00F50# => romdata <= X"02020202";
    when 16#00F51# => romdata <= X"02020202";
    when 16#00F52# => romdata <= X"02020202";
    when 16#00F53# => romdata <= X"02020202";
    when 16#00F54# => romdata <= X"10101010";
    when 16#00F55# => romdata <= X"20000000";
    when 16#00F56# => romdata <= X"00000000";
    when 16#00F57# => romdata <= X"00000000";
    when 16#00F58# => romdata <= X"00000000";
    when 16#00F59# => romdata <= X"00000000";
    when 16#00F5A# => romdata <= X"00000000";
    when 16#00F5B# => romdata <= X"00000000";
    when 16#00F5C# => romdata <= X"00000000";
    when 16#00F5D# => romdata <= X"00000000";
    when 16#00F5E# => romdata <= X"00000000";
    when 16#00F5F# => romdata <= X"00000000";
    when 16#00F60# => romdata <= X"00000000";
    when 16#00F61# => romdata <= X"00000000";
    when 16#00F62# => romdata <= X"00000000";
    when 16#00F63# => romdata <= X"00000000";
    when 16#00F64# => romdata <= X"00000000";
    when 16#00F65# => romdata <= X"00000000";
    when 16#00F66# => romdata <= X"00000000";
    when 16#00F67# => romdata <= X"00000000";
    when 16#00F68# => romdata <= X"00000000";
    when 16#00F69# => romdata <= X"00000000";
    when 16#00F6A# => romdata <= X"00000000";
    when 16#00F6B# => romdata <= X"00000000";
    when 16#00F6C# => romdata <= X"00000000";
    when 16#00F6D# => romdata <= X"00000000";
    when 16#00F6E# => romdata <= X"00000000";
    when 16#00F6F# => romdata <= X"00000000";
    when 16#00F70# => romdata <= X"00000000";
    when 16#00F71# => romdata <= X"00000000";
    when 16#00F72# => romdata <= X"00000000";
    when 16#00F73# => romdata <= X"00000000";
    when 16#00F74# => romdata <= X"00000000";
    when 16#00F75# => romdata <= X"00000000";
    when 16#00F76# => romdata <= X"43000000";
    when 16#00F77# => romdata <= X"00000000";
    when 16#00F78# => romdata <= X"00000000";
    when 16#00F79# => romdata <= X"80000B00";
    when 16#00F7A# => romdata <= X"10000000";
    when 16#00F7B# => romdata <= X"80000D00";
    when 16#00F7C# => romdata <= X"00FFFFFF";
    when 16#00F7D# => romdata <= X"FF00FFFF";
    when 16#00F7E# => romdata <= X"FFFF00FF";
    when 16#00F7F# => romdata <= X"FFFFFF00";
    when 16#00F80# => romdata <= X"00000000";
    when 16#00F81# => romdata <= X"00000000";
    when 16#00F82# => romdata <= X"80000A00";
    when 16#00F83# => romdata <= X"80000400";
    when 16#00F84# => romdata <= X"80000200";
    when 16#00F85# => romdata <= X"80000100";
    when 16#00F86# => romdata <= X"80000004";
    when 16#00F87# => romdata <= X"80000000";
    when 16#00F88# => romdata <= X"00003E24";
    when 16#00F89# => romdata <= X"00000000";
    when 16#00F8A# => romdata <= X"0000408C";
    when 16#00F8B# => romdata <= X"000040E8";
    when 16#00F8C# => romdata <= X"00004144";
    when 16#00F8D# => romdata <= X"00000000";
    when 16#00F8E# => romdata <= X"00000000";
    when 16#00F8F# => romdata <= X"00000000";
    when 16#00F90# => romdata <= X"00000000";
    when 16#00F91# => romdata <= X"00000000";
    when 16#00F92# => romdata <= X"00000000";
    when 16#00F93# => romdata <= X"00000000";
    when 16#00F94# => romdata <= X"00000000";
    when 16#00F95# => romdata <= X"00000000";
    when 16#00F96# => romdata <= X"00003DD8";
    when 16#00F97# => romdata <= X"00000000";
    when 16#00F98# => romdata <= X"00000000";
    when 16#00F99# => romdata <= X"00000000";
    when 16#00F9A# => romdata <= X"00000000";
    when 16#00F9B# => romdata <= X"00000000";
    when 16#00F9C# => romdata <= X"00000000";
    when 16#00F9D# => romdata <= X"00000000";
    when 16#00F9E# => romdata <= X"00000000";
    when 16#00F9F# => romdata <= X"00000000";
    when 16#00FA0# => romdata <= X"00000000";
    when 16#00FA1# => romdata <= X"00000000";
    when 16#00FA2# => romdata <= X"00000000";
    when 16#00FA3# => romdata <= X"00000000";
    when 16#00FA4# => romdata <= X"00000000";
    when 16#00FA5# => romdata <= X"00000000";
    when 16#00FA6# => romdata <= X"00000000";
    when 16#00FA7# => romdata <= X"00000000";
    when 16#00FA8# => romdata <= X"00000000";
    when 16#00FA9# => romdata <= X"00000000";
    when 16#00FAA# => romdata <= X"00000000";
    when 16#00FAB# => romdata <= X"00000000";
    when 16#00FAC# => romdata <= X"00000000";
    when 16#00FAD# => romdata <= X"00000000";
    when 16#00FAE# => romdata <= X"00000000";
    when 16#00FAF# => romdata <= X"00000000";
    when 16#00FB0# => romdata <= X"00000000";
    when 16#00FB1# => romdata <= X"00000000";
    when 16#00FB2# => romdata <= X"00000000";
    when 16#00FB3# => romdata <= X"00000001";
    when 16#00FB4# => romdata <= X"330EABCD";
    when 16#00FB5# => romdata <= X"1234E66D";
    when 16#00FB6# => romdata <= X"DEEC0005";
    when 16#00FB7# => romdata <= X"000B0000";
    when 16#00FB8# => romdata <= X"00000000";
    when 16#00FB9# => romdata <= X"00000000";
    when 16#00FBA# => romdata <= X"00000000";
    when 16#00FBB# => romdata <= X"00000000";
    when 16#00FBC# => romdata <= X"00000000";
    when 16#00FBD# => romdata <= X"00000000";
    when 16#00FBE# => romdata <= X"00000000";
    when 16#00FBF# => romdata <= X"00000000";
    when 16#00FC0# => romdata <= X"00000000";
    when 16#00FC1# => romdata <= X"00000000";
    when 16#00FC2# => romdata <= X"00000000";
    when 16#00FC3# => romdata <= X"00000000";
    when 16#00FC4# => romdata <= X"00000000";
    when 16#00FC5# => romdata <= X"00000000";
    when 16#00FC6# => romdata <= X"00000000";
    when 16#00FC7# => romdata <= X"00000000";
    when 16#00FC8# => romdata <= X"00000000";
    when 16#00FC9# => romdata <= X"00000000";
    when 16#00FCA# => romdata <= X"00000000";
    when 16#00FCB# => romdata <= X"00000000";
    when 16#00FCC# => romdata <= X"00000000";
    when 16#00FCD# => romdata <= X"00000000";
    when 16#00FCE# => romdata <= X"00000000";
    when 16#00FCF# => romdata <= X"00000000";
    when 16#00FD0# => romdata <= X"00000000";
    when 16#00FD1# => romdata <= X"00000000";
    when 16#00FD2# => romdata <= X"00000000";
    when 16#00FD3# => romdata <= X"00000000";
    when 16#00FD4# => romdata <= X"00000000";
    when 16#00FD5# => romdata <= X"00000000";
    when 16#00FD6# => romdata <= X"00000000";
    when 16#00FD7# => romdata <= X"00000000";
    when 16#00FD8# => romdata <= X"00000000";
    when 16#00FD9# => romdata <= X"00000000";
    when 16#00FDA# => romdata <= X"00000000";
    when 16#00FDB# => romdata <= X"00000000";
    when 16#00FDC# => romdata <= X"00000000";
    when 16#00FDD# => romdata <= X"00000000";
    when 16#00FDE# => romdata <= X"00000000";
    when 16#00FDF# => romdata <= X"00000000";
    when 16#00FE0# => romdata <= X"00000000";
    when 16#00FE1# => romdata <= X"00000000";
    when 16#00FE2# => romdata <= X"00000000";
    when 16#00FE3# => romdata <= X"00000000";
    when 16#00FE4# => romdata <= X"00000000";
    when 16#00FE5# => romdata <= X"00000000";
    when 16#00FE6# => romdata <= X"00000000";
    when 16#00FE7# => romdata <= X"00000000";
    when 16#00FE8# => romdata <= X"00000000";
    when 16#00FE9# => romdata <= X"00000000";
    when 16#00FEA# => romdata <= X"00000000";
    when 16#00FEB# => romdata <= X"00000000";
    when 16#00FEC# => romdata <= X"00000000";
    when 16#00FED# => romdata <= X"00000000";
    when 16#00FEE# => romdata <= X"00000000";
    when 16#00FEF# => romdata <= X"00000000";
    when 16#00FF0# => romdata <= X"00000000";
    when 16#00FF1# => romdata <= X"00000000";
    when 16#00FF2# => romdata <= X"00000000";
    when 16#00FF3# => romdata <= X"00000000";
    when 16#00FF4# => romdata <= X"00000000";
    when 16#00FF5# => romdata <= X"00000000";
    when 16#00FF6# => romdata <= X"00000000";
    when 16#00FF7# => romdata <= X"00000000";
    when 16#00FF8# => romdata <= X"00000000";
    when 16#00FF9# => romdata <= X"00000000";
    when 16#00FFA# => romdata <= X"00000000";
    when 16#00FFB# => romdata <= X"00000000";
    when 16#00FFC# => romdata <= X"00000000";
    when 16#00FFD# => romdata <= X"00000000";
    when 16#00FFE# => romdata <= X"00000000";
    when 16#00FFF# => romdata <= X"00000000";
    when 16#01000# => romdata <= X"00000000";
    when 16#01001# => romdata <= X"00000000";
    when 16#01002# => romdata <= X"00000000";
    when 16#01003# => romdata <= X"00000000";
    when 16#01004# => romdata <= X"00000000";
    when 16#01005# => romdata <= X"00000000";
    when 16#01006# => romdata <= X"00000000";
    when 16#01007# => romdata <= X"00000000";
    when 16#01008# => romdata <= X"00000000";
    when 16#01009# => romdata <= X"00000000";
    when 16#0100A# => romdata <= X"00000000";
    when 16#0100B# => romdata <= X"00000000";
    when 16#0100C# => romdata <= X"00000000";
    when 16#0100D# => romdata <= X"00000000";
    when 16#0100E# => romdata <= X"00000000";
    when 16#0100F# => romdata <= X"00000000";
    when 16#01010# => romdata <= X"00000000";
    when 16#01011# => romdata <= X"00000000";
    when 16#01012# => romdata <= X"00000000";
    when 16#01013# => romdata <= X"00000000";
    when 16#01014# => romdata <= X"00000000";
    when 16#01015# => romdata <= X"00000000";
    when 16#01016# => romdata <= X"00000000";
    when 16#01017# => romdata <= X"00000000";
    when 16#01018# => romdata <= X"00000000";
    when 16#01019# => romdata <= X"00000000";
    when 16#0101A# => romdata <= X"00000000";
    when 16#0101B# => romdata <= X"00000000";
    when 16#0101C# => romdata <= X"00000000";
    when 16#0101D# => romdata <= X"00000000";
    when 16#0101E# => romdata <= X"00000000";
    when 16#0101F# => romdata <= X"00000000";
    when 16#01020# => romdata <= X"00000000";
    when 16#01021# => romdata <= X"00000000";
    when 16#01022# => romdata <= X"00000000";
    when 16#01023# => romdata <= X"00000000";
    when 16#01024# => romdata <= X"00000000";
    when 16#01025# => romdata <= X"00000000";
    when 16#01026# => romdata <= X"00000000";
    when 16#01027# => romdata <= X"00000000";
    when 16#01028# => romdata <= X"00000000";
    when 16#01029# => romdata <= X"00000000";
    when 16#0102A# => romdata <= X"00000000";
    when 16#0102B# => romdata <= X"00000000";
    when 16#0102C# => romdata <= X"00000000";
    when 16#0102D# => romdata <= X"00000000";
    when 16#0102E# => romdata <= X"00000000";
    when 16#0102F# => romdata <= X"00000000";
    when 16#01030# => romdata <= X"00000000";
    when 16#01031# => romdata <= X"00000000";
    when 16#01032# => romdata <= X"00000000";
    when 16#01033# => romdata <= X"00000000";
    when 16#01034# => romdata <= X"00000000";
    when 16#01035# => romdata <= X"00000000";
    when 16#01036# => romdata <= X"00000000";
    when 16#01037# => romdata <= X"00000000";
    when 16#01038# => romdata <= X"00000000";
    when 16#01039# => romdata <= X"00000000";
    when 16#0103A# => romdata <= X"00000000";
    when 16#0103B# => romdata <= X"00000000";
    when 16#0103C# => romdata <= X"00000000";
    when 16#0103D# => romdata <= X"00000000";
    when 16#0103E# => romdata <= X"00000000";
    when 16#0103F# => romdata <= X"00000000";
    when 16#01040# => romdata <= X"00000000";
    when 16#01041# => romdata <= X"00000000";
    when 16#01042# => romdata <= X"00000000";
    when 16#01043# => romdata <= X"00000000";
    when 16#01044# => romdata <= X"00000000";
    when 16#01045# => romdata <= X"00000000";
    when 16#01046# => romdata <= X"00000000";
    when 16#01047# => romdata <= X"00000000";
    when 16#01048# => romdata <= X"00000000";
    when 16#01049# => romdata <= X"00000000";
    when 16#0104A# => romdata <= X"00000000";
    when 16#0104B# => romdata <= X"00000000";
    when 16#0104C# => romdata <= X"00000000";
    when 16#0104D# => romdata <= X"00000000";
    when 16#0104E# => romdata <= X"00000000";
    when 16#0104F# => romdata <= X"00000000";
    when 16#01050# => romdata <= X"00000000";
    when 16#01051# => romdata <= X"00000000";
    when 16#01052# => romdata <= X"00000000";
    when 16#01053# => romdata <= X"00000000";
    when 16#01054# => romdata <= X"00000000";
    when 16#01055# => romdata <= X"00000000";
    when 16#01056# => romdata <= X"00000000";
    when 16#01057# => romdata <= X"00000000";
    when 16#01058# => romdata <= X"00000000";
    when 16#01059# => romdata <= X"00000000";
    when 16#0105A# => romdata <= X"00000000";
    when 16#0105B# => romdata <= X"00000000";
    when 16#0105C# => romdata <= X"00000000";
    when 16#0105D# => romdata <= X"00000000";
    when 16#0105E# => romdata <= X"00000000";
    when 16#0105F# => romdata <= X"00000000";
    when 16#01060# => romdata <= X"00000000";
    when 16#01061# => romdata <= X"00000000";
    when 16#01062# => romdata <= X"00000000";
    when 16#01063# => romdata <= X"00000000";
    when 16#01064# => romdata <= X"00000000";
    when 16#01065# => romdata <= X"00000000";
    when 16#01066# => romdata <= X"00000000";
    when 16#01067# => romdata <= X"00000000";
    when 16#01068# => romdata <= X"00000000";
    when 16#01069# => romdata <= X"00000000";
    when 16#0106A# => romdata <= X"00000000";
    when 16#0106B# => romdata <= X"00000000";
    when 16#0106C# => romdata <= X"00000000";
    when 16#0106D# => romdata <= X"00000000";
    when 16#0106E# => romdata <= X"00000000";
    when 16#0106F# => romdata <= X"00000000";
    when 16#01070# => romdata <= X"00000000";
    when 16#01071# => romdata <= X"00000000";
    when 16#01072# => romdata <= X"00000000";
    when 16#01073# => romdata <= X"00000000";
    when 16#01074# => romdata <= X"FFFFFFFF";
    when 16#01075# => romdata <= X"00000000";
    when 16#01076# => romdata <= X"00020000";
    when 16#01077# => romdata <= X"00000000";
    when 16#01078# => romdata <= X"00000000";
    when 16#01079# => romdata <= X"000041DC";
    when 16#0107A# => romdata <= X"000041DC";
    when 16#0107B# => romdata <= X"000041E4";
    when 16#0107C# => romdata <= X"000041E4";
    when 16#0107D# => romdata <= X"000041EC";
    when 16#0107E# => romdata <= X"000041EC";
    when 16#0107F# => romdata <= X"000041F4";
    when 16#01080# => romdata <= X"000041F4";
    when 16#01081# => romdata <= X"000041FC";
    when 16#01082# => romdata <= X"000041FC";
    when 16#01083# => romdata <= X"00004204";
    when 16#01084# => romdata <= X"00004204";
    when 16#01085# => romdata <= X"0000420C";
    when 16#01086# => romdata <= X"0000420C";
    when 16#01087# => romdata <= X"00004214";
    when 16#01088# => romdata <= X"00004214";
    when 16#01089# => romdata <= X"0000421C";
    when 16#0108A# => romdata <= X"0000421C";
    when 16#0108B# => romdata <= X"00004224";
    when 16#0108C# => romdata <= X"00004224";
    when 16#0108D# => romdata <= X"0000422C";
    when 16#0108E# => romdata <= X"0000422C";
    when 16#0108F# => romdata <= X"00004234";
    when 16#01090# => romdata <= X"00004234";
    when 16#01091# => romdata <= X"0000423C";
    when 16#01092# => romdata <= X"0000423C";
    when 16#01093# => romdata <= X"00004244";
    when 16#01094# => romdata <= X"00004244";
    when 16#01095# => romdata <= X"0000424C";
    when 16#01096# => romdata <= X"0000424C";
    when 16#01097# => romdata <= X"00004254";
    when 16#01098# => romdata <= X"00004254";
    when 16#01099# => romdata <= X"0000425C";
    when 16#0109A# => romdata <= X"0000425C";
    when 16#0109B# => romdata <= X"00004264";
    when 16#0109C# => romdata <= X"00004264";
    when 16#0109D# => romdata <= X"0000426C";
    when 16#0109E# => romdata <= X"0000426C";
    when 16#0109F# => romdata <= X"00004274";
    when 16#010A0# => romdata <= X"00004274";
    when 16#010A1# => romdata <= X"0000427C";
    when 16#010A2# => romdata <= X"0000427C";
    when 16#010A3# => romdata <= X"00004284";
    when 16#010A4# => romdata <= X"00004284";
    when 16#010A5# => romdata <= X"0000428C";
    when 16#010A6# => romdata <= X"0000428C";
    when 16#010A7# => romdata <= X"00004294";
    when 16#010A8# => romdata <= X"00004294";
    when 16#010A9# => romdata <= X"0000429C";
    when 16#010AA# => romdata <= X"0000429C";
    when 16#010AB# => romdata <= X"000042A4";
    when 16#010AC# => romdata <= X"000042A4";
    when 16#010AD# => romdata <= X"000042AC";
    when 16#010AE# => romdata <= X"000042AC";
    when 16#010AF# => romdata <= X"000042B4";
    when 16#010B0# => romdata <= X"000042B4";
    when 16#010B1# => romdata <= X"000042BC";
    when 16#010B2# => romdata <= X"000042BC";
    when 16#010B3# => romdata <= X"000042C4";
    when 16#010B4# => romdata <= X"000042C4";
    when 16#010B5# => romdata <= X"000042CC";
    when 16#010B6# => romdata <= X"000042CC";
    when 16#010B7# => romdata <= X"000042D4";
    when 16#010B8# => romdata <= X"000042D4";
    when 16#010B9# => romdata <= X"000042DC";
    when 16#010BA# => romdata <= X"000042DC";
    when 16#010BB# => romdata <= X"000042E4";
    when 16#010BC# => romdata <= X"000042E4";
    when 16#010BD# => romdata <= X"000042EC";
    when 16#010BE# => romdata <= X"000042EC";
    when 16#010BF# => romdata <= X"000042F4";
    when 16#010C0# => romdata <= X"000042F4";
    when 16#010C1# => romdata <= X"000042FC";
    when 16#010C2# => romdata <= X"000042FC";
    when 16#010C3# => romdata <= X"00004304";
    when 16#010C4# => romdata <= X"00004304";
    when 16#010C5# => romdata <= X"0000430C";
    when 16#010C6# => romdata <= X"0000430C";
    when 16#010C7# => romdata <= X"00004314";
    when 16#010C8# => romdata <= X"00004314";
    when 16#010C9# => romdata <= X"0000431C";
    when 16#010CA# => romdata <= X"0000431C";
    when 16#010CB# => romdata <= X"00004324";
    when 16#010CC# => romdata <= X"00004324";
    when 16#010CD# => romdata <= X"0000432C";
    when 16#010CE# => romdata <= X"0000432C";
    when 16#010CF# => romdata <= X"00004334";
    when 16#010D0# => romdata <= X"00004334";
    when 16#010D1# => romdata <= X"0000433C";
    when 16#010D2# => romdata <= X"0000433C";
    when 16#010D3# => romdata <= X"00004344";
    when 16#010D4# => romdata <= X"00004344";
    when 16#010D5# => romdata <= X"0000434C";
    when 16#010D6# => romdata <= X"0000434C";
    when 16#010D7# => romdata <= X"00004354";
    when 16#010D8# => romdata <= X"00004354";
    when 16#010D9# => romdata <= X"0000435C";
    when 16#010DA# => romdata <= X"0000435C";
    when 16#010DB# => romdata <= X"00004364";
    when 16#010DC# => romdata <= X"00004364";
    when 16#010DD# => romdata <= X"0000436C";
    when 16#010DE# => romdata <= X"0000436C";
    when 16#010DF# => romdata <= X"00004374";
    when 16#010E0# => romdata <= X"00004374";
    when 16#010E1# => romdata <= X"0000437C";
    when 16#010E2# => romdata <= X"0000437C";
    when 16#010E3# => romdata <= X"00004384";
    when 16#010E4# => romdata <= X"00004384";
    when 16#010E5# => romdata <= X"0000438C";
    when 16#010E6# => romdata <= X"0000438C";
    when 16#010E7# => romdata <= X"00004394";
    when 16#010E8# => romdata <= X"00004394";
    when 16#010E9# => romdata <= X"0000439C";
    when 16#010EA# => romdata <= X"0000439C";
    when 16#010EB# => romdata <= X"000043A4";
    when 16#010EC# => romdata <= X"000043A4";
    when 16#010ED# => romdata <= X"000043AC";
    when 16#010EE# => romdata <= X"000043AC";
    when 16#010EF# => romdata <= X"000043B4";
    when 16#010F0# => romdata <= X"000043B4";
    when 16#010F1# => romdata <= X"000043BC";
    when 16#010F2# => romdata <= X"000043BC";
    when 16#010F3# => romdata <= X"000043C4";
    when 16#010F4# => romdata <= X"000043C4";
    when 16#010F5# => romdata <= X"000043CC";
    when 16#010F6# => romdata <= X"000043CC";
    when 16#010F7# => romdata <= X"000043D4";
    when 16#010F8# => romdata <= X"000043D4";
    when 16#010F9# => romdata <= X"000043DC";
    when 16#010FA# => romdata <= X"000043DC";
    when 16#010FB# => romdata <= X"000043E4";
    when 16#010FC# => romdata <= X"000043E4";
    when 16#010FD# => romdata <= X"000043EC";
    when 16#010FE# => romdata <= X"000043EC";
    when 16#010FF# => romdata <= X"000043F4";
    when 16#01100# => romdata <= X"000043F4";
    when 16#01101# => romdata <= X"000043FC";
    when 16#01102# => romdata <= X"000043FC";
    when 16#01103# => romdata <= X"00004404";
    when 16#01104# => romdata <= X"00004404";
    when 16#01105# => romdata <= X"0000440C";
    when 16#01106# => romdata <= X"0000440C";
    when 16#01107# => romdata <= X"00004414";
    when 16#01108# => romdata <= X"00004414";
    when 16#01109# => romdata <= X"0000441C";
    when 16#0110A# => romdata <= X"0000441C";
    when 16#0110B# => romdata <= X"00004424";
    when 16#0110C# => romdata <= X"00004424";
    when 16#0110D# => romdata <= X"0000442C";
    when 16#0110E# => romdata <= X"0000442C";
    when 16#0110F# => romdata <= X"00004434";
    when 16#01110# => romdata <= X"00004434";
    when 16#01111# => romdata <= X"0000443C";
    when 16#01112# => romdata <= X"0000443C";
    when 16#01113# => romdata <= X"00004444";
    when 16#01114# => romdata <= X"00004444";
    when 16#01115# => romdata <= X"0000444C";
    when 16#01116# => romdata <= X"0000444C";
    when 16#01117# => romdata <= X"00004454";
    when 16#01118# => romdata <= X"00004454";
    when 16#01119# => romdata <= X"0000445C";
    when 16#0111A# => romdata <= X"0000445C";
    when 16#0111B# => romdata <= X"00004464";
    when 16#0111C# => romdata <= X"00004464";
    when 16#0111D# => romdata <= X"0000446C";
    when 16#0111E# => romdata <= X"0000446C";
    when 16#0111F# => romdata <= X"00004474";
    when 16#01120# => romdata <= X"00004474";
    when 16#01121# => romdata <= X"0000447C";
    when 16#01122# => romdata <= X"0000447C";
    when 16#01123# => romdata <= X"00004484";
    when 16#01124# => romdata <= X"00004484";
    when 16#01125# => romdata <= X"0000448C";
    when 16#01126# => romdata <= X"0000448C";
    when 16#01127# => romdata <= X"00004494";
    when 16#01128# => romdata <= X"00004494";
    when 16#01129# => romdata <= X"0000449C";
    when 16#0112A# => romdata <= X"0000449C";
    when 16#0112B# => romdata <= X"000044A4";
    when 16#0112C# => romdata <= X"000044A4";
    when 16#0112D# => romdata <= X"000044AC";
    when 16#0112E# => romdata <= X"000044AC";
    when 16#0112F# => romdata <= X"000044B4";
    when 16#01130# => romdata <= X"000044B4";
    when 16#01131# => romdata <= X"000044BC";
    when 16#01132# => romdata <= X"000044BC";
    when 16#01133# => romdata <= X"000044C4";
    when 16#01134# => romdata <= X"000044C4";
    when 16#01135# => romdata <= X"000044CC";
    when 16#01136# => romdata <= X"000044CC";
    when 16#01137# => romdata <= X"000044D4";
    when 16#01138# => romdata <= X"000044D4";
    when 16#01139# => romdata <= X"000044DC";
    when 16#0113A# => romdata <= X"000044DC";
    when 16#0113B# => romdata <= X"000044E4";
    when 16#0113C# => romdata <= X"000044E4";
    when 16#0113D# => romdata <= X"000044EC";
    when 16#0113E# => romdata <= X"000044EC";
    when 16#0113F# => romdata <= X"000044F4";
    when 16#01140# => romdata <= X"000044F4";
    when 16#01141# => romdata <= X"000044FC";
    when 16#01142# => romdata <= X"000044FC";
    when 16#01143# => romdata <= X"00004504";
    when 16#01144# => romdata <= X"00004504";
    when 16#01145# => romdata <= X"0000450C";
    when 16#01146# => romdata <= X"0000450C";
    when 16#01147# => romdata <= X"00004514";
    when 16#01148# => romdata <= X"00004514";
    when 16#01149# => romdata <= X"0000451C";
    when 16#0114A# => romdata <= X"0000451C";
    when 16#0114B# => romdata <= X"00004524";
    when 16#0114C# => romdata <= X"00004524";
    when 16#0114D# => romdata <= X"0000452C";
    when 16#0114E# => romdata <= X"0000452C";
    when 16#0114F# => romdata <= X"00004534";
    when 16#01150# => romdata <= X"00004534";
    when 16#01151# => romdata <= X"0000453C";
    when 16#01152# => romdata <= X"0000453C";
    when 16#01153# => romdata <= X"00004544";
    when 16#01154# => romdata <= X"00004544";
    when 16#01155# => romdata <= X"0000454C";
    when 16#01156# => romdata <= X"0000454C";
    when 16#01157# => romdata <= X"00004554";
    when 16#01158# => romdata <= X"00004554";
    when 16#01159# => romdata <= X"0000455C";
    when 16#0115A# => romdata <= X"0000455C";
    when 16#0115B# => romdata <= X"00004564";
    when 16#0115C# => romdata <= X"00004564";
    when 16#0115D# => romdata <= X"0000456C";
    when 16#0115E# => romdata <= X"0000456C";
    when 16#0115F# => romdata <= X"00004574";
    when 16#01160# => romdata <= X"00004574";
    when 16#01161# => romdata <= X"0000457C";
    when 16#01162# => romdata <= X"0000457C";
    when 16#01163# => romdata <= X"00004584";
    when 16#01164# => romdata <= X"00004584";
    when 16#01165# => romdata <= X"0000458C";
    when 16#01166# => romdata <= X"0000458C";
    when 16#01167# => romdata <= X"00004594";
    when 16#01168# => romdata <= X"00004594";
    when 16#01169# => romdata <= X"0000459C";
    when 16#0116A# => romdata <= X"0000459C";
    when 16#0116B# => romdata <= X"000045A4";
    when 16#0116C# => romdata <= X"000045A4";
    when 16#0116D# => romdata <= X"000045AC";
    when 16#0116E# => romdata <= X"000045AC";
    when 16#0116F# => romdata <= X"000045B4";
    when 16#01170# => romdata <= X"000045B4";
    when 16#01171# => romdata <= X"000045BC";
    when 16#01172# => romdata <= X"000045BC";
    when 16#01173# => romdata <= X"000045C4";
    when 16#01174# => romdata <= X"000045C4";
    when 16#01175# => romdata <= X"000045CC";
    when 16#01176# => romdata <= X"000045CC";
    when 16#01177# => romdata <= X"000045D4";
    when 16#01178# => romdata <= X"000045D4";
    when 16#01179# => romdata <= X"000045D4";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
