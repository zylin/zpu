
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 16;
constant bytes : integer := 33508;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B8191";
    when 16#00001# => romdata <= X"FF040000";
    when 16#00002# => romdata <= X"00000000";
    when 16#00003# => romdata <= X"00000000";
    when 16#00004# => romdata <= X"00000000";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"0B0B8194";
    when 16#00009# => romdata <= X"E7040000";
    when 16#0000A# => romdata <= X"00000000";
    when 16#0000B# => romdata <= X"00000000";
    when 16#0000C# => romdata <= X"00000000";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B8194";
    when 16#00049# => romdata <= X"99040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B8193FC";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B81F5";
    when 16#000A2# => romdata <= X"E4738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B81";
    when 16#000A5# => romdata <= X"93FF0400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"0B0B8194";
    when 16#000A9# => romdata <= X"CE040000";
    when 16#000AA# => romdata <= X"00000000";
    when 16#000AB# => romdata <= X"00000000";
    when 16#000AC# => romdata <= X"00000000";
    when 16#000AD# => romdata <= X"00000000";
    when 16#000AE# => romdata <= X"00000000";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"0B0B8194";
    when 16#000B1# => romdata <= X"B5040000";
    when 16#000B2# => romdata <= X"00000000";
    when 16#000B3# => romdata <= X"00000000";
    when 16#000B4# => romdata <= X"00000000";
    when 16#000B5# => romdata <= X"00000000";
    when 16#000B6# => romdata <= X"00000000";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"81F5F40C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"FF3D0D02";
    when 16#00101# => romdata <= X"8F053370";
    when 16#00102# => romdata <= X"52528191";
    when 16#00103# => romdata <= X"E43F7151";
    when 16#00104# => romdata <= X"8192D23F";
    when 16#00105# => romdata <= X"71B00C83";
    when 16#00106# => romdata <= X"3D0D04FF";
    when 16#00107# => romdata <= X"3D0D028F";
    when 16#00108# => romdata <= X"05337052";
    when 16#00109# => romdata <= X"528191C9";
    when 16#0010A# => romdata <= X"3F715181";
    when 16#0010B# => romdata <= X"92B73F71";
    when 16#0010C# => romdata <= X"5180CAC3";
    when 16#0010D# => romdata <= X"3F71B00C";
    when 16#0010E# => romdata <= X"833D0D04";
    when 16#0010F# => romdata <= X"FF3D0D81";
    when 16#00110# => romdata <= X"F5CC08B8";
    when 16#00111# => romdata <= X"11085351";
    when 16#00112# => romdata <= X"800BB812";
    when 16#00113# => romdata <= X"0C71B00C";
    when 16#00114# => romdata <= X"833D0D04";
    when 16#00115# => romdata <= X"FA3D0D8A";
    when 16#00116# => romdata <= X"51818CB1";
    when 16#00117# => romdata <= X"3F96BC3F";
    when 16#00118# => romdata <= X"80E0EB53";
    when 16#00119# => romdata <= X"81C48C52";
    when 16#0011A# => romdata <= X"81C4A051";
    when 16#0011B# => romdata <= X"96C03F80";
    when 16#0011C# => romdata <= X"F4AF5381";
    when 16#0011D# => romdata <= X"C4A45281";
    when 16#0011E# => romdata <= X"C4B85196";
    when 16#0011F# => romdata <= X"B13F80F4";
    when 16#00120# => romdata <= X"855381C4";
    when 16#00121# => romdata <= X"BC5281C4";
    when 16#00122# => romdata <= X"E45196A2";
    when 16#00123# => romdata <= X"3F80FCF0";
    when 16#00124# => romdata <= X"5381C4EC";
    when 16#00125# => romdata <= X"5281C4FC";
    when 16#00126# => romdata <= X"5196933F";
    when 16#00127# => romdata <= X"80FD8753";
    when 16#00128# => romdata <= X"81C58452";
    when 16#00129# => romdata <= X"81C5A051";
    when 16#0012A# => romdata <= X"96843F80";
    when 16#0012B# => romdata <= X"F6E15381";
    when 16#0012C# => romdata <= X"C5A85281";
    when 16#0012D# => romdata <= X"C5C05195";
    when 16#0012E# => romdata <= X"F53F8180";
    when 16#0012F# => romdata <= X"E85381C5";
    when 16#00130# => romdata <= X"C85281C5";
    when 16#00131# => romdata <= X"EC5195E6";
    when 16#00132# => romdata <= X"3F90B453";
    when 16#00133# => romdata <= X"81C5F452";
    when 16#00134# => romdata <= X"81C69051";
    when 16#00135# => romdata <= X"95D83F91";
    when 16#00136# => romdata <= X"CF5381C6";
    when 16#00137# => romdata <= X"945281C6";
    when 16#00138# => romdata <= X"B85195CA";
    when 16#00139# => romdata <= X"3F8FD253";
    when 16#0013A# => romdata <= X"81C6C052";
    when 16#0013B# => romdata <= X"81C6E451";
    when 16#0013C# => romdata <= X"95BC3F81";
    when 16#0013D# => romdata <= X"8FDA5381";
    when 16#0013E# => romdata <= X"C6EC5281";
    when 16#0013F# => romdata <= X"C7945195";
    when 16#00140# => romdata <= X"AD3F8191";
    when 16#00141# => romdata <= X"875381C7";
    when 16#00142# => romdata <= X"9C5281C7";
    when 16#00143# => romdata <= X"BC51959E";
    when 16#00144# => romdata <= X"3F88BC53";
    when 16#00145# => romdata <= X"81C7C452";
    when 16#00146# => romdata <= X"81C7E451";
    when 16#00147# => romdata <= X"95903F80";
    when 16#00148# => romdata <= X"F78C5381";
    when 16#00149# => romdata <= X"C7EC5281";
    when 16#0014A# => romdata <= X"C8805195";
    when 16#0014B# => romdata <= X"813F80FD";
    when 16#0014C# => romdata <= X"A25381C8";
    when 16#0014D# => romdata <= X"885281C7";
    when 16#0014E# => romdata <= X"B45194F2";
    when 16#0014F# => romdata <= X"3F8180B4";
    when 16#00150# => romdata <= X"5381C8A4";
    when 16#00151# => romdata <= X"5281C8B8";
    when 16#00152# => romdata <= X"5194E33F";
    when 16#00153# => romdata <= X"80FEB253";
    when 16#00154# => romdata <= X"81C8C052";
    when 16#00155# => romdata <= X"81C8E051";
    when 16#00156# => romdata <= X"94D43F80";
    when 16#00157# => romdata <= X"FF945381";
    when 16#00158# => romdata <= X"C8E85281";
    when 16#00159# => romdata <= X"C9885194";
    when 16#0015A# => romdata <= X"C53F818F";
    when 16#0015B# => romdata <= X"B25381C9";
    when 16#0015C# => romdata <= X"905281C9";
    when 16#0015D# => romdata <= X"AC5194B6";
    when 16#0015E# => romdata <= X"3F818694";
    when 16#0015F# => romdata <= X"5381C9B4";
    when 16#00160# => romdata <= X"5281C9C8";
    when 16#00161# => romdata <= X"5194A73F";
    when 16#00162# => romdata <= X"81828153";
    when 16#00163# => romdata <= X"81C9D052";
    when 16#00164# => romdata <= X"81C9F451";
    when 16#00165# => romdata <= X"94983F96";
    when 16#00166# => romdata <= X"8C5381C9";
    when 16#00167# => romdata <= X"FC5281CA";
    when 16#00168# => romdata <= X"8C51948A";
    when 16#00169# => romdata <= X"3F93BC53";
    when 16#0016A# => romdata <= X"81CA9052";
    when 16#0016B# => romdata <= X"81CAAC51";
    when 16#0016C# => romdata <= X"93FC3F8F";
    when 16#0016D# => romdata <= X"B65381CA";
    when 16#0016E# => romdata <= X"B45281CA";
    when 16#0016F# => romdata <= X"CC5193EE";
    when 16#00170# => romdata <= X"3F93C453";
    when 16#00171# => romdata <= X"81CAD452";
    when 16#00172# => romdata <= X"81CAE851";
    when 16#00173# => romdata <= X"93E03F80";
    when 16#00174# => romdata <= X"D3975381";
    when 16#00175# => romdata <= X"CAF05281";
    when 16#00176# => romdata <= X"CB845193";
    when 16#00177# => romdata <= X"D13F80D7";
    when 16#00178# => romdata <= X"965381CB";
    when 16#00179# => romdata <= X"885281CB";
    when 16#0017A# => romdata <= X"B05193C2";
    when 16#0017B# => romdata <= X"3F80FABC";
    when 16#0017C# => romdata <= X"5381CBB8";
    when 16#0017D# => romdata <= X"5281CBD8";
    when 16#0017E# => romdata <= X"5193B33F";
    when 16#0017F# => romdata <= X"80F9E053";
    when 16#00180# => romdata <= X"81CBE052";
    when 16#00181# => romdata <= X"81CBF451";
    when 16#00182# => romdata <= X"93A43F80";
    when 16#00183# => romdata <= X"D9835381";
    when 16#00184# => romdata <= X"CBFC5281";
    when 16#00185# => romdata <= X"CC945193";
    when 16#00186# => romdata <= X"953FBBC5";
    when 16#00187# => romdata <= X"5381CC9C";
    when 16#00188# => romdata <= X"5281CCB4";
    when 16#00189# => romdata <= X"5193873F";
    when 16#0018A# => romdata <= X"80D9E753";
    when 16#0018B# => romdata <= X"81CCBC52";
    when 16#0018C# => romdata <= X"81CCE451";
    when 16#0018D# => romdata <= X"92F83F80";
    when 16#0018E# => romdata <= X"FAE65381";
    when 16#0018F# => romdata <= X"CCEC5281";
    when 16#00190# => romdata <= X"CCF85192";
    when 16#00191# => romdata <= X"E93F80FC";
    when 16#00192# => romdata <= X"975381CC";
    when 16#00193# => romdata <= X"FC5281CD";
    when 16#00194# => romdata <= X"A45192DA";
    when 16#00195# => romdata <= X"3F80FAE6";
    when 16#00196# => romdata <= X"5381CDAC";
    when 16#00197# => romdata <= X"5281F0D8";
    when 16#00198# => romdata <= X"5192CB3F";
    when 16#00199# => romdata <= X"80FCE053";
    when 16#0019A# => romdata <= X"81CDCC52";
    when 16#0019B# => romdata <= X"81CDDC51";
    when 16#0019C# => romdata <= X"92BC3F80";
    when 16#0019D# => romdata <= X"FADB5381";
    when 16#0019E# => romdata <= X"DEFC5281";
    when 16#0019F# => romdata <= X"C3FC5192";
    when 16#001A0# => romdata <= X"AD3FA6AD";
    when 16#001A1# => romdata <= X"5381DEFC";
    when 16#001A2# => romdata <= X"5281C484";
    when 16#001A3# => romdata <= X"51929F3F";
    when 16#001A4# => romdata <= X"999B3F92";
    when 16#001A5# => romdata <= X"F93F810B";
    when 16#001A6# => romdata <= X"829DD834";
    when 16#001A7# => romdata <= X"8285E833";
    when 16#001A8# => romdata <= X"7081FF06";
    when 16#001A9# => romdata <= X"555573B2";
    when 16#001AA# => romdata <= X"38818BED";
    when 16#001AB# => romdata <= X"3FB00890";
    when 16#001AC# => romdata <= X"3892EA3F";
    when 16#001AD# => romdata <= X"829DD833";
    when 16#001AE# => romdata <= X"5675E138";
    when 16#001AF# => romdata <= X"883D0D04";
    when 16#001B0# => romdata <= X"818BE93F";
    when 16#001B1# => romdata <= X"B00881FF";
    when 16#001B2# => romdata <= X"065193C8";
    when 16#001B3# => romdata <= X"3F92CE3F";
    when 16#001B4# => romdata <= X"829DD833";
    when 16#001B5# => romdata <= X"5675C538";
    when 16#001B6# => romdata <= X"E339800B";
    when 16#001B7# => romdata <= X"8285E834";
    when 16#001B8# => romdata <= X"99F43F81";
    when 16#001B9# => romdata <= X"F68C0870";
    when 16#001BA# => romdata <= X"0870872A";
    when 16#001BB# => romdata <= X"81065257";
    when 16#001BC# => romdata <= X"5473802E";
    when 16#001BD# => romdata <= X"8F387680";
    when 16#001BE# => romdata <= X"2E819738";
    when 16#001BF# => romdata <= X"FF177081";
    when 16#001C0# => romdata <= X"FF065854";
    when 16#001C1# => romdata <= X"75862A81";
    when 16#001C2# => romdata <= X"06557480";
    when 16#001C3# => romdata <= X"2E8F3876";
    when 16#001C4# => romdata <= X"802E8190";
    when 16#001C5# => romdata <= X"38FF1770";
    when 16#001C6# => romdata <= X"81FF0658";
    when 16#001C7# => romdata <= X"5575852A";
    when 16#001C8# => romdata <= X"81065473";
    when 16#001C9# => romdata <= X"802E9638";
    when 16#001CA# => romdata <= X"76BA3881";
    when 16#001CB# => romdata <= X"960B81F5";
    when 16#001CC# => romdata <= X"CC08B811";
    when 16#001CD# => romdata <= X"08575557";
    when 16#001CE# => romdata <= X"800BB815";
    when 16#001CF# => romdata <= X"0C75842A";
    when 16#001D0# => romdata <= X"81065675";
    when 16#001D1# => romdata <= X"802EFEE1";
    when 16#001D2# => romdata <= X"3876802E";
    when 16#001D3# => romdata <= X"A138FF17";
    when 16#001D4# => romdata <= X"7081FF06";
    when 16#001D5# => romdata <= X"5855818A";
    when 16#001D6# => romdata <= X"C03FB008";
    when 16#001D7# => romdata <= X"802EFED1";
    when 16#001D8# => romdata <= X"38FEDD39";
    when 16#001D9# => romdata <= X"FF177081";
    when 16#001DA# => romdata <= X"FF065855";
    when 16#001DB# => romdata <= X"D0398196";
    when 16#001DC# => romdata <= X"0B81F68C";
    when 16#001DD# => romdata <= X"08841108";
    when 16#001DE# => romdata <= X"840A0784";
    when 16#001DF# => romdata <= X"120C5657";
    when 16#001E0# => romdata <= X"80E4DA3F";
    when 16#001E1# => romdata <= X"818A923F";
    when 16#001E2# => romdata <= X"B008802E";
    when 16#001E3# => romdata <= X"FEA338FE";
    when 16#001E4# => romdata <= X"AF398196";
    when 16#001E5# => romdata <= X"76822A83";
    when 16#001E6# => romdata <= X"06535780";
    when 16#001E7# => romdata <= X"5180FADB";
    when 16#001E8# => romdata <= X"3FFEE139";
    when 16#001E9# => romdata <= X"81965780";
    when 16#001EA# => romdata <= X"5181829F";
    when 16#001EB# => romdata <= X"3F815181";
    when 16#001EC# => romdata <= X"82993FFE";
    when 16#001ED# => romdata <= X"E839FE3D";
    when 16#001EE# => romdata <= X"0D815194";
    when 16#001EF# => romdata <= X"8A3FB008";
    when 16#001F0# => romdata <= X"81FF0681";
    when 16#001F1# => romdata <= X"F5C00871";
    when 16#001F2# => romdata <= X"88120C53";
    when 16#001F3# => romdata <= X"B00C843D";
    when 16#001F4# => romdata <= X"0D04FC3D";
    when 16#001F5# => romdata <= X"0D815193";
    when 16#001F6# => romdata <= X"EE3FB008";
    when 16#001F7# => romdata <= X"81FF0654";
    when 16#001F8# => romdata <= X"825193E3";
    when 16#001F9# => romdata <= X"3FB00881";
    when 16#001FA# => romdata <= X"FF0681F6";
    when 16#001FB# => romdata <= X"8C088411";
    when 16#001FC# => romdata <= X"0870FE8F";
    when 16#001FD# => romdata <= X"0A067798";
    when 16#001FE# => romdata <= X"2B075154";
    when 16#001FF# => romdata <= X"56537280";
    when 16#00200# => romdata <= X"2E863871";
    when 16#00201# => romdata <= X"810A0752";
    when 16#00202# => romdata <= X"7184160C";
    when 16#00203# => romdata <= X"71B00C86";
    when 16#00204# => romdata <= X"3D0D04FF";
    when 16#00205# => romdata <= X"3D0D81F6";
    when 16#00206# => romdata <= X"8C087008";
    when 16#00207# => romdata <= X"709E2A70";
    when 16#00208# => romdata <= X"81065152";
    when 16#00209# => romdata <= X"53518152";
    when 16#0020A# => romdata <= X"70833870";
    when 16#0020B# => romdata <= X"5271B00C";
    when 16#0020C# => romdata <= X"833D0D04";
    when 16#0020D# => romdata <= X"FC3D0D81";
    when 16#0020E# => romdata <= X"51938C3F";
    when 16#0020F# => romdata <= X"B00881FF";
    when 16#00210# => romdata <= X"0681CDE4";
    when 16#00211# => romdata <= X"52558184";
    when 16#00212# => romdata <= X"DE3F81F6";
    when 16#00213# => romdata <= X"8C087008";
    when 16#00214# => romdata <= X"709E2A70";
    when 16#00215# => romdata <= X"81065154";
    when 16#00216# => romdata <= X"54548153";
    when 16#00217# => romdata <= X"71833871";
    when 16#00218# => romdata <= X"5372802E";
    when 16#00219# => romdata <= X"80CB3881";
    when 16#0021A# => romdata <= X"CDF45181";
    when 16#0021B# => romdata <= X"84B93F81";
    when 16#0021C# => romdata <= X"CDE45181";
    when 16#0021D# => romdata <= X"84B13F74";
    when 16#0021E# => romdata <= X"802EAC38";
    when 16#0021F# => romdata <= X"81CDFC51";
    when 16#00220# => romdata <= X"8184A43F";
    when 16#00221# => romdata <= X"81F68C08";
    when 16#00222# => romdata <= X"84110870";
    when 16#00223# => romdata <= X"FD0A0655";
    when 16#00224# => romdata <= X"53547480";
    when 16#00225# => romdata <= X"2E863871";
    when 16#00226# => romdata <= X"820A0753";
    when 16#00227# => romdata <= X"7284150C";
    when 16#00228# => romdata <= X"71B00C86";
    when 16#00229# => romdata <= X"3D0D0481";
    when 16#0022A# => romdata <= X"CE885181";
    when 16#0022B# => romdata <= X"83F93FCC";
    when 16#0022C# => romdata <= X"3981CE88";
    when 16#0022D# => romdata <= X"518183EF";
    when 16#0022E# => romdata <= X"3F81CDF4";
    when 16#0022F# => romdata <= X"518183E7";
    when 16#00230# => romdata <= X"3F81CDE4";
    when 16#00231# => romdata <= X"518183DF";
    when 16#00232# => romdata <= X"3F74FFB0";
    when 16#00233# => romdata <= X"38D939FD";
    when 16#00234# => romdata <= X"3D0D8151";
    when 16#00235# => romdata <= X"91F13FB0";
    when 16#00236# => romdata <= X"0881FF06";
    when 16#00237# => romdata <= X"81CE9052";
    when 16#00238# => romdata <= X"548183C3";
    when 16#00239# => romdata <= X"3F73A638";
    when 16#0023A# => romdata <= X"81C6E451";
    when 16#0023B# => romdata <= X"8183B83F";
    when 16#0023C# => romdata <= X"81F68C08";
    when 16#0023D# => romdata <= X"84110870";
    when 16#0023E# => romdata <= X"FB0A0684";
    when 16#0023F# => romdata <= X"130C5353";
    when 16#00240# => romdata <= X"8A518183";
    when 16#00241# => romdata <= X"883F73B0";
    when 16#00242# => romdata <= X"0C853D0D";
    when 16#00243# => romdata <= X"0481CEA4";
    when 16#00244# => romdata <= X"51818393";
    when 16#00245# => romdata <= X"3F81F68C";
    when 16#00246# => romdata <= X"08841108";
    when 16#00247# => romdata <= X"70840A07";
    when 16#00248# => romdata <= X"84130C53";
    when 16#00249# => romdata <= X"538A5181";
    when 16#0024A# => romdata <= X"82E33F73";
    when 16#0024B# => romdata <= X"B00C853D";
    when 16#0024C# => romdata <= X"0D04F73D";
    when 16#0024D# => romdata <= X"0D853D54";
    when 16#0024E# => romdata <= X"965381CE";
    when 16#0024F# => romdata <= X"B0527351";
    when 16#00250# => romdata <= X"8189FC3F";
    when 16#00251# => romdata <= X"AD8B3F81";
    when 16#00252# => romdata <= X"5190FC3F";
    when 16#00253# => romdata <= X"80528051";
    when 16#00254# => romdata <= X"AAEB3F73";
    when 16#00255# => romdata <= X"53805281";
    when 16#00256# => romdata <= X"D68451BF";
    when 16#00257# => romdata <= X"AA3F8052";
    when 16#00258# => romdata <= X"8151AAD9";
    when 16#00259# => romdata <= X"3F735382";
    when 16#0025A# => romdata <= X"5281D684";
    when 16#0025B# => romdata <= X"51BF983F";
    when 16#0025C# => romdata <= X"80528251";
    when 16#0025D# => romdata <= X"AAC73F73";
    when 16#0025E# => romdata <= X"53815281";
    when 16#0025F# => romdata <= X"D68451BF";
    when 16#00260# => romdata <= X"863F8052";
    when 16#00261# => romdata <= X"8451AAB5";
    when 16#00262# => romdata <= X"3F735384";
    when 16#00263# => romdata <= X"5281D684";
    when 16#00264# => romdata <= X"51BEF43F";
    when 16#00265# => romdata <= X"80528551";
    when 16#00266# => romdata <= X"AAA33F73";
    when 16#00267# => romdata <= X"53905281";
    when 16#00268# => romdata <= X"D68451BE";
    when 16#00269# => romdata <= X"E23F8052";
    when 16#0026A# => romdata <= X"8651AA91";
    when 16#0026B# => romdata <= X"3F735383";
    when 16#0026C# => romdata <= X"5281D684";
    when 16#0026D# => romdata <= X"51BED03F";
    when 16#0026E# => romdata <= X"8B3D0D04";
    when 16#0026F# => romdata <= X"FEF43F80";
    when 16#00270# => romdata <= X"0BB00C04";
    when 16#00271# => romdata <= X"FC3D0DAB";
    when 16#00272# => romdata <= X"973F81BE";
    when 16#00273# => romdata <= X"94548055";
    when 16#00274# => romdata <= X"84527451";
    when 16#00275# => romdata <= X"A9E73F80";
    when 16#00276# => romdata <= X"53737081";
    when 16#00277# => romdata <= X"05553351";
    when 16#00278# => romdata <= X"AAE13F81";
    when 16#00279# => romdata <= X"137081FF";
    when 16#0027A# => romdata <= X"06515380";
    when 16#0027B# => romdata <= X"DC7327E9";
    when 16#0027C# => romdata <= X"38811570";
    when 16#0027D# => romdata <= X"81FF0656";
    when 16#0027E# => romdata <= X"53877527";
    when 16#0027F# => romdata <= X"D338800B";
    when 16#00280# => romdata <= X"B00C863D";
    when 16#00281# => romdata <= X"0D04FD3D";
    when 16#00282# => romdata <= X"0D81F5DC";
    when 16#00283# => romdata <= X"337081FF";
    when 16#00284# => romdata <= X"06545472";
    when 16#00285# => romdata <= X"BF26AB38";
    when 16#00286# => romdata <= X"81F5DC33";
    when 16#00287# => romdata <= X"7081FF06";
    when 16#00288# => romdata <= X"81F5C008";
    when 16#00289# => romdata <= X"5288120C";
    when 16#0028A# => romdata <= X"5480E452";
    when 16#0028B# => romdata <= X"94865194";
    when 16#0028C# => romdata <= X"853F81F5";
    when 16#0028D# => romdata <= X"DC338105";
    when 16#0028E# => romdata <= X"537281F5";
    when 16#0028F# => romdata <= X"DC34853D";
    when 16#00290# => romdata <= X"0D0480E4";
    when 16#00291# => romdata <= X"5294DB51";
    when 16#00292# => romdata <= X"93EC3F81";
    when 16#00293# => romdata <= X"F5DC3381";
    when 16#00294# => romdata <= X"05537281";
    when 16#00295# => romdata <= X"F5DC3485";
    when 16#00296# => romdata <= X"3D0D04FD";
    when 16#00297# => romdata <= X"3D0D81F5";
    when 16#00298# => romdata <= X"DC337081";
    when 16#00299# => romdata <= X"FF065454";
    when 16#0029A# => romdata <= X"72BF2680";
    when 16#0029B# => romdata <= X"C83881F5";
    when 16#0029C# => romdata <= X"DC337081";
    when 16#0029D# => romdata <= X"FF0681F5";
    when 16#0029E# => romdata <= X"C0085688";
    when 16#0029F# => romdata <= X"160C5381";
    when 16#002A0# => romdata <= X"F5DC3370";
    when 16#002A1# => romdata <= X"81FF0655";
    when 16#002A2# => romdata <= X"5373BF2E";
    when 16#002A3# => romdata <= X"80D03880";
    when 16#002A4# => romdata <= X"E45294DB";
    when 16#002A5# => romdata <= X"51939F3F";
    when 16#002A6# => romdata <= X"81F5DC33";
    when 16#002A7# => romdata <= X"81055372";
    when 16#002A8# => romdata <= X"81F5DC34";
    when 16#002A9# => romdata <= X"81F5DC33";
    when 16#002AA# => romdata <= X"80FF0653";
    when 16#002AB# => romdata <= X"7281F5DC";
    when 16#002AC# => romdata <= X"34853D0D";
    when 16#002AD# => romdata <= X"0481F5DC";
    when 16#002AE# => romdata <= X"337081FF";
    when 16#002AF# => romdata <= X"0680FF71";
    when 16#002B0# => romdata <= X"3181F5C0";
    when 16#002B1# => romdata <= X"08528812";
    when 16#002B2# => romdata <= X"0C555381";
    when 16#002B3# => romdata <= X"F5DC3370";
    when 16#002B4# => romdata <= X"81FF0655";
    when 16#002B5# => romdata <= X"5373BF2E";
    when 16#002B6# => romdata <= X"098106FF";
    when 16#002B7# => romdata <= X"B23880CE";
    when 16#002B8# => romdata <= X"905294DB";
    when 16#002B9# => romdata <= X"5192CF3F";
    when 16#002BA# => romdata <= X"81F5DC33";
    when 16#002BB# => romdata <= X"81055372";
    when 16#002BC# => romdata <= X"81F5DC34";
    when 16#002BD# => romdata <= X"81F5DC33";
    when 16#002BE# => romdata <= X"80FF0653";
    when 16#002BF# => romdata <= X"7281F5DC";
    when 16#002C0# => romdata <= X"34853D0D";
    when 16#002C1# => romdata <= X"04810B81";
    when 16#002C2# => romdata <= X"F5C43404";
    when 16#002C3# => romdata <= X"FD3D0D82";
    when 16#002C4# => romdata <= X"85E40852";
    when 16#002C5# => romdata <= X"F881C08E";
    when 16#002C6# => romdata <= X"800B81F6";
    when 16#002C7# => romdata <= X"8C085553";
    when 16#002C8# => romdata <= X"71802E80";
    when 16#002C9# => romdata <= X"F8387281";
    when 16#002CA# => romdata <= X"FF068415";
    when 16#002CB# => romdata <= X"0C81F5DC";
    when 16#002CC# => romdata <= X"337081FF";
    when 16#002CD# => romdata <= X"06515271";
    when 16#002CE# => romdata <= X"802E80C2";
    when 16#002CF# => romdata <= X"38729F2A";
    when 16#002D0# => romdata <= X"73100753";
    when 16#002D1# => romdata <= X"8285E833";
    when 16#002D2# => romdata <= X"7081FF06";
    when 16#002D3# => romdata <= X"51527180";
    when 16#002D4# => romdata <= X"2ED43880";
    when 16#002D5# => romdata <= X"0B8285E8";
    when 16#002D6# => romdata <= X"3490FB3F";
    when 16#002D7# => romdata <= X"81F5C433";
    when 16#002D8# => romdata <= X"547380E4";
    when 16#002D9# => romdata <= X"3881F68C";
    when 16#002DA# => romdata <= X"087381FF";
    when 16#002DB# => romdata <= X"0684120C";
    when 16#002DC# => romdata <= X"81F5DC33";
    when 16#002DD# => romdata <= X"7081FF06";
    when 16#002DE# => romdata <= X"51535471";
    when 16#002DF# => romdata <= X"C0387281";
    when 16#002E0# => romdata <= X"2A739F2B";
    when 16#002E1# => romdata <= X"0753FFBC";
    when 16#002E2# => romdata <= X"3972812A";
    when 16#002E3# => romdata <= X"739F2B07";
    when 16#002E4# => romdata <= X"5380FD51";
    when 16#002E5# => romdata <= X"8181A33F";
    when 16#002E6# => romdata <= X"81F68C08";
    when 16#002E7# => romdata <= X"547281FF";
    when 16#002E8# => romdata <= X"0684150C";
    when 16#002E9# => romdata <= X"81F5DC33";
    when 16#002EA# => romdata <= X"7081FF06";
    when 16#002EB# => romdata <= X"53547180";
    when 16#002EC# => romdata <= X"2ED73872";
    when 16#002ED# => romdata <= X"9F2A7310";
    when 16#002EE# => romdata <= X"075380FD";
    when 16#002EF# => romdata <= X"518180FA";
    when 16#002F0# => romdata <= X"3F81F68C";
    when 16#002F1# => romdata <= X"0854D639";
    when 16#002F2# => romdata <= X"800BB00C";
    when 16#002F3# => romdata <= X"853D0D04";
    when 16#002F4# => romdata <= X"FE3D0D81";
    when 16#002F5# => romdata <= X"F6900898";
    when 16#002F6# => romdata <= X"11087084";
    when 16#002F7# => romdata <= X"2A708106";
    when 16#002F8# => romdata <= X"51535353";
    when 16#002F9# => romdata <= X"70802E8D";
    when 16#002FA# => romdata <= X"3871EF06";
    when 16#002FB# => romdata <= X"98140C81";
    when 16#002FC# => romdata <= X"0B8285E8";
    when 16#002FD# => romdata <= X"34843D0D";
    when 16#002FE# => romdata <= X"04FB3D0D";
    when 16#002FF# => romdata <= X"81F68C08";
    when 16#00300# => romdata <= X"7008810A";
    when 16#00301# => romdata <= X"068285E4";
    when 16#00302# => romdata <= X"0C548180";
    when 16#00303# => romdata <= X"D03F8180";
    when 16#00304# => romdata <= X"F23F91DF";
    when 16#00305# => romdata <= X"3F81F690";
    when 16#00306# => romdata <= X"08981108";
    when 16#00307# => romdata <= X"88079812";
    when 16#00308# => romdata <= X"0C548285";
    when 16#00309# => romdata <= X"E4085372";
    when 16#0030A# => romdata <= X"802E85A9";
    when 16#0030B# => romdata <= X"388194F7";
    when 16#0030C# => romdata <= X"0B829EBC";
    when 16#0030D# => romdata <= X"0C81CEC8";
    when 16#0030E# => romdata <= X"5180FCEB";
    when 16#0030F# => romdata <= X"3F8C5180";
    when 16#00310# => romdata <= X"FCCB3F81";
    when 16#00311# => romdata <= X"CEB05180";
    when 16#00312# => romdata <= X"FCDD3F82";
    when 16#00313# => romdata <= X"85E40880";
    when 16#00314# => romdata <= X"2E81EE38";
    when 16#00315# => romdata <= X"81CECC51";
    when 16#00316# => romdata <= X"80FCCC3F";
    when 16#00317# => romdata <= X"8285E408";
    when 16#00318# => romdata <= X"5473802E";
    when 16#00319# => romdata <= X"82F33881";
    when 16#0031A# => romdata <= X"F5E00854";
    when 16#0031B# => romdata <= X"81740C81";
    when 16#0031C# => romdata <= X"F68C0884";
    when 16#0031D# => romdata <= X"11087056";
    when 16#0031E# => romdata <= X"57558053";
    when 16#0031F# => romdata <= X"73FE8F0A";
    when 16#00320# => romdata <= X"0673982B";
    when 16#00321# => romdata <= X"07708417";
    when 16#00322# => romdata <= X"0C811470";
    when 16#00323# => romdata <= X"81FF0651";
    when 16#00324# => romdata <= X"54548F73";
    when 16#00325# => romdata <= X"27E63875";
    when 16#00326# => romdata <= X"84160C81";
    when 16#00327# => romdata <= X"F5CC0853";
    when 16#00328# => romdata <= X"800BB814";
    when 16#00329# => romdata <= X"0C81F5FC";
    when 16#0032A# => romdata <= X"087008FE";
    when 16#0032B# => romdata <= X"8006710C";
    when 16#0032C# => romdata <= X"54A0808D";
    when 16#0032D# => romdata <= X"0A085180";
    when 16#0032E# => romdata <= X"FDB73F8A";
    when 16#0032F# => romdata <= X"5180FBCD";
    when 16#00330# => romdata <= X"3F825296";
    when 16#00331# => romdata <= X"85518EEE";
    when 16#00332# => romdata <= X"3FF881C0";
    when 16#00333# => romdata <= X"8E800B81";
    when 16#00334# => romdata <= X"F68C0856";
    when 16#00335# => romdata <= X"548285E4";
    when 16#00336# => romdata <= X"08802E81";
    when 16#00337# => romdata <= X"D1387381";
    when 16#00338# => romdata <= X"FF068416";
    when 16#00339# => romdata <= X"0C81F5DC";
    when 16#0033A# => romdata <= X"337081FF";
    when 16#0033B# => romdata <= X"06545672";
    when 16#0033C# => romdata <= X"802E80C2";
    when 16#0033D# => romdata <= X"38739F2A";
    when 16#0033E# => romdata <= X"74100754";
    when 16#0033F# => romdata <= X"8285E833";
    when 16#00340# => romdata <= X"7081FF06";
    when 16#00341# => romdata <= X"57537580";
    when 16#00342# => romdata <= X"2ED43880";
    when 16#00343# => romdata <= X"0B8285E8";
    when 16#00344# => romdata <= X"348DC33F";
    when 16#00345# => romdata <= X"81F5C433";
    when 16#00346# => romdata <= X"557484FB";
    when 16#00347# => romdata <= X"3881F68C";
    when 16#00348# => romdata <= X"087481FF";
    when 16#00349# => romdata <= X"0684120C";
    when 16#0034A# => romdata <= X"81F5DC33";
    when 16#0034B# => romdata <= X"7081FF06";
    when 16#0034C# => romdata <= X"55575572";
    when 16#0034D# => romdata <= X"C0387381";
    when 16#0034E# => romdata <= X"2A749F2B";
    when 16#0034F# => romdata <= X"0754FFBC";
    when 16#00350# => romdata <= X"3981CED8";
    when 16#00351# => romdata <= X"5180FADF";
    when 16#00352# => romdata <= X"3F810A51";
    when 16#00353# => romdata <= X"80FAD83F";
    when 16#00354# => romdata <= X"81CEEC51";
    when 16#00355# => romdata <= X"80FAD03F";
    when 16#00356# => romdata <= X"81CF9451";
    when 16#00357# => romdata <= X"80FAC83F";
    when 16#00358# => romdata <= X"B45180FC";
    when 16#00359# => romdata <= X"8C3F81CF";
    when 16#0035A# => romdata <= X"A85180FA";
    when 16#0035B# => romdata <= X"BA3F81CF";
    when 16#0035C# => romdata <= X"B05180FA";
    when 16#0035D# => romdata <= X"B23F81CF";
    when 16#0035E# => romdata <= X"BC5180FA";
    when 16#0035F# => romdata <= X"AA3F81CF";
    when 16#00360# => romdata <= X"C45180FA";
    when 16#00361# => romdata <= X"A23F81CF";
    when 16#00362# => romdata <= X"E05180FA";
    when 16#00363# => romdata <= X"9A3F8285";
    when 16#00364# => romdata <= X"E4085473";
    when 16#00365# => romdata <= X"FDD13880";
    when 16#00366# => romdata <= X"C0397381";
    when 16#00367# => romdata <= X"2A749F2B";
    when 16#00368# => romdata <= X"075480FD";
    when 16#00369# => romdata <= X"5180FD92";
    when 16#0036A# => romdata <= X"3F81F68C";
    when 16#0036B# => romdata <= X"08557381";
    when 16#0036C# => romdata <= X"FF068416";
    when 16#0036D# => romdata <= X"0C81F5DC";
    when 16#0036E# => romdata <= X"337081FF";
    when 16#0036F# => romdata <= X"06565674";
    when 16#00370# => romdata <= X"802ED738";
    when 16#00371# => romdata <= X"739F2A74";
    when 16#00372# => romdata <= X"10075480";
    when 16#00373# => romdata <= X"FD5180FC";
    when 16#00374# => romdata <= X"E93F81F6";
    when 16#00375# => romdata <= X"8C0855D6";
    when 16#00376# => romdata <= X"39889B0B";
    when 16#00377# => romdata <= X"829EBC0C";
    when 16#00378# => romdata <= X"81CFE851";
    when 16#00379# => romdata <= X"80F9C03F";
    when 16#0037A# => romdata <= X"810A5180";
    when 16#0037B# => romdata <= X"F9B93F81";
    when 16#0037C# => romdata <= X"D0805180";
    when 16#0037D# => romdata <= X"F9B13F81";
    when 16#0037E# => romdata <= X"F5CC0874";
    when 16#0037F# => romdata <= X"B4120C74";
    when 16#00380# => romdata <= X"B8120C55";
    when 16#00381# => romdata <= X"81D09851";
    when 16#00382# => romdata <= X"80F99C3F";
    when 16#00383# => romdata <= X"735180DD";
    when 16#00384# => romdata <= X"823FB008";
    when 16#00385# => romdata <= X"982B5372";
    when 16#00386# => romdata <= X"82C83881";
    when 16#00387# => romdata <= X"D0A45180";
    when 16#00388# => romdata <= X"F9853F81";
    when 16#00389# => romdata <= X"F68C0870";
    when 16#0038A# => romdata <= X"08709E2A";
    when 16#0038B# => romdata <= X"81065557";
    when 16#0038C# => romdata <= X"54815572";
    when 16#0038D# => romdata <= X"802E81BA";
    when 16#0038E# => romdata <= X"387481FF";
    when 16#0038F# => romdata <= X"06841508";
    when 16#00390# => romdata <= X"70FD0A06";
    when 16#00391# => romdata <= X"58565372";
    when 16#00392# => romdata <= X"802E8638";
    when 16#00393# => romdata <= X"74820A07";
    when 16#00394# => romdata <= X"56758415";
    when 16#00395# => romdata <= X"0C730870";
    when 16#00396# => romdata <= X"9E2A8106";
    when 16#00397# => romdata <= X"54558154";
    when 16#00398# => romdata <= X"72833872";
    when 16#00399# => romdata <= X"5473802E";
    when 16#0039A# => romdata <= X"818D3881";
    when 16#0039B# => romdata <= X"D0B05180";
    when 16#0039C# => romdata <= X"F8B53F81";
    when 16#0039D# => romdata <= X"5180F4D3";
    when 16#0039E# => romdata <= X"3F81F68C";
    when 16#0039F# => romdata <= X"08841108";
    when 16#003A0# => romdata <= X"840A0784";
    when 16#003A1# => romdata <= X"120C5581";
    when 16#003A2# => romdata <= X"D0BC5180";
    when 16#003A3# => romdata <= X"F8993F81";
    when 16#003A4# => romdata <= X"F5CC0854";
    when 16#003A5# => romdata <= X"800BB815";
    when 16#003A6# => romdata <= X"0C81F5E0";
    when 16#003A7# => romdata <= X"08568176";
    when 16#003A8# => romdata <= X"0C88800B";
    when 16#003A9# => romdata <= X"829EBC0C";
    when 16#003AA# => romdata <= X"A7885293";
    when 16#003AB# => romdata <= X"C4518B86";
    when 16#003AC# => romdata <= X"3F87E852";
    when 16#003AD# => romdata <= X"9486518A";
    when 16#003AE# => romdata <= X"FD3FEB98";
    when 16#003AF# => romdata <= X"3F81F5E0";
    when 16#003B0# => romdata <= X"08548174";
    when 16#003B1# => romdata <= X"0C81F68C";
    when 16#003B2# => romdata <= X"08841108";
    when 16#003B3# => romdata <= X"70565755";
    when 16#003B4# => romdata <= X"8053FBA8";
    when 16#003B5# => romdata <= X"3980FCE9";
    when 16#003B6# => romdata <= X"3F9DEA3F";
    when 16#003B7# => romdata <= X"A1F33F72";
    when 16#003B8# => romdata <= X"5281D684";
    when 16#003B9# => romdata <= X"51A3CC3F";
    when 16#003BA# => romdata <= X"88800B82";
    when 16#003BB# => romdata <= X"9EBC0CFA";
    when 16#003BC# => romdata <= X"C4397255";
    when 16#003BD# => romdata <= X"FEC33981";
    when 16#003BE# => romdata <= X"D0C85180";
    when 16#003BF# => romdata <= X"F7A93F81";
    when 16#003C0# => romdata <= X"F5CC08B8";
    when 16#003C1# => romdata <= X"1108810A";
    when 16#003C2# => romdata <= X"07B8120C";
    when 16#003C3# => romdata <= X"5481D0B0";
    when 16#003C4# => romdata <= X"5180F793";
    when 16#003C5# => romdata <= X"3F815180";
    when 16#003C6# => romdata <= X"F3B13F81";
    when 16#003C7# => romdata <= X"F68C0884";
    when 16#003C8# => romdata <= X"1108840A";
    when 16#003C9# => romdata <= X"0784120C";
    when 16#003CA# => romdata <= X"5581D0BC";
    when 16#003CB# => romdata <= X"5180F6F7";
    when 16#003CC# => romdata <= X"3F81F5CC";
    when 16#003CD# => romdata <= X"0854800B";
    when 16#003CE# => romdata <= X"B8150C81";
    when 16#003CF# => romdata <= X"F5E00856";
    when 16#003D0# => romdata <= X"81760C88";
    when 16#003D1# => romdata <= X"800B829E";
    when 16#003D2# => romdata <= X"BC0CA788";
    when 16#003D3# => romdata <= X"5293C451";
    when 16#003D4# => romdata <= X"89E43F87";
    when 16#003D5# => romdata <= X"E8529486";
    when 16#003D6# => romdata <= X"5189DB3F";
    when 16#003D7# => romdata <= X"E9F63FFE";
    when 16#003D8# => romdata <= X"DC3981D0";
    when 16#003D9# => romdata <= X"C85180F6";
    when 16#003DA# => romdata <= X"BE3F81F5";
    when 16#003DB# => romdata <= X"CC08B811";
    when 16#003DC# => romdata <= X"08810A07";
    when 16#003DD# => romdata <= X"B8120C56";
    when 16#003DE# => romdata <= X"81D0A451";
    when 16#003DF# => romdata <= X"80F6A83F";
    when 16#003E0# => romdata <= X"81F68C08";
    when 16#003E1# => romdata <= X"7008709E";
    when 16#003E2# => romdata <= X"2A810655";
    when 16#003E3# => romdata <= X"57548155";
    when 16#003E4# => romdata <= X"72FDA638";
    when 16#003E5# => romdata <= X"FEDC3980";
    when 16#003E6# => romdata <= X"FD983F80";
    when 16#003E7# => romdata <= X"0B829DD0";
    when 16#003E8# => romdata <= X"34800B82";
    when 16#003E9# => romdata <= X"9DCC3480";
    when 16#003EA# => romdata <= X"0B829DD4";
    when 16#003EB# => romdata <= X"0C04FC3D";
    when 16#003EC# => romdata <= X"0D829DCC";
    when 16#003ED# => romdata <= X"335372A7";
    when 16#003EE# => romdata <= X"2680C738";
    when 16#003EF# => romdata <= X"76527210";
    when 16#003F0# => romdata <= X"10107310";
    when 16#003F1# => romdata <= X"058285EC";
    when 16#003F2# => romdata <= X"05518182";
    when 16#003F3# => romdata <= X"803F7752";
    when 16#003F4# => romdata <= X"829DCC33";
    when 16#003F5# => romdata <= X"70902971";
    when 16#003F6# => romdata <= X"31701010";
    when 16#003F7# => romdata <= X"8288FC05";
    when 16#003F8# => romdata <= X"53565481";
    when 16#003F9# => romdata <= X"81E73F82";
    when 16#003FA# => romdata <= X"9DCC3370";
    when 16#003FB# => romdata <= X"1010829B";
    when 16#003FC# => romdata <= X"DC057A71";
    when 16#003FD# => romdata <= X"0C548105";
    when 16#003FE# => romdata <= X"5372829D";
    when 16#003FF# => romdata <= X"CC34863D";
    when 16#00400# => romdata <= X"0D0481D0";
    when 16#00401# => romdata <= X"D45180F5";
    when 16#00402# => romdata <= X"9E3F863D";
    when 16#00403# => romdata <= X"0D04803D";
    when 16#00404# => romdata <= X"0D81D0F0";
    when 16#00405# => romdata <= X"5180F58F";
    when 16#00406# => romdata <= X"3F823D0D";
    when 16#00407# => romdata <= X"04FE3D0D";
    when 16#00408# => romdata <= X"829DD408";
    when 16#00409# => romdata <= X"53728538";
    when 16#0040A# => romdata <= X"843D0D04";
    when 16#0040B# => romdata <= X"722DB008";
    when 16#0040C# => romdata <= X"53800B82";
    when 16#0040D# => romdata <= X"9DD40CB0";
    when 16#0040E# => romdata <= X"088D3881";
    when 16#0040F# => romdata <= X"D0F05180";
    when 16#00410# => romdata <= X"F4E53F84";
    when 16#00411# => romdata <= X"3D0D0481";
    when 16#00412# => romdata <= X"D5AC5180";
    when 16#00413# => romdata <= X"F4D93F72";
    when 16#00414# => romdata <= X"83FFFF26";
    when 16#00415# => romdata <= X"AF3881FF";
    when 16#00416# => romdata <= X"73279938";
    when 16#00417# => romdata <= X"72529051";
    when 16#00418# => romdata <= X"80F4E73F";
    when 16#00419# => romdata <= X"8A5180F4";
    when 16#0041A# => romdata <= X"A43F81D0";
    when 16#0041B# => romdata <= X"F05180F4";
    when 16#0041C# => romdata <= X"B63FD039";
    when 16#0041D# => romdata <= X"72528851";
    when 16#0041E# => romdata <= X"80F4CF3F";
    when 16#0041F# => romdata <= X"8A5180F4";
    when 16#00420# => romdata <= X"8C3FE739";
    when 16#00421# => romdata <= X"7252A051";
    when 16#00422# => romdata <= X"80F4BF3F";
    when 16#00423# => romdata <= X"8A5180F3";
    when 16#00424# => romdata <= X"FC3FD739";
    when 16#00425# => romdata <= X"FA3D0D02";
    when 16#00426# => romdata <= X"A3053356";
    when 16#00427# => romdata <= X"758D2E80";
    when 16#00428# => romdata <= X"F8387588";
    when 16#00429# => romdata <= X"32703077";
    when 16#0042A# => romdata <= X"80FF3270";
    when 16#0042B# => romdata <= X"30728025";
    when 16#0042C# => romdata <= X"71802507";
    when 16#0042D# => romdata <= X"54515658";
    when 16#0042E# => romdata <= X"55749538";
    when 16#0042F# => romdata <= X"9F76278C";
    when 16#00430# => romdata <= X"38829DD0";
    when 16#00431# => romdata <= X"335580CE";
    when 16#00432# => romdata <= X"7527B138";
    when 16#00433# => romdata <= X"883D0D04";
    when 16#00434# => romdata <= X"829DD033";
    when 16#00435# => romdata <= X"5675802E";
    when 16#00436# => romdata <= X"F3388851";
    when 16#00437# => romdata <= X"80F3AE3F";
    when 16#00438# => romdata <= X"A05180F3";
    when 16#00439# => romdata <= X"A83F8851";
    when 16#0043A# => romdata <= X"80F3A23F";
    when 16#0043B# => romdata <= X"829DD033";
    when 16#0043C# => romdata <= X"FF055776";
    when 16#0043D# => romdata <= X"829DD034";
    when 16#0043E# => romdata <= X"883D0D04";
    when 16#0043F# => romdata <= X"755180F3";
    when 16#00440# => romdata <= X"8C3F829D";
    when 16#00441# => romdata <= X"D0338111";
    when 16#00442# => romdata <= X"55577382";
    when 16#00443# => romdata <= X"9DD03475";
    when 16#00444# => romdata <= X"829CFC18";
    when 16#00445# => romdata <= X"34883D0D";
    when 16#00446# => romdata <= X"048A5180";
    when 16#00447# => romdata <= X"F2EF3F82";
    when 16#00448# => romdata <= X"9DD03381";
    when 16#00449# => romdata <= X"11565474";
    when 16#0044A# => romdata <= X"829DD034";
    when 16#0044B# => romdata <= X"800B829C";
    when 16#0044C# => romdata <= X"FC153480";
    when 16#0044D# => romdata <= X"56800B82";
    when 16#0044E# => romdata <= X"9CFC1733";
    when 16#0044F# => romdata <= X"565474A0";
    when 16#00450# => romdata <= X"2E833881";
    when 16#00451# => romdata <= X"5474802E";
    when 16#00452# => romdata <= X"90387380";
    when 16#00453# => romdata <= X"2E8B3881";
    when 16#00454# => romdata <= X"167081FF";
    when 16#00455# => romdata <= X"065757DD";
    when 16#00456# => romdata <= X"3975802E";
    when 16#00457# => romdata <= X"80C13880";
    when 16#00458# => romdata <= X"0B829DCC";
    when 16#00459# => romdata <= X"33555574";
    when 16#0045A# => romdata <= X"7427AC38";
    when 16#0045B# => romdata <= X"73577410";
    when 16#0045C# => romdata <= X"10107510";
    when 16#0045D# => romdata <= X"05765482";
    when 16#0045E# => romdata <= X"9CFC5382";
    when 16#0045F# => romdata <= X"85EC0551";
    when 16#00460# => romdata <= X"8180963F";
    when 16#00461# => romdata <= X"B008802E";
    when 16#00462# => romdata <= X"A8388115";
    when 16#00463# => romdata <= X"7081FF06";
    when 16#00464# => romdata <= X"56547675";
    when 16#00465# => romdata <= X"26D83881";
    when 16#00466# => romdata <= X"D0F45180";
    when 16#00467# => romdata <= X"F2893F81";
    when 16#00468# => romdata <= X"D0F05180";
    when 16#00469# => romdata <= X"F2813F80";
    when 16#0046A# => romdata <= X"0B829DD0";
    when 16#0046B# => romdata <= X"34883D0D";
    when 16#0046C# => romdata <= X"04741010";
    when 16#0046D# => romdata <= X"829BDC05";
    when 16#0046E# => romdata <= X"7008829D";
    when 16#0046F# => romdata <= X"D40C5680";
    when 16#00470# => romdata <= X"0B829DD0";
    when 16#00471# => romdata <= X"34E739F7";
    when 16#00472# => romdata <= X"3D0D02AF";
    when 16#00473# => romdata <= X"05335980";
    when 16#00474# => romdata <= X"0B829CFC";
    when 16#00475# => romdata <= X"33829CFC";
    when 16#00476# => romdata <= X"59555673";
    when 16#00477# => romdata <= X"A02E0981";
    when 16#00478# => romdata <= X"06963881";
    when 16#00479# => romdata <= X"167081FF";
    when 16#0047A# => romdata <= X"06829CFC";
    when 16#0047B# => romdata <= X"11703353";
    when 16#0047C# => romdata <= X"59575473";
    when 16#0047D# => romdata <= X"A02EEC38";
    when 16#0047E# => romdata <= X"80587779";
    when 16#0047F# => romdata <= X"2780EA38";
    when 16#00480# => romdata <= X"80773356";
    when 16#00481# => romdata <= X"5474742E";
    when 16#00482# => romdata <= X"83388154";
    when 16#00483# => romdata <= X"74A02E9A";
    when 16#00484# => romdata <= X"387380C5";
    when 16#00485# => romdata <= X"3874A02E";
    when 16#00486# => romdata <= X"91388118";
    when 16#00487# => romdata <= X"7081FF06";
    when 16#00488# => romdata <= X"59557878";
    when 16#00489# => romdata <= X"26DA3880";
    when 16#0048A# => romdata <= X"C0398116";
    when 16#0048B# => romdata <= X"7081FF06";
    when 16#0048C# => romdata <= X"829CFC11";
    when 16#0048D# => romdata <= X"70335752";
    when 16#0048E# => romdata <= X"575773A0";
    when 16#0048F# => romdata <= X"2E098106";
    when 16#00490# => romdata <= X"D9388116";
    when 16#00491# => romdata <= X"7081FF06";
    when 16#00492# => romdata <= X"829CFC11";
    when 16#00493# => romdata <= X"70335752";
    when 16#00494# => romdata <= X"575773A0";
    when 16#00495# => romdata <= X"2ED438C2";
    when 16#00496# => romdata <= X"39811670";
    when 16#00497# => romdata <= X"81FF0682";
    when 16#00498# => romdata <= X"9CFC1159";
    when 16#00499# => romdata <= X"5755FF98";
    when 16#0049A# => romdata <= X"3980538B";
    when 16#0049B# => romdata <= X"3DFC0552";
    when 16#0049C# => romdata <= X"76518182";
    when 16#0049D# => romdata <= X"E93F8B3D";
    when 16#0049E# => romdata <= X"0D04F73D";
    when 16#0049F# => romdata <= X"0D02AF05";
    when 16#004A0# => romdata <= X"3359800B";
    when 16#004A1# => romdata <= X"829CFC33";
    when 16#004A2# => romdata <= X"829CFC59";
    when 16#004A3# => romdata <= X"555673A0";
    when 16#004A4# => romdata <= X"2E098106";
    when 16#004A5# => romdata <= X"96388116";
    when 16#004A6# => romdata <= X"7081FF06";
    when 16#004A7# => romdata <= X"829CFC11";
    when 16#004A8# => romdata <= X"70335359";
    when 16#004A9# => romdata <= X"575473A0";
    when 16#004AA# => romdata <= X"2EEC3880";
    when 16#004AB# => romdata <= X"58777927";
    when 16#004AC# => romdata <= X"80EA3880";
    when 16#004AD# => romdata <= X"77335654";
    when 16#004AE# => romdata <= X"74742E83";
    when 16#004AF# => romdata <= X"38815474";
    when 16#004B0# => romdata <= X"A02E9A38";
    when 16#004B1# => romdata <= X"7380C538";
    when 16#004B2# => romdata <= X"74A02E91";
    when 16#004B3# => romdata <= X"38811870";
    when 16#004B4# => romdata <= X"81FF0659";
    when 16#004B5# => romdata <= X"55787826";
    when 16#004B6# => romdata <= X"DA3880C0";
    when 16#004B7# => romdata <= X"39811670";
    when 16#004B8# => romdata <= X"81FF0682";
    when 16#004B9# => romdata <= X"9CFC1170";
    when 16#004BA# => romdata <= X"33575257";
    when 16#004BB# => romdata <= X"5773A02E";
    when 16#004BC# => romdata <= X"098106D9";
    when 16#004BD# => romdata <= X"38811670";
    when 16#004BE# => romdata <= X"81FF0682";
    when 16#004BF# => romdata <= X"9CFC1170";
    when 16#004C0# => romdata <= X"33575257";
    when 16#004C1# => romdata <= X"5773A02E";
    when 16#004C2# => romdata <= X"D438C239";
    when 16#004C3# => romdata <= X"81167081";
    when 16#004C4# => romdata <= X"FF06829C";
    when 16#004C5# => romdata <= X"FC115957";
    when 16#004C6# => romdata <= X"55FF9839";
    when 16#004C7# => romdata <= X"90538B3D";
    when 16#004C8# => romdata <= X"FC055276";
    when 16#004C9# => romdata <= X"518184D3";
    when 16#004CA# => romdata <= X"3F8B3D0D";
    when 16#004CB# => romdata <= X"04FC3D0D";
    when 16#004CC# => romdata <= X"8A5180EE";
    when 16#004CD# => romdata <= X"D83F81D1";
    when 16#004CE# => romdata <= X"885180EE";
    when 16#004CF# => romdata <= X"EA3F800B";
    when 16#004D0# => romdata <= X"829DCC33";
    when 16#004D1# => romdata <= X"53537272";
    when 16#004D2# => romdata <= X"2780FB38";
    when 16#004D3# => romdata <= X"72101010";
    when 16#004D4# => romdata <= X"73100582";
    when 16#004D5# => romdata <= X"85EC0570";
    when 16#004D6# => romdata <= X"525480EE";
    when 16#004D7# => romdata <= X"CA3F7284";
    when 16#004D8# => romdata <= X"2B707431";
    when 16#004D9# => romdata <= X"822B8288";
    when 16#004DA# => romdata <= X"FC113351";
    when 16#004DB# => romdata <= X"53557180";
    when 16#004DC# => romdata <= X"2EBB3873";
    when 16#004DD# => romdata <= X"5180FBC2";
    when 16#004DE# => romdata <= X"3FB00881";
    when 16#004DF# => romdata <= X"FF065271";
    when 16#004E0# => romdata <= X"89269438";
    when 16#004E1# => romdata <= X"A05180EE";
    when 16#004E2# => romdata <= X"843F8112";
    when 16#004E3# => romdata <= X"7081FF06";
    when 16#004E4# => romdata <= X"53548972";
    when 16#004E5# => romdata <= X"27EE3881";
    when 16#004E6# => romdata <= X"D1A05180";
    when 16#004E7# => romdata <= X"EE893F74";
    when 16#004E8# => romdata <= X"7331822B";
    when 16#004E9# => romdata <= X"8288FC05";
    when 16#004EA# => romdata <= X"5180EDFB";
    when 16#004EB# => romdata <= X"3F8A5180";
    when 16#004EC# => romdata <= X"EDDB3F81";
    when 16#004ED# => romdata <= X"137081FF";
    when 16#004EE# => romdata <= X"06829DCC";
    when 16#004EF# => romdata <= X"33545455";
    when 16#004F0# => romdata <= X"717326FF";
    when 16#004F1# => romdata <= X"87388A51";
    when 16#004F2# => romdata <= X"80EDC23F";
    when 16#004F3# => romdata <= X"829DCC33";
    when 16#004F4# => romdata <= X"B00C863D";
    when 16#004F5# => romdata <= X"0D04FE3D";
    when 16#004F6# => romdata <= X"0D829EAC";
    when 16#004F7# => romdata <= X"22FF0551";
    when 16#004F8# => romdata <= X"70829EAC";
    when 16#004F9# => romdata <= X"237083FF";
    when 16#004FA# => romdata <= X"FF065170";
    when 16#004FB# => romdata <= X"80C43882";
    when 16#004FC# => romdata <= X"9EB03351";
    when 16#004FD# => romdata <= X"7081FF2E";
    when 16#004FE# => romdata <= X"B9387010";
    when 16#004FF# => romdata <= X"1010829D";
    when 16#00500# => romdata <= X"DC055271";
    when 16#00501# => romdata <= X"33829EB0";
    when 16#00502# => romdata <= X"34FE7234";
    when 16#00503# => romdata <= X"829EB033";
    when 16#00504# => romdata <= X"70101010";
    when 16#00505# => romdata <= X"829DDC05";
    when 16#00506# => romdata <= X"52538211";
    when 16#00507# => romdata <= X"22829EAC";
    when 16#00508# => romdata <= X"23841208";
    when 16#00509# => romdata <= X"53722D82";
    when 16#0050A# => romdata <= X"9EAC2251";
    when 16#0050B# => romdata <= X"70802EFF";
    when 16#0050C# => romdata <= X"BE38843D";
    when 16#0050D# => romdata <= X"0D04F93D";
    when 16#0050E# => romdata <= X"0D02AA05";
    when 16#0050F# => romdata <= X"22568055";
    when 16#00510# => romdata <= X"74101010";
    when 16#00511# => romdata <= X"829DDC05";
    when 16#00512# => romdata <= X"70335252";
    when 16#00513# => romdata <= X"7081FE2E";
    when 16#00514# => romdata <= X"99388115";
    when 16#00515# => romdata <= X"7081FF06";
    when 16#00516# => romdata <= X"5652748A";
    when 16#00517# => romdata <= X"2E098106";
    when 16#00518# => romdata <= X"DF38810B";
    when 16#00519# => romdata <= X"B00C893D";
    when 16#0051A# => romdata <= X"0D04829E";
    when 16#0051B# => romdata <= X"B0337081";
    when 16#0051C# => romdata <= X"FF06829E";
    when 16#0051D# => romdata <= X"AC225354";
    when 16#0051E# => romdata <= X"587281FF";
    when 16#0051F# => romdata <= X"2EB03872";
    when 16#00520# => romdata <= X"832B5470";
    when 16#00521# => romdata <= X"762780DE";
    when 16#00522# => romdata <= X"38757131";
    when 16#00523# => romdata <= X"7083FFFF";
    when 16#00524# => romdata <= X"0674829D";
    when 16#00525# => romdata <= X"DC173370";
    when 16#00526# => romdata <= X"832B829D";
    when 16#00527# => romdata <= X"DE112256";
    when 16#00528# => romdata <= X"58565257";
    when 16#00529# => romdata <= X"577281FF";
    when 16#0052A# => romdata <= X"2E098106";
    when 16#0052B# => romdata <= X"D6387272";
    when 16#0052C# => romdata <= X"34758213";
    when 16#0052D# => romdata <= X"23798413";
    when 16#0052E# => romdata <= X"0C7781FF";
    when 16#0052F# => romdata <= X"06547373";
    when 16#00530# => romdata <= X"2E963876";
    when 16#00531# => romdata <= X"10101082";
    when 16#00532# => romdata <= X"9DDC0553";
    when 16#00533# => romdata <= X"74733480";
    when 16#00534# => romdata <= X"5170B00C";
    when 16#00535# => romdata <= X"893D0D04";
    when 16#00536# => romdata <= X"74829EB0";
    when 16#00537# => romdata <= X"3475829E";
    when 16#00538# => romdata <= X"AC238051";
    when 16#00539# => romdata <= X"EC397076";
    when 16#0053A# => romdata <= X"31517082";
    when 16#0053B# => romdata <= X"9DDE1523";
    when 16#0053C# => romdata <= X"FFBC39FF";
    when 16#0053D# => romdata <= X"3D0D8A52";
    when 16#0053E# => romdata <= X"71101010";
    when 16#0053F# => romdata <= X"829DD405";
    when 16#00540# => romdata <= X"51FE7134";
    when 16#00541# => romdata <= X"FF127081";
    when 16#00542# => romdata <= X"FF065351";
    when 16#00543# => romdata <= X"71EA38FF";
    when 16#00544# => romdata <= X"0B829EB0";
    when 16#00545# => romdata <= X"34833D0D";
    when 16#00546# => romdata <= X"04F53D0D";
    when 16#00547# => romdata <= X"7D598A54";
    when 16#00548# => romdata <= X"81028405";
    when 16#00549# => romdata <= X"BA052257";
    when 16#0054A# => romdata <= X"5C80E453";
    when 16#0054B# => romdata <= X"805280EE";
    when 16#0054C# => romdata <= X"E83FB008";
    when 16#0054D# => romdata <= X"722E0981";
    when 16#0054E# => romdata <= X"06833881";
    when 16#0054F# => romdata <= X"5272802E";
    when 16#00550# => romdata <= X"B3387180";
    when 16#00551# => romdata <= X"2E923880";
    when 16#00552# => romdata <= X"E45180ED";
    when 16#00553# => romdata <= X"ED3FFF13";
    when 16#00554# => romdata <= X"7081FF06";
    when 16#00555# => romdata <= X"5452D539";
    when 16#00556# => romdata <= X"72802E98";
    when 16#00557# => romdata <= X"3880EECC";
    when 16#00558# => romdata <= X"3FB00881";
    when 16#00559# => romdata <= X"FF065271";
    when 16#0055A# => romdata <= X"952E82A7";
    when 16#0055B# => romdata <= X"387180C3";
    when 16#0055C# => romdata <= X"2E81F838";
    when 16#0055D# => romdata <= X"FF147081";
    when 16#0055E# => romdata <= X"FF065553";
    when 16#0055F# => romdata <= X"73FFAA38";
    when 16#00560# => romdata <= X"75802E81";
    when 16#00561# => romdata <= X"D6388A7C";
    when 16#00562# => romdata <= X"095C5A81";
    when 16#00563# => romdata <= X"5180EEBE";
    when 16#00564# => romdata <= X"3F7B5180";
    when 16#00565# => romdata <= X"EEB83F7A";
    when 16#00566# => romdata <= X"5180EEB2";
    when 16#00567# => romdata <= X"3F807055";
    when 16#00568# => romdata <= X"57818055";
    when 16#00569# => romdata <= X"FF157081";
    when 16#0056A# => romdata <= X"FF065652";
    when 16#0056B# => romdata <= X"9A537580";
    when 16#0056C# => romdata <= X"2E913878";
    when 16#0056D# => romdata <= X"7081055A";
    when 16#0056E# => romdata <= X"33FF1770";
    when 16#0056F# => romdata <= X"83FFFF06";
    when 16#00570# => romdata <= X"58535372";
    when 16#00571# => romdata <= X"5180EE86";
    when 16#00572# => romdata <= X"3F77802E";
    when 16#00573# => romdata <= X"81B13872";
    when 16#00574# => romdata <= X"882B7432";
    when 16#00575# => romdata <= X"53875472";
    when 16#00576# => romdata <= X"902B5280";
    when 16#00577# => romdata <= X"72248190";
    when 16#00578# => romdata <= X"38721083";
    when 16#00579# => romdata <= X"FFFE0653";
    when 16#0057A# => romdata <= X"FF145473";
    when 16#0057B# => romdata <= X"8025E838";
    when 16#0057C# => romdata <= X"7283FFFF";
    when 16#0057D# => romdata <= X"065474FF";
    when 16#0057E# => romdata <= X"AB387780";
    when 16#0057F# => romdata <= X"2E818B38";
    when 16#00580# => romdata <= X"73882A51";
    when 16#00581# => romdata <= X"80EDC73F";
    when 16#00582# => romdata <= X"7381FF06";
    when 16#00583# => romdata <= X"5180EDBE";
    when 16#00584# => romdata <= X"3F80ED85";
    when 16#00585# => romdata <= X"3FB008F9";
    when 16#00586# => romdata <= X"3880ED90";
    when 16#00587# => romdata <= X"3FB00881";
    when 16#00588# => romdata <= X"FF065271";
    when 16#00589# => romdata <= X"862E80F0";
    when 16#0058A# => romdata <= X"3871982E";
    when 16#0058B# => romdata <= X"80F538FF";
    when 16#0058C# => romdata <= X"1A7081FF";
    when 16#0058D# => romdata <= X"065B5479";
    when 16#0058E# => romdata <= X"FED138FE";
    when 16#0058F# => romdata <= X"5271B00C";
    when 16#00590# => romdata <= X"8D3D0D04";
    when 16#00591# => romdata <= X"80ECD23F";
    when 16#00592# => romdata <= X"B008F938";
    when 16#00593# => romdata <= X"80ECDD3F";
    when 16#00594# => romdata <= X"B00881FF";
    when 16#00595# => romdata <= X"06527186";
    when 16#00596# => romdata <= X"2EE33884";
    when 16#00597# => romdata <= X"5180ECEE";
    when 16#00598# => romdata <= X"3F80ECB5";
    when 16#00599# => romdata <= X"3FB008DC";
    when 16#0059A# => romdata <= X"38E23981";
    when 16#0059B# => romdata <= X"58FE9139";
    when 16#0059C# => romdata <= X"7210A0A1";
    when 16#0059D# => romdata <= X"327083FF";
    when 16#0059E# => romdata <= X"FF065452";
    when 16#0059F# => romdata <= X"FEEA3972";
    when 16#005A0# => romdata <= X"177081FF";
    when 16#005A1# => romdata <= X"065852FE";
    when 16#005A2# => romdata <= X"ED397651";
    when 16#005A3# => romdata <= X"80ECBF3F";
    when 16#005A4# => romdata <= X"FEFF3980";
    when 16#005A5# => romdata <= X"58FDE939";
    when 16#005A6# => romdata <= X"811C7081";
    when 16#005A7# => romdata <= X"FF065D55";
    when 16#005A8# => romdata <= X"FDDE39FF";
    when 16#005A9# => romdata <= X"0BB00C8D";
    when 16#005AA# => romdata <= X"3D0D04F6";
    when 16#005AB# => romdata <= X"3D0D7C7E";
    when 16#005AC# => romdata <= X"5B5980C3";
    when 16#005AD# => romdata <= X"578A5581";
    when 16#005AE# => romdata <= X"5B805880";
    when 16#005AF# => romdata <= X"E4538054";
    when 16#005B0# => romdata <= X"777A2482";
    when 16#005B1# => romdata <= X"B4387651";
    when 16#005B2# => romdata <= X"80EC833F";
    when 16#005B3# => romdata <= X"805280EB";
    when 16#005B4# => romdata <= X"C83FB008";
    when 16#005B5# => romdata <= X"722E0981";
    when 16#005B6# => romdata <= X"06833881";
    when 16#005B7# => romdata <= X"5272802E";
    when 16#005B8# => romdata <= X"81ED3871";
    when 16#005B9# => romdata <= X"802E9238";
    when 16#005BA# => romdata <= X"80E45180";
    when 16#005BB# => romdata <= X"EACC3FFF";
    when 16#005BC# => romdata <= X"137081FF";
    when 16#005BD# => romdata <= X"065452D4";
    when 16#005BE# => romdata <= X"3972802E";
    when 16#005BF# => romdata <= X"81D13880";
    when 16#005C0# => romdata <= X"EBAA3FB0";
    when 16#005C1# => romdata <= X"0881FF06";
    when 16#005C2# => romdata <= X"5271842E";
    when 16#005C3# => romdata <= X"82883871";
    when 16#005C4# => romdata <= X"842481CF";
    when 16#005C5# => romdata <= X"3871812E";
    when 16#005C6# => romdata <= X"09810681";
    when 16#005C7# => romdata <= X"B2388657";
    when 16#005C8# => romdata <= X"80EB893F";
    when 16#005C9# => romdata <= X"B00881FF";
    when 16#005CA# => romdata <= X"06537A73";
    when 16#005CB# => romdata <= X"2E833895";
    when 16#005CC# => romdata <= X"5780EAF8";
    when 16#005CD# => romdata <= X"3FB00809";
    when 16#005CE# => romdata <= X"7081FF06";
    when 16#005CF# => romdata <= X"57527A76";
    when 16#005D0# => romdata <= X"2E833895";
    when 16#005D1# => romdata <= X"57805380";
    when 16#005D2# => romdata <= X"EAE23F78";
    when 16#005D3# => romdata <= X"1356B008";
    when 16#005D4# => romdata <= X"76348113";
    when 16#005D5# => romdata <= X"7081FF06";
    when 16#005D6# => romdata <= X"70982B58";
    when 16#005D7# => romdata <= X"54527580";
    when 16#005D8# => romdata <= X"25E53880";
    when 16#005D9# => romdata <= X"56781670";
    when 16#005DA# => romdata <= X"3370882B";
    when 16#005DB# => romdata <= X"76325253";
    when 16#005DC# => romdata <= X"53875472";
    when 16#005DD# => romdata <= X"902B5280";
    when 16#005DE# => romdata <= X"7224818B";
    when 16#005DF# => romdata <= X"38721083";
    when 16#005E0# => romdata <= X"FFFE0653";
    when 16#005E1# => romdata <= X"FF145473";
    when 16#005E2# => romdata <= X"8025E838";
    when 16#005E3# => romdata <= X"7283FFFF";
    when 16#005E4# => romdata <= X"06811770";
    when 16#005E5# => romdata <= X"81FF0670";
    when 16#005E6# => romdata <= X"982B5658";
    when 16#005E7# => romdata <= X"53547280";
    when 16#005E8# => romdata <= X"25C33880";
    when 16#005E9# => romdata <= X"EA863FB0";
    when 16#005EA# => romdata <= X"0881FF06";
    when 16#005EB# => romdata <= X"74882A57";
    when 16#005EC# => romdata <= X"5372762E";
    when 16#005ED# => romdata <= X"83389557";
    when 16#005EE# => romdata <= X"80E9F13F";
    when 16#005EF# => romdata <= X"B00881FF";
    when 16#005F0# => romdata <= X"067481FF";
    when 16#005F1# => romdata <= X"06535675";
    when 16#005F2# => romdata <= X"722E80D7";
    when 16#005F3# => romdata <= X"389557FF";
    when 16#005F4# => romdata <= X"157081FF";
    when 16#005F5# => romdata <= X"06565274";
    when 16#005F6# => romdata <= X"FDE138FE";
    when 16#005F7# => romdata <= X"0BB00C8C";
    when 16#005F8# => romdata <= X"3D0D0471";
    when 16#005F9# => romdata <= X"982E0981";
    when 16#005FA# => romdata <= X"06E53886";
    when 16#005FB# => romdata <= X"5180E9DE";
    when 16#005FC# => romdata <= X"3FFF0BB0";
    when 16#005FD# => romdata <= X"0C8C3D0D";
    when 16#005FE# => romdata <= X"04985180";
    when 16#005FF# => romdata <= X"E9D03FFD";
    when 16#00600# => romdata <= X"0BB00C8C";
    when 16#00601# => romdata <= X"3D0D0472";
    when 16#00602# => romdata <= X"10A0A132";
    when 16#00603# => romdata <= X"7083FFFF";
    when 16#00604# => romdata <= X"065452FE";
    when 16#00605# => romdata <= X"EF398651";
    when 16#00606# => romdata <= X"80E9B33F";
    when 16#00607# => romdata <= X"77B00C8C";
    when 16#00608# => romdata <= X"3D0D0476";
    when 16#00609# => romdata <= X"862E0981";
    when 16#0060A# => romdata <= X"06FFA438";
    when 16#0060B# => romdata <= X"77848080";
    when 16#0060C# => romdata <= X"2982800A";
    when 16#0060D# => romdata <= X"0570902C";
    when 16#0060E# => romdata <= X"81801B81";
    when 16#0060F# => romdata <= X"1E7081FF";
    when 16#00610# => romdata <= X"065F575B";
    when 16#00611# => romdata <= X"595374FC";
    when 16#00612# => romdata <= X"F238FF8F";
    when 16#00613# => romdata <= X"39FE3D0D";
    when 16#00614# => romdata <= X"02930533";
    when 16#00615# => romdata <= X"02840597";
    when 16#00616# => romdata <= X"05335452";
    when 16#00617# => romdata <= X"71842E80";
    when 16#00618# => romdata <= X"ED387184";
    when 16#00619# => romdata <= X"24923871";
    when 16#0061A# => romdata <= X"812EAF38";
    when 16#0061B# => romdata <= X"81D1A451";
    when 16#0061C# => romdata <= X"80E4B43F";
    when 16#0061D# => romdata <= X"843D0D04";
    when 16#0061E# => romdata <= X"7180D52E";
    when 16#0061F# => romdata <= X"098106EC";
    when 16#00620# => romdata <= X"3881D1B0";
    when 16#00621# => romdata <= X"5180E49F";
    when 16#00622# => romdata <= X"3F728A26";
    when 16#00623# => romdata <= X"80CD3872";
    when 16#00624# => romdata <= X"101081D5";
    when 16#00625# => romdata <= X"D8055271";
    when 16#00626# => romdata <= X"080481D1";
    when 16#00627# => romdata <= X"BC5180E4";
    when 16#00628# => romdata <= X"863F729A";
    when 16#00629# => romdata <= X"2E829C38";
    when 16#0062A# => romdata <= X"729A2480";
    when 16#0062B# => romdata <= X"C638728C";
    when 16#0062C# => romdata <= X"2E829C38";
    when 16#0062D# => romdata <= X"728C2481";
    when 16#0062E# => romdata <= X"EF387286";
    when 16#0062F# => romdata <= X"2E098106";
    when 16#00630# => romdata <= X"9A3881D1";
    when 16#00631# => romdata <= X"C85180E3";
    when 16#00632# => romdata <= X"DE3F843D";
    when 16#00633# => romdata <= X"0D0481D1";
    when 16#00634# => romdata <= X"D85180E3";
    when 16#00635# => romdata <= X"D23F728F";
    when 16#00636# => romdata <= X"2E8D3881";
    when 16#00637# => romdata <= X"D1E45180";
    when 16#00638# => romdata <= X"E3C53F84";
    when 16#00639# => romdata <= X"3D0D0481";
    when 16#0063A# => romdata <= X"D1F45180";
    when 16#0063B# => romdata <= X"E3B93F84";
    when 16#0063C# => romdata <= X"3D0D0472";
    when 16#0063D# => romdata <= X"A82E81E3";
    when 16#0063E# => romdata <= X"3872A824";
    when 16#0063F# => romdata <= X"818D3872";
    when 16#00640# => romdata <= X"9D2E0981";
    when 16#00641# => romdata <= X"06D53881";
    when 16#00642# => romdata <= X"D28C5180";
    when 16#00643# => romdata <= X"E3993F84";
    when 16#00644# => romdata <= X"3D0D0481";
    when 16#00645# => romdata <= X"D2A85180";
    when 16#00646# => romdata <= X"E38D3F84";
    when 16#00647# => romdata <= X"3D0D0481";
    when 16#00648# => romdata <= X"D2C85180";
    when 16#00649# => romdata <= X"E3813F84";
    when 16#0064A# => romdata <= X"3D0D0481";
    when 16#0064B# => romdata <= X"D2DC5180";
    when 16#0064C# => romdata <= X"E2F53F84";
    when 16#0064D# => romdata <= X"3D0D0481";
    when 16#0064E# => romdata <= X"D2F85180";
    when 16#0064F# => romdata <= X"E2E93F84";
    when 16#00650# => romdata <= X"3D0D0481";
    when 16#00651# => romdata <= X"CEB05180";
    when 16#00652# => romdata <= X"E2DD3F84";
    when 16#00653# => romdata <= X"3D0D0481";
    when 16#00654# => romdata <= X"D3905180";
    when 16#00655# => romdata <= X"E2D13F84";
    when 16#00656# => romdata <= X"3D0D0481";
    when 16#00657# => romdata <= X"D3A45180";
    when 16#00658# => romdata <= X"E2C53F84";
    when 16#00659# => romdata <= X"3D0D0481";
    when 16#0065A# => romdata <= X"D3B45180";
    when 16#0065B# => romdata <= X"E2B93F84";
    when 16#0065C# => romdata <= X"3D0D0481";
    when 16#0065D# => romdata <= X"D3CC5180";
    when 16#0065E# => romdata <= X"E2AD3F84";
    when 16#0065F# => romdata <= X"3D0D0481";
    when 16#00660# => romdata <= X"D3E05180";
    when 16#00661# => romdata <= X"E2A13F84";
    when 16#00662# => romdata <= X"3D0D0472";
    when 16#00663# => romdata <= X"80C52E80";
    when 16#00664# => romdata <= X"D6387280";
    when 16#00665# => romdata <= X"E12E0981";
    when 16#00666# => romdata <= X"06FEC038";
    when 16#00667# => romdata <= X"81D3F051";
    when 16#00668# => romdata <= X"80E2843F";
    when 16#00669# => romdata <= X"843D0D04";
    when 16#0066A# => romdata <= X"728F2E80";
    when 16#0066B# => romdata <= X"C6387291";
    when 16#0066C# => romdata <= X"2E098106";
    when 16#0066D# => romdata <= X"FEA53881";
    when 16#0066E# => romdata <= X"D4805180";
    when 16#0066F# => romdata <= X"E1E93F84";
    when 16#00670# => romdata <= X"3D0D0481";
    when 16#00671# => romdata <= X"D4945180";
    when 16#00672# => romdata <= X"E1DD3F84";
    when 16#00673# => romdata <= X"3D0D0481";
    when 16#00674# => romdata <= X"D4B05180";
    when 16#00675# => romdata <= X"E1D13F84";
    when 16#00676# => romdata <= X"3D0D0481";
    when 16#00677# => romdata <= X"D4C05180";
    when 16#00678# => romdata <= X"E1C53F84";
    when 16#00679# => romdata <= X"3D0D0481";
    when 16#0067A# => romdata <= X"D4E05180";
    when 16#0067B# => romdata <= X"E1B93F84";
    when 16#0067C# => romdata <= X"3D0D0481";
    when 16#0067D# => romdata <= X"D4F85180";
    when 16#0067E# => romdata <= X"E1AD3F84";
    when 16#0067F# => romdata <= X"3D0D04F7";
    when 16#00680# => romdata <= X"3D0D02B3";
    when 16#00681# => romdata <= X"05337C70";
    when 16#00682# => romdata <= X"08C08080";
    when 16#00683# => romdata <= X"0659545A";
    when 16#00684# => romdata <= X"80567583";
    when 16#00685# => romdata <= X"2B7707BF";
    when 16#00686# => romdata <= X"E0800770";
    when 16#00687# => romdata <= X"70840552";
    when 16#00688# => romdata <= X"0871088C";
    when 16#00689# => romdata <= X"2ABFFE80";
    when 16#0068A# => romdata <= X"06790771";
    when 16#0068B# => romdata <= X"982A728C";
    when 16#0068C# => romdata <= X"2A9FFF06";
    when 16#0068D# => romdata <= X"73852A70";
    when 16#0068E# => romdata <= X"8F06759F";
    when 16#0068F# => romdata <= X"06565158";
    when 16#00690# => romdata <= X"5D585255";
    when 16#00691# => romdata <= X"58748D38";
    when 16#00692# => romdata <= X"8116568F";
    when 16#00693# => romdata <= X"7627C338";
    when 16#00694# => romdata <= X"8B3D0D04";
    when 16#00695# => romdata <= X"81D59451";
    when 16#00696# => romdata <= X"80E0CC3F";
    when 16#00697# => romdata <= X"755180E2";
    when 16#00698# => romdata <= X"903F8452";
    when 16#00699# => romdata <= X"B00851A5";
    when 16#0069A# => romdata <= X"CB3F81D5";
    when 16#0069B# => romdata <= X"A05180E0";
    when 16#0069C# => romdata <= X"B63F7452";
    when 16#0069D# => romdata <= X"885180E0";
    when 16#0069E# => romdata <= X"D13F8452";
    when 16#0069F# => romdata <= X"B00851A5";
    when 16#006A0# => romdata <= X"B33F81D5";
    when 16#006A1# => romdata <= X"A85180E0";
    when 16#006A2# => romdata <= X"9E3F7852";
    when 16#006A3# => romdata <= X"905180E0";
    when 16#006A4# => romdata <= X"B93F8652";
    when 16#006A5# => romdata <= X"B00851A5";
    when 16#006A6# => romdata <= X"9B3F81D5";
    when 16#006A7# => romdata <= X"B05180E0";
    when 16#006A8# => romdata <= X"863F7251";
    when 16#006A9# => romdata <= X"80E1CA3F";
    when 16#006AA# => romdata <= X"8452B008";
    when 16#006AB# => romdata <= X"51A5853F";
    when 16#006AC# => romdata <= X"81D5B851";
    when 16#006AD# => romdata <= X"80DFF03F";
    when 16#006AE# => romdata <= X"735180E1";
    when 16#006AF# => romdata <= X"B43F8452";
    when 16#006B0# => romdata <= X"B00851A4";
    when 16#006B1# => romdata <= X"EF3F81D5";
    when 16#006B2# => romdata <= X"C05180DF";
    when 16#006B3# => romdata <= X"DA3F7752";
    when 16#006B4# => romdata <= X"A05180DF";
    when 16#006B5# => romdata <= X"F53F8A52";
    when 16#006B6# => romdata <= X"B00851A4";
    when 16#006B7# => romdata <= X"D73F7993";
    when 16#006B8# => romdata <= X"388A5180";
    when 16#006B9# => romdata <= X"DFA73F81";
    when 16#006BA# => romdata <= X"16568F76";
    when 16#006BB# => romdata <= X"27FEA338";
    when 16#006BC# => romdata <= X"FEDE3978";
    when 16#006BD# => romdata <= X"81FF0652";
    when 16#006BE# => romdata <= X"7451FAD1";
    when 16#006BF# => romdata <= X"3F8A5180";
    when 16#006C0# => romdata <= X"DF8B3FE3";
    when 16#006C1# => romdata <= X"39F83D0D";
    when 16#006C2# => romdata <= X"02AB0533";
    when 16#006C3# => romdata <= X"59805675";
    when 16#006C4# => romdata <= X"852BE090";
    when 16#006C5# => romdata <= X"11E08012";
    when 16#006C6# => romdata <= X"0870982A";
    when 16#006C7# => romdata <= X"718C2A9F";
    when 16#006C8# => romdata <= X"FF067285";
    when 16#006C9# => romdata <= X"2A708F06";
    when 16#006CA# => romdata <= X"749F0655";
    when 16#006CB# => romdata <= X"51585B53";
    when 16#006CC# => romdata <= X"56595574";
    when 16#006CD# => romdata <= X"802E81AE";
    when 16#006CE# => romdata <= X"3875BF26";
    when 16#006CF# => romdata <= X"81B63881";
    when 16#006D0# => romdata <= X"D5C85180";
    when 16#006D1# => romdata <= X"DEE13F75";
    when 16#006D2# => romdata <= X"5180E0A5";
    when 16#006D3# => romdata <= X"3F8652B0";
    when 16#006D4# => romdata <= X"0851A3E0";
    when 16#006D5# => romdata <= X"3F81D5A0";
    when 16#006D6# => romdata <= X"5180DECB";
    when 16#006D7# => romdata <= X"3F745288";
    when 16#006D8# => romdata <= X"5180DEE6";
    when 16#006D9# => romdata <= X"3F8452B0";
    when 16#006DA# => romdata <= X"0851A3C8";
    when 16#006DB# => romdata <= X"3F81D5A8";
    when 16#006DC# => romdata <= X"5180DEB3";
    when 16#006DD# => romdata <= X"3F765290";
    when 16#006DE# => romdata <= X"5180DECE";
    when 16#006DF# => romdata <= X"3F8652B0";
    when 16#006E0# => romdata <= X"0851A3B0";
    when 16#006E1# => romdata <= X"3F81D5B0";
    when 16#006E2# => romdata <= X"5180DE9B";
    when 16#006E3# => romdata <= X"3F725180";
    when 16#006E4# => romdata <= X"DFDF3F84";
    when 16#006E5# => romdata <= X"52B00851";
    when 16#006E6# => romdata <= X"A39A3F81";
    when 16#006E7# => romdata <= X"D5B85180";
    when 16#006E8# => romdata <= X"DE853F73";
    when 16#006E9# => romdata <= X"5180DFC9";
    when 16#006EA# => romdata <= X"3F8452B0";
    when 16#006EB# => romdata <= X"0851A384";
    when 16#006EC# => romdata <= X"3F81D5C0";
    when 16#006ED# => romdata <= X"5180DDEF";
    when 16#006EE# => romdata <= X"3F7708C0";
    when 16#006EF# => romdata <= X"80800652";
    when 16#006F0# => romdata <= X"A05180DE";
    when 16#006F1# => romdata <= X"853F8A52";
    when 16#006F2# => romdata <= X"B00851A2";
    when 16#006F3# => romdata <= X"E73F7881";
    when 16#006F4# => romdata <= X"B9388A51";
    when 16#006F5# => romdata <= X"80DDB63F";
    when 16#006F6# => romdata <= X"80537481";
    when 16#006F7# => romdata <= X"2E81E638";
    when 16#006F8# => romdata <= X"76862E81";
    when 16#006F9# => romdata <= X"C2388116";
    when 16#006FA# => romdata <= X"5680FF76";
    when 16#006FB# => romdata <= X"27FEA038";
    when 16#006FC# => romdata <= X"8A3D0D04";
    when 16#006FD# => romdata <= X"81D5D051";
    when 16#006FE# => romdata <= X"80DDAC3F";
    when 16#006FF# => romdata <= X"C0165180";
    when 16#00700# => romdata <= X"DEEF3F86";
    when 16#00701# => romdata <= X"52B00851";
    when 16#00702# => romdata <= X"A2AA3F81";
    when 16#00703# => romdata <= X"D5A05180";
    when 16#00704# => romdata <= X"DD953F74";
    when 16#00705# => romdata <= X"52885180";
    when 16#00706# => romdata <= X"DDB03F84";
    when 16#00707# => romdata <= X"52B00851";
    when 16#00708# => romdata <= X"A2923F81";
    when 16#00709# => romdata <= X"D5A85180";
    when 16#0070A# => romdata <= X"DCFD3F76";
    when 16#0070B# => romdata <= X"52905180";
    when 16#0070C# => romdata <= X"DD983F86";
    when 16#0070D# => romdata <= X"52B00851";
    when 16#0070E# => romdata <= X"A1FA3F81";
    when 16#0070F# => romdata <= X"D5B05180";
    when 16#00710# => romdata <= X"DCE53F72";
    when 16#00711# => romdata <= X"5180DEA9";
    when 16#00712# => romdata <= X"3F8452B0";
    when 16#00713# => romdata <= X"0851A1E4";
    when 16#00714# => romdata <= X"3F81D5B8";
    when 16#00715# => romdata <= X"5180DCCF";
    when 16#00716# => romdata <= X"3F735180";
    when 16#00717# => romdata <= X"DE933F84";
    when 16#00718# => romdata <= X"52B00851";
    when 16#00719# => romdata <= X"A1CE3F81";
    when 16#0071A# => romdata <= X"D5C05180";
    when 16#0071B# => romdata <= X"DCB93F77";
    when 16#0071C# => romdata <= X"08C08080";
    when 16#0071D# => romdata <= X"0652A051";
    when 16#0071E# => romdata <= X"80DCCF3F";
    when 16#0071F# => romdata <= X"8A52B008";
    when 16#00720# => romdata <= X"51A1B13F";
    when 16#00721# => romdata <= X"78802EFE";
    when 16#00722# => romdata <= X"C9387681";
    when 16#00723# => romdata <= X"FF065274";
    when 16#00724# => romdata <= X"51F7BA3F";
    when 16#00725# => romdata <= X"8A5180DB";
    when 16#00726# => romdata <= X"F43F8053";
    when 16#00727# => romdata <= X"74812E09";
    when 16#00728# => romdata <= X"8106FEBC";
    when 16#00729# => romdata <= X"389F3972";
    when 16#0072A# => romdata <= X"81065776";
    when 16#0072B# => romdata <= X"802EFEB6";
    when 16#0072C# => romdata <= X"38785277";
    when 16#0072D# => romdata <= X"51FAC83F";
    when 16#0072E# => romdata <= X"81165680";
    when 16#0072F# => romdata <= X"FF7627FC";
    when 16#00730# => romdata <= X"CE38FEAC";
    when 16#00731# => romdata <= X"39745376";
    when 16#00732# => romdata <= X"862E0981";
    when 16#00733# => romdata <= X"06FE9738";
    when 16#00734# => romdata <= X"D639803D";
    when 16#00735# => romdata <= X"0D81F684";
    when 16#00736# => romdata <= X"08519971";
    when 16#00737# => romdata <= X"0C81800B";
    when 16#00738# => romdata <= X"84120C81";
    when 16#00739# => romdata <= X"F6800851";
    when 16#0073A# => romdata <= X"99710C81";
    when 16#0073B# => romdata <= X"800B8412";
    when 16#0073C# => romdata <= X"0C823D0D";
    when 16#0073D# => romdata <= X"04FE3D0D";
    when 16#0073E# => romdata <= X"74028405";
    when 16#0073F# => romdata <= X"97053302";
    when 16#00740# => romdata <= X"88059B05";
    when 16#00741# => romdata <= X"3388130C";
    when 16#00742# => romdata <= X"8C120C53";
    when 16#00743# => romdata <= X"8C130870";
    when 16#00744# => romdata <= X"812A8106";
    when 16#00745# => romdata <= X"515271F4";
    when 16#00746# => romdata <= X"388C1308";
    when 16#00747# => romdata <= X"7081FF06";
    when 16#00748# => romdata <= X"B00C5184";
    when 16#00749# => romdata <= X"3D0D0480";
    when 16#0074A# => romdata <= X"3D0D728C";
    when 16#0074B# => romdata <= X"11087087";
    when 16#0074C# => romdata <= X"2A813281";
    when 16#0074D# => romdata <= X"06B00C51";
    when 16#0074E# => romdata <= X"51823D0D";
    when 16#0074F# => romdata <= X"04FD3D0D";
    when 16#00750# => romdata <= X"02970533";
    when 16#00751# => romdata <= X"5481EC53";
    when 16#00752# => romdata <= X"81905281";
    when 16#00753# => romdata <= X"F6840851";
    when 16#00754# => romdata <= X"FFA33F73";
    when 16#00755# => romdata <= X"53905281";
    when 16#00756# => romdata <= X"F6840851";
    when 16#00757# => romdata <= X"FF973F81";
    when 16#00758# => romdata <= X"ED538190";
    when 16#00759# => romdata <= X"5281F684";
    when 16#0075A# => romdata <= X"0851FF89";
    when 16#0075B# => romdata <= X"3F805380";
    when 16#0075C# => romdata <= X"E05281F6";
    when 16#0075D# => romdata <= X"840851FE";
    when 16#0075E# => romdata <= X"FC3F81F6";
    when 16#0075F# => romdata <= X"84088811";
    when 16#00760# => romdata <= X"08B00C54";
    when 16#00761# => romdata <= X"853D0D04";
    when 16#00762# => romdata <= X"FC3D0D02";
    when 16#00763# => romdata <= X"9B053302";
    when 16#00764# => romdata <= X"84059F05";
    when 16#00765# => romdata <= X"33565481";
    when 16#00766# => romdata <= X"EC538190";
    when 16#00767# => romdata <= X"5281F684";
    when 16#00768# => romdata <= X"0851FED1";
    when 16#00769# => romdata <= X"3F735390";
    when 16#0076A# => romdata <= X"5281F684";
    when 16#0076B# => romdata <= X"0851FEC5";
    when 16#0076C# => romdata <= X"3F745380";
    when 16#0076D# => romdata <= X"D05281F6";
    when 16#0076E# => romdata <= X"840851FE";
    when 16#0076F# => romdata <= X"B83F73B0";
    when 16#00770# => romdata <= X"0C863D0D";
    when 16#00771# => romdata <= X"04FE3D0D";
    when 16#00772# => romdata <= X"FE883F81";
    when 16#00773# => romdata <= X"EC538190";
    when 16#00774# => romdata <= X"5281F684";
    when 16#00775# => romdata <= X"0851FE9D";
    when 16#00776# => romdata <= X"3F9D5390";
    when 16#00777# => romdata <= X"5281F684";
    when 16#00778# => romdata <= X"0851FE91";
    when 16#00779# => romdata <= X"3F80C553";
    when 16#0077A# => romdata <= X"80D05281";
    when 16#0077B# => romdata <= X"F6840851";
    when 16#0077C# => romdata <= X"FE833F81";
    when 16#0077D# => romdata <= X"EC538190";
    when 16#0077E# => romdata <= X"5281F684";
    when 16#0077F# => romdata <= X"0851FDF5";
    when 16#00780# => romdata <= X"3FA15390";
    when 16#00781# => romdata <= X"5281F684";
    when 16#00782# => romdata <= X"0851FDE9";
    when 16#00783# => romdata <= X"3F895380";
    when 16#00784# => romdata <= X"D05281F6";
    when 16#00785# => romdata <= X"840851FD";
    when 16#00786# => romdata <= X"DC3F81EC";
    when 16#00787# => romdata <= X"53819052";
    when 16#00788# => romdata <= X"81F68408";
    when 16#00789# => romdata <= X"51FDCE3F";
    when 16#0078A# => romdata <= X"B3539052";
    when 16#0078B# => romdata <= X"81F68408";
    when 16#0078C# => romdata <= X"51FDC23F";
    when 16#0078D# => romdata <= X"885380D0";
    when 16#0078E# => romdata <= X"5281F684";
    when 16#0078F# => romdata <= X"0851FDB5";
    when 16#00790# => romdata <= X"3F81EC53";
    when 16#00791# => romdata <= X"81905281";
    when 16#00792# => romdata <= X"F6840851";
    when 16#00793# => romdata <= X"FDA73FB4";
    when 16#00794# => romdata <= X"53905281";
    when 16#00795# => romdata <= X"F6840851";
    when 16#00796# => romdata <= X"FD9B3F96";
    when 16#00797# => romdata <= X"5380D052";
    when 16#00798# => romdata <= X"81F68408";
    when 16#00799# => romdata <= X"51FD8E3F";
    when 16#0079A# => romdata <= X"81EC5381";
    when 16#0079B# => romdata <= X"905281F6";
    when 16#0079C# => romdata <= X"840851FD";
    when 16#0079D# => romdata <= X"803FB653";
    when 16#0079E# => romdata <= X"905281F6";
    when 16#0079F# => romdata <= X"840851FC";
    when 16#007A0# => romdata <= X"F43F80E0";
    when 16#007A1# => romdata <= X"5380D052";
    when 16#007A2# => romdata <= X"81F68408";
    when 16#007A3# => romdata <= X"51FCE63F";
    when 16#007A4# => romdata <= X"81EC5381";
    when 16#007A5# => romdata <= X"905281F6";
    when 16#007A6# => romdata <= X"840851FC";
    when 16#007A7# => romdata <= X"D83F80C9";
    when 16#007A8# => romdata <= X"53905281";
    when 16#007A9# => romdata <= X"F6840851";
    when 16#007AA# => romdata <= X"FCCB3F81";
    when 16#007AB# => romdata <= X"C05380D0";
    when 16#007AC# => romdata <= X"5281F684";
    when 16#007AD# => romdata <= X"0851FCBD";
    when 16#007AE# => romdata <= X"3F843D0D";
    when 16#007AF# => romdata <= X"04FD3D0D";
    when 16#007B0# => romdata <= X"02970533";
    when 16#007B1# => romdata <= X"0284059B";
    when 16#007B2# => romdata <= X"05337181";
    when 16#007B3# => romdata <= X"B00781BF";
    when 16#007B4# => romdata <= X"06535454";
    when 16#007B5# => romdata <= X"F8808098";
    when 16#007B6# => romdata <= X"8071710C";
    when 16#007B7# => romdata <= X"73842A90";
    when 16#007B8# => romdata <= X"07710C73";
    when 16#007B9# => romdata <= X"8F06710C";
    when 16#007BA# => romdata <= X"527281F5";
    when 16#007BB# => romdata <= X"D0347381";
    when 16#007BC# => romdata <= X"F5D43485";
    when 16#007BD# => romdata <= X"3D0D04FD";
    when 16#007BE# => romdata <= X"3D0D0297";
    when 16#007BF# => romdata <= X"053381F5";
    when 16#007C0# => romdata <= X"D4335473";
    when 16#007C1# => romdata <= X"05870602";
    when 16#007C2# => romdata <= X"84059A05";
    when 16#007C3# => romdata <= X"2281F5D0";
    when 16#007C4# => romdata <= X"33547305";
    when 16#007C5# => romdata <= X"7081FF06";
    when 16#007C6# => romdata <= X"7281B007";
    when 16#007C7# => romdata <= X"54515454";
    when 16#007C8# => romdata <= X"F8808098";
    when 16#007C9# => romdata <= X"8071710C";
    when 16#007CA# => romdata <= X"73842A90";
    when 16#007CB# => romdata <= X"07710C73";
    when 16#007CC# => romdata <= X"8F06710C";
    when 16#007CD# => romdata <= X"527281F5";
    when 16#007CE# => romdata <= X"D0347381";
    when 16#007CF# => romdata <= X"F5D43485";
    when 16#007D0# => romdata <= X"3D0D04FF";
    when 16#007D1# => romdata <= X"3D0D028F";
    when 16#007D2# => romdata <= X"0533F880";
    when 16#007D3# => romdata <= X"8098840C";
    when 16#007D4# => romdata <= X"81F5D033";
    when 16#007D5# => romdata <= X"81055170";
    when 16#007D6# => romdata <= X"81F5D034";
    when 16#007D7# => romdata <= X"833D0D04";
    when 16#007D8# => romdata <= X"FF3D0D80";
    when 16#007D9# => romdata <= X"527181B0";
    when 16#007DA# => romdata <= X"0781BF06";
    when 16#007DB# => romdata <= X"F8808098";
    when 16#007DC# => romdata <= X"800C900B";
    when 16#007DD# => romdata <= X"F8808098";
    when 16#007DE# => romdata <= X"800C800B";
    when 16#007DF# => romdata <= X"F8808098";
    when 16#007E0# => romdata <= X"800C8051";
    when 16#007E1# => romdata <= X"800BF880";
    when 16#007E2# => romdata <= X"8098840C";
    when 16#007E3# => romdata <= X"81117081";
    when 16#007E4# => romdata <= X"FF065151";
    when 16#007E5# => romdata <= X"80E57127";
    when 16#007E6# => romdata <= X"EB388112";
    when 16#007E7# => romdata <= X"7081FF06";
    when 16#007E8# => romdata <= X"53518772";
    when 16#007E9# => romdata <= X"27FFBE38";
    when 16#007EA# => romdata <= X"81B00BF8";
    when 16#007EB# => romdata <= X"80809880";
    when 16#007EC# => romdata <= X"0C900BF8";
    when 16#007ED# => romdata <= X"80809880";
    when 16#007EE# => romdata <= X"0C800BF8";
    when 16#007EF# => romdata <= X"80809880";
    when 16#007F0# => romdata <= X"0C800B81";
    when 16#007F1# => romdata <= X"F5D03480";
    when 16#007F2# => romdata <= X"0B81F5D4";
    when 16#007F3# => romdata <= X"34833D0D";
    when 16#007F4# => romdata <= X"04FF3D0D";
    when 16#007F5# => romdata <= X"80C00BF8";
    when 16#007F6# => romdata <= X"80809880";
    when 16#007F7# => romdata <= X"0C81A10B";
    when 16#007F8# => romdata <= X"F8808098";
    when 16#007F9# => romdata <= X"800C81C0";
    when 16#007FA# => romdata <= X"0BF88080";
    when 16#007FB# => romdata <= X"98800C81";
    when 16#007FC# => romdata <= X"A40BF880";
    when 16#007FD# => romdata <= X"8098800C";
    when 16#007FE# => romdata <= X"81A60BF8";
    when 16#007FF# => romdata <= X"80809880";
    when 16#00800# => romdata <= X"0C81A20B";
    when 16#00801# => romdata <= X"F8808098";
    when 16#00802# => romdata <= X"800CAF0B";
    when 16#00803# => romdata <= X"F8808098";
    when 16#00804# => romdata <= X"800CA50B";
    when 16#00805# => romdata <= X"F8808098";
    when 16#00806# => romdata <= X"800C8181";
    when 16#00807# => romdata <= X"0BF88080";
    when 16#00808# => romdata <= X"98800C9D";
    when 16#00809# => romdata <= X"0BF88080";
    when 16#0080A# => romdata <= X"98800C81";
    when 16#0080B# => romdata <= X"FA0BF880";
    when 16#0080C# => romdata <= X"8098800C";
    when 16#0080D# => romdata <= X"800BF880";
    when 16#0080E# => romdata <= X"8098800C";
    when 16#0080F# => romdata <= X"80527181";
    when 16#00810# => romdata <= X"B00781BF";
    when 16#00811# => romdata <= X"06F88080";
    when 16#00812# => romdata <= X"98800C90";
    when 16#00813# => romdata <= X"0BF88080";
    when 16#00814# => romdata <= X"98800C80";
    when 16#00815# => romdata <= X"0BF88080";
    when 16#00816# => romdata <= X"98800C80";
    when 16#00817# => romdata <= X"51800BF8";
    when 16#00818# => romdata <= X"80809884";
    when 16#00819# => romdata <= X"0C811170";
    when 16#0081A# => romdata <= X"81FF0651";
    when 16#0081B# => romdata <= X"5180E571";
    when 16#0081C# => romdata <= X"27EB3881";
    when 16#0081D# => romdata <= X"127081FF";
    when 16#0081E# => romdata <= X"06535187";
    when 16#0081F# => romdata <= X"7227FFBE";
    when 16#00820# => romdata <= X"3881B00B";
    when 16#00821# => romdata <= X"F8808098";
    when 16#00822# => romdata <= X"800C900B";
    when 16#00823# => romdata <= X"F8808098";
    when 16#00824# => romdata <= X"800C800B";
    when 16#00825# => romdata <= X"F8808098";
    when 16#00826# => romdata <= X"800C800B";
    when 16#00827# => romdata <= X"81F5D034";
    when 16#00828# => romdata <= X"800B81F5";
    when 16#00829# => romdata <= X"D43481AF";
    when 16#0082A# => romdata <= X"0BF88080";
    when 16#0082B# => romdata <= X"98800C83";
    when 16#0082C# => romdata <= X"3D0D0480";
    when 16#0082D# => romdata <= X"3D0D028F";
    when 16#0082E# => romdata <= X"05337382";
    when 16#0082F# => romdata <= X"9EB40C51";
    when 16#00830# => romdata <= X"70829EB8";
    when 16#00831# => romdata <= X"34823D0D";
    when 16#00832# => romdata <= X"04EE3D0D";
    when 16#00833# => romdata <= X"64028405";
    when 16#00834# => romdata <= X"80D70533";
    when 16#00835# => romdata <= X"02880580";
    when 16#00836# => romdata <= X"DB053359";
    when 16#00837# => romdata <= X"57598076";
    when 16#00838# => romdata <= X"81067781";
    when 16#00839# => romdata <= X"2A810678";
    when 16#0083A# => romdata <= X"832B8180";
    when 16#0083B# => romdata <= X"0679822A";
    when 16#0083C# => romdata <= X"8106575E";
    when 16#0083D# => romdata <= X"415F5D81";
    when 16#0083E# => romdata <= X"FF42727D";
    when 16#0083F# => romdata <= X"2E098106";
    when 16#00840# => romdata <= X"83387C42";
    when 16#00841# => romdata <= X"768A2E83";
    when 16#00842# => romdata <= X"B9388819";
    when 16#00843# => romdata <= X"08557480";
    when 16#00844# => romdata <= X"2E83A438";
    when 16#00845# => romdata <= X"8519335A";
    when 16#00846# => romdata <= X"FF53767A";
    when 16#00847# => romdata <= X"268E3884";
    when 16#00848# => romdata <= X"19335473";
    when 16#00849# => romdata <= X"77268538";
    when 16#0084A# => romdata <= X"76743153";
    when 16#0084B# => romdata <= X"74137033";
    when 16#0084C# => romdata <= X"54587281";
    when 16#0084D# => romdata <= X"FF06831A";
    when 16#0084E# => romdata <= X"3370982B";
    when 16#0084F# => romdata <= X"81FF0A11";
    when 16#00850# => romdata <= X"9B2A8105";
    when 16#00851# => romdata <= X"5B454240";
    when 16#00852# => romdata <= X"81537483";
    when 16#00853# => romdata <= X"38745372";
    when 16#00854# => romdata <= X"81FF0643";
    when 16#00855# => romdata <= X"807A81FF";
    when 16#00856# => romdata <= X"06545CFF";
    when 16#00857# => romdata <= X"54767326";
    when 16#00858# => romdata <= X"8B388419";
    when 16#00859# => romdata <= X"33537673";
    when 16#0085A# => romdata <= X"2783F438";
    when 16#0085B# => romdata <= X"737481FF";
    when 16#0085C# => romdata <= X"06555380";
    when 16#0085D# => romdata <= X"5A797324";
    when 16#0085E# => romdata <= X"AB38747A";
    when 16#0085F# => romdata <= X"2E098106";
    when 16#00860# => romdata <= X"82E13860";
    when 16#00861# => romdata <= X"982B81FF";
    when 16#00862# => romdata <= X"0A119B2A";
    when 16#00863# => romdata <= X"821B3371";
    when 16#00864# => romdata <= X"71291170";
    when 16#00865# => romdata <= X"81FF0678";
    when 16#00866# => romdata <= X"71298C1F";
    when 16#00867# => romdata <= X"08055245";
    when 16#00868# => romdata <= X"5D575D53";
    when 16#00869# => romdata <= X"7F630570";
    when 16#0086A# => romdata <= X"81FF0670";
    when 16#0086B# => romdata <= X"612B7081";
    when 16#0086C# => romdata <= X"FF067B62";
    when 16#0086D# => romdata <= X"2B7081FF";
    when 16#0086E# => romdata <= X"067B832A";
    when 16#0086F# => romdata <= X"81065F53";
    when 16#00870# => romdata <= X"58525E42";
    when 16#00871# => romdata <= X"5578802E";
    when 16#00872# => romdata <= X"8F3881F5";
    when 16#00873# => romdata <= X"D0336105";
    when 16#00874# => romdata <= X"567580E6";
    when 16#00875# => romdata <= X"2483C538";
    when 16#00876# => romdata <= X"7F782961";
    when 16#00877# => romdata <= X"3041577C";
    when 16#00878# => romdata <= X"7E2C982B";
    when 16#00879# => romdata <= X"70982C55";
    when 16#0087A# => romdata <= X"55737725";
    when 16#0087B# => romdata <= X"818238FF";
    when 16#0087C# => romdata <= X"1C7D8106";
    when 16#0087D# => romdata <= X"5A537C73";
    when 16#0087E# => romdata <= X"2E83C438";
    when 16#0087F# => romdata <= X"7E86A638";
    when 16#00880# => romdata <= X"6184EB38";
    when 16#00881# => romdata <= X"7D802E82";
    when 16#00882# => romdata <= X"A4387914";
    when 16#00883# => romdata <= X"70337058";
    when 16#00884# => romdata <= X"54558055";
    when 16#00885# => romdata <= X"78752E85";
    when 16#00886# => romdata <= X"3872842A";
    when 16#00887# => romdata <= X"5675832A";
    when 16#00888# => romdata <= X"70810651";
    when 16#00889# => romdata <= X"5372802E";
    when 16#0088A# => romdata <= X"843881C0";
    when 16#0088B# => romdata <= X"5575822A";
    when 16#0088C# => romdata <= X"70810651";
    when 16#0088D# => romdata <= X"5372802E";
    when 16#0088E# => romdata <= X"853874B0";
    when 16#0088F# => romdata <= X"07557581";
    when 16#00890# => romdata <= X"2A708106";
    when 16#00891# => romdata <= X"51537280";
    when 16#00892# => romdata <= X"2E853874";
    when 16#00893# => romdata <= X"8C075575";
    when 16#00894# => romdata <= X"81065372";
    when 16#00895# => romdata <= X"802E8538";
    when 16#00896# => romdata <= X"74830755";
    when 16#00897# => romdata <= X"7451F9E3";
    when 16#00898# => romdata <= X"3F771498";
    when 16#00899# => romdata <= X"2B70982C";
    when 16#0089A# => romdata <= X"55567674";
    when 16#0089B# => romdata <= X"24FF9B38";
    when 16#0089C# => romdata <= X"62802E95";
    when 16#0089D# => romdata <= X"3861FF1D";
    when 16#0089E# => romdata <= X"54547C73";
    when 16#0089F# => romdata <= X"2E81FB38";
    when 16#008A0# => romdata <= X"7351F9BF";
    when 16#008A1# => romdata <= X"3F7E81EA";
    when 16#008A2# => romdata <= X"387F5281";
    when 16#008A3# => romdata <= X"51F8E83F";
    when 16#008A4# => romdata <= X"811D7081";
    when 16#008A5# => romdata <= X"FF065E54";
    when 16#008A6# => romdata <= X"7B7D26FE";
    when 16#008A7# => romdata <= X"C2386052";
    when 16#008A8# => romdata <= X"7B307098";
    when 16#008A9# => romdata <= X"2B70982C";
    when 16#008AA# => romdata <= X"53585BF8";
    when 16#008AB# => romdata <= X"CA3F6053";
    when 16#008AC# => romdata <= X"72B00C94";
    when 16#008AD# => romdata <= X"3D0D0482";
    when 16#008AE# => romdata <= X"1933851A";
    when 16#008AF# => romdata <= X"335B53FC";
    when 16#008B0# => romdata <= X"F13981F5";
    when 16#008B1# => romdata <= X"D4335372";
    when 16#008B2# => romdata <= X"8726819A";
    when 16#008B3# => romdata <= X"38811356";
    when 16#008B4# => romdata <= X"80527581";
    when 16#008B5# => romdata <= X"FF0651F7";
    when 16#008B6# => romdata <= X"E43F8053";
    when 16#008B7# => romdata <= X"72B00C94";
    when 16#008B8# => romdata <= X"3D0D0473";
    when 16#008B9# => romdata <= X"802EAF38";
    when 16#008BA# => romdata <= X"FF147081";
    when 16#008BB# => romdata <= X"FF06555A";
    when 16#008BC# => romdata <= X"7381FF2E";
    when 16#008BD# => romdata <= X"A1387470";
    when 16#008BE# => romdata <= X"81055633";
    when 16#008BF# => romdata <= X"7C057083";
    when 16#008C0# => romdata <= X"FFFF06FF";
    when 16#008C1# => romdata <= X"167081FF";
    when 16#008C2# => romdata <= X"06575C5D";
    when 16#008C3# => romdata <= X"537381FF";
    when 16#008C4# => romdata <= X"2E098106";
    when 16#008C5# => romdata <= X"E1386098";
    when 16#008C6# => romdata <= X"2B81FF0A";
    when 16#008C7# => romdata <= X"119B2A70";
    when 16#008C8# => romdata <= X"7E291E8C";
    when 16#008C9# => romdata <= X"1C08055C";
    when 16#008CA# => romdata <= X"4255FCF8";
    when 16#008CB# => romdata <= X"39791470";
    when 16#008CC# => romdata <= X"335259F8";
    when 16#008CD# => romdata <= X"8E3F7714";
    when 16#008CE# => romdata <= X"982B7098";
    when 16#008CF# => romdata <= X"2C555673";
    when 16#008D0# => romdata <= X"7725FEAC";
    when 16#008D1# => romdata <= X"38791470";
    when 16#008D2# => romdata <= X"335259F7";
    when 16#008D3# => romdata <= X"F63F7714";
    when 16#008D4# => romdata <= X"982B7098";
    when 16#008D5# => romdata <= X"2C555676";
    when 16#008D6# => romdata <= X"7424D238";
    when 16#008D7# => romdata <= X"FE923976";
    when 16#008D8# => romdata <= X"733154FC";
    when 16#008D9# => romdata <= X"87398052";
    when 16#008DA# => romdata <= X"8051F6D1";
    when 16#008DB# => romdata <= X"3F8053FE";
    when 16#008DC# => romdata <= X"EB397351";
    when 16#008DD# => romdata <= X"F7CD3FFE";
    when 16#008DE# => romdata <= X"9039617B";
    when 16#008DF# => romdata <= X"327081FF";
    when 16#008E0# => romdata <= X"0655557D";
    when 16#008E1# => romdata <= X"802EFDF8";
    when 16#008E2# => romdata <= X"387A812A";
    when 16#008E3# => romdata <= X"74327052";
    when 16#008E4# => romdata <= X"54F7B03F";
    when 16#008E5# => romdata <= X"7E802EFD";
    when 16#008E6# => romdata <= X"F038D739";
    when 16#008E7# => romdata <= X"81F5D433";
    when 16#008E8# => romdata <= X"7C055380";
    when 16#008E9# => romdata <= X"527281FF";
    when 16#008EA# => romdata <= X"0651F691";
    when 16#008EB# => romdata <= X"3F805376";
    when 16#008EC# => romdata <= X"A02EFDFC";
    when 16#008ED# => romdata <= X"387F7829";
    when 16#008EE# => romdata <= X"61304157";
    when 16#008EF# => romdata <= X"FCA1397E";
    when 16#008F0# => romdata <= X"87AD3861";
    when 16#008F1# => romdata <= X"85EB387D";
    when 16#008F2# => romdata <= X"802E80EC";
    when 16#008F3# => romdata <= X"38791470";
    when 16#008F4# => romdata <= X"337C0770";
    when 16#008F5# => romdata <= X"52545680";
    when 16#008F6# => romdata <= X"5578752E";
    when 16#008F7# => romdata <= X"85387284";
    when 16#008F8# => romdata <= X"2A567583";
    when 16#008F9# => romdata <= X"2A708106";
    when 16#008FA# => romdata <= X"51537280";
    when 16#008FB# => romdata <= X"2E843881";
    when 16#008FC# => romdata <= X"C0557582";
    when 16#008FD# => romdata <= X"2A708106";
    when 16#008FE# => romdata <= X"51537280";
    when 16#008FF# => romdata <= X"2E853874";
    when 16#00900# => romdata <= X"B0075575";
    when 16#00901# => romdata <= X"812A7081";
    when 16#00902# => romdata <= X"06515372";
    when 16#00903# => romdata <= X"802E8538";
    when 16#00904# => romdata <= X"748C0755";
    when 16#00905# => romdata <= X"75810653";
    when 16#00906# => romdata <= X"72802E85";
    when 16#00907# => romdata <= X"38748307";
    when 16#00908# => romdata <= X"557451F6";
    when 16#00909# => romdata <= X"9E3F7714";
    when 16#0090A# => romdata <= X"982B7098";
    when 16#0090B# => romdata <= X"2C555376";
    when 16#0090C# => romdata <= X"7424FF99";
    when 16#0090D# => romdata <= X"38FCB939";
    when 16#0090E# => romdata <= X"79147033";
    when 16#0090F# => romdata <= X"7C075256";
    when 16#00910# => romdata <= X"F6813F77";
    when 16#00911# => romdata <= X"14982B70";
    when 16#00912# => romdata <= X"982C5559";
    when 16#00913# => romdata <= X"737725FC";
    when 16#00914# => romdata <= X"9F387914";
    when 16#00915# => romdata <= X"70337C07";
    when 16#00916# => romdata <= X"5256F5E7";
    when 16#00917# => romdata <= X"3F771498";
    when 16#00918# => romdata <= X"2B70982C";
    when 16#00919# => romdata <= X"55597674";
    when 16#0091A# => romdata <= X"24CE38FC";
    when 16#0091B# => romdata <= X"83397D80";
    when 16#0091C# => romdata <= X"2E80F038";
    when 16#0091D# => romdata <= X"79147033";
    when 16#0091E# => romdata <= X"70585455";
    when 16#0091F# => romdata <= X"80557875";
    when 16#00920# => romdata <= X"2E853872";
    when 16#00921# => romdata <= X"842A5675";
    when 16#00922# => romdata <= X"832A7081";
    when 16#00923# => romdata <= X"06515372";
    when 16#00924# => romdata <= X"802E8438";
    when 16#00925# => romdata <= X"81C05575";
    when 16#00926# => romdata <= X"822A7081";
    when 16#00927# => romdata <= X"06515372";
    when 16#00928# => romdata <= X"802E8538";
    when 16#00929# => romdata <= X"74B00755";
    when 16#0092A# => romdata <= X"75812A70";
    when 16#0092B# => romdata <= X"81065153";
    when 16#0092C# => romdata <= X"72802E85";
    when 16#0092D# => romdata <= X"38748C07";
    when 16#0092E# => romdata <= X"55758106";
    when 16#0092F# => romdata <= X"5372802E";
    when 16#00930# => romdata <= X"85387483";
    when 16#00931# => romdata <= X"07557409";
    when 16#00932# => romdata <= X"7081FF06";
    when 16#00933# => romdata <= X"5253F4F3";
    when 16#00934# => romdata <= X"3F771498";
    when 16#00935# => romdata <= X"2B70982C";
    when 16#00936# => romdata <= X"55567674";
    when 16#00937# => romdata <= X"24FF9538";
    when 16#00938# => romdata <= X"FB8E3979";
    when 16#00939# => romdata <= X"14703370";
    when 16#0093A# => romdata <= X"097081FF";
    when 16#0093B# => romdata <= X"06545854";
    when 16#0093C# => romdata <= X"55F4D03F";
    when 16#0093D# => romdata <= X"7714982B";
    when 16#0093E# => romdata <= X"70982C55";
    when 16#0093F# => romdata <= X"59737725";
    when 16#00940# => romdata <= X"FAEE3879";
    when 16#00941# => romdata <= X"14703370";
    when 16#00942# => romdata <= X"097081FF";
    when 16#00943# => romdata <= X"06545854";
    when 16#00944# => romdata <= X"55F4B03F";
    when 16#00945# => romdata <= X"7714982B";
    when 16#00946# => romdata <= X"70982C55";
    when 16#00947# => romdata <= X"59767424";
    when 16#00948# => romdata <= X"C238FACC";
    when 16#00949# => romdata <= X"3961802E";
    when 16#0094A# => romdata <= X"81CE387D";
    when 16#0094B# => romdata <= X"802E80F7";
    when 16#0094C# => romdata <= X"38791470";
    when 16#0094D# => romdata <= X"33705854";
    when 16#0094E# => romdata <= X"55805578";
    when 16#0094F# => romdata <= X"752E8538";
    when 16#00950# => romdata <= X"72842A56";
    when 16#00951# => romdata <= X"75832A70";
    when 16#00952# => romdata <= X"81065153";
    when 16#00953# => romdata <= X"72802E84";
    when 16#00954# => romdata <= X"3881C055";
    when 16#00955# => romdata <= X"75822A70";
    when 16#00956# => romdata <= X"81065153";
    when 16#00957# => romdata <= X"72802E85";
    when 16#00958# => romdata <= X"3874B007";
    when 16#00959# => romdata <= X"5575812A";
    when 16#0095A# => romdata <= X"70810651";
    when 16#0095B# => romdata <= X"5372802E";
    when 16#0095C# => romdata <= X"8538748C";
    when 16#0095D# => romdata <= X"07557581";
    when 16#0095E# => romdata <= X"06537280";
    when 16#0095F# => romdata <= X"2E853874";
    when 16#00960# => romdata <= X"83075574";
    when 16#00961# => romdata <= X"097081FF";
    when 16#00962# => romdata <= X"06705357";
    when 16#00963# => romdata <= X"53F3B43F";
    when 16#00964# => romdata <= X"7551F3AF";
    when 16#00965# => romdata <= X"3F771498";
    when 16#00966# => romdata <= X"2B70982C";
    when 16#00967# => romdata <= X"55557674";
    when 16#00968# => romdata <= X"24FF8E38";
    when 16#00969# => romdata <= X"F9CA3979";
    when 16#0096A# => romdata <= X"14703370";
    when 16#0096B# => romdata <= X"097081FF";
    when 16#0096C# => romdata <= X"06705559";
    when 16#0096D# => romdata <= X"555659F3";
    when 16#0096E# => romdata <= X"8A3F7551";
    when 16#0096F# => romdata <= X"F3853F77";
    when 16#00970# => romdata <= X"14982B70";
    when 16#00971# => romdata <= X"982C5559";
    when 16#00972# => romdata <= X"737725F9";
    when 16#00973# => romdata <= X"A3387914";
    when 16#00974# => romdata <= X"70337009";
    when 16#00975# => romdata <= X"7081FF06";
    when 16#00976# => romdata <= X"70555955";
    when 16#00977# => romdata <= X"5659F2E3";
    when 16#00978# => romdata <= X"3F7551F2";
    when 16#00979# => romdata <= X"DE3F7714";
    when 16#0097A# => romdata <= X"982B7098";
    when 16#0097B# => romdata <= X"2C555976";
    when 16#0097C# => romdata <= X"7424FFB3";
    when 16#0097D# => romdata <= X"38F8F939";
    when 16#0097E# => romdata <= X"7D802E80";
    when 16#0097F# => romdata <= X"F4387914";
    when 16#00980# => romdata <= X"70337058";
    when 16#00981# => romdata <= X"54558055";
    when 16#00982# => romdata <= X"78752E85";
    when 16#00983# => romdata <= X"3872842A";
    when 16#00984# => romdata <= X"5675832A";
    when 16#00985# => romdata <= X"70810651";
    when 16#00986# => romdata <= X"5372802E";
    when 16#00987# => romdata <= X"843881C0";
    when 16#00988# => romdata <= X"5575822A";
    when 16#00989# => romdata <= X"70810651";
    when 16#0098A# => romdata <= X"5372802E";
    when 16#0098B# => romdata <= X"853874B0";
    when 16#0098C# => romdata <= X"07557581";
    when 16#0098D# => romdata <= X"2A708106";
    when 16#0098E# => romdata <= X"51537280";
    when 16#0098F# => romdata <= X"2E853874";
    when 16#00990# => romdata <= X"8C075575";
    when 16#00991# => romdata <= X"81065372";
    when 16#00992# => romdata <= X"802E8538";
    when 16#00993# => romdata <= X"74830755";
    when 16#00994# => romdata <= X"7481FF06";
    when 16#00995# => romdata <= X"705256F1";
    when 16#00996# => romdata <= X"EA3F7551";
    when 16#00997# => romdata <= X"F1E53F77";
    when 16#00998# => romdata <= X"14982B70";
    when 16#00999# => romdata <= X"982C5555";
    when 16#0099A# => romdata <= X"767424FF";
    when 16#0099B# => romdata <= X"9138F880";
    when 16#0099C# => romdata <= X"39791470";
    when 16#0099D# => romdata <= X"33705357";
    when 16#0099E# => romdata <= X"53F1C83F";
    when 16#0099F# => romdata <= X"7551F1C3";
    when 16#009A0# => romdata <= X"3F771498";
    when 16#009A1# => romdata <= X"2B70982C";
    when 16#009A2# => romdata <= X"55597377";
    when 16#009A3# => romdata <= X"25F7E138";
    when 16#009A4# => romdata <= X"79147033";
    when 16#009A5# => romdata <= X"70535753";
    when 16#009A6# => romdata <= X"F1A93F75";
    when 16#009A7# => romdata <= X"51F1A43F";
    when 16#009A8# => romdata <= X"7714982B";
    when 16#009A9# => romdata <= X"70982C55";
    when 16#009AA# => romdata <= X"59767424";
    when 16#009AB# => romdata <= X"C438F7C0";
    when 16#009AC# => romdata <= X"397D802E";
    when 16#009AD# => romdata <= X"80F23879";
    when 16#009AE# => romdata <= X"1470337C";
    when 16#009AF# => romdata <= X"07705254";
    when 16#009B0# => romdata <= X"56805578";
    when 16#009B1# => romdata <= X"752E8538";
    when 16#009B2# => romdata <= X"72842A56";
    when 16#009B3# => romdata <= X"75832A70";
    when 16#009B4# => romdata <= X"81065153";
    when 16#009B5# => romdata <= X"72802E84";
    when 16#009B6# => romdata <= X"3881C055";
    when 16#009B7# => romdata <= X"75822A70";
    when 16#009B8# => romdata <= X"81065153";
    when 16#009B9# => romdata <= X"72802E85";
    when 16#009BA# => romdata <= X"3874B007";
    when 16#009BB# => romdata <= X"5575812A";
    when 16#009BC# => romdata <= X"70810651";
    when 16#009BD# => romdata <= X"5372802E";
    when 16#009BE# => romdata <= X"8538748C";
    when 16#009BF# => romdata <= X"07557581";
    when 16#009C0# => romdata <= X"06537280";
    when 16#009C1# => romdata <= X"2E853874";
    when 16#009C2# => romdata <= X"83075574";
    when 16#009C3# => romdata <= X"097081FF";
    when 16#009C4# => romdata <= X"065256F0";
    when 16#009C5# => romdata <= X"AE3F7714";
    when 16#009C6# => romdata <= X"982B7098";
    when 16#009C7# => romdata <= X"2C555376";
    when 16#009C8# => romdata <= X"7424FF93";
    when 16#009C9# => romdata <= X"38F6C939";
    when 16#009CA# => romdata <= X"79147033";
    when 16#009CB# => romdata <= X"7C077009";
    when 16#009CC# => romdata <= X"7081FF06";
    when 16#009CD# => romdata <= X"54555659";
    when 16#009CE# => romdata <= X"F0893F77";
    when 16#009CF# => romdata <= X"14982B70";
    when 16#009D0# => romdata <= X"982C5559";
    when 16#009D1# => romdata <= X"737725F6";
    when 16#009D2# => romdata <= X"A7387914";
    when 16#009D3# => romdata <= X"70337C07";
    when 16#009D4# => romdata <= X"70097081";
    when 16#009D5# => romdata <= X"FF065455";
    when 16#009D6# => romdata <= X"5659EFE7";
    when 16#009D7# => romdata <= X"3F771498";
    when 16#009D8# => romdata <= X"2B70982C";
    when 16#009D9# => romdata <= X"55597674";
    when 16#009DA# => romdata <= X"24FFBD38";
    when 16#009DB# => romdata <= X"F6823961";
    when 16#009DC# => romdata <= X"802E81D4";
    when 16#009DD# => romdata <= X"387D802E";
    when 16#009DE# => romdata <= X"80F93879";
    when 16#009DF# => romdata <= X"1470337C";
    when 16#009E0# => romdata <= X"07705254";
    when 16#009E1# => romdata <= X"56805578";
    when 16#009E2# => romdata <= X"752E8538";
    when 16#009E3# => romdata <= X"72842A56";
    when 16#009E4# => romdata <= X"75832A70";
    when 16#009E5# => romdata <= X"81065153";
    when 16#009E6# => romdata <= X"72802E84";
    when 16#009E7# => romdata <= X"3881C055";
    when 16#009E8# => romdata <= X"75822A70";
    when 16#009E9# => romdata <= X"81065153";
    when 16#009EA# => romdata <= X"72802E85";
    when 16#009EB# => romdata <= X"3874B007";
    when 16#009EC# => romdata <= X"5575812A";
    when 16#009ED# => romdata <= X"70810651";
    when 16#009EE# => romdata <= X"5372802E";
    when 16#009EF# => romdata <= X"8538748C";
    when 16#009F0# => romdata <= X"07557581";
    when 16#009F1# => romdata <= X"06537280";
    when 16#009F2# => romdata <= X"2E853874";
    when 16#009F3# => romdata <= X"83075574";
    when 16#009F4# => romdata <= X"097081FF";
    when 16#009F5# => romdata <= X"06705354";
    when 16#009F6# => romdata <= X"56EEE83F";
    when 16#009F7# => romdata <= X"7251EEE3";
    when 16#009F8# => romdata <= X"3F771498";
    when 16#009F9# => romdata <= X"2B70982C";
    when 16#009FA# => romdata <= X"55567674";
    when 16#009FB# => romdata <= X"24FF8C38";
    when 16#009FC# => romdata <= X"F4FE3979";
    when 16#009FD# => romdata <= X"1470337C";
    when 16#009FE# => romdata <= X"07700970";
    when 16#009FF# => romdata <= X"81FF0670";
    when 16#00A00# => romdata <= X"55535757";
    when 16#00A01# => romdata <= X"53EEBC3F";
    when 16#00A02# => romdata <= X"7251EEB7";
    when 16#00A03# => romdata <= X"3F771498";
    when 16#00A04# => romdata <= X"2B70982C";
    when 16#00A05# => romdata <= X"55597377";
    when 16#00A06# => romdata <= X"25F4D538";
    when 16#00A07# => romdata <= X"79147033";
    when 16#00A08# => romdata <= X"7C077009";
    when 16#00A09# => romdata <= X"7081FF06";
    when 16#00A0A# => romdata <= X"70555357";
    when 16#00A0B# => romdata <= X"5753EE93";
    when 16#00A0C# => romdata <= X"3F7251EE";
    when 16#00A0D# => romdata <= X"8E3F7714";
    when 16#00A0E# => romdata <= X"982B7098";
    when 16#00A0F# => romdata <= X"2C555976";
    when 16#00A10# => romdata <= X"7424FFAF";
    when 16#00A11# => romdata <= X"38F4A939";
    when 16#00A12# => romdata <= X"7D802E80";
    when 16#00A13# => romdata <= X"F6387914";
    when 16#00A14# => romdata <= X"70337C07";
    when 16#00A15# => romdata <= X"70525456";
    when 16#00A16# => romdata <= X"80557875";
    when 16#00A17# => romdata <= X"2E853872";
    when 16#00A18# => romdata <= X"842A5675";
    when 16#00A19# => romdata <= X"832A7081";
    when 16#00A1A# => romdata <= X"06515372";
    when 16#00A1B# => romdata <= X"802E8438";
    when 16#00A1C# => romdata <= X"81C05575";
    when 16#00A1D# => romdata <= X"822A7081";
    when 16#00A1E# => romdata <= X"06515372";
    when 16#00A1F# => romdata <= X"802E8538";
    when 16#00A20# => romdata <= X"74B00755";
    when 16#00A21# => romdata <= X"75812A70";
    when 16#00A22# => romdata <= X"81065153";
    when 16#00A23# => romdata <= X"72802E85";
    when 16#00A24# => romdata <= X"38748C07";
    when 16#00A25# => romdata <= X"55758106";
    when 16#00A26# => romdata <= X"5372802E";
    when 16#00A27# => romdata <= X"85387483";
    when 16#00A28# => romdata <= X"07557481";
    when 16#00A29# => romdata <= X"FF067052";
    when 16#00A2A# => romdata <= X"56ED983F";
    when 16#00A2B# => romdata <= X"7551ED93";
    when 16#00A2C# => romdata <= X"3F771498";
    when 16#00A2D# => romdata <= X"2B70982C";
    when 16#00A2E# => romdata <= X"55537674";
    when 16#00A2F# => romdata <= X"24FF8F38";
    when 16#00A30# => romdata <= X"F3AE3979";
    when 16#00A31# => romdata <= X"1470337C";
    when 16#00A32# => romdata <= X"07705354";
    when 16#00A33# => romdata <= X"56ECF43F";
    when 16#00A34# => romdata <= X"7251ECEF";
    when 16#00A35# => romdata <= X"3F771498";
    when 16#00A36# => romdata <= X"2B70982C";
    when 16#00A37# => romdata <= X"55597377";
    when 16#00A38# => romdata <= X"25F38D38";
    when 16#00A39# => romdata <= X"79147033";
    when 16#00A3A# => romdata <= X"7C077053";
    when 16#00A3B# => romdata <= X"5456ECD3";
    when 16#00A3C# => romdata <= X"3F7251EC";
    when 16#00A3D# => romdata <= X"CE3F7714";
    when 16#00A3E# => romdata <= X"982B7098";
    when 16#00A3F# => romdata <= X"2C555976";
    when 16#00A40# => romdata <= X"7424C038";
    when 16#00A41# => romdata <= X"F2EA39F8";
    when 16#00A42# => romdata <= X"3D0D7A7D";
    when 16#00A43# => romdata <= X"028805AF";
    when 16#00A44# => romdata <= X"05335A55";
    when 16#00A45# => romdata <= X"59807470";
    when 16#00A46# => romdata <= X"81055633";
    when 16#00A47# => romdata <= X"75585657";
    when 16#00A48# => romdata <= X"74772E09";
    when 16#00A49# => romdata <= X"81068838";
    when 16#00A4A# => romdata <= X"76B00C8A";
    when 16#00A4B# => romdata <= X"3D0D0474";
    when 16#00A4C# => romdata <= X"53775278";
    when 16#00A4D# => romdata <= X"51EF923F";
    when 16#00A4E# => romdata <= X"B00881FF";
    when 16#00A4F# => romdata <= X"06770570";
    when 16#00A50# => romdata <= X"83FFFF06";
    when 16#00A51# => romdata <= X"77708105";
    when 16#00A52# => romdata <= X"59335258";
    when 16#00A53# => romdata <= X"5574802E";
    when 16#00A54# => romdata <= X"D7387453";
    when 16#00A55# => romdata <= X"77527851";
    when 16#00A56# => romdata <= X"EEEF3FB0";
    when 16#00A57# => romdata <= X"0881FF06";
    when 16#00A58# => romdata <= X"77057083";
    when 16#00A59# => romdata <= X"FFFF0677";
    when 16#00A5A# => romdata <= X"70810559";
    when 16#00A5B# => romdata <= X"33525855";
    when 16#00A5C# => romdata <= X"74FFBC38";
    when 16#00A5D# => romdata <= X"FFB239FE";
    when 16#00A5E# => romdata <= X"3D0D0293";
    when 16#00A5F# => romdata <= X"05335382";
    when 16#00A60# => romdata <= X"9EB83352";
    when 16#00A61# => romdata <= X"829EB408";
    when 16#00A62# => romdata <= X"51EEBE3F";
    when 16#00A63# => romdata <= X"B00881FF";
    when 16#00A64# => romdata <= X"06B00C84";
    when 16#00A65# => romdata <= X"3D0D04FB";
    when 16#00A66# => romdata <= X"3D0D800B";
    when 16#00A67# => romdata <= X"81DEE852";
    when 16#00A68# => romdata <= X"5680C283";
    when 16#00A69# => romdata <= X"3F755574";
    when 16#00A6A# => romdata <= X"105381D0";
    when 16#00A6B# => romdata <= X"5281F684";
    when 16#00A6C# => romdata <= X"0851E6C1";
    when 16#00A6D# => romdata <= X"3FB00887";
    when 16#00A6E# => romdata <= X"2A708106";
    when 16#00A6F# => romdata <= X"51547380";
    when 16#00A70# => romdata <= X"2E80D138";
    when 16#00A71# => romdata <= X"81157081";
    when 16#00A72# => romdata <= X"FF067098";
    when 16#00A73# => romdata <= X"2B525654";
    when 16#00A74# => romdata <= X"738025D3";
    when 16#00A75# => romdata <= X"3881DEF4";
    when 16#00A76# => romdata <= X"5180C1CB";
    when 16#00A77# => romdata <= X"3F805574";
    when 16#00A78# => romdata <= X"105381D0";
    when 16#00A79# => romdata <= X"5281F680";
    when 16#00A7A# => romdata <= X"0851E689";
    when 16#00A7B# => romdata <= X"3FB00887";
    when 16#00A7C# => romdata <= X"2A708106";
    when 16#00A7D# => romdata <= X"51547380";
    when 16#00A7E# => romdata <= X"2E80CF38";
    when 16#00A7F# => romdata <= X"81157081";
    when 16#00A80# => romdata <= X"FF067098";
    when 16#00A81# => romdata <= X"2B525654";
    when 16#00A82# => romdata <= X"738025D3";
    when 16#00A83# => romdata <= X"3875B00C";
    when 16#00A84# => romdata <= X"873D0D04";
    when 16#00A85# => romdata <= X"81DF8051";
    when 16#00A86# => romdata <= X"80C18C3F";
    when 16#00A87# => romdata <= X"74528851";
    when 16#00A88# => romdata <= X"80C1A73F";
    when 16#00A89# => romdata <= X"81DF8C51";
    when 16#00A8A# => romdata <= X"80C0FC3F";
    when 16#00A8B# => romdata <= X"81167083";
    when 16#00A8C# => romdata <= X"FFFF0681";
    when 16#00A8D# => romdata <= X"177081FF";
    when 16#00A8E# => romdata <= X"0670982B";
    when 16#00A8F# => romdata <= X"52585257";
    when 16#00A90# => romdata <= X"54738025";
    when 16#00A91# => romdata <= X"FEE138FF";
    when 16#00A92# => romdata <= X"8C3981DF";
    when 16#00A93# => romdata <= X"805180C0";
    when 16#00A94# => romdata <= X"D63F7452";
    when 16#00A95# => romdata <= X"885180C0";
    when 16#00A96# => romdata <= X"F13F81DF";
    when 16#00A97# => romdata <= X"8C5180C0";
    when 16#00A98# => romdata <= X"C63F8116";
    when 16#00A99# => romdata <= X"7083FFFF";
    when 16#00A9A# => romdata <= X"06811770";
    when 16#00A9B# => romdata <= X"81FF0670";
    when 16#00A9C# => romdata <= X"982B5258";
    when 16#00A9D# => romdata <= X"52575473";
    when 16#00A9E# => romdata <= X"8025FEE3";
    when 16#00A9F# => romdata <= X"38FF8E39";
    when 16#00AA0# => romdata <= X"F33D0D7F";
    when 16#00AA1# => romdata <= X"02840580";
    when 16#00AA2# => romdata <= X"C3053302";
    when 16#00AA3# => romdata <= X"880580C6";
    when 16#00AA4# => romdata <= X"052281DF";
    when 16#00AA5# => romdata <= X"9C545B55";
    when 16#00AA6# => romdata <= X"5880C08B";
    when 16#00AA7# => romdata <= X"3F785180";
    when 16#00AA8# => romdata <= X"C1CF3F81";
    when 16#00AA9# => romdata <= X"DFA851BF";
    when 16#00AAA# => romdata <= X"FE3F7352";
    when 16#00AAB# => romdata <= X"885180C0";
    when 16#00AAC# => romdata <= X"993F81CE";
    when 16#00AAD# => romdata <= X"C851BFEF";
    when 16#00AAE# => romdata <= X"3F805776";
    when 16#00AAF# => romdata <= X"79278191";
    when 16#00AB0# => romdata <= X"3873108E";
    when 16#00AB1# => romdata <= X"3D5C5A79";
    when 16#00AB2# => romdata <= X"53819052";
    when 16#00AB3# => romdata <= X"7751E4A5";
    when 16#00AB4# => romdata <= X"3F76882A";
    when 16#00AB5# => romdata <= X"53905277";
    when 16#00AB6# => romdata <= X"51E49A3F";
    when 16#00AB7# => romdata <= X"7681FF06";
    when 16#00AB8# => romdata <= X"53905277";
    when 16#00AB9# => romdata <= X"51E48E3F";
    when 16#00ABA# => romdata <= X"811A5381";
    when 16#00ABB# => romdata <= X"90527751";
    when 16#00ABC# => romdata <= X"E4833F80";
    when 16#00ABD# => romdata <= X"5380E052";
    when 16#00ABE# => romdata <= X"7751E3F9";
    when 16#00ABF# => romdata <= X"3FB00887";
    when 16#00AC0# => romdata <= X"2A810654";
    when 16#00AC1# => romdata <= X"738A3888";
    when 16#00AC2# => romdata <= X"18087081";
    when 16#00AC3# => romdata <= X"FF065D56";
    when 16#00AC4# => romdata <= X"7B81FF06";
    when 16#00AC5# => romdata <= X"81D5AC52";
    when 16#00AC6# => romdata <= X"56BF8C3F";
    when 16#00AC7# => romdata <= X"75528851";
    when 16#00AC8# => romdata <= X"BFA83F81";
    when 16#00AC9# => romdata <= X"E9E051BE";
    when 16#00ACA# => romdata <= X"FE3FE016";
    when 16#00ACB# => romdata <= X"5480DF74";
    when 16#00ACC# => romdata <= X"27B63876";
    when 16#00ACD# => romdata <= X"8706701C";
    when 16#00ACE# => romdata <= X"5755A076";
    when 16#00ACF# => romdata <= X"3474872E";
    when 16#00AD0# => romdata <= X"B9388117";
    when 16#00AD1# => romdata <= X"7083FFFF";
    when 16#00AD2# => romdata <= X"06585578";
    when 16#00AD3# => romdata <= X"7726FEF7";
    when 16#00AD4# => romdata <= X"3880E00B";
    when 16#00AD5# => romdata <= X"8C190C8C";
    when 16#00AD6# => romdata <= X"18087081";
    when 16#00AD7# => romdata <= X"2A810658";
    when 16#00AD8# => romdata <= X"5A76F438";
    when 16#00AD9# => romdata <= X"8F3D0D04";
    when 16#00ADA# => romdata <= X"76870670";
    when 16#00ADB# => romdata <= X"1C555575";
    when 16#00ADC# => romdata <= X"74347487";
    when 16#00ADD# => romdata <= X"2E098106";
    when 16#00ADE# => romdata <= X"C9387A51";
    when 16#00ADF# => romdata <= X"BEA93F8A";
    when 16#00AE0# => romdata <= X"51BE8A3F";
    when 16#00AE1# => romdata <= X"81177083";
    when 16#00AE2# => romdata <= X"FFFF0658";
    when 16#00AE3# => romdata <= X"55787726";
    when 16#00AE4# => romdata <= X"FEB538FF";
    when 16#00AE5# => romdata <= X"BC39FB3D";
    when 16#00AE6# => romdata <= X"0D8151CC";
    when 16#00AE7# => romdata <= X"AA3FB008";
    when 16#00AE8# => romdata <= X"81FF0654";
    when 16#00AE9# => romdata <= X"8251CDD2";
    when 16#00AEA# => romdata <= X"3FB00881";
    when 16#00AEB# => romdata <= X"FF065683";
    when 16#00AEC# => romdata <= X"51CC943F";
    when 16#00AED# => romdata <= X"B00883FF";
    when 16#00AEE# => romdata <= X"FF065573";
    when 16#00AEF# => romdata <= X"9C3881F6";
    when 16#00AF0# => romdata <= X"80085474";
    when 16#00AF1# => romdata <= X"84388180";
    when 16#00AF2# => romdata <= X"55745375";
    when 16#00AF3# => romdata <= X"527351FD";
    when 16#00AF4# => romdata <= X"AF3F74B0";
    when 16#00AF5# => romdata <= X"0C873D0D";
    when 16#00AF6# => romdata <= X"0481F684";
    when 16#00AF7# => romdata <= X"0854E439";
    when 16#00AF8# => romdata <= X"FB3D0D77";
    when 16#00AF9# => romdata <= X"028405A7";
    when 16#00AFA# => romdata <= X"05330288";
    when 16#00AFB# => romdata <= X"05A30533";
    when 16#00AFC# => romdata <= X"70105658";
    when 16#00AFD# => romdata <= X"56548190";
    when 16#00AFE# => romdata <= X"527351E1";
    when 16#00AFF# => romdata <= X"F83F7351";
    when 16#00B00# => romdata <= X"E2A53FB0";
    when 16#00B01# => romdata <= X"08802E93";
    when 16#00B02# => romdata <= X"38745380";
    when 16#00B03# => romdata <= X"D0527351";
    when 16#00B04# => romdata <= X"E1E33F80";
    when 16#00B05# => romdata <= X"0BB00C87";
    when 16#00B06# => romdata <= X"3D0D0481";
    when 16#00B07# => romdata <= X"DFC451BD";
    when 16#00B08# => romdata <= X"863FFF0B";
    when 16#00B09# => romdata <= X"B00C873D";
    when 16#00B0A# => romdata <= X"0D04FC3D";
    when 16#00B0B# => romdata <= X"0D760284";
    when 16#00B0C# => romdata <= X"059F0533";
    when 16#00B0D# => romdata <= X"70108105";
    when 16#00B0E# => romdata <= X"55565481";
    when 16#00B0F# => romdata <= X"90527351";
    when 16#00B10# => romdata <= X"E1B33F73";
    when 16#00B11# => romdata <= X"51E1E03F";
    when 16#00B12# => romdata <= X"B008802E";
    when 16#00B13# => romdata <= X"A7388053";
    when 16#00B14# => romdata <= X"80E05273";
    when 16#00B15# => romdata <= X"51E19E3F";
    when 16#00B16# => romdata <= X"7351E1CB";
    when 16#00B17# => romdata <= X"3FB00880";
    when 16#00B18# => romdata <= X"2E923888";
    when 16#00B19# => romdata <= X"14087090";
    when 16#00B1A# => romdata <= X"2B70902C";
    when 16#00B1B# => romdata <= X"B00C5555";
    when 16#00B1C# => romdata <= X"863D0D04";
    when 16#00B1D# => romdata <= X"81DFC451";
    when 16#00B1E# => romdata <= X"BCAD3FFF";
    when 16#00B1F# => romdata <= X"0BB00C86";
    when 16#00B20# => romdata <= X"3D0D04FD";
    when 16#00B21# => romdata <= X"3D0D9C54";
    when 16#00B22# => romdata <= X"81DFCC51";
    when 16#00B23# => romdata <= X"BC993F73";
    when 16#00B24# => romdata <= X"528851BC";
    when 16#00B25# => romdata <= X"B53F7351";
    when 16#00B26# => romdata <= X"E1A33FB0";
    when 16#00B27# => romdata <= X"0881FF06";
    when 16#00B28# => romdata <= X"81F68408";
    when 16#00B29# => romdata <= X"5253E0FF";
    when 16#00B2A# => romdata <= X"3FB00880";
    when 16#00B2B# => romdata <= X"2EAA3881";
    when 16#00B2C# => romdata <= X"DFDC51BB";
    when 16#00B2D# => romdata <= X"F23F7252";
    when 16#00B2E# => romdata <= X"8851BC8E";
    when 16#00B2F# => romdata <= X"3F8A51BB";
    when 16#00B30# => romdata <= X"CC3F8114";
    when 16#00B31# => romdata <= X"7081FF06";
    when 16#00B32# => romdata <= X"555380D5";
    when 16#00B33# => romdata <= X"7427FFB8";
    when 16#00B34# => romdata <= X"3872B00C";
    when 16#00B35# => romdata <= X"853D0D04";
    when 16#00B36# => romdata <= X"81DFE451";
    when 16#00B37# => romdata <= X"BBC93FFF";
    when 16#00B38# => romdata <= X"0BB00C85";
    when 16#00B39# => romdata <= X"3D0D04FE";
    when 16#00B3A# => romdata <= X"3D0D8151";
    when 16#00B3B# => romdata <= X"CB8C3FB0";
    when 16#00B3C# => romdata <= X"0881FF06";
    when 16#00B3D# => romdata <= X"538251CB";
    when 16#00B3E# => romdata <= X"813FB008";
    when 16#00B3F# => romdata <= X"81FF0652";
    when 16#00B40# => romdata <= X"7251E184";
    when 16#00B41# => romdata <= X"3F7251E0";
    when 16#00B42# => romdata <= X"B43FB008";
    when 16#00B43# => romdata <= X"81FF0681";
    when 16#00B44# => romdata <= X"F6840852";
    when 16#00B45# => romdata <= X"53E0903F";
    when 16#00B46# => romdata <= X"B008802E";
    when 16#00B47# => romdata <= X"883872B0";
    when 16#00B48# => romdata <= X"0C843D0D";
    when 16#00B49# => romdata <= X"0481DFEC";
    when 16#00B4A# => romdata <= X"51BAFC3F";
    when 16#00B4B# => romdata <= X"FF0BB00C";
    when 16#00B4C# => romdata <= X"843D0D04";
    when 16#00B4D# => romdata <= X"FE3D0D02";
    when 16#00B4E# => romdata <= X"93053302";
    when 16#00B4F# => romdata <= X"84059705";
    when 16#00B50# => romdata <= X"33545271";
    when 16#00B51# => romdata <= X"73279338";
    when 16#00B52# => romdata <= X"A051BAC1";
    when 16#00B53# => romdata <= X"3F811270";
    when 16#00B54# => romdata <= X"81FF0651";
    when 16#00B55# => romdata <= X"52727226";
    when 16#00B56# => romdata <= X"EF38843D";
    when 16#00B57# => romdata <= X"0D04FE3D";
    when 16#00B58# => romdata <= X"0D747081";
    when 16#00B59# => romdata <= X"06535371";
    when 16#00B5A# => romdata <= X"85DF3872";
    when 16#00B5B# => romdata <= X"812A7081";
    when 16#00B5C# => romdata <= X"06515271";
    when 16#00B5D# => romdata <= X"85BC3872";
    when 16#00B5E# => romdata <= X"822A7081";
    when 16#00B5F# => romdata <= X"06515271";
    when 16#00B60# => romdata <= X"85993872";
    when 16#00B61# => romdata <= X"832A7081";
    when 16#00B62# => romdata <= X"06515271";
    when 16#00B63# => romdata <= X"84F63872";
    when 16#00B64# => romdata <= X"842A7081";
    when 16#00B65# => romdata <= X"06515271";
    when 16#00B66# => romdata <= X"84D33872";
    when 16#00B67# => romdata <= X"852A7081";
    when 16#00B68# => romdata <= X"06515271";
    when 16#00B69# => romdata <= X"84B03872";
    when 16#00B6A# => romdata <= X"862A7081";
    when 16#00B6B# => romdata <= X"06515271";
    when 16#00B6C# => romdata <= X"848D3872";
    when 16#00B6D# => romdata <= X"872A7081";
    when 16#00B6E# => romdata <= X"06515271";
    when 16#00B6F# => romdata <= X"83EA3872";
    when 16#00B70# => romdata <= X"882A7081";
    when 16#00B71# => romdata <= X"06515271";
    when 16#00B72# => romdata <= X"83C73872";
    when 16#00B73# => romdata <= X"892A7081";
    when 16#00B74# => romdata <= X"06515271";
    when 16#00B75# => romdata <= X"83A43872";
    when 16#00B76# => romdata <= X"8A2A7081";
    when 16#00B77# => romdata <= X"06515271";
    when 16#00B78# => romdata <= X"83813872";
    when 16#00B79# => romdata <= X"8B2A7081";
    when 16#00B7A# => romdata <= X"06515271";
    when 16#00B7B# => romdata <= X"82DE3872";
    when 16#00B7C# => romdata <= X"8C2A7081";
    when 16#00B7D# => romdata <= X"06515271";
    when 16#00B7E# => romdata <= X"82BB3872";
    when 16#00B7F# => romdata <= X"8D2A7081";
    when 16#00B80# => romdata <= X"06515271";
    when 16#00B81# => romdata <= X"82983872";
    when 16#00B82# => romdata <= X"8E2A7081";
    when 16#00B83# => romdata <= X"06515271";
    when 16#00B84# => romdata <= X"81F53872";
    when 16#00B85# => romdata <= X"8F2A7081";
    when 16#00B86# => romdata <= X"06515271";
    when 16#00B87# => romdata <= X"81D23872";
    when 16#00B88# => romdata <= X"902A7081";
    when 16#00B89# => romdata <= X"06515271";
    when 16#00B8A# => romdata <= X"81AF3872";
    when 16#00B8B# => romdata <= X"912A7081";
    when 16#00B8C# => romdata <= X"06515271";
    when 16#00B8D# => romdata <= X"818C3872";
    when 16#00B8E# => romdata <= X"922A7081";
    when 16#00B8F# => romdata <= X"06515271";
    when 16#00B90# => romdata <= X"80E93872";
    when 16#00B91# => romdata <= X"932A7081";
    when 16#00B92# => romdata <= X"06515271";
    when 16#00B93# => romdata <= X"80C63872";
    when 16#00B94# => romdata <= X"942A7081";
    when 16#00B95# => romdata <= X"06515271";
    when 16#00B96# => romdata <= X"A5387295";
    when 16#00B97# => romdata <= X"2A708106";
    when 16#00B98# => romdata <= X"5152718B";
    when 16#00B99# => romdata <= X"38807324";
    when 16#00B9A# => romdata <= X"83F63884";
    when 16#00B9B# => romdata <= X"3D0D0481";
    when 16#00B9C# => romdata <= X"DFFC51B8";
    when 16#00B9D# => romdata <= X"B23F7280";
    when 16#00B9E# => romdata <= X"25F13883";
    when 16#00B9F# => romdata <= X"E33981E0";
    when 16#00BA0# => romdata <= X"9851B8A3";
    when 16#00BA1# => romdata <= X"3F72952A";
    when 16#00BA2# => romdata <= X"70810651";
    when 16#00BA3# => romdata <= X"5271802E";
    when 16#00BA4# => romdata <= X"D438DC39";
    when 16#00BA5# => romdata <= X"81E0B451";
    when 16#00BA6# => romdata <= X"B88D3F72";
    when 16#00BA7# => romdata <= X"942A7081";
    when 16#00BA8# => romdata <= X"06515271";
    when 16#00BA9# => romdata <= X"802EFFB2";
    when 16#00BAA# => romdata <= X"38D43981";
    when 16#00BAB# => romdata <= X"E0D051B7";
    when 16#00BAC# => romdata <= X"F63F7293";
    when 16#00BAD# => romdata <= X"2A708106";
    when 16#00BAE# => romdata <= X"51527180";
    when 16#00BAF# => romdata <= X"2EFF9038";
    when 16#00BB0# => romdata <= X"D33981E0";
    when 16#00BB1# => romdata <= X"EC51B7DF";
    when 16#00BB2# => romdata <= X"3F72922A";
    when 16#00BB3# => romdata <= X"70810651";
    when 16#00BB4# => romdata <= X"5271802E";
    when 16#00BB5# => romdata <= X"FEED38D3";
    when 16#00BB6# => romdata <= X"3981E18C";
    when 16#00BB7# => romdata <= X"51B7C83F";
    when 16#00BB8# => romdata <= X"72912A70";
    when 16#00BB9# => romdata <= X"81065152";
    when 16#00BBA# => romdata <= X"71802EFE";
    when 16#00BBB# => romdata <= X"CA38D339";
    when 16#00BBC# => romdata <= X"81E1AC51";
    when 16#00BBD# => romdata <= X"B7B13F72";
    when 16#00BBE# => romdata <= X"902A7081";
    when 16#00BBF# => romdata <= X"06515271";
    when 16#00BC0# => romdata <= X"802EFEA7";
    when 16#00BC1# => romdata <= X"38D33981";
    when 16#00BC2# => romdata <= X"E1CC51B7";
    when 16#00BC3# => romdata <= X"9A3F728F";
    when 16#00BC4# => romdata <= X"2A708106";
    when 16#00BC5# => romdata <= X"51527180";
    when 16#00BC6# => romdata <= X"2EFE8438";
    when 16#00BC7# => romdata <= X"D33981E1";
    when 16#00BC8# => romdata <= X"EC51B783";
    when 16#00BC9# => romdata <= X"3F728E2A";
    when 16#00BCA# => romdata <= X"70810651";
    when 16#00BCB# => romdata <= X"5271802E";
    when 16#00BCC# => romdata <= X"FDE138D3";
    when 16#00BCD# => romdata <= X"3981E284";
    when 16#00BCE# => romdata <= X"51B6EC3F";
    when 16#00BCF# => romdata <= X"728D2A70";
    when 16#00BD0# => romdata <= X"81065152";
    when 16#00BD1# => romdata <= X"71802EFD";
    when 16#00BD2# => romdata <= X"BE38D339";
    when 16#00BD3# => romdata <= X"81E29851";
    when 16#00BD4# => romdata <= X"B6D53F72";
    when 16#00BD5# => romdata <= X"8C2A7081";
    when 16#00BD6# => romdata <= X"06515271";
    when 16#00BD7# => romdata <= X"802EFD9B";
    when 16#00BD8# => romdata <= X"38D33981";
    when 16#00BD9# => romdata <= X"E2B851B6";
    when 16#00BDA# => romdata <= X"BE3F728B";
    when 16#00BDB# => romdata <= X"2A708106";
    when 16#00BDC# => romdata <= X"51527180";
    when 16#00BDD# => romdata <= X"2EFCF838";
    when 16#00BDE# => romdata <= X"D33981E2";
    when 16#00BDF# => romdata <= X"E051B6A7";
    when 16#00BE0# => romdata <= X"3F728A2A";
    when 16#00BE1# => romdata <= X"70810651";
    when 16#00BE2# => romdata <= X"5271802E";
    when 16#00BE3# => romdata <= X"FCD538D3";
    when 16#00BE4# => romdata <= X"3981E380";
    when 16#00BE5# => romdata <= X"51B6903F";
    when 16#00BE6# => romdata <= X"72892A70";
    when 16#00BE7# => romdata <= X"81065152";
    when 16#00BE8# => romdata <= X"71802EFC";
    when 16#00BE9# => romdata <= X"B238D339";
    when 16#00BEA# => romdata <= X"81E3A051";
    when 16#00BEB# => romdata <= X"B5F93F72";
    when 16#00BEC# => romdata <= X"882A7081";
    when 16#00BED# => romdata <= X"06515271";
    when 16#00BEE# => romdata <= X"802EFC8F";
    when 16#00BEF# => romdata <= X"38D33981";
    when 16#00BF0# => romdata <= X"E3C851B5";
    when 16#00BF1# => romdata <= X"E23F7287";
    when 16#00BF2# => romdata <= X"2A708106";
    when 16#00BF3# => romdata <= X"51527180";
    when 16#00BF4# => romdata <= X"2EFBEC38";
    when 16#00BF5# => romdata <= X"D33981E3";
    when 16#00BF6# => romdata <= X"E851B5CB";
    when 16#00BF7# => romdata <= X"3F72862A";
    when 16#00BF8# => romdata <= X"70810651";
    when 16#00BF9# => romdata <= X"5271802E";
    when 16#00BFA# => romdata <= X"FBC938D3";
    when 16#00BFB# => romdata <= X"3981E488";
    when 16#00BFC# => romdata <= X"51B5B43F";
    when 16#00BFD# => romdata <= X"72852A70";
    when 16#00BFE# => romdata <= X"81065152";
    when 16#00BFF# => romdata <= X"71802EFB";
    when 16#00C00# => romdata <= X"A638D339";
    when 16#00C01# => romdata <= X"81E4B051";
    when 16#00C02# => romdata <= X"B59D3F72";
    when 16#00C03# => romdata <= X"842A7081";
    when 16#00C04# => romdata <= X"06515271";
    when 16#00C05# => romdata <= X"802EFB83";
    when 16#00C06# => romdata <= X"38D33981";
    when 16#00C07# => romdata <= X"E4D051B5";
    when 16#00C08# => romdata <= X"863F7283";
    when 16#00C09# => romdata <= X"2A708106";
    when 16#00C0A# => romdata <= X"51527180";
    when 16#00C0B# => romdata <= X"2EFAE038";
    when 16#00C0C# => romdata <= X"D33981E4";
    when 16#00C0D# => romdata <= X"F051B4EF";
    when 16#00C0E# => romdata <= X"3F72822A";
    when 16#00C0F# => romdata <= X"70810651";
    when 16#00C10# => romdata <= X"5271802E";
    when 16#00C11# => romdata <= X"FABD38D3";
    when 16#00C12# => romdata <= X"3981E598";
    when 16#00C13# => romdata <= X"51B4D83F";
    when 16#00C14# => romdata <= X"72812A70";
    when 16#00C15# => romdata <= X"81065152";
    when 16#00C16# => romdata <= X"71802EFA";
    when 16#00C17# => romdata <= X"9A38D339";
    when 16#00C18# => romdata <= X"81E5B851";
    when 16#00C19# => romdata <= X"B4C13F84";
    when 16#00C1A# => romdata <= X"3D0D04FD";
    when 16#00C1B# => romdata <= X"3D0D81E5";
    when 16#00C1C# => romdata <= X"CC51B4B3";
    when 16#00C1D# => romdata <= X"3FFFAF9B";
    when 16#00C1E# => romdata <= X"3FB00880";
    when 16#00C1F# => romdata <= X"2E889A38";
    when 16#00C20# => romdata <= X"81E5E851";
    when 16#00C21# => romdata <= X"B4A13F81";
    when 16#00C22# => romdata <= X"E5F051B4";
    when 16#00C23# => romdata <= X"9A3F81F6";
    when 16#00C24# => romdata <= X"8C088411";
    when 16#00C25# => romdata <= X"08709D2A";
    when 16#00C26# => romdata <= X"81065154";
    when 16#00C27# => romdata <= X"5472802E";
    when 16#00C28# => romdata <= X"87933881";
    when 16#00C29# => romdata <= X"CEA451B3";
    when 16#00C2A# => romdata <= X"FE3F81E6";
    when 16#00C2B# => romdata <= X"8C51B3F7";
    when 16#00C2C# => romdata <= X"3F81F5CC";
    when 16#00C2D# => romdata <= X"0880D411";
    when 16#00C2E# => romdata <= X"085253B5";
    when 16#00C2F# => romdata <= X"B43F81E6";
    when 16#00C30# => romdata <= X"A851B3E3";
    when 16#00C31# => romdata <= X"3F81F5CC";
    when 16#00C32# => romdata <= X"0880D011";
    when 16#00C33# => romdata <= X"085254B5";
    when 16#00C34# => romdata <= X"A03F8A51";
    when 16#00C35# => romdata <= X"B3B73F81";
    when 16#00C36# => romdata <= X"E6C451B3";
    when 16#00C37# => romdata <= X"CA3F81E6";
    when 16#00C38# => romdata <= X"E851B3C3";
    when 16#00C39# => romdata <= X"3F81E7B0";
    when 16#00C3A# => romdata <= X"51B3BC3F";
    when 16#00C3B# => romdata <= X"81E7F851";
    when 16#00C3C# => romdata <= X"B3B53F81";
    when 16#00C3D# => romdata <= X"F5CC0870";
    when 16#00C3E# => romdata <= X"085253B4";
    when 16#00C3F# => romdata <= X"F43FB008";
    when 16#00C40# => romdata <= X"81FF0653";
    when 16#00C41# => romdata <= X"728C2793";
    when 16#00C42# => romdata <= X"38A051B3";
    when 16#00C43# => romdata <= X"803F8113";
    when 16#00C44# => romdata <= X"7081FF06";
    when 16#00C45# => romdata <= X"54548C73";
    when 16#00C46# => romdata <= X"26EF3881";
    when 16#00C47# => romdata <= X"F5CC0884";
    when 16#00C48# => romdata <= X"11085253";
    when 16#00C49# => romdata <= X"B4CB3FB0";
    when 16#00C4A# => romdata <= X"0881FF06";
    when 16#00C4B# => romdata <= X"53728C27";
    when 16#00C4C# => romdata <= X"9338A051";
    when 16#00C4D# => romdata <= X"B2D73F81";
    when 16#00C4E# => romdata <= X"137081FF";
    when 16#00C4F# => romdata <= X"0654548C";
    when 16#00C50# => romdata <= X"7326EF38";
    when 16#00C51# => romdata <= X"81F5CC08";
    when 16#00C52# => romdata <= X"88110852";
    when 16#00C53# => romdata <= X"53B4A23F";
    when 16#00C54# => romdata <= X"B00881FF";
    when 16#00C55# => romdata <= X"0653728C";
    when 16#00C56# => romdata <= X"279338A0";
    when 16#00C57# => romdata <= X"51B2AE3F";
    when 16#00C58# => romdata <= X"81137081";
    when 16#00C59# => romdata <= X"FF065454";
    when 16#00C5A# => romdata <= X"8C7326EF";
    when 16#00C5B# => romdata <= X"3881F5CC";
    when 16#00C5C# => romdata <= X"088C1108";
    when 16#00C5D# => romdata <= X"5253B3F9";
    when 16#00C5E# => romdata <= X"3FB00881";
    when 16#00C5F# => romdata <= X"FF065372";
    when 16#00C60# => romdata <= X"8C279338";
    when 16#00C61# => romdata <= X"A051B285";
    when 16#00C62# => romdata <= X"3F811370";
    when 16#00C63# => romdata <= X"81FF0654";
    when 16#00C64# => romdata <= X"548C7326";
    when 16#00C65# => romdata <= X"EF3881E8";
    when 16#00C66# => romdata <= X"9451B28B";
    when 16#00C67# => romdata <= X"3F81F5CC";
    when 16#00C68# => romdata <= X"08901108";
    when 16#00C69# => romdata <= X"5253B3C9";
    when 16#00C6A# => romdata <= X"3FB00881";
    when 16#00C6B# => romdata <= X"FF065372";
    when 16#00C6C# => romdata <= X"8C279338";
    when 16#00C6D# => romdata <= X"A051B1D5";
    when 16#00C6E# => romdata <= X"3F811370";
    when 16#00C6F# => romdata <= X"81FF0654";
    when 16#00C70# => romdata <= X"548C7326";
    when 16#00C71# => romdata <= X"EF3881F5";
    when 16#00C72# => romdata <= X"CC089411";
    when 16#00C73# => romdata <= X"085253B3";
    when 16#00C74# => romdata <= X"A03FB008";
    when 16#00C75# => romdata <= X"81FF0653";
    when 16#00C76# => romdata <= X"728C2793";
    when 16#00C77# => romdata <= X"38A051B1";
    when 16#00C78# => romdata <= X"AC3F8113";
    when 16#00C79# => romdata <= X"7081FF06";
    when 16#00C7A# => romdata <= X"54548C73";
    when 16#00C7B# => romdata <= X"26EF3881";
    when 16#00C7C# => romdata <= X"F5CC0898";
    when 16#00C7D# => romdata <= X"11085253";
    when 16#00C7E# => romdata <= X"B2F73FB0";
    when 16#00C7F# => romdata <= X"0881FF06";
    when 16#00C80# => romdata <= X"53728C27";
    when 16#00C81# => romdata <= X"9338A051";
    when 16#00C82# => romdata <= X"B1833F81";
    when 16#00C83# => romdata <= X"137081FF";
    when 16#00C84# => romdata <= X"0654548C";
    when 16#00C85# => romdata <= X"7326EF38";
    when 16#00C86# => romdata <= X"81F5CC08";
    when 16#00C87# => romdata <= X"9C110852";
    when 16#00C88# => romdata <= X"53B2CE3F";
    when 16#00C89# => romdata <= X"B00881FF";
    when 16#00C8A# => romdata <= X"0653728C";
    when 16#00C8B# => romdata <= X"279338A0";
    when 16#00C8C# => romdata <= X"51B0DA3F";
    when 16#00C8D# => romdata <= X"81137081";
    when 16#00C8E# => romdata <= X"FF065454";
    when 16#00C8F# => romdata <= X"8C7326EF";
    when 16#00C90# => romdata <= X"3881E8B0";
    when 16#00C91# => romdata <= X"51B0E03F";
    when 16#00C92# => romdata <= X"81F5CC08";
    when 16#00C93# => romdata <= X"54810BB0";
    when 16#00C94# => romdata <= X"150CB014";
    when 16#00C95# => romdata <= X"08537280";
    when 16#00C96# => romdata <= X"25F838A0";
    when 16#00C97# => romdata <= X"140851B2";
    when 16#00C98# => romdata <= X"903FB008";
    when 16#00C99# => romdata <= X"81FF0653";
    when 16#00C9A# => romdata <= X"728C2793";
    when 16#00C9B# => romdata <= X"38A051B0";
    when 16#00C9C# => romdata <= X"9C3F8113";
    when 16#00C9D# => romdata <= X"7081FF06";
    when 16#00C9E# => romdata <= X"54548C73";
    when 16#00C9F# => romdata <= X"26EF3881";
    when 16#00CA0# => romdata <= X"F5CC08A4";
    when 16#00CA1# => romdata <= X"11085253";
    when 16#00CA2# => romdata <= X"B1E73FB0";
    when 16#00CA3# => romdata <= X"0881FF06";
    when 16#00CA4# => romdata <= X"53728C27";
    when 16#00CA5# => romdata <= X"9338A051";
    when 16#00CA6# => romdata <= X"AFF33F81";
    when 16#00CA7# => romdata <= X"137081FF";
    when 16#00CA8# => romdata <= X"0654548C";
    when 16#00CA9# => romdata <= X"7326EF38";
    when 16#00CAA# => romdata <= X"81F5CC08";
    when 16#00CAB# => romdata <= X"A8110852";
    when 16#00CAC# => romdata <= X"53B1BE3F";
    when 16#00CAD# => romdata <= X"B00881FF";
    when 16#00CAE# => romdata <= X"0653728C";
    when 16#00CAF# => romdata <= X"279338A0";
    when 16#00CB0# => romdata <= X"51AFCA3F";
    when 16#00CB1# => romdata <= X"81137081";
    when 16#00CB2# => romdata <= X"FF065454";
    when 16#00CB3# => romdata <= X"8C7326EF";
    when 16#00CB4# => romdata <= X"3881F5CC";
    when 16#00CB5# => romdata <= X"08AC1108";
    when 16#00CB6# => romdata <= X"5253B195";
    when 16#00CB7# => romdata <= X"3FB00881";
    when 16#00CB8# => romdata <= X"FF065372";
    when 16#00CB9# => romdata <= X"8C279338";
    when 16#00CBA# => romdata <= X"A051AFA1";
    when 16#00CBB# => romdata <= X"3F811370";
    when 16#00CBC# => romdata <= X"81FF0654";
    when 16#00CBD# => romdata <= X"548C7326";
    when 16#00CBE# => romdata <= X"EF3881E8";
    when 16#00CBF# => romdata <= X"CC51AFA7";
    when 16#00CC0# => romdata <= X"3F81F5CC";
    when 16#00CC1# => romdata <= X"0880E011";
    when 16#00CC2# => romdata <= X"085254B0";
    when 16#00CC3# => romdata <= X"E43F81E8";
    when 16#00CC4# => romdata <= X"E451AF93";
    when 16#00CC5# => romdata <= X"3F81F5CC";
    when 16#00CC6# => romdata <= X"0880D811";
    when 16#00CC7# => romdata <= X"085253B0";
    when 16#00CC8# => romdata <= X"D03F81E8";
    when 16#00CC9# => romdata <= X"FC51AEFF";
    when 16#00CCA# => romdata <= X"3F81F5CC";
    when 16#00CCB# => romdata <= X"08B01108";
    when 16#00CCC# => romdata <= X"FE0A0652";
    when 16#00CCD# => romdata <= X"54B0BA3F";
    when 16#00CCE# => romdata <= X"81F5CC08";
    when 16#00CCF# => romdata <= X"54800BB0";
    when 16#00CD0# => romdata <= X"150C81E9";
    when 16#00CD1# => romdata <= X"9451AEDF";
    when 16#00CD2# => romdata <= X"3F81E9AC";
    when 16#00CD3# => romdata <= X"51AED83F";
    when 16#00CD4# => romdata <= X"81F5CC08";
    when 16#00CD5# => romdata <= X"80C01108";
    when 16#00CD6# => romdata <= X"5253B095";
    when 16#00CD7# => romdata <= X"3FB00881";
    when 16#00CD8# => romdata <= X"FF065372";
    when 16#00CD9# => romdata <= X"98279338";
    when 16#00CDA# => romdata <= X"A051AEA1";
    when 16#00CDB# => romdata <= X"3F811370";
    when 16#00CDC# => romdata <= X"81FF0651";
    when 16#00CDD# => romdata <= X"53987326";
    when 16#00CDE# => romdata <= X"EF3881F5";
    when 16#00CDF# => romdata <= X"CC0880C8";
    when 16#00CE0# => romdata <= X"11085254";
    when 16#00CE1# => romdata <= X"AFEB3FB0";
    when 16#00CE2# => romdata <= X"0881FF06";
    when 16#00CE3# => romdata <= X"53729827";
    when 16#00CE4# => romdata <= X"9338A051";
    when 16#00CE5# => romdata <= X"ADF73F81";
    when 16#00CE6# => romdata <= X"137081FF";
    when 16#00CE7# => romdata <= X"06515398";
    when 16#00CE8# => romdata <= X"7326EF38";
    when 16#00CE9# => romdata <= X"81E9C851";
    when 16#00CEA# => romdata <= X"ADFD3F81";
    when 16#00CEB# => romdata <= X"F5CC0880";
    when 16#00CEC# => romdata <= X"C4110852";
    when 16#00CED# => romdata <= X"54AFBA3F";
    when 16#00CEE# => romdata <= X"B00881FF";
    when 16#00CEF# => romdata <= X"06537298";
    when 16#00CF0# => romdata <= X"279338A0";
    when 16#00CF1# => romdata <= X"51ADC63F";
    when 16#00CF2# => romdata <= X"81137081";
    when 16#00CF3# => romdata <= X"FF065153";
    when 16#00CF4# => romdata <= X"987326EF";
    when 16#00CF5# => romdata <= X"3881F5CC";
    when 16#00CF6# => romdata <= X"0880CC11";
    when 16#00CF7# => romdata <= X"085254AF";
    when 16#00CF8# => romdata <= X"903FB008";
    when 16#00CF9# => romdata <= X"81FF0653";
    when 16#00CFA# => romdata <= X"72982793";
    when 16#00CFB# => romdata <= X"38A051AD";
    when 16#00CFC# => romdata <= X"9C3F8113";
    when 16#00CFD# => romdata <= X"7081FF06";
    when 16#00CFE# => romdata <= X"51539873";
    when 16#00CFF# => romdata <= X"26EF388A";
    when 16#00D00# => romdata <= X"51AD8A3F";
    when 16#00D01# => romdata <= X"81F5CC08";
    when 16#00D02# => romdata <= X"B4110881";
    when 16#00D03# => romdata <= X"E9E45354";
    when 16#00D04# => romdata <= X"54AD943F";
    when 16#00D05# => romdata <= X"80732481";
    when 16#00D06# => romdata <= X"8A387251";
    when 16#00D07# => romdata <= X"AED33FA0";
    when 16#00D08# => romdata <= X"51ACEA3F";
    when 16#00D09# => romdata <= X"72862681";
    when 16#00D0A# => romdata <= X"81387210";
    when 16#00D0B# => romdata <= X"1081EEC8";
    when 16#00D0C# => romdata <= X"05537208";
    when 16#00D0D# => romdata <= X"0481C6E4";
    when 16#00D0E# => romdata <= X"51ACEC3F";
    when 16#00D0F# => romdata <= X"81E68C51";
    when 16#00D10# => romdata <= X"ACE53F81";
    when 16#00D11# => romdata <= X"F5CC0880";
    when 16#00D12# => romdata <= X"D4110852";
    when 16#00D13# => romdata <= X"53AEA23F";
    when 16#00D14# => romdata <= X"81E6A851";
    when 16#00D15# => romdata <= X"ACD13F81";
    when 16#00D16# => romdata <= X"F5CC0880";
    when 16#00D17# => romdata <= X"D0110852";
    when 16#00D18# => romdata <= X"54AE8E3F";
    when 16#00D19# => romdata <= X"8A51ACA5";
    when 16#00D1A# => romdata <= X"3F81E6C4";
    when 16#00D1B# => romdata <= X"51ACB83F";
    when 16#00D1C# => romdata <= X"81E6E851";
    when 16#00D1D# => romdata <= X"ACB13F81";
    when 16#00D1E# => romdata <= X"E7B051AC";
    when 16#00D1F# => romdata <= X"AA3F81E7";
    when 16#00D20# => romdata <= X"F851ACA3";
    when 16#00D21# => romdata <= X"3F81F5CC";
    when 16#00D22# => romdata <= X"08700852";
    when 16#00D23# => romdata <= X"53ADE23F";
    when 16#00D24# => romdata <= X"B00881FF";
    when 16#00D25# => romdata <= X"0653F8EC";
    when 16#00D26# => romdata <= X"3981CE88";
    when 16#00D27# => romdata <= X"51AC883F";
    when 16#00D28# => romdata <= X"F7DE3981";
    when 16#00D29# => romdata <= X"E9F851AB";
    when 16#00D2A# => romdata <= X"FE3F81F5";
    when 16#00D2B# => romdata <= X"CC08B811";
    when 16#00D2C# => romdata <= X"0881EA84";
    when 16#00D2D# => romdata <= X"535553AB";
    when 16#00D2E# => romdata <= X"EE3F7352";
    when 16#00D2F# => romdata <= X"A051AC8A";
    when 16#00D30# => romdata <= X"3F7351F1";
    when 16#00D31# => romdata <= X"993F8A51";
    when 16#00D32# => romdata <= X"ABC33F80";
    when 16#00D33# => romdata <= X"0BB00C85";
    when 16#00D34# => romdata <= X"3D0D0481";
    when 16#00D35# => romdata <= X"EA9851AB";
    when 16#00D36# => romdata <= X"CE3FCF39";
    when 16#00D37# => romdata <= X"81EAA451";
    when 16#00D38# => romdata <= X"ABC53FC6";
    when 16#00D39# => romdata <= X"3981EAB0";
    when 16#00D3A# => romdata <= X"51ABBC3F";
    when 16#00D3B# => romdata <= X"FFBC3981";
    when 16#00D3C# => romdata <= X"EAB451AB";
    when 16#00D3D# => romdata <= X"B23FFFB2";
    when 16#00D3E# => romdata <= X"3981EAC0";
    when 16#00D3F# => romdata <= X"51ABA83F";
    when 16#00D40# => romdata <= X"FFA83981";
    when 16#00D41# => romdata <= X"EACC51AB";
    when 16#00D42# => romdata <= X"9E3FFF9E";
    when 16#00D43# => romdata <= X"3981EAD8";
    when 16#00D44# => romdata <= X"51AB943F";
    when 16#00D45# => romdata <= X"FF9439FD";
    when 16#00D46# => romdata <= X"3D0D81EA";
    when 16#00D47# => romdata <= X"E451AB87";
    when 16#00D48# => romdata <= X"3FFFA5EF";
    when 16#00D49# => romdata <= X"3FB00882";
    when 16#00D4A# => romdata <= X"C63881EA";
    when 16#00D4B# => romdata <= X"EC51AAF7";
    when 16#00D4C# => romdata <= X"3F81F5D4";
    when 16#00D4D# => romdata <= X"3353B352";
    when 16#00D4E# => romdata <= X"7251D381";
    when 16#00D4F# => romdata <= X"3F81EAF0";
    when 16#00D50# => romdata <= X"51AAE43F";
    when 16#00D51# => romdata <= X"81F68C08";
    when 16#00D52# => romdata <= X"84110870";
    when 16#00D53# => romdata <= X"9D2A8106";
    when 16#00D54# => romdata <= X"51545472";
    when 16#00D55# => romdata <= X"802E81EF";
    when 16#00D56# => romdata <= X"3881EAF8";
    when 16#00D57# => romdata <= X"51AAC83F";
    when 16#00D58# => romdata <= X"81EAFC51";
    when 16#00D59# => romdata <= X"AAC13F81";
    when 16#00D5A# => romdata <= X"F5CC0880";
    when 16#00D5B# => romdata <= X"D0110852";
    when 16#00D5C# => romdata <= X"54ABFE3F";
    when 16#00D5D# => romdata <= X"81F5CC08";
    when 16#00D5E# => romdata <= X"54810BB0";
    when 16#00D5F# => romdata <= X"150CB014";
    when 16#00D60# => romdata <= X"08537280";
    when 16#00D61# => romdata <= X"25F83881";
    when 16#00D62# => romdata <= X"EB8C51AA";
    when 16#00D63# => romdata <= X"9A3F81F5";
    when 16#00D64# => romdata <= X"CC08A011";
    when 16#00D65# => romdata <= X"085254AB";
    when 16#00D66# => romdata <= X"D83F81F5";
    when 16#00D67# => romdata <= X"D43353B3";
    when 16#00D68# => romdata <= X"527251D2";
    when 16#00D69# => romdata <= X"983F81EB";
    when 16#00D6A# => romdata <= X"9451A9FB";
    when 16#00D6B# => romdata <= X"3F81F5CC";
    when 16#00D6C# => romdata <= X"08A41108";
    when 16#00D6D# => romdata <= X"5254ABB9";
    when 16#00D6E# => romdata <= X"3F81EB9C";
    when 16#00D6F# => romdata <= X"51A9E83F";
    when 16#00D70# => romdata <= X"81F5CC08";
    when 16#00D71# => romdata <= X"A8110852";
    when 16#00D72# => romdata <= X"53ABA63F";
    when 16#00D73# => romdata <= X"81F5D433";
    when 16#00D74# => romdata <= X"54B35273";
    when 16#00D75# => romdata <= X"51D1E63F";
    when 16#00D76# => romdata <= X"81EBA451";
    when 16#00D77# => romdata <= X"A9C93F81";
    when 16#00D78# => romdata <= X"F5CC08AC";
    when 16#00D79# => romdata <= X"11085253";
    when 16#00D7A# => romdata <= X"AB873F81";
    when 16#00D7B# => romdata <= X"EBAC51A9";
    when 16#00D7C# => romdata <= X"B63F81F5";
    when 16#00D7D# => romdata <= X"CC0880E0";
    when 16#00D7E# => romdata <= X"11085254";
    when 16#00D7F# => romdata <= X"AAF33F81";
    when 16#00D80# => romdata <= X"F5D43353";
    when 16#00D81# => romdata <= X"B3527251";
    when 16#00D82# => romdata <= X"D1B33F81";
    when 16#00D83# => romdata <= X"EBB451A9";
    when 16#00D84# => romdata <= X"963F81F5";
    when 16#00D85# => romdata <= X"CC08B011";
    when 16#00D86# => romdata <= X"08FE0A06";
    when 16#00D87# => romdata <= X"5254AAD1";
    when 16#00D88# => romdata <= X"3F81F5CC";
    when 16#00D89# => romdata <= X"0854800B";
    when 16#00D8A# => romdata <= X"B0150CB4";
    when 16#00D8B# => romdata <= X"140881EB";
    when 16#00D8C# => romdata <= X"BC5253A8";
    when 16#00D8D# => romdata <= X"F23F7286";
    when 16#00D8E# => romdata <= X"2680C238";
    when 16#00D8F# => romdata <= X"72101081";
    when 16#00D90# => romdata <= X"EEE40553";
    when 16#00D91# => romdata <= X"72080481";
    when 16#00D92# => romdata <= X"EBC851A8";
    when 16#00D93# => romdata <= X"DA3F81EA";
    when 16#00D94# => romdata <= X"FC51A8D3";
    when 16#00D95# => romdata <= X"3F81F5CC";
    when 16#00D96# => romdata <= X"0880D011";
    when 16#00D97# => romdata <= X"085254AA";
    when 16#00D98# => romdata <= X"903F81F5";
    when 16#00D99# => romdata <= X"CC085481";
    when 16#00D9A# => romdata <= X"0BB0150C";
    when 16#00D9B# => romdata <= X"FE903981";
    when 16#00D9C# => romdata <= X"EAF851FD";
    when 16#00D9D# => romdata <= X"B93981EA";
    when 16#00D9E# => romdata <= X"D851A8AB";
    when 16#00D9F# => romdata <= X"3F81F5CC";
    when 16#00DA0# => romdata <= X"08B81108";
    when 16#00DA1# => romdata <= X"81EBD053";
    when 16#00DA2# => romdata <= X"5553A89B";
    when 16#00DA3# => romdata <= X"3F7352A0";
    when 16#00DA4# => romdata <= X"51A8B73F";
    when 16#00DA5# => romdata <= X"8A51A7F5";
    when 16#00DA6# => romdata <= X"3F738106";
    when 16#00DA7# => romdata <= X"537285DF";
    when 16#00DA8# => romdata <= X"3873812A";
    when 16#00DA9# => romdata <= X"70810651";
    when 16#00DAA# => romdata <= X"537285BC";
    when 16#00DAB# => romdata <= X"3873822A";
    when 16#00DAC# => romdata <= X"70810651";
    when 16#00DAD# => romdata <= X"53728599";
    when 16#00DAE# => romdata <= X"3873832A";
    when 16#00DAF# => romdata <= X"70810651";
    when 16#00DB0# => romdata <= X"537284F6";
    when 16#00DB1# => romdata <= X"3873842A";
    when 16#00DB2# => romdata <= X"70810651";
    when 16#00DB3# => romdata <= X"537284D3";
    when 16#00DB4# => romdata <= X"3873852A";
    when 16#00DB5# => romdata <= X"70810651";
    when 16#00DB6# => romdata <= X"537284B0";
    when 16#00DB7# => romdata <= X"3873862A";
    when 16#00DB8# => romdata <= X"70810651";
    when 16#00DB9# => romdata <= X"5372848D";
    when 16#00DBA# => romdata <= X"3873872A";
    when 16#00DBB# => romdata <= X"70810651";
    when 16#00DBC# => romdata <= X"537283EA";
    when 16#00DBD# => romdata <= X"3873882A";
    when 16#00DBE# => romdata <= X"70810651";
    when 16#00DBF# => romdata <= X"537283C7";
    when 16#00DC0# => romdata <= X"3873892A";
    when 16#00DC1# => romdata <= X"70810651";
    when 16#00DC2# => romdata <= X"537283A4";
    when 16#00DC3# => romdata <= X"38738A2A";
    when 16#00DC4# => romdata <= X"70810651";
    when 16#00DC5# => romdata <= X"53728381";
    when 16#00DC6# => romdata <= X"38738B2A";
    when 16#00DC7# => romdata <= X"70810651";
    when 16#00DC8# => romdata <= X"537282DE";
    when 16#00DC9# => romdata <= X"38738C2A";
    when 16#00DCA# => romdata <= X"70810651";
    when 16#00DCB# => romdata <= X"537282BB";
    when 16#00DCC# => romdata <= X"38738D2A";
    when 16#00DCD# => romdata <= X"70810651";
    when 16#00DCE# => romdata <= X"53728298";
    when 16#00DCF# => romdata <= X"38738E2A";
    when 16#00DD0# => romdata <= X"70810651";
    when 16#00DD1# => romdata <= X"537281F5";
    when 16#00DD2# => romdata <= X"38738F2A";
    when 16#00DD3# => romdata <= X"70810651";
    when 16#00DD4# => romdata <= X"537281D2";
    when 16#00DD5# => romdata <= X"3873902A";
    when 16#00DD6# => romdata <= X"70810651";
    when 16#00DD7# => romdata <= X"537281AF";
    when 16#00DD8# => romdata <= X"3873912A";
    when 16#00DD9# => romdata <= X"70810651";
    when 16#00DDA# => romdata <= X"5372818C";
    when 16#00DDB# => romdata <= X"3873922A";
    when 16#00DDC# => romdata <= X"70810651";
    when 16#00DDD# => romdata <= X"537280E9";
    when 16#00DDE# => romdata <= X"3873932A";
    when 16#00DDF# => romdata <= X"70810651";
    when 16#00DE0# => romdata <= X"537280C6";
    when 16#00DE1# => romdata <= X"3873942A";
    when 16#00DE2# => romdata <= X"70810651";
    when 16#00DE3# => romdata <= X"5372A538";
    when 16#00DE4# => romdata <= X"73952A70";
    when 16#00DE5# => romdata <= X"81065153";
    when 16#00DE6# => romdata <= X"728B3880";
    when 16#00DE7# => romdata <= X"742483F6";
    when 16#00DE8# => romdata <= X"38853D0D";
    when 16#00DE9# => romdata <= X"0481EBE0";
    when 16#00DEA# => romdata <= X"51A5FC3F";
    when 16#00DEB# => romdata <= X"738025F1";
    when 16#00DEC# => romdata <= X"3883E339";
    when 16#00DED# => romdata <= X"81EBF051";
    when 16#00DEE# => romdata <= X"A5ED3F73";
    when 16#00DEF# => romdata <= X"952A7081";
    when 16#00DF0# => romdata <= X"06515372";
    when 16#00DF1# => romdata <= X"802ED438";
    when 16#00DF2# => romdata <= X"DC3981EC";
    when 16#00DF3# => romdata <= X"8051A5D7";
    when 16#00DF4# => romdata <= X"3F73942A";
    when 16#00DF5# => romdata <= X"70810651";
    when 16#00DF6# => romdata <= X"5372802E";
    when 16#00DF7# => romdata <= X"FFB238D4";
    when 16#00DF8# => romdata <= X"3981EC90";
    when 16#00DF9# => romdata <= X"51A5C03F";
    when 16#00DFA# => romdata <= X"73932A70";
    when 16#00DFB# => romdata <= X"81065153";
    when 16#00DFC# => romdata <= X"72802EFF";
    when 16#00DFD# => romdata <= X"9038D339";
    when 16#00DFE# => romdata <= X"81ECA051";
    when 16#00DFF# => romdata <= X"A5A93F73";
    when 16#00E00# => romdata <= X"922A7081";
    when 16#00E01# => romdata <= X"06515372";
    when 16#00E02# => romdata <= X"802EFEED";
    when 16#00E03# => romdata <= X"38D33981";
    when 16#00E04# => romdata <= X"ECB051A5";
    when 16#00E05# => romdata <= X"923F7391";
    when 16#00E06# => romdata <= X"2A708106";
    when 16#00E07# => romdata <= X"51537280";
    when 16#00E08# => romdata <= X"2EFECA38";
    when 16#00E09# => romdata <= X"D33981EC";
    when 16#00E0A# => romdata <= X"C051A4FB";
    when 16#00E0B# => romdata <= X"3F73902A";
    when 16#00E0C# => romdata <= X"70810651";
    when 16#00E0D# => romdata <= X"5372802E";
    when 16#00E0E# => romdata <= X"FEA738D3";
    when 16#00E0F# => romdata <= X"3981ECD0";
    when 16#00E10# => romdata <= X"51A4E43F";
    when 16#00E11# => romdata <= X"738F2A70";
    when 16#00E12# => romdata <= X"81065153";
    when 16#00E13# => romdata <= X"72802EFE";
    when 16#00E14# => romdata <= X"8438D339";
    when 16#00E15# => romdata <= X"81ECE051";
    when 16#00E16# => romdata <= X"A4CD3F73";
    when 16#00E17# => romdata <= X"8E2A7081";
    when 16#00E18# => romdata <= X"06515372";
    when 16#00E19# => romdata <= X"802EFDE1";
    when 16#00E1A# => romdata <= X"38D33981";
    when 16#00E1B# => romdata <= X"ECF051A4";
    when 16#00E1C# => romdata <= X"B63F738D";
    when 16#00E1D# => romdata <= X"2A708106";
    when 16#00E1E# => romdata <= X"51537280";
    when 16#00E1F# => romdata <= X"2EFDBE38";
    when 16#00E20# => romdata <= X"D33981EC";
    when 16#00E21# => romdata <= X"FC51A49F";
    when 16#00E22# => romdata <= X"3F738C2A";
    when 16#00E23# => romdata <= X"70810651";
    when 16#00E24# => romdata <= X"5372802E";
    when 16#00E25# => romdata <= X"FD9B38D3";
    when 16#00E26# => romdata <= X"3981ED8C";
    when 16#00E27# => romdata <= X"51A4883F";
    when 16#00E28# => romdata <= X"738B2A70";
    when 16#00E29# => romdata <= X"81065153";
    when 16#00E2A# => romdata <= X"72802EFC";
    when 16#00E2B# => romdata <= X"F838D339";
    when 16#00E2C# => romdata <= X"81ED9C51";
    when 16#00E2D# => romdata <= X"A3F13F73";
    when 16#00E2E# => romdata <= X"8A2A7081";
    when 16#00E2F# => romdata <= X"06515372";
    when 16#00E30# => romdata <= X"802EFCD5";
    when 16#00E31# => romdata <= X"38D33981";
    when 16#00E32# => romdata <= X"EDAC51A3";
    when 16#00E33# => romdata <= X"DA3F7389";
    when 16#00E34# => romdata <= X"2A708106";
    when 16#00E35# => romdata <= X"51537280";
    when 16#00E36# => romdata <= X"2EFCB238";
    when 16#00E37# => romdata <= X"D33981ED";
    when 16#00E38# => romdata <= X"BC51A3C3";
    when 16#00E39# => romdata <= X"3F73882A";
    when 16#00E3A# => romdata <= X"70810651";
    when 16#00E3B# => romdata <= X"5372802E";
    when 16#00E3C# => romdata <= X"FC8F38D3";
    when 16#00E3D# => romdata <= X"3981EDCC";
    when 16#00E3E# => romdata <= X"51A3AC3F";
    when 16#00E3F# => romdata <= X"73872A70";
    when 16#00E40# => romdata <= X"81065153";
    when 16#00E41# => romdata <= X"72802EFB";
    when 16#00E42# => romdata <= X"EC38D339";
    when 16#00E43# => romdata <= X"81EDDC51";
    when 16#00E44# => romdata <= X"A3953F73";
    when 16#00E45# => romdata <= X"862A7081";
    when 16#00E46# => romdata <= X"06515372";
    when 16#00E47# => romdata <= X"802EFBC9";
    when 16#00E48# => romdata <= X"38D33981";
    when 16#00E49# => romdata <= X"EDEC51A2";
    when 16#00E4A# => romdata <= X"FE3F7385";
    when 16#00E4B# => romdata <= X"2A708106";
    when 16#00E4C# => romdata <= X"51537280";
    when 16#00E4D# => romdata <= X"2EFBA638";
    when 16#00E4E# => romdata <= X"D33981ED";
    when 16#00E4F# => romdata <= X"FC51A2E7";
    when 16#00E50# => romdata <= X"3F73842A";
    when 16#00E51# => romdata <= X"70810651";
    when 16#00E52# => romdata <= X"5372802E";
    when 16#00E53# => romdata <= X"FB8338D3";
    when 16#00E54# => romdata <= X"3981EE8C";
    when 16#00E55# => romdata <= X"51A2D03F";
    when 16#00E56# => romdata <= X"73832A70";
    when 16#00E57# => romdata <= X"81065153";
    when 16#00E58# => romdata <= X"72802EFA";
    when 16#00E59# => romdata <= X"E038D339";
    when 16#00E5A# => romdata <= X"81EE9C51";
    when 16#00E5B# => romdata <= X"A2B93F73";
    when 16#00E5C# => romdata <= X"822A7081";
    when 16#00E5D# => romdata <= X"06515372";
    when 16#00E5E# => romdata <= X"802EFABD";
    when 16#00E5F# => romdata <= X"38D33981";
    when 16#00E60# => romdata <= X"EEAC51A2";
    when 16#00E61# => romdata <= X"A23F7381";
    when 16#00E62# => romdata <= X"2A708106";
    when 16#00E63# => romdata <= X"51537280";
    when 16#00E64# => romdata <= X"2EFA9A38";
    when 16#00E65# => romdata <= X"D33981EE";
    when 16#00E66# => romdata <= X"BC51A28B";
    when 16#00E67# => romdata <= X"3F853D0D";
    when 16#00E68# => romdata <= X"0481EA98";
    when 16#00E69# => romdata <= X"51A2803F";
    when 16#00E6A# => romdata <= X"F9D33981";
    when 16#00E6B# => romdata <= X"EAA451A1";
    when 16#00E6C# => romdata <= X"F63FF9C9";
    when 16#00E6D# => romdata <= X"3981EAB0";
    when 16#00E6E# => romdata <= X"51A1EC3F";
    when 16#00E6F# => romdata <= X"F9BF3981";
    when 16#00E70# => romdata <= X"EAB451A1";
    when 16#00E71# => romdata <= X"E23FF9B5";
    when 16#00E72# => romdata <= X"3981EAC0";
    when 16#00E73# => romdata <= X"51A1D83F";
    when 16#00E74# => romdata <= X"F9AB3981";
    when 16#00E75# => romdata <= X"EACC51A1";
    when 16#00E76# => romdata <= X"CE3FF9A1";
    when 16#00E77# => romdata <= X"39FE3D0D";
    when 16#00E78# => romdata <= X"CAFE3F80";
    when 16#00E79# => romdata <= X"5281D684";
    when 16#00E7A# => romdata <= X"51CDC83F";
    when 16#00E7B# => romdata <= X"829EBC08";
    when 16#00E7C# => romdata <= X"80D2F70B";
    when 16#00E7D# => romdata <= X"829EBC0C";
    when 16#00E7E# => romdata <= X"53F69C3F";
    when 16#00E7F# => romdata <= X"72829EBC";
    when 16#00E80# => romdata <= X"0C843D0D";
    when 16#00E81# => romdata <= X"04FD3D0D";
    when 16#00E82# => romdata <= X"8151FFAF";
    when 16#00E83# => romdata <= X"BA3FB008";
    when 16#00E84# => romdata <= X"81FF0654";
    when 16#00E85# => romdata <= X"8251FFAF";
    when 16#00E86# => romdata <= X"AE3FB008";
    when 16#00E87# => romdata <= X"9F2B7407";
    when 16#00E88# => romdata <= X"81F5CC08";
    when 16#00E89# => romdata <= X"53B4130C";
    when 16#00E8A# => romdata <= X"73B00C85";
    when 16#00E8B# => romdata <= X"3D0D04FD";
    when 16#00E8C# => romdata <= X"3D0D81EF";
    when 16#00E8D# => romdata <= X"F851A0EF";
    when 16#00E8E# => romdata <= X"3F81F5C8";
    when 16#00E8F# => romdata <= X"08841108";
    when 16#00E90# => romdata <= X"5254A2AD";
    when 16#00E91# => romdata <= X"3F81F088";
    when 16#00E92# => romdata <= X"51A0DC3F";
    when 16#00E93# => romdata <= X"81F5C808";
    when 16#00E94# => romdata <= X"88110852";
    when 16#00E95# => romdata <= X"53A29A3F";
    when 16#00E96# => romdata <= X"81F09851";
    when 16#00E97# => romdata <= X"A0C93F81";
    when 16#00E98# => romdata <= X"F5C8088C";
    when 16#00E99# => romdata <= X"11085254";
    when 16#00E9A# => romdata <= X"A2873F81";
    when 16#00E9B# => romdata <= X"F0A851A0";
    when 16#00E9C# => romdata <= X"B63F81F5";
    when 16#00E9D# => romdata <= X"C8089011";
    when 16#00E9E# => romdata <= X"085253A1";
    when 16#00E9F# => romdata <= X"F43F81F0";
    when 16#00EA0# => romdata <= X"B851A0A3";
    when 16#00EA1# => romdata <= X"3F81F5C8";
    when 16#00EA2# => romdata <= X"08941108";
    when 16#00EA3# => romdata <= X"5254A1E1";
    when 16#00EA4# => romdata <= X"3F81F5C8";
    when 16#00EA5# => romdata <= X"08700881";
    when 16#00EA6# => romdata <= X"F0C85355";
    when 16#00EA7# => romdata <= X"53A0883F";
    when 16#00EA8# => romdata <= X"73528851";
    when 16#00EA9# => romdata <= X"A0A43F73";
    when 16#00EAA# => romdata <= X"81065372";
    when 16#00EAB# => romdata <= X"802E80C2";
    when 16#00EAC# => romdata <= X"3881EF80";
    when 16#00EAD# => romdata <= X"519FF03F";
    when 16#00EAE# => romdata <= X"73812A70";
    when 16#00EAF# => romdata <= X"81065153";
    when 16#00EB0# => romdata <= X"72818738";
    when 16#00EB1# => romdata <= X"73822A70";
    when 16#00EB2# => romdata <= X"81065153";
    when 16#00EB3# => romdata <= X"7280E438";
    when 16#00EB4# => romdata <= X"73832A70";
    when 16#00EB5# => romdata <= X"81065153";
    when 16#00EB6# => romdata <= X"7280C338";
    when 16#00EB7# => romdata <= X"73842A81";
    when 16#00EB8# => romdata <= X"065473A6";
    when 16#00EB9# => romdata <= X"388A519F";
    when 16#00EBA# => romdata <= X"A43F800B";
    when 16#00EBB# => romdata <= X"B00C853D";
    when 16#00EBC# => romdata <= X"0D0481EF";
    when 16#00EBD# => romdata <= X"90519FAF";
    when 16#00EBE# => romdata <= X"3F73812A";
    when 16#00EBF# => romdata <= X"70810651";
    when 16#00EC0# => romdata <= X"5372802E";
    when 16#00EC1# => romdata <= X"FFBE3880";
    when 16#00EC2# => romdata <= X"C13981EF";
    when 16#00EC3# => romdata <= X"A4519F97";
    when 16#00EC4# => romdata <= X"3F8A519E";
    when 16#00EC5# => romdata <= X"F83F800B";
    when 16#00EC6# => romdata <= X"B00C853D";
    when 16#00EC7# => romdata <= X"0D0481EF";
    when 16#00EC8# => romdata <= X"BC519F83";
    when 16#00EC9# => romdata <= X"3F73842A";
    when 16#00ECA# => romdata <= X"81065473";
    when 16#00ECB# => romdata <= X"802EFFB5";
    when 16#00ECC# => romdata <= X"38D83981";
    when 16#00ECD# => romdata <= X"EFD8519E";
    when 16#00ECE# => romdata <= X"EE3F7383";
    when 16#00ECF# => romdata <= X"2A708106";
    when 16#00ED0# => romdata <= X"51537280";
    when 16#00ED1# => romdata <= X"2EFF9538";
    when 16#00ED2# => romdata <= X"D53981EF";
    when 16#00ED3# => romdata <= X"EC519ED7";
    when 16#00ED4# => romdata <= X"3F73822A";
    when 16#00ED5# => romdata <= X"70810651";
    when 16#00ED6# => romdata <= X"5372802E";
    when 16#00ED7# => romdata <= X"FEF238D3";
    when 16#00ED8# => romdata <= X"39FF3D0D";
    when 16#00ED9# => romdata <= X"8151FFAC";
    when 16#00EDA# => romdata <= X"DE3F81F5";
    when 16#00EDB# => romdata <= X"C808B008";
    when 16#00EDC# => romdata <= X"90120C52";
    when 16#00EDD# => romdata <= X"8251FFAC";
    when 16#00EDE# => romdata <= X"CE3F81F5";
    when 16#00EDF# => romdata <= X"C808B008";
    when 16#00EE0# => romdata <= X"94120C52";
    when 16#00EE1# => romdata <= X"800BB00C";
    when 16#00EE2# => romdata <= X"833D0D04";
    when 16#00EE3# => romdata <= X"FF3D0D81";
    when 16#00EE4# => romdata <= X"F5C80870";
    when 16#00EE5# => romdata <= X"08535180";
    when 16#00EE6# => romdata <= X"710C71B0";
    when 16#00EE7# => romdata <= X"0C833D0D";
    when 16#00EE8# => romdata <= X"04F93D0D";
    when 16#00EE9# => romdata <= X"02A60522";
    when 16#00EEA# => romdata <= X"81F5D833";
    when 16#00EEB# => romdata <= X"81F70655";
    when 16#00EEC# => romdata <= X"567381F5";
    when 16#00EED# => romdata <= X"D8347353";
    when 16#00EEE# => romdata <= X"A05281F6";
    when 16#00EEF# => romdata <= X"800851E0";
    when 16#00EF0# => romdata <= X"9F3F8057";
    when 16#00EF1# => romdata <= X"8F5581F5";
    when 16#00EF2# => romdata <= X"D83381FE";
    when 16#00EF3# => romdata <= X"06547381";
    when 16#00EF4# => romdata <= X"F5D83473";
    when 16#00EF5# => romdata <= X"53A05281";
    when 16#00EF6# => romdata <= X"F6800851";
    when 16#00EF7# => romdata <= X"E0823F75";
    when 16#00EF8# => romdata <= X"752C8106";
    when 16#00EF9# => romdata <= X"5877802E";
    when 16#00EFA# => romdata <= X"819E3881";
    when 16#00EFB# => romdata <= X"F5D83382";
    when 16#00EFC# => romdata <= X"07547381";
    when 16#00EFD# => romdata <= X"F5D83473";
    when 16#00EFE# => romdata <= X"53A05281";
    when 16#00EFF# => romdata <= X"F6800851";
    when 16#00F00# => romdata <= X"DFDE3FA0";
    when 16#00F01# => romdata <= X"5281F680";
    when 16#00F02# => romdata <= X"0851E09E";
    when 16#00F03# => romdata <= X"3FB00882";
    when 16#00F04# => romdata <= X"2A810654";
    when 16#00F05# => romdata <= X"73802E8D";
    when 16#00F06# => romdata <= X"3881752B";
    when 16#00F07# => romdata <= X"77077083";
    when 16#00F08# => romdata <= X"FFFF0658";
    when 16#00F09# => romdata <= X"5481F5D8";
    when 16#00F0A# => romdata <= X"33810754";
    when 16#00F0B# => romdata <= X"7381F5D8";
    when 16#00F0C# => romdata <= X"347353A0";
    when 16#00F0D# => romdata <= X"5281F680";
    when 16#00F0E# => romdata <= X"0851DFA4";
    when 16#00F0F# => romdata <= X"3F748180";
    when 16#00F10# => romdata <= X"0A2981FF";
    when 16#00F11# => romdata <= X"0A057098";
    when 16#00F12# => romdata <= X"2C565874";
    when 16#00F13# => romdata <= X"8025FEF6";
    when 16#00F14# => romdata <= X"3881F5D8";
    when 16#00F15# => romdata <= X"33820754";
    when 16#00F16# => romdata <= X"7381F5D8";
    when 16#00F17# => romdata <= X"347353A0";
    when 16#00F18# => romdata <= X"5281F680";
    when 16#00F19# => romdata <= X"0851DEF8";
    when 16#00F1A# => romdata <= X"3F81F5D8";
    when 16#00F1B# => romdata <= X"33880756";
    when 16#00F1C# => romdata <= X"7581F5D8";
    when 16#00F1D# => romdata <= X"347553A0";
    when 16#00F1E# => romdata <= X"5281F680";
    when 16#00F1F# => romdata <= X"0851DEE0";
    when 16#00F20# => romdata <= X"3F76B00C";
    when 16#00F21# => romdata <= X"893D0D04";
    when 16#00F22# => romdata <= X"81F5D833";
    when 16#00F23# => romdata <= X"81FD0654";
    when 16#00F24# => romdata <= X"FEE039FB";
    when 16#00F25# => romdata <= X"3D0D029F";
    when 16#00F26# => romdata <= X"05335680";
    when 16#00F27# => romdata <= X"C05381D0";
    when 16#00F28# => romdata <= X"5281F680";
    when 16#00F29# => romdata <= X"0851C0CD";
    when 16#00F2A# => romdata <= X"3FB00887";
    when 16#00F2B# => romdata <= X"2A810655";
    when 16#00F2C# => romdata <= X"FF5474A5";
    when 16#00F2D# => romdata <= X"38818051";
    when 16#00F2E# => romdata <= X"FDE73F82";
    when 16#00F2F# => romdata <= X"8051FDE1";
    when 16#00F30# => romdata <= X"3F848351";
    when 16#00F31# => romdata <= X"FDDB3F86";
    when 16#00F32# => romdata <= X"F151FDD5";
    when 16#00F33# => romdata <= X"3F75832B";
    when 16#00F34# => romdata <= X"88830751";
    when 16#00F35# => romdata <= X"FDCB3F74";
    when 16#00F36# => romdata <= X"5473B00C";
    when 16#00F37# => romdata <= X"873D0D04";
    when 16#00F38# => romdata <= X"FC3D0D81";
    when 16#00F39# => romdata <= X"51FFA9DF";
    when 16#00F3A# => romdata <= X"3FB00881";
    when 16#00F3B# => romdata <= X"FF065580";
    when 16#00F3C# => romdata <= X"C05381D0";
    when 16#00F3D# => romdata <= X"5281F680";
    when 16#00F3E# => romdata <= X"0851FFBF";
    when 16#00F3F# => romdata <= X"F83FB008";
    when 16#00F40# => romdata <= X"872A7081";
    when 16#00F41# => romdata <= X"06515473";
    when 16#00F42# => romdata <= X"802E8838";
    when 16#00F43# => romdata <= X"74B00C86";
    when 16#00F44# => romdata <= X"3D0D0481";
    when 16#00F45# => romdata <= X"8051FD89";
    when 16#00F46# => romdata <= X"3F828051";
    when 16#00F47# => romdata <= X"FD833F84";
    when 16#00F48# => romdata <= X"8351FCFD";
    when 16#00F49# => romdata <= X"3F86F151";
    when 16#00F4A# => romdata <= X"FCF73F74";
    when 16#00F4B# => romdata <= X"832B8883";
    when 16#00F4C# => romdata <= X"0751FCED";
    when 16#00F4D# => romdata <= X"3F74B00C";
    when 16#00F4E# => romdata <= X"863D0D04";
    when 16#00F4F# => romdata <= X"803D0D81";
    when 16#00F50# => romdata <= X"51FFAAB6";
    when 16#00F51# => romdata <= X"3FB00883";
    when 16#00F52# => romdata <= X"FFFF0651";
    when 16#00F53# => romdata <= X"FCD33FB0";
    when 16#00F54# => romdata <= X"0883FFFF";
    when 16#00F55# => romdata <= X"06B00C82";
    when 16#00F56# => romdata <= X"3D0D0480";
    when 16#00F57# => romdata <= X"0B829DD8";
    when 16#00F58# => romdata <= X"34800BB0";
    when 16#00F59# => romdata <= X"0C04FB3D";
    when 16#00F5A# => romdata <= X"0D8151FF";
    when 16#00F5B# => romdata <= X"AA8C3FB0";
    when 16#00F5C# => romdata <= X"08538251";
    when 16#00F5D# => romdata <= X"FFAA833F";
    when 16#00F5E# => romdata <= X"B00856B0";
    when 16#00F5F# => romdata <= X"08833890";
    when 16#00F60# => romdata <= X"5672FC06";
    when 16#00F61# => romdata <= X"5575812E";
    when 16#00F62# => romdata <= X"80F13880";
    when 16#00F63# => romdata <= X"54737627";
    when 16#00F64# => romdata <= X"AA387383";
    when 16#00F65# => romdata <= X"06537280";
    when 16#00F66# => romdata <= X"2EAE3881";
    when 16#00F67# => romdata <= X"D5AC519A";
    when 16#00F68# => romdata <= X"863F7470";
    when 16#00F69# => romdata <= X"84055608";
    when 16#00F6A# => romdata <= X"52A0519A";
    when 16#00F6B# => romdata <= X"9D3FA051";
    when 16#00F6C# => romdata <= X"99DB3F81";
    when 16#00F6D# => romdata <= X"14547574";
    when 16#00F6E# => romdata <= X"26D8388A";
    when 16#00F6F# => romdata <= X"5199CE3F";
    when 16#00F70# => romdata <= X"800BB00C";
    when 16#00F71# => romdata <= X"873D0D04";
    when 16#00F72# => romdata <= X"81F0DC51";
    when 16#00F73# => romdata <= X"99D93F74";
    when 16#00F74# => romdata <= X"52A05199";
    when 16#00F75# => romdata <= X"F53F81F1";
    when 16#00F76# => romdata <= X"FC5199CB";
    when 16#00F77# => romdata <= X"3F81D5AC";
    when 16#00F78# => romdata <= X"5199C43F";
    when 16#00F79# => romdata <= X"74708405";
    when 16#00F7A# => romdata <= X"560852A0";
    when 16#00F7B# => romdata <= X"5199DB3F";
    when 16#00F7C# => romdata <= X"A0519999";
    when 16#00F7D# => romdata <= X"3F811454";
    when 16#00F7E# => romdata <= X"FFBC3981";
    when 16#00F7F# => romdata <= X"D5AC5199";
    when 16#00F80# => romdata <= X"A63F7408";
    when 16#00F81# => romdata <= X"52A05199";
    when 16#00F82# => romdata <= X"C13F8A51";
    when 16#00F83# => romdata <= X"98FF3F80";
    when 16#00F84# => romdata <= X"0BB00C87";
    when 16#00F85# => romdata <= X"3D0D04FC";
    when 16#00F86# => romdata <= X"3D0D8151";
    when 16#00F87# => romdata <= X"FFA8DB3F";
    when 16#00F88# => romdata <= X"B0085282";
    when 16#00F89# => romdata <= X"51FFA79F";
    when 16#00F8A# => romdata <= X"3FB00881";
    when 16#00F8B# => romdata <= X"FF067256";
    when 16#00F8C# => romdata <= X"53835472";
    when 16#00F8D# => romdata <= X"802EA238";
    when 16#00F8E# => romdata <= X"7351FFA8";
    when 16#00F8F# => romdata <= X"BD3F8114";
    when 16#00F90# => romdata <= X"7081FF06";
    when 16#00F91# => romdata <= X"FF157081";
    when 16#00F92# => romdata <= X"FF06B008";
    when 16#00F93# => romdata <= X"79708405";
    when 16#00F94# => romdata <= X"5B0C5652";
    when 16#00F95# => romdata <= X"555272E0";
    when 16#00F96# => romdata <= X"3872B00C";
    when 16#00F97# => romdata <= X"863D0D04";
    when 16#00F98# => romdata <= X"803D0D8C";
    when 16#00F99# => romdata <= X"5198A63F";
    when 16#00F9A# => romdata <= X"800BB00C";
    when 16#00F9B# => romdata <= X"823D0D04";
    when 16#00F9C# => romdata <= X"803D0D81";
    when 16#00F9D# => romdata <= X"F6980851";
    when 16#00F9E# => romdata <= X"F8BB9586";
    when 16#00F9F# => romdata <= X"A1710C81";
    when 16#00FA0# => romdata <= X"0BB00C82";
    when 16#00FA1# => romdata <= X"3D0D0480";
    when 16#00FA2# => romdata <= X"3D0D8151";
    when 16#00FA3# => romdata <= X"FFA6B83F";
    when 16#00FA4# => romdata <= X"B00881FF";
    when 16#00FA5# => romdata <= X"0651FFB8";
    when 16#00FA6# => romdata <= X"EC3F800B";
    when 16#00FA7# => romdata <= X"B00C823D";
    when 16#00FA8# => romdata <= X"0D04FA3D";
    when 16#00FA9# => romdata <= X"0D880A57";
    when 16#00FAA# => romdata <= X"840A5681";
    when 16#00FAB# => romdata <= X"51FFA697";
    when 16#00FAC# => romdata <= X"3FB00883";
    when 16#00FAD# => romdata <= X"FFFF0654";
    when 16#00FAE# => romdata <= X"73833890";
    when 16#00FAF# => romdata <= X"54805574";
    when 16#00FB0# => romdata <= X"742780E7";
    when 16#00FB1# => romdata <= X"38757084";
    when 16#00FB2# => romdata <= X"05570870";
    when 16#00FB3# => romdata <= X"902C5253";
    when 16#00FB4# => romdata <= X"999F3F8A";
    when 16#00FB5# => romdata <= X"52B00851";
    when 16#00FB6# => romdata <= X"DCDA3F72";
    when 16#00FB7# => romdata <= X"902B7090";
    when 16#00FB8# => romdata <= X"2C525399";
    when 16#00FB9# => romdata <= X"8C3F8A52";
    when 16#00FBA# => romdata <= X"B00851DC";
    when 16#00FBB# => romdata <= X"C73F7670";
    when 16#00FBC# => romdata <= X"84055808";
    when 16#00FBD# => romdata <= X"70902C52";
    when 16#00FBE# => romdata <= X"5398F63F";
    when 16#00FBF# => romdata <= X"8A52B008";
    when 16#00FC0# => romdata <= X"51DCB13F";
    when 16#00FC1# => romdata <= X"72902B70";
    when 16#00FC2# => romdata <= X"902C5253";
    when 16#00FC3# => romdata <= X"98E33F8A";
    when 16#00FC4# => romdata <= X"52B00851";
    when 16#00FC5# => romdata <= X"DC9E3F8A";
    when 16#00FC6# => romdata <= X"5196F23F";
    when 16#00FC7# => romdata <= X"81157083";
    when 16#00FC8# => romdata <= X"FFFF0656";
    when 16#00FC9# => romdata <= X"53737526";
    when 16#00FCA# => romdata <= X"FF9B3873";
    when 16#00FCB# => romdata <= X"B00C883D";
    when 16#00FCC# => romdata <= X"0D04FD3D";
    when 16#00FCD# => romdata <= X"0D81F5E0";
    when 16#00FCE# => romdata <= X"088C1108";
    when 16#00FCF# => romdata <= X"70822B83";
    when 16#00FD0# => romdata <= X"FFFC0681";
    when 16#00FD1# => romdata <= X"F0E05451";
    when 16#00FD2# => romdata <= X"545496DB";
    when 16#00FD3# => romdata <= X"3F725288";
    when 16#00FD4# => romdata <= X"0A51FFAB";
    when 16#00FD5# => romdata <= X"C43FB008";
    when 16#00FD6# => romdata <= X"54B008FE";
    when 16#00FD7# => romdata <= X"2EA838B0";
    when 16#00FD8# => romdata <= X"08FF2E94";
    when 16#00FD9# => romdata <= X"38725198";
    when 16#00FDA# => romdata <= X"883F81F0";
    when 16#00FDB# => romdata <= X"F45196B7";
    when 16#00FDC# => romdata <= X"3F73B00C";
    when 16#00FDD# => romdata <= X"853D0D04";
    when 16#00FDE# => romdata <= X"81F18851";
    when 16#00FDF# => romdata <= X"96A93F73";
    when 16#00FE0# => romdata <= X"B00C853D";
    when 16#00FE1# => romdata <= X"0D0481F1";
    when 16#00FE2# => romdata <= X"9051969B";
    when 16#00FE3# => romdata <= X"3F73B00C";
    when 16#00FE4# => romdata <= X"853D0D04";
    when 16#00FE5# => romdata <= X"FC3D0D81";
    when 16#00FE6# => romdata <= X"F5E0088C";
    when 16#00FE7# => romdata <= X"11087082";
    when 16#00FE8# => romdata <= X"2B83FFFC";
    when 16#00FE9# => romdata <= X"0681F19C";
    when 16#00FEA# => romdata <= X"54515555";
    when 16#00FEB# => romdata <= X"95F93F81";
    when 16#00FEC# => romdata <= X"F6940888";
    when 16#00FED# => romdata <= X"11087080";
    when 16#00FEE# => romdata <= X"C0078813";
    when 16#00FEF# => romdata <= X"0C545573";
    when 16#00FF0# => romdata <= X"52880A51";
    when 16#00FF1# => romdata <= X"FFADE43F";
    when 16#00FF2# => romdata <= X"B00881F6";
    when 16#00FF3# => romdata <= X"94088811";
    when 16#00FF4# => romdata <= X"0870FFBF";
    when 16#00FF5# => romdata <= X"0688130C";
    when 16#00FF6# => romdata <= X"555555B0";
    when 16#00FF7# => romdata <= X"08FE2E80";
    when 16#00FF8# => romdata <= X"C538B008";
    when 16#00FF9# => romdata <= X"FE249A38";
    when 16#00FFA# => romdata <= X"B008FD2E";
    when 16#00FFB# => romdata <= X"AB387451";
    when 16#00FFC# => romdata <= X"96FF3F81";
    when 16#00FFD# => romdata <= X"F1B05195";
    when 16#00FFE# => romdata <= X"AE3F74B0";
    when 16#00FFF# => romdata <= X"0C863D0D";
    when 16#01000# => romdata <= X"04B008FF";
    when 16#01001# => romdata <= X"2E098106";
    when 16#01002# => romdata <= X"E53881F1";
    when 16#01003# => romdata <= X"88519597";
    when 16#01004# => romdata <= X"3F74B00C";
    when 16#01005# => romdata <= X"863D0D04";
    when 16#01006# => romdata <= X"81F1C451";
    when 16#01007# => romdata <= X"95893F74";
    when 16#01008# => romdata <= X"B00C863D";
    when 16#01009# => romdata <= X"0D0481F1";
    when 16#0100A# => romdata <= X"D45194FB";
    when 16#0100B# => romdata <= X"3F74B00C";
    when 16#0100C# => romdata <= X"863D0D04";
    when 16#0100D# => romdata <= X"FE3D0D88";
    when 16#0100E# => romdata <= X"0A53840A";
    when 16#0100F# => romdata <= X"0B81F5E0";
    when 16#01010# => romdata <= X"088C1108";
    when 16#01011# => romdata <= X"51525280";
    when 16#01012# => romdata <= X"71279538";
    when 16#01013# => romdata <= X"80737084";
    when 16#01014# => romdata <= X"05550C80";
    when 16#01015# => romdata <= X"72708405";
    when 16#01016# => romdata <= X"540CFF11";
    when 16#01017# => romdata <= X"5170ED38";
    when 16#01018# => romdata <= X"800BB00C";
    when 16#01019# => romdata <= X"843D0D04";
    when 16#0101A# => romdata <= X"FD3D0D81";
    when 16#0101B# => romdata <= X"51FFA2D7";
    when 16#0101C# => romdata <= X"3FB00881";
    when 16#0101D# => romdata <= X"FF065473";
    when 16#0101E# => romdata <= X"802EA438";
    when 16#0101F# => romdata <= X"73842690";
    when 16#01020# => romdata <= X"3881F5E0";
    when 16#01021# => romdata <= X"0874710C";
    when 16#01022# => romdata <= X"5373B00C";
    when 16#01023# => romdata <= X"853D0D04";
    when 16#01024# => romdata <= X"81F5E008";
    when 16#01025# => romdata <= X"5380730C";
    when 16#01026# => romdata <= X"73B00C85";
    when 16#01027# => romdata <= X"3D0D0481";
    when 16#01028# => romdata <= X"F1E05194";
    when 16#01029# => romdata <= X"823F81F1";
    when 16#0102A# => romdata <= X"F05193FB";
    when 16#0102B# => romdata <= X"3F81F5E0";
    when 16#0102C# => romdata <= X"08700852";
    when 16#0102D# => romdata <= X"5395BA3F";
    when 16#0102E# => romdata <= X"81F28051";
    when 16#0102F# => romdata <= X"93E93F81";
    when 16#01030# => romdata <= X"F5E00884";
    when 16#01031# => romdata <= X"11085353";
    when 16#01032# => romdata <= X"A05193FE";
    when 16#01033# => romdata <= X"3F81F294";
    when 16#01034# => romdata <= X"5193D43F";
    when 16#01035# => romdata <= X"81F5E008";
    when 16#01036# => romdata <= X"88110853";
    when 16#01037# => romdata <= X"53A05193";
    when 16#01038# => romdata <= X"E93F81F2";
    when 16#01039# => romdata <= X"A85193BF";
    when 16#0103A# => romdata <= X"3F81F5E0";
    when 16#0103B# => romdata <= X"088C1108";
    when 16#0103C# => romdata <= X"525394FD";
    when 16#0103D# => romdata <= X"3F8A5193";
    when 16#0103E# => romdata <= X"943F73B0";
    when 16#0103F# => romdata <= X"0C853D0D";
    when 16#01040# => romdata <= X"04BC0802";
    when 16#01041# => romdata <= X"BC0CF93D";
    when 16#01042# => romdata <= X"0D02BC08";
    when 16#01043# => romdata <= X"FC050C88";
    when 16#01044# => romdata <= X"0A0BBC08";
    when 16#01045# => romdata <= X"F4050CFC";
    when 16#01046# => romdata <= X"3D0D823D";
    when 16#01047# => romdata <= X"BC08F005";
    when 16#01048# => romdata <= X"0C8151FF";
    when 16#01049# => romdata <= X"A1A13FB0";
    when 16#0104A# => romdata <= X"0881FF06";
    when 16#0104B# => romdata <= X"BC08F805";
    when 16#0104C# => romdata <= X"0C8251FF";
    when 16#0104D# => romdata <= X"A1913FB0";
    when 16#0104E# => romdata <= X"08BC08F0";
    when 16#0104F# => romdata <= X"05082383";
    when 16#01050# => romdata <= X"51FFA183";
    when 16#01051# => romdata <= X"3FB008BC";
    when 16#01052# => romdata <= X"08F00508";
    when 16#01053# => romdata <= X"82052384";
    when 16#01054# => romdata <= X"51FFA0F3";
    when 16#01055# => romdata <= X"3FB008BC";
    when 16#01056# => romdata <= X"08F00508";
    when 16#01057# => romdata <= X"84052385";
    when 16#01058# => romdata <= X"51FFA0E3";
    when 16#01059# => romdata <= X"3FB008BC";
    when 16#0105A# => romdata <= X"08F00508";
    when 16#0105B# => romdata <= X"86052386";
    when 16#0105C# => romdata <= X"51FFA0D3";
    when 16#0105D# => romdata <= X"3FB008BC";
    when 16#0105E# => romdata <= X"08F00508";
    when 16#0105F# => romdata <= X"88052387";
    when 16#01060# => romdata <= X"51FFA0C3";
    when 16#01061# => romdata <= X"3FB008BC";
    when 16#01062# => romdata <= X"08F00508";
    when 16#01063# => romdata <= X"8A052388";
    when 16#01064# => romdata <= X"51FFA0B3";
    when 16#01065# => romdata <= X"3FB008BC";
    when 16#01066# => romdata <= X"08F00508";
    when 16#01067# => romdata <= X"8C052389";
    when 16#01068# => romdata <= X"51FFA0A3";
    when 16#01069# => romdata <= X"3FB008BC";
    when 16#0106A# => romdata <= X"08F00508";
    when 16#0106B# => romdata <= X"8E052380";
    when 16#0106C# => romdata <= X"0B81F5E0";
    when 16#0106D# => romdata <= X"08708C05";
    when 16#0106E# => romdata <= X"0851BC08";
    when 16#0106F# => romdata <= X"E4050CBC";
    when 16#01070# => romdata <= X"08EC050C";
    when 16#01071# => romdata <= X"BC08EC05";
    when 16#01072# => romdata <= X"08BC08E4";
    when 16#01073# => romdata <= X"05082781";
    when 16#01074# => romdata <= X"8F38BC08";
    when 16#01075# => romdata <= X"E40508BC";
    when 16#01076# => romdata <= X"08E8050C";
    when 16#01077# => romdata <= X"BC08F805";
    when 16#01078# => romdata <= X"08802E81";
    when 16#01079# => romdata <= X"B638BC08";
    when 16#0107A# => romdata <= X"EC050810";
    when 16#0107B# => romdata <= X"BC08F005";
    when 16#0107C# => romdata <= X"08057022";
    when 16#0107D# => romdata <= X"BC08F405";
    when 16#0107E# => romdata <= X"08820522";
    when 16#0107F# => romdata <= X"71902B07";
    when 16#01080# => romdata <= X"BC08F405";
    when 16#01081# => romdata <= X"080CBC08";
    when 16#01082# => romdata <= X"E4050CBC";
    when 16#01083# => romdata <= X"08F8050C";
    when 16#01084# => romdata <= X"BC08EC05";
    when 16#01085# => romdata <= X"08810570";
    when 16#01086# => romdata <= X"81FF06BC";
    when 16#01087# => romdata <= X"08E4050C";
    when 16#01088# => romdata <= X"BC08F805";
    when 16#01089# => romdata <= X"0C860BBC";
    when 16#0108A# => romdata <= X"08EC0508";
    when 16#0108B# => romdata <= X"27883880";
    when 16#0108C# => romdata <= X"0BBC08E4";
    when 16#0108D# => romdata <= X"050CBC08";
    when 16#0108E# => romdata <= X"E40508BC";
    when 16#0108F# => romdata <= X"08F40508";
    when 16#01090# => romdata <= X"8405BC08";
    when 16#01091# => romdata <= X"E80508FF";
    when 16#01092# => romdata <= X"05BC08E8";
    when 16#01093# => romdata <= X"050CBC08";
    when 16#01094# => romdata <= X"F4050CBC";
    when 16#01095# => romdata <= X"08EC050C";
    when 16#01096# => romdata <= X"BC08E805";
    when 16#01097# => romdata <= X"08FF8738";
    when 16#01098# => romdata <= X"BC08FC05";
    when 16#01099# => romdata <= X"080D800B";
    when 16#0109A# => romdata <= X"B00C893D";
    when 16#0109B# => romdata <= X"0DBC0C04";
    when 16#0109C# => romdata <= X"BC08E405";
    when 16#0109D# => romdata <= X"08BC08F4";
    when 16#0109E# => romdata <= X"05088405";
    when 16#0109F# => romdata <= X"BC08E805";
    when 16#010A0# => romdata <= X"08FF05BC";
    when 16#010A1# => romdata <= X"08E8050C";
    when 16#010A2# => romdata <= X"BC08F405";
    when 16#010A3# => romdata <= X"0CBC08EC";
    when 16#010A4# => romdata <= X"050CBC08";
    when 16#010A5# => romdata <= X"E8050880";
    when 16#010A6# => romdata <= X"2EC638BC";
    when 16#010A7# => romdata <= X"08EC0508";
    when 16#010A8# => romdata <= X"10BC08F0";
    when 16#010A9# => romdata <= X"05080570";
    when 16#010AA# => romdata <= X"2270902B";
    when 16#010AB# => romdata <= X"BC08F405";
    when 16#010AC# => romdata <= X"0808FC80";
    when 16#010AD# => romdata <= X"80067190";
    when 16#010AE# => romdata <= X"2C07BC08";
    when 16#010AF# => romdata <= X"F405080C";
    when 16#010B0# => romdata <= X"52BC08E4";
    when 16#010B1# => romdata <= X"050CBC08";
    when 16#010B2# => romdata <= X"F8050C80";
    when 16#010B3# => romdata <= X"0BBC08E4";
    when 16#010B4# => romdata <= X"050CBC08";
    when 16#010B5# => romdata <= X"EC050886";
    when 16#010B6# => romdata <= X"26FF9538";
    when 16#010B7# => romdata <= X"BC08EC05";
    when 16#010B8# => romdata <= X"08810570";
    when 16#010B9# => romdata <= X"81FF06BC";
    when 16#010BA# => romdata <= X"08F40508";
    when 16#010BB# => romdata <= X"8405BC08";
    when 16#010BC# => romdata <= X"E80508FF";
    when 16#010BD# => romdata <= X"05BC08E8";
    when 16#010BE# => romdata <= X"050CBC08";
    when 16#010BF# => romdata <= X"F4050CBC";
    when 16#010C0# => romdata <= X"08EC050C";
    when 16#010C1# => romdata <= X"BC08E405";
    when 16#010C2# => romdata <= X"0CBC08E8";
    when 16#010C3# => romdata <= X"0508FF8B";
    when 16#010C4# => romdata <= X"38FECD39";
    when 16#010C5# => romdata <= X"F93D0D81";
    when 16#010C6# => romdata <= X"51FF9DAB";
    when 16#010C7# => romdata <= X"3FB00881";
    when 16#010C8# => romdata <= X"FF0681F2";
    when 16#010C9# => romdata <= X"B852578E";
    when 16#010CA# => romdata <= X"FE3F81F2";
    when 16#010CB# => romdata <= X"CC518EF7";
    when 16#010CC# => romdata <= X"3FF88080";
    when 16#010CD# => romdata <= X"9A805480";
    when 16#010CE# => romdata <= X"55737084";
    when 16#010CF# => romdata <= X"05550874";
    when 16#010D0# => romdata <= X"70840556";
    when 16#010D1# => romdata <= X"08545672";
    when 16#010D2# => romdata <= X"A0388115";
    when 16#010D3# => romdata <= X"7081FF06";
    when 16#010D4# => romdata <= X"56538775";
    when 16#010D5# => romdata <= X"27E33876";
    when 16#010D6# => romdata <= X"812E80C3";
    when 16#010D7# => romdata <= X"388A518E";
    when 16#010D8# => romdata <= X"AC3F76B0";
    when 16#010D9# => romdata <= X"0C893D0D";
    when 16#010DA# => romdata <= X"048A518E";
    when 16#010DB# => romdata <= X"A03F7251";
    when 16#010DC# => romdata <= X"8FFF3F8C";
    when 16#010DD# => romdata <= X"52B00851";
    when 16#010DE# => romdata <= X"D3BA3F81";
    when 16#010DF# => romdata <= X"F2E4518E";
    when 16#010E0# => romdata <= X"A63F7552";
    when 16#010E1# => romdata <= X"A0518EC2";
    when 16#010E2# => romdata <= X"3F7551D3";
    when 16#010E3# => romdata <= X"D13F8115";
    when 16#010E4# => romdata <= X"7081FF06";
    when 16#010E5# => romdata <= X"56538775";
    when 16#010E6# => romdata <= X"27FF9E38";
    when 16#010E7# => romdata <= X"FFB939F8";
    when 16#010E8# => romdata <= X"80809A80";
    when 16#010E9# => romdata <= X"54805380";
    when 16#010EA# => romdata <= X"74708405";
    when 16#010EB# => romdata <= X"560C8074";
    when 16#010EC# => romdata <= X"70840556";
    when 16#010ED# => romdata <= X"0C811370";
    when 16#010EE# => romdata <= X"81FF0654";
    when 16#010EF# => romdata <= X"55728726";
    when 16#010F0# => romdata <= X"FF9B3880";
    when 16#010F1# => romdata <= X"74708405";
    when 16#010F2# => romdata <= X"560C8074";
    when 16#010F3# => romdata <= X"70840556";
    when 16#010F4# => romdata <= X"0C811370";
    when 16#010F5# => romdata <= X"81FF0654";
    when 16#010F6# => romdata <= X"55877327";
    when 16#010F7# => romdata <= X"CA38FEFD";
    when 16#010F8# => romdata <= X"39FB3D0D";
    when 16#010F9# => romdata <= X"029F0533";
    when 16#010FA# => romdata <= X"79982B70";
    when 16#010FB# => romdata <= X"982C5154";
    when 16#010FC# => romdata <= X"55810A54";
    when 16#010FD# => romdata <= X"805672E8";
    when 16#010FE# => romdata <= X"25BD38E8";
    when 16#010FF# => romdata <= X"53751081";
    when 16#01100# => romdata <= X"07738180";
    when 16#01101# => romdata <= X"0A298180";
    when 16#01102# => romdata <= X"0A057098";
    when 16#01103# => romdata <= X"2C515456";
    when 16#01104# => romdata <= X"807324E9";
    when 16#01105# => romdata <= X"38807325";
    when 16#01106# => romdata <= X"80C73873";
    when 16#01107# => romdata <= X"812A810A";
    when 16#01108# => romdata <= X"07738180";
    when 16#01109# => romdata <= X"0A2981FF";
    when 16#0110A# => romdata <= X"0A057098";
    when 16#0110B# => romdata <= X"2C515454";
    when 16#0110C# => romdata <= X"728024E7";
    when 16#0110D# => romdata <= X"38AB3997";
    when 16#0110E# => romdata <= X"73259A38";
    when 16#0110F# => romdata <= X"9774812A";
    when 16#01110# => romdata <= X"810A0771";
    when 16#01111# => romdata <= X"81800A29";
    when 16#01112# => romdata <= X"81FF0A05";
    when 16#01113# => romdata <= X"70982C51";
    when 16#01114# => romdata <= X"525553DC";
    when 16#01115# => romdata <= X"39807324";
    when 16#01116# => romdata <= X"FFA33872";
    when 16#01117# => romdata <= X"8024FFBB";
    when 16#01118# => romdata <= X"38745280";
    when 16#01119# => romdata <= X"51FFB4D5";
    when 16#0111A# => romdata <= X"3F7381FF";
    when 16#0111B# => romdata <= X"0651FFB5";
    when 16#0111C# => romdata <= X"D23F7452";
    when 16#0111D# => romdata <= X"8151FFB4";
    when 16#0111E# => romdata <= X"C43F7388";
    when 16#0111F# => romdata <= X"2A7081FF";
    when 16#01120# => romdata <= X"065253FF";
    when 16#01121# => romdata <= X"B5BD3F74";
    when 16#01122# => romdata <= X"528251FF";
    when 16#01123# => romdata <= X"B4AF3F73";
    when 16#01124# => romdata <= X"902A7081";
    when 16#01125# => romdata <= X"FF065253";
    when 16#01126# => romdata <= X"FFB5A83F";
    when 16#01127# => romdata <= X"74528351";
    when 16#01128# => romdata <= X"FFB49A3F";
    when 16#01129# => romdata <= X"73982A51";
    when 16#0112A# => romdata <= X"FFB5983F";
    when 16#0112B# => romdata <= X"74528451";
    when 16#0112C# => romdata <= X"FFB48A3F";
    when 16#0112D# => romdata <= X"7581FF06";
    when 16#0112E# => romdata <= X"51FFB587";
    when 16#0112F# => romdata <= X"3F745285";
    when 16#01130# => romdata <= X"51FFB3F9";
    when 16#01131# => romdata <= X"3F75882A";
    when 16#01132# => romdata <= X"7081FF06";
    when 16#01133# => romdata <= X"5253FFB4";
    when 16#01134# => romdata <= X"F23F7452";
    when 16#01135# => romdata <= X"8651FFB3";
    when 16#01136# => romdata <= X"E43F7590";
    when 16#01137# => romdata <= X"2A7081FF";
    when 16#01138# => romdata <= X"065254FF";
    when 16#01139# => romdata <= X"B4DD3F74";
    when 16#0113A# => romdata <= X"528751FF";
    when 16#0113B# => romdata <= X"B3CF3F75";
    when 16#0113C# => romdata <= X"982A51FF";
    when 16#0113D# => romdata <= X"B4CD3F87";
    when 16#0113E# => romdata <= X"3D0D04F2";
    when 16#0113F# => romdata <= X"3D0D0280";
    when 16#01140# => romdata <= X"C3053302";
    when 16#01141# => romdata <= X"840580C7";
    when 16#01142# => romdata <= X"05338180";
    when 16#01143# => romdata <= X"0A712B98";
    when 16#01144# => romdata <= X"2A81F5E0";
    when 16#01145# => romdata <= X"088C1108";
    when 16#01146# => romdata <= X"71084453";
    when 16#01147# => romdata <= X"565C5557";
    when 16#01148# => romdata <= X"80730C80";
    when 16#01149# => romdata <= X"7071725C";
    when 16#0114A# => romdata <= X"5A5E5B80";
    when 16#0114B# => romdata <= X"56757A27";
    when 16#0114C# => romdata <= X"80D73881";
    when 16#0114D# => romdata <= X"772783CB";
    when 16#0114E# => romdata <= X"387783FF";
    when 16#0114F# => romdata <= X"FF068119";
    when 16#01150# => romdata <= X"71101084";
    when 16#01151# => romdata <= X"0A057930";
    when 16#01152# => romdata <= X"7A823270";
    when 16#01153# => romdata <= X"30728025";
    when 16#01154# => romdata <= X"71802507";
    when 16#01155# => romdata <= X"56585841";
    when 16#01156# => romdata <= X"57595C7B";
    when 16#01157# => romdata <= X"802E83D2";
    when 16#01158# => romdata <= X"38821522";
    when 16#01159# => romdata <= X"5372902B";
    when 16#0115A# => romdata <= X"70902C54";
    when 16#0115B# => romdata <= X"55727B25";
    when 16#0115C# => romdata <= X"8338725B";
    when 16#0115D# => romdata <= X"7C732583";
    when 16#0115E# => romdata <= X"38725D81";
    when 16#0115F# => romdata <= X"167081FF";
    when 16#01160# => romdata <= X"06575E79";
    when 16#01161# => romdata <= X"7626FFB1";
    when 16#01162# => romdata <= X"38811970";
    when 16#01163# => romdata <= X"81FF065A";
    when 16#01164# => romdata <= X"5680E579";
    when 16#01165# => romdata <= X"27FF9438";
    when 16#01166# => romdata <= X"987D3590";
    when 16#01167# => romdata <= X"2B70902C";
    when 16#01168# => romdata <= X"7C309871";
    when 16#01169# => romdata <= X"35902B70";
    when 16#0116A# => romdata <= X"902C5C5C";
    when 16#0116B# => romdata <= X"55565477";
    when 16#0116C# => romdata <= X"54777525";
    when 16#0116D# => romdata <= X"83387454";
    when 16#0116E# => romdata <= X"73902B70";
    when 16#0116F# => romdata <= X"902C5D55";
    when 16#01170# => romdata <= X"7B54807C";
    when 16#01171# => romdata <= X"2583D438";
    when 16#01172# => romdata <= X"73902B70";
    when 16#01173# => romdata <= X"902C5F56";
    when 16#01174# => romdata <= X"80705D58";
    when 16#01175# => romdata <= X"80705A56";
    when 16#01176# => romdata <= X"757A2780";
    when 16#01177# => romdata <= X"E4388177";
    when 16#01178# => romdata <= X"27838938";
    when 16#01179# => romdata <= X"7783FFFF";
    when 16#0117A# => romdata <= X"06811971";
    when 16#0117B# => romdata <= X"1010840A";
    when 16#0117C# => romdata <= X"0579307A";
    when 16#0117D# => romdata <= X"82327030";
    when 16#0117E# => romdata <= X"72802571";
    when 16#0117F# => romdata <= X"80250753";
    when 16#01180# => romdata <= X"51575357";
    when 16#01181# => romdata <= X"59547380";
    when 16#01182# => romdata <= X"2E83A138";
    when 16#01183# => romdata <= X"82152254";
    when 16#01184# => romdata <= X"73902B70";
    when 16#01185# => romdata <= X"902C719F";
    when 16#01186# => romdata <= X"2C707232";
    when 16#01187# => romdata <= X"7131799F";
    when 16#01188# => romdata <= X"2C707B32";
    when 16#01189# => romdata <= X"71315154";
    when 16#0118A# => romdata <= X"51565653";
    when 16#0118B# => romdata <= X"72742583";
    when 16#0118C# => romdata <= X"38745681";
    when 16#0118D# => romdata <= X"197081FF";
    when 16#0118E# => romdata <= X"065A5579";
    when 16#0118F# => romdata <= X"7926FFA4";
    when 16#01190# => romdata <= X"387D7635";
    when 16#01191# => romdata <= X"982B7098";
    when 16#01192# => romdata <= X"2C53547B";
    when 16#01193# => romdata <= X"51FB923F";
    when 16#01194# => romdata <= X"811C7081";
    when 16#01195# => romdata <= X"FF065D59";
    when 16#01196# => romdata <= X"80E57C27";
    when 16#01197# => romdata <= X"FEF63881";
    when 16#01198# => romdata <= X"F5E0087F";
    when 16#01199# => romdata <= X"710C5880";
    when 16#0119A# => romdata <= X"5281D684";
    when 16#0119B# => romdata <= X"51FFB4C3";
    when 16#0119C# => romdata <= X"3F829EBC";
    when 16#0119D# => romdata <= X"0880D2F7";
    when 16#0119E# => romdata <= X"0B829EBC";
    when 16#0119F# => romdata <= X"0C5F8052";
    when 16#011A0# => romdata <= X"8051FFB0";
    when 16#011A1# => romdata <= X"B83F81F2";
    when 16#011A2# => romdata <= X"EC51889B";
    when 16#011A3# => romdata <= X"3F7C5189";
    when 16#011A4# => romdata <= X"E03F8052";
    when 16#011A5# => romdata <= X"8751FFB0";
    when 16#011A6# => romdata <= X"A43F81F2";
    when 16#011A7# => romdata <= X"F4518887";
    when 16#011A8# => romdata <= X"3F7A5189";
    when 16#011A9# => romdata <= X"CC3F80D2";
    when 16#011AA# => romdata <= X"528051FF";
    when 16#011AB# => romdata <= X"B08F3F81";
    when 16#011AC# => romdata <= X"F2FC5187";
    when 16#011AD# => romdata <= X"F23F7651";
    when 16#011AE# => romdata <= X"89B73F80";
    when 16#011AF# => romdata <= X"C0528751";
    when 16#011B0# => romdata <= X"FFAFFA3F";
    when 16#011B1# => romdata <= X"81F38451";
    when 16#011B2# => romdata <= X"87DD3F79";
    when 16#011B3# => romdata <= X"80E62951";
    when 16#011B4# => romdata <= X"899F3F7E";
    when 16#011B5# => romdata <= X"829EBC0C";
    when 16#011B6# => romdata <= X"903D0D04";
    when 16#011B7# => romdata <= X"74225372";
    when 16#011B8# => romdata <= X"902B7090";
    when 16#011B9# => romdata <= X"2C545C72";
    when 16#011BA# => romdata <= X"7B258338";
    when 16#011BB# => romdata <= X"725B7C73";
    when 16#011BC# => romdata <= X"25833872";
    when 16#011BD# => romdata <= X"5D811670";
    when 16#011BE# => romdata <= X"81FF0657";
    when 16#011BF# => romdata <= X"5E757A27";
    when 16#011C0# => romdata <= X"FD873877";
    when 16#011C1# => romdata <= X"83FFFF06";
    when 16#011C2# => romdata <= X"81197110";
    when 16#011C3# => romdata <= X"10880A05";
    when 16#011C4# => romdata <= X"79307A82";
    when 16#011C5# => romdata <= X"32703072";
    when 16#011C6# => romdata <= X"80257180";
    when 16#011C7# => romdata <= X"25075658";
    when 16#011C8# => romdata <= X"40415759";
    when 16#011C9# => romdata <= X"5473802E";
    when 16#011CA# => romdata <= X"FFB23882";
    when 16#011CB# => romdata <= X"152253FF";
    when 16#011CC# => romdata <= X"AE397422";
    when 16#011CD# => romdata <= X"53FCAE39";
    when 16#011CE# => romdata <= X"74225473";
    when 16#011CF# => romdata <= X"902B7090";
    when 16#011D0# => romdata <= X"2C719F2C";
    when 16#011D1# => romdata <= X"70723271";
    when 16#011D2# => romdata <= X"31799F2C";
    when 16#011D3# => romdata <= X"707B3271";
    when 16#011D4# => romdata <= X"31515451";
    when 16#011D5# => romdata <= X"56565372";
    when 16#011D6# => romdata <= X"74258338";
    when 16#011D7# => romdata <= X"74568119";
    when 16#011D8# => romdata <= X"7081FF06";
    when 16#011D9# => romdata <= X"5A55787A";
    when 16#011DA# => romdata <= X"27FDD638";
    when 16#011DB# => romdata <= X"7783FFFF";
    when 16#011DC# => romdata <= X"06811971";
    when 16#011DD# => romdata <= X"1010880A";
    when 16#011DE# => romdata <= X"0579307A";
    when 16#011DF# => romdata <= X"82327030";
    when 16#011E0# => romdata <= X"72802571";
    when 16#011E1# => romdata <= X"80250753";
    when 16#011E2# => romdata <= X"51575357";
    when 16#011E3# => romdata <= X"59547380";
    when 16#011E4# => romdata <= X"2EFFA538";
    when 16#011E5# => romdata <= X"82152254";
    when 16#011E6# => romdata <= X"FFA13981";
    when 16#011E7# => romdata <= X"70902B70";
    when 16#011E8# => romdata <= X"902C4057";
    when 16#011E9# => romdata <= X"5480705D";
    when 16#011EA# => romdata <= X"58FCA939";
    when 16#011EB# => romdata <= X"742254FC";
    when 16#011EC# => romdata <= X"DF39FE3D";
    when 16#011ED# => romdata <= X"0D8151FF";
    when 16#011EE# => romdata <= X"948D3FB0";
    when 16#011EF# => romdata <= X"0881FF06";
    when 16#011F0# => romdata <= X"538251FF";
    when 16#011F1# => romdata <= X"94813FB0";
    when 16#011F2# => romdata <= X"0881FF06";
    when 16#011F3# => romdata <= X"527251FA";
    when 16#011F4# => romdata <= X"AA3F800B";
    when 16#011F5# => romdata <= X"B00C843D";
    when 16#011F6# => romdata <= X"0D04FD3D";
    when 16#011F7# => romdata <= X"0D81F68C";
    when 16#011F8# => romdata <= X"08841108";
    when 16#011F9# => romdata <= X"55538151";
    when 16#011FA# => romdata <= X"FF93DC3F";
    when 16#011FB# => romdata <= X"B00881FF";
    when 16#011FC# => romdata <= X"0674DFFF";
    when 16#011FD# => romdata <= X"FF065452";
    when 16#011FE# => romdata <= X"71802E87";
    when 16#011FF# => romdata <= X"3873A080";
    when 16#01200# => romdata <= X"80075382";
    when 16#01201# => romdata <= X"51FF93BF";
    when 16#01202# => romdata <= X"3FB00881";
    when 16#01203# => romdata <= X"FF0673EF";
    when 16#01204# => romdata <= X"FF0A0655";
    when 16#01205# => romdata <= X"5271802E";
    when 16#01206# => romdata <= X"87387290";
    when 16#01207# => romdata <= X"800A0754";
    when 16#01208# => romdata <= X"8351FF93";
    when 16#01209# => romdata <= X"A23FB008";
    when 16#0120A# => romdata <= X"81FF0674";
    when 16#0120B# => romdata <= X"F7FF0A06";
    when 16#0120C# => romdata <= X"54527180";
    when 16#0120D# => romdata <= X"2E873873";
    when 16#0120E# => romdata <= X"88800A07";
    when 16#0120F# => romdata <= X"538451FF";
    when 16#01210# => romdata <= X"93853FB0";
    when 16#01211# => romdata <= X"0881FF06";
    when 16#01212# => romdata <= X"73FBFF0A";
    when 16#01213# => romdata <= X"06555271";
    when 16#01214# => romdata <= X"802E8738";
    when 16#01215# => romdata <= X"7284800A";
    when 16#01216# => romdata <= X"07548551";
    when 16#01217# => romdata <= X"FF92E83F";
    when 16#01218# => romdata <= X"B00881FF";
    when 16#01219# => romdata <= X"0674FDFF";
    when 16#0121A# => romdata <= X"0A065452";
    when 16#0121B# => romdata <= X"71802E87";
    when 16#0121C# => romdata <= X"38738280";
    when 16#0121D# => romdata <= X"0A075381";
    when 16#0121E# => romdata <= X"F68C0873";
    when 16#0121F# => romdata <= X"84120C54";
    when 16#01220# => romdata <= X"72B00C85";
    when 16#01221# => romdata <= X"3D0D04FA";
    when 16#01222# => romdata <= X"3D0D880A";
    when 16#01223# => romdata <= X"0B81F5E0";
    when 16#01224# => romdata <= X"088C1108";
    when 16#01225# => romdata <= X"59555681";
    when 16#01226# => romdata <= X"51FF92AB";
    when 16#01227# => romdata <= X"3FB00890";
    when 16#01228# => romdata <= X"2B70902C";
    when 16#01229# => romdata <= X"56538077";
    when 16#0122A# => romdata <= X"27993880";
    when 16#0122B# => romdata <= X"77545473";
    when 16#0122C# => romdata <= X"83FFFF06";
    when 16#0122D# => romdata <= X"76708405";
    when 16#0122E# => romdata <= X"580CFF13";
    when 16#0122F# => romdata <= X"75155553";
    when 16#01230# => romdata <= X"72ED3880";
    when 16#01231# => romdata <= X"0BB00C88";
    when 16#01232# => romdata <= X"3D0D04FD";
    when 16#01233# => romdata <= X"3D0D0297";
    when 16#01234# => romdata <= X"053381F6";
    when 16#01235# => romdata <= X"8C088411";
    when 16#01236# => romdata <= X"0870B080";
    when 16#01237# => romdata <= X"0A0770EF";
    when 16#01238# => romdata <= X"FF0A0651";
    when 16#01239# => romdata <= X"54555552";
    when 16#0123A# => romdata <= X"71802E87";
    when 16#0123B# => romdata <= X"3872B080";
    when 16#0123C# => romdata <= X"0A075170";
    when 16#0123D# => romdata <= X"8E800A07";
    when 16#0123E# => romdata <= X"84150C85";
    when 16#0123F# => romdata <= X"3D0D04FF";
    when 16#01240# => romdata <= X"85F73F04";
    when 16#01241# => romdata <= X"FB3D0D77";
    when 16#01242# => romdata <= X"79555580";
    when 16#01243# => romdata <= X"56757524";
    when 16#01244# => romdata <= X"AB388074";
    when 16#01245# => romdata <= X"249D3880";
    when 16#01246# => romdata <= X"53735274";
    when 16#01247# => romdata <= X"5180E13F";
    when 16#01248# => romdata <= X"B0085475";
    when 16#01249# => romdata <= X"802E8538";
    when 16#0124A# => romdata <= X"B0083054";
    when 16#0124B# => romdata <= X"73B00C87";
    when 16#0124C# => romdata <= X"3D0D0473";
    when 16#0124D# => romdata <= X"30768132";
    when 16#0124E# => romdata <= X"5754DC39";
    when 16#0124F# => romdata <= X"74305581";
    when 16#01250# => romdata <= X"56738025";
    when 16#01251# => romdata <= X"D238EC39";
    when 16#01252# => romdata <= X"FA3D0D78";
    when 16#01253# => romdata <= X"7A575580";
    when 16#01254# => romdata <= X"57767524";
    when 16#01255# => romdata <= X"A438759F";
    when 16#01256# => romdata <= X"2C548153";
    when 16#01257# => romdata <= X"75743274";
    when 16#01258# => romdata <= X"31527451";
    when 16#01259# => romdata <= X"9B3FB008";
    when 16#0125A# => romdata <= X"5476802E";
    when 16#0125B# => romdata <= X"8538B008";
    when 16#0125C# => romdata <= X"305473B0";
    when 16#0125D# => romdata <= X"0C883D0D";
    when 16#0125E# => romdata <= X"04743055";
    when 16#0125F# => romdata <= X"8157D739";
    when 16#01260# => romdata <= X"FC3D0D76";
    when 16#01261# => romdata <= X"78535481";
    when 16#01262# => romdata <= X"53807473";
    when 16#01263# => romdata <= X"26525572";
    when 16#01264# => romdata <= X"802E9838";
    when 16#01265# => romdata <= X"70802EA9";
    when 16#01266# => romdata <= X"38807224";
    when 16#01267# => romdata <= X"A4387110";
    when 16#01268# => romdata <= X"73107572";
    when 16#01269# => romdata <= X"26535452";
    when 16#0126A# => romdata <= X"72EA3873";
    when 16#0126B# => romdata <= X"51788338";
    when 16#0126C# => romdata <= X"745170B0";
    when 16#0126D# => romdata <= X"0C863D0D";
    when 16#0126E# => romdata <= X"0472812A";
    when 16#0126F# => romdata <= X"72812A53";
    when 16#01270# => romdata <= X"5372802E";
    when 16#01271# => romdata <= X"E6387174";
    when 16#01272# => romdata <= X"26EF3873";
    when 16#01273# => romdata <= X"72317574";
    when 16#01274# => romdata <= X"0774812A";
    when 16#01275# => romdata <= X"74812A55";
    when 16#01276# => romdata <= X"555654E5";
    when 16#01277# => romdata <= X"39101010";
    when 16#01278# => romdata <= X"10101010";
    when 16#01279# => romdata <= X"10101010";
    when 16#0127A# => romdata <= X"10101010";
    when 16#0127B# => romdata <= X"10101010";
    when 16#0127C# => romdata <= X"10101010";
    when 16#0127D# => romdata <= X"10101010";
    when 16#0127E# => romdata <= X"10101010";
    when 16#0127F# => romdata <= X"53510473";
    when 16#01280# => romdata <= X"81FF0673";
    when 16#01281# => romdata <= X"83060981";
    when 16#01282# => romdata <= X"05830510";
    when 16#01283# => romdata <= X"10102B07";
    when 16#01284# => romdata <= X"72FC060C";
    when 16#01285# => romdata <= X"5151043C";
    when 16#01286# => romdata <= X"04727280";
    when 16#01287# => romdata <= X"728106FF";
    when 16#01288# => romdata <= X"05097206";
    when 16#01289# => romdata <= X"05711052";
    when 16#0128A# => romdata <= X"720A100A";
    when 16#0128B# => romdata <= X"5372ED38";
    when 16#0128C# => romdata <= X"51515351";
    when 16#0128D# => romdata <= X"04B008B4";
    when 16#0128E# => romdata <= X"08B80875";
    when 16#0128F# => romdata <= X"758192C8";
    when 16#01290# => romdata <= X"2D5050B0";
    when 16#01291# => romdata <= X"0856B80C";
    when 16#01292# => romdata <= X"B40CB00C";
    when 16#01293# => romdata <= X"5104B008";
    when 16#01294# => romdata <= X"B408B808";
    when 16#01295# => romdata <= X"75758192";
    when 16#01296# => romdata <= X"842D5050";
    when 16#01297# => romdata <= X"B00856B8";
    when 16#01298# => romdata <= X"0CB40CB0";
    when 16#01299# => romdata <= X"0C5104B0";
    when 16#0129A# => romdata <= X"08B408B8";
    when 16#0129B# => romdata <= X"0897D02D";
    when 16#0129C# => romdata <= X"B80CB40C";
    when 16#0129D# => romdata <= X"B00C04FF";
    when 16#0129E# => romdata <= X"3D0D028F";
    when 16#0129F# => romdata <= X"053381F6";
    when 16#012A0# => romdata <= X"9C085271";
    when 16#012A1# => romdata <= X"0C800BB0";
    when 16#012A2# => romdata <= X"0C833D0D";
    when 16#012A3# => romdata <= X"04FF3D0D";
    when 16#012A4# => romdata <= X"028F0533";
    when 16#012A5# => romdata <= X"51829EBC";
    when 16#012A6# => romdata <= X"0852712D";
    when 16#012A7# => romdata <= X"B00881FF";
    when 16#012A8# => romdata <= X"06B00C83";
    when 16#012A9# => romdata <= X"3D0D04FE";
    when 16#012AA# => romdata <= X"3D0D7470";
    when 16#012AB# => romdata <= X"33535371";
    when 16#012AC# => romdata <= X"802E9338";
    when 16#012AD# => romdata <= X"81137252";
    when 16#012AE# => romdata <= X"829EBC08";
    when 16#012AF# => romdata <= X"5353712D";
    when 16#012B0# => romdata <= X"72335271";
    when 16#012B1# => romdata <= X"EF38843D";
    when 16#012B2# => romdata <= X"0D04F43D";
    when 16#012B3# => romdata <= X"0D7F0284";
    when 16#012B4# => romdata <= X"05BB0533";
    when 16#012B5# => romdata <= X"5557880B";
    when 16#012B6# => romdata <= X"8C3D5B59";
    when 16#012B7# => romdata <= X"895381F3";
    when 16#012B8# => romdata <= X"B0527951";
    when 16#012B9# => romdata <= X"86D93F73";
    when 16#012BA# => romdata <= X"792E80FF";
    when 16#012BB# => romdata <= X"38785673";
    when 16#012BC# => romdata <= X"902E80EC";
    when 16#012BD# => romdata <= X"3802A705";
    when 16#012BE# => romdata <= X"58768F06";
    when 16#012BF# => romdata <= X"54738926";
    when 16#012C0# => romdata <= X"80C23875";
    when 16#012C1# => romdata <= X"18B01555";
    when 16#012C2# => romdata <= X"55737534";
    when 16#012C3# => romdata <= X"76842AFF";
    when 16#012C4# => romdata <= X"177081FF";
    when 16#012C5# => romdata <= X"06585557";
    when 16#012C6# => romdata <= X"75DF3878";
    when 16#012C7# => romdata <= X"1A557575";
    when 16#012C8# => romdata <= X"34797033";
    when 16#012C9# => romdata <= X"55557380";
    when 16#012CA# => romdata <= X"2E933881";
    when 16#012CB# => romdata <= X"15745282";
    when 16#012CC# => romdata <= X"9EBC0857";
    when 16#012CD# => romdata <= X"55752D74";
    when 16#012CE# => romdata <= X"335473EF";
    when 16#012CF# => romdata <= X"3878B00C";
    when 16#012D0# => romdata <= X"8E3D0D04";
    when 16#012D1# => romdata <= X"7518B715";
    when 16#012D2# => romdata <= X"55557375";
    when 16#012D3# => romdata <= X"3476842A";
    when 16#012D4# => romdata <= X"FF177081";
    when 16#012D5# => romdata <= X"FF065855";
    when 16#012D6# => romdata <= X"5775FF9D";
    when 16#012D7# => romdata <= X"38FFBC39";
    when 16#012D8# => romdata <= X"84705759";
    when 16#012D9# => romdata <= X"02A70558";
    when 16#012DA# => romdata <= X"FF8F3982";
    when 16#012DB# => romdata <= X"705759F4";
    when 16#012DC# => romdata <= X"39F13D0D";
    when 16#012DD# => romdata <= X"618D3D70";
    when 16#012DE# => romdata <= X"5B5C5A80";
    when 16#012DF# => romdata <= X"7A565776";
    when 16#012E0# => romdata <= X"7A248185";
    when 16#012E1# => romdata <= X"38781754";
    when 16#012E2# => romdata <= X"8A527451";
    when 16#012E3# => romdata <= X"84FF3FB0";
    when 16#012E4# => romdata <= X"08B00553";
    when 16#012E5# => romdata <= X"72743481";
    when 16#012E6# => romdata <= X"17578A52";
    when 16#012E7# => romdata <= X"745184C8";
    when 16#012E8# => romdata <= X"3FB00855";
    when 16#012E9# => romdata <= X"B008DE38";
    when 16#012EA# => romdata <= X"B008779F";
    when 16#012EB# => romdata <= X"2A187081";
    when 16#012EC# => romdata <= X"2C5A5656";
    when 16#012ED# => romdata <= X"8078259E";
    when 16#012EE# => romdata <= X"387817FF";
    when 16#012EF# => romdata <= X"05557519";
    when 16#012F0# => romdata <= X"70335553";
    when 16#012F1# => romdata <= X"74337334";
    when 16#012F2# => romdata <= X"73753481";
    when 16#012F3# => romdata <= X"16FF1656";
    when 16#012F4# => romdata <= X"56777624";
    when 16#012F5# => romdata <= X"E9387619";
    when 16#012F6# => romdata <= X"58807834";
    when 16#012F7# => romdata <= X"807A2417";
    when 16#012F8# => romdata <= X"7081FF06";
    when 16#012F9# => romdata <= X"7C703356";
    when 16#012FA# => romdata <= X"57555672";
    when 16#012FB# => romdata <= X"802E9338";
    when 16#012FC# => romdata <= X"81157352";
    when 16#012FD# => romdata <= X"829EBC08";
    when 16#012FE# => romdata <= X"5855762D";
    when 16#012FF# => romdata <= X"74335372";
    when 16#01300# => romdata <= X"EF3873B0";
    when 16#01301# => romdata <= X"0C913D0D";
    when 16#01302# => romdata <= X"04AD7B34";
    when 16#01303# => romdata <= X"02AD057A";
    when 16#01304# => romdata <= X"30711956";
    when 16#01305# => romdata <= X"56598A52";
    when 16#01306# => romdata <= X"745183F1";
    when 16#01307# => romdata <= X"3FB008B0";
    when 16#01308# => romdata <= X"05537274";
    when 16#01309# => romdata <= X"34811757";
    when 16#0130A# => romdata <= X"8A527451";
    when 16#0130B# => romdata <= X"83BA3FB0";
    when 16#0130C# => romdata <= X"0855B008";
    when 16#0130D# => romdata <= X"FECF38FE";
    when 16#0130E# => romdata <= X"EF39FD3D";
    when 16#0130F# => romdata <= X"0D81F690";
    when 16#01310# => romdata <= X"0876B2E4";
    when 16#01311# => romdata <= X"2994120C";
    when 16#01312# => romdata <= X"54850B98";
    when 16#01313# => romdata <= X"150C9814";
    when 16#01314# => romdata <= X"08708106";
    when 16#01315# => romdata <= X"515372F6";
    when 16#01316# => romdata <= X"38853D0D";
    when 16#01317# => romdata <= X"04803D0D";
    when 16#01318# => romdata <= X"81F69008";
    when 16#01319# => romdata <= X"51870B84";
    when 16#0131A# => romdata <= X"120CFF0B";
    when 16#0131B# => romdata <= X"A4120CA7";
    when 16#0131C# => romdata <= X"0BA8120C";
    when 16#0131D# => romdata <= X"B2E40B94";
    when 16#0131E# => romdata <= X"120C870B";
    when 16#0131F# => romdata <= X"98120C82";
    when 16#01320# => romdata <= X"3D0D0480";
    when 16#01321# => romdata <= X"3D0D81F6";
    when 16#01322# => romdata <= X"940851B8";
    when 16#01323# => romdata <= X"0B8C120C";
    when 16#01324# => romdata <= X"830B8812";
    when 16#01325# => romdata <= X"0C823D0D";
    when 16#01326# => romdata <= X"04803D0D";
    when 16#01327# => romdata <= X"81F69408";
    when 16#01328# => romdata <= X"84110881";
    when 16#01329# => romdata <= X"06B00C51";
    when 16#0132A# => romdata <= X"823D0D04";
    when 16#0132B# => romdata <= X"FF3D0D81";
    when 16#0132C# => romdata <= X"F6940852";
    when 16#0132D# => romdata <= X"84120870";
    when 16#0132E# => romdata <= X"81065151";
    when 16#0132F# => romdata <= X"70802EF4";
    when 16#01330# => romdata <= X"38710870";
    when 16#01331# => romdata <= X"81FF06B0";
    when 16#01332# => romdata <= X"0C51833D";
    when 16#01333# => romdata <= X"0D04FE3D";
    when 16#01334# => romdata <= X"0D029305";
    when 16#01335# => romdata <= X"3381F694";
    when 16#01336# => romdata <= X"08535384";
    when 16#01337# => romdata <= X"12087089";
    when 16#01338# => romdata <= X"2A708106";
    when 16#01339# => romdata <= X"51515170";
    when 16#0133A# => romdata <= X"F2387272";
    when 16#0133B# => romdata <= X"0C843D0D";
    when 16#0133C# => romdata <= X"04FE3D0D";
    when 16#0133D# => romdata <= X"02930533";
    when 16#0133E# => romdata <= X"53728A2E";
    when 16#0133F# => romdata <= X"9C3881F6";
    when 16#01340# => romdata <= X"94085284";
    when 16#01341# => romdata <= X"12087089";
    when 16#01342# => romdata <= X"2A708106";
    when 16#01343# => romdata <= X"51515170";
    when 16#01344# => romdata <= X"F2387272";
    when 16#01345# => romdata <= X"0C843D0D";
    when 16#01346# => romdata <= X"0481F694";
    when 16#01347# => romdata <= X"08528412";
    when 16#01348# => romdata <= X"0870892A";
    when 16#01349# => romdata <= X"70810651";
    when 16#0134A# => romdata <= X"515170F2";
    when 16#0134B# => romdata <= X"388D720C";
    when 16#0134C# => romdata <= X"84120870";
    when 16#0134D# => romdata <= X"892A7081";
    when 16#0134E# => romdata <= X"06515151";
    when 16#0134F# => romdata <= X"70C538D2";
    when 16#01350# => romdata <= X"39803D0D";
    when 16#01351# => romdata <= X"81F68808";
    when 16#01352# => romdata <= X"51800B84";
    when 16#01353# => romdata <= X"120C83FE";
    when 16#01354# => romdata <= X"800B8812";
    when 16#01355# => romdata <= X"0C800B82";
    when 16#01356# => romdata <= X"9EC03480";
    when 16#01357# => romdata <= X"0B829EC4";
    when 16#01358# => romdata <= X"34823D0D";
    when 16#01359# => romdata <= X"04FA3D0D";
    when 16#0135A# => romdata <= X"02A30533";
    when 16#0135B# => romdata <= X"81F68808";
    when 16#0135C# => romdata <= X"829EC033";
    when 16#0135D# => romdata <= X"7081FF06";
    when 16#0135E# => romdata <= X"70101011";
    when 16#0135F# => romdata <= X"829EC433";
    when 16#01360# => romdata <= X"7081FF06";
    when 16#01361# => romdata <= X"72902911";
    when 16#01362# => romdata <= X"70882B78";
    when 16#01363# => romdata <= X"07770C53";
    when 16#01364# => romdata <= X"5B5B5555";
    when 16#01365# => romdata <= X"59545473";
    when 16#01366# => romdata <= X"8A2E9838";
    when 16#01367# => romdata <= X"7480CF2E";
    when 16#01368# => romdata <= X"9238738C";
    when 16#01369# => romdata <= X"2EA43881";
    when 16#0136A# => romdata <= X"16537282";
    when 16#0136B# => romdata <= X"9EC43488";
    when 16#0136C# => romdata <= X"3D0D0471";
    when 16#0136D# => romdata <= X"A326A338";
    when 16#0136E# => romdata <= X"81175271";
    when 16#0136F# => romdata <= X"829EC034";
    when 16#01370# => romdata <= X"800B829E";
    when 16#01371# => romdata <= X"C434883D";
    when 16#01372# => romdata <= X"0D048052";
    when 16#01373# => romdata <= X"71882B73";
    when 16#01374# => romdata <= X"0C811252";
    when 16#01375# => romdata <= X"97907226";
    when 16#01376# => romdata <= X"F338800B";
    when 16#01377# => romdata <= X"829EC034";
    when 16#01378# => romdata <= X"800B829E";
    when 16#01379# => romdata <= X"C434DF39";
    when 16#0137A# => romdata <= X"BC0802BC";
    when 16#0137B# => romdata <= X"0CFD3D0D";
    when 16#0137C# => romdata <= X"8053BC08";
    when 16#0137D# => romdata <= X"8C050852";
    when 16#0137E# => romdata <= X"BC088805";
    when 16#0137F# => romdata <= X"0851F780";
    when 16#01380# => romdata <= X"3FB00870";
    when 16#01381# => romdata <= X"B00C5485";
    when 16#01382# => romdata <= X"3D0DBC0C";
    when 16#01383# => romdata <= X"04BC0802";
    when 16#01384# => romdata <= X"BC0CFD3D";
    when 16#01385# => romdata <= X"0D8153BC";
    when 16#01386# => romdata <= X"088C0508";
    when 16#01387# => romdata <= X"52BC0888";
    when 16#01388# => romdata <= X"050851F6";
    when 16#01389# => romdata <= X"DB3FB008";
    when 16#0138A# => romdata <= X"70B00C54";
    when 16#0138B# => romdata <= X"853D0DBC";
    when 16#0138C# => romdata <= X"0C04803D";
    when 16#0138D# => romdata <= X"0D865184";
    when 16#0138E# => romdata <= X"963F8151";
    when 16#0138F# => romdata <= X"A1D33FFC";
    when 16#01390# => romdata <= X"3D0D7670";
    when 16#01391# => romdata <= X"797B5555";
    when 16#01392# => romdata <= X"55558F72";
    when 16#01393# => romdata <= X"278C3872";
    when 16#01394# => romdata <= X"75078306";
    when 16#01395# => romdata <= X"5170802E";
    when 16#01396# => romdata <= X"A738FF12";
    when 16#01397# => romdata <= X"5271FF2E";
    when 16#01398# => romdata <= X"98387270";
    when 16#01399# => romdata <= X"81055433";
    when 16#0139A# => romdata <= X"74708105";
    when 16#0139B# => romdata <= X"5634FF12";
    when 16#0139C# => romdata <= X"5271FF2E";
    when 16#0139D# => romdata <= X"098106EA";
    when 16#0139E# => romdata <= X"3874B00C";
    when 16#0139F# => romdata <= X"863D0D04";
    when 16#013A0# => romdata <= X"74517270";
    when 16#013A1# => romdata <= X"84055408";
    when 16#013A2# => romdata <= X"71708405";
    when 16#013A3# => romdata <= X"530C7270";
    when 16#013A4# => romdata <= X"84055408";
    when 16#013A5# => romdata <= X"71708405";
    when 16#013A6# => romdata <= X"530C7270";
    when 16#013A7# => romdata <= X"84055408";
    when 16#013A8# => romdata <= X"71708405";
    when 16#013A9# => romdata <= X"530C7270";
    when 16#013AA# => romdata <= X"84055408";
    when 16#013AB# => romdata <= X"71708405";
    when 16#013AC# => romdata <= X"530CF012";
    when 16#013AD# => romdata <= X"52718F26";
    when 16#013AE# => romdata <= X"C9388372";
    when 16#013AF# => romdata <= X"27953872";
    when 16#013B0# => romdata <= X"70840554";
    when 16#013B1# => romdata <= X"08717084";
    when 16#013B2# => romdata <= X"05530CFC";
    when 16#013B3# => romdata <= X"12527183";
    when 16#013B4# => romdata <= X"26ED3870";
    when 16#013B5# => romdata <= X"54FF8339";
    when 16#013B6# => romdata <= X"FD3D0D75";
    when 16#013B7# => romdata <= X"5384D813";
    when 16#013B8# => romdata <= X"08802E8A";
    when 16#013B9# => romdata <= X"38805372";
    when 16#013BA# => romdata <= X"B00C853D";
    when 16#013BB# => romdata <= X"0D048180";
    when 16#013BC# => romdata <= X"5272518D";
    when 16#013BD# => romdata <= X"9B3FB008";
    when 16#013BE# => romdata <= X"84D8140C";
    when 16#013BF# => romdata <= X"FF53B008";
    when 16#013C0# => romdata <= X"802EE438";
    when 16#013C1# => romdata <= X"B008549F";
    when 16#013C2# => romdata <= X"53807470";
    when 16#013C3# => romdata <= X"8405560C";
    when 16#013C4# => romdata <= X"FF135380";
    when 16#013C5# => romdata <= X"7324CE38";
    when 16#013C6# => romdata <= X"80747084";
    when 16#013C7# => romdata <= X"05560CFF";
    when 16#013C8# => romdata <= X"13537280";
    when 16#013C9# => romdata <= X"25E338FF";
    when 16#013CA# => romdata <= X"BC39FD3D";
    when 16#013CB# => romdata <= X"0D757755";
    when 16#013CC# => romdata <= X"539F7427";
    when 16#013CD# => romdata <= X"8D389673";
    when 16#013CE# => romdata <= X"0CFF5271";
    when 16#013CF# => romdata <= X"B00C853D";
    when 16#013D0# => romdata <= X"0D0484D8";
    when 16#013D1# => romdata <= X"13085271";
    when 16#013D2# => romdata <= X"802E9338";
    when 16#013D3# => romdata <= X"73101012";
    when 16#013D4# => romdata <= X"70087972";
    when 16#013D5# => romdata <= X"0C515271";
    when 16#013D6# => romdata <= X"B00C853D";
    when 16#013D7# => romdata <= X"0D047251";
    when 16#013D8# => romdata <= X"FEF63FFF";
    when 16#013D9# => romdata <= X"52B008D3";
    when 16#013DA# => romdata <= X"3884D813";
    when 16#013DB# => romdata <= X"08741010";
    when 16#013DC# => romdata <= X"1170087A";
    when 16#013DD# => romdata <= X"720C5151";
    when 16#013DE# => romdata <= X"52DD39F9";
    when 16#013DF# => romdata <= X"3D0D797B";
    when 16#013E0# => romdata <= X"5856769F";
    when 16#013E1# => romdata <= X"2680E838";
    when 16#013E2# => romdata <= X"84D81608";
    when 16#013E3# => romdata <= X"5473802E";
    when 16#013E4# => romdata <= X"AA387610";
    when 16#013E5# => romdata <= X"10147008";
    when 16#013E6# => romdata <= X"55557380";
    when 16#013E7# => romdata <= X"2EBA3880";
    when 16#013E8# => romdata <= X"5873812E";
    when 16#013E9# => romdata <= X"8F3873FF";
    when 16#013EA# => romdata <= X"2EA33880";
    when 16#013EB# => romdata <= X"750C7651";
    when 16#013EC# => romdata <= X"732D8058";
    when 16#013ED# => romdata <= X"77B00C89";
    when 16#013EE# => romdata <= X"3D0D0475";
    when 16#013EF# => romdata <= X"51FE993F";
    when 16#013F0# => romdata <= X"FF58B008";
    when 16#013F1# => romdata <= X"EF3884D8";
    when 16#013F2# => romdata <= X"160854C6";
    when 16#013F3# => romdata <= X"3996760C";
    when 16#013F4# => romdata <= X"810BB00C";
    when 16#013F5# => romdata <= X"893D0D04";
    when 16#013F6# => romdata <= X"755181ED";
    when 16#013F7# => romdata <= X"3F7653B0";
    when 16#013F8# => romdata <= X"08527551";
    when 16#013F9# => romdata <= X"81AD3FB0";
    when 16#013FA# => romdata <= X"08B00C89";
    when 16#013FB# => romdata <= X"3D0D0496";
    when 16#013FC# => romdata <= X"760CFF0B";
    when 16#013FD# => romdata <= X"B00C893D";
    when 16#013FE# => romdata <= X"0D04FC3D";
    when 16#013FF# => romdata <= X"0D767856";
    when 16#01400# => romdata <= X"53FF5474";
    when 16#01401# => romdata <= X"9F26B138";
    when 16#01402# => romdata <= X"84D81308";
    when 16#01403# => romdata <= X"5271802E";
    when 16#01404# => romdata <= X"AE387410";
    when 16#01405# => romdata <= X"10127008";
    when 16#01406# => romdata <= X"53538154";
    when 16#01407# => romdata <= X"71802E98";
    when 16#01408# => romdata <= X"38825471";
    when 16#01409# => romdata <= X"FF2E9138";
    when 16#0140A# => romdata <= X"83547181";
    when 16#0140B# => romdata <= X"2E8A3880";
    when 16#0140C# => romdata <= X"730C7451";
    when 16#0140D# => romdata <= X"712D8054";
    when 16#0140E# => romdata <= X"73B00C86";
    when 16#0140F# => romdata <= X"3D0D0472";
    when 16#01410# => romdata <= X"51FD953F";
    when 16#01411# => romdata <= X"B008F138";
    when 16#01412# => romdata <= X"84D81308";
    when 16#01413# => romdata <= X"52C439FF";
    when 16#01414# => romdata <= X"3D0D7352";
    when 16#01415# => romdata <= X"81F6A008";
    when 16#01416# => romdata <= X"51FEA03F";
    when 16#01417# => romdata <= X"833D0D04";
    when 16#01418# => romdata <= X"FE3D0D75";
    when 16#01419# => romdata <= X"53745281";
    when 16#0141A# => romdata <= X"F6A00851";
    when 16#0141B# => romdata <= X"FDBC3F84";
    when 16#0141C# => romdata <= X"3D0D0480";
    when 16#0141D# => romdata <= X"3D0D81F6";
    when 16#0141E# => romdata <= X"A00851FC";
    when 16#0141F# => romdata <= X"DB3F823D";
    when 16#01420# => romdata <= X"0D04FF3D";
    when 16#01421# => romdata <= X"0D735281";
    when 16#01422# => romdata <= X"F6A00851";
    when 16#01423# => romdata <= X"FEEC3F83";
    when 16#01424# => romdata <= X"3D0D04FC";
    when 16#01425# => romdata <= X"3D0D800B";
    when 16#01426# => romdata <= X"829ECC0C";
    when 16#01427# => romdata <= X"78527751";
    when 16#01428# => romdata <= X"9CAA3FB0";
    when 16#01429# => romdata <= X"0854B008";
    when 16#0142A# => romdata <= X"FF2E8838";
    when 16#0142B# => romdata <= X"73B00C86";
    when 16#0142C# => romdata <= X"3D0D0482";
    when 16#0142D# => romdata <= X"9ECC0855";
    when 16#0142E# => romdata <= X"74802EF0";
    when 16#0142F# => romdata <= X"38767571";
    when 16#01430# => romdata <= X"0C5373B0";
    when 16#01431# => romdata <= X"0C863D0D";
    when 16#01432# => romdata <= X"049BFC3F";
    when 16#01433# => romdata <= X"04FC3D0D";
    when 16#01434# => romdata <= X"76707970";
    when 16#01435# => romdata <= X"73078306";
    when 16#01436# => romdata <= X"54545455";
    when 16#01437# => romdata <= X"7080C338";
    when 16#01438# => romdata <= X"71700870";
    when 16#01439# => romdata <= X"0970F7FB";
    when 16#0143A# => romdata <= X"FDFF1306";
    when 16#0143B# => romdata <= X"70F88482";
    when 16#0143C# => romdata <= X"81800651";
    when 16#0143D# => romdata <= X"51535354";
    when 16#0143E# => romdata <= X"70A63884";
    when 16#0143F# => romdata <= X"14727470";
    when 16#01440# => romdata <= X"8405560C";
    when 16#01441# => romdata <= X"70087009";
    when 16#01442# => romdata <= X"70F7FBFD";
    when 16#01443# => romdata <= X"FF130670";
    when 16#01444# => romdata <= X"F8848281";
    when 16#01445# => romdata <= X"80065151";
    when 16#01446# => romdata <= X"53535470";
    when 16#01447# => romdata <= X"802EDC38";
    when 16#01448# => romdata <= X"73527170";
    when 16#01449# => romdata <= X"81055333";
    when 16#0144A# => romdata <= X"51707370";
    when 16#0144B# => romdata <= X"81055534";
    when 16#0144C# => romdata <= X"70F03874";
    when 16#0144D# => romdata <= X"B00C863D";
    when 16#0144E# => romdata <= X"0D04FD3D";
    when 16#0144F# => romdata <= X"0D757071";
    when 16#01450# => romdata <= X"83065355";
    when 16#01451# => romdata <= X"5270B838";
    when 16#01452# => romdata <= X"71700870";
    when 16#01453# => romdata <= X"09F7FBFD";
    when 16#01454# => romdata <= X"FF120670";
    when 16#01455# => romdata <= X"F8848281";
    when 16#01456# => romdata <= X"80065151";
    when 16#01457# => romdata <= X"5253709D";
    when 16#01458# => romdata <= X"38841370";
    when 16#01459# => romdata <= X"087009F7";
    when 16#0145A# => romdata <= X"FBFDFF12";
    when 16#0145B# => romdata <= X"0670F884";
    when 16#0145C# => romdata <= X"82818006";
    when 16#0145D# => romdata <= X"51515253";
    when 16#0145E# => romdata <= X"70802EE5";
    when 16#0145F# => romdata <= X"38725271";
    when 16#01460# => romdata <= X"33517080";
    when 16#01461# => romdata <= X"2E8A3881";
    when 16#01462# => romdata <= X"12703352";
    when 16#01463# => romdata <= X"5270F838";
    when 16#01464# => romdata <= X"717431B0";
    when 16#01465# => romdata <= X"0C853D0D";
    when 16#01466# => romdata <= X"04FA3D0D";
    when 16#01467# => romdata <= X"787A7C70";
    when 16#01468# => romdata <= X"54555552";
    when 16#01469# => romdata <= X"72802E80";
    when 16#0146A# => romdata <= X"D9387174";
    when 16#0146B# => romdata <= X"07830651";
    when 16#0146C# => romdata <= X"70802E80";
    when 16#0146D# => romdata <= X"D438FF13";
    when 16#0146E# => romdata <= X"5372FF2E";
    when 16#0146F# => romdata <= X"B1387133";
    when 16#01470# => romdata <= X"74335651";
    when 16#01471# => romdata <= X"74712E09";
    when 16#01472# => romdata <= X"8106A938";
    when 16#01473# => romdata <= X"72802E81";
    when 16#01474# => romdata <= X"87387081";
    when 16#01475# => romdata <= X"FF065170";
    when 16#01476# => romdata <= X"802E80FC";
    when 16#01477# => romdata <= X"38811281";
    when 16#01478# => romdata <= X"15FF1555";
    when 16#01479# => romdata <= X"555272FF";
    when 16#0147A# => romdata <= X"2E098106";
    when 16#0147B# => romdata <= X"D1387133";
    when 16#0147C# => romdata <= X"74335651";
    when 16#0147D# => romdata <= X"7081FF06";
    when 16#0147E# => romdata <= X"7581FF06";
    when 16#0147F# => romdata <= X"71713151";
    when 16#01480# => romdata <= X"525270B0";
    when 16#01481# => romdata <= X"0C883D0D";
    when 16#01482# => romdata <= X"04717457";
    when 16#01483# => romdata <= X"55837327";
    when 16#01484# => romdata <= X"88387108";
    when 16#01485# => romdata <= X"74082E88";
    when 16#01486# => romdata <= X"38747655";
    when 16#01487# => romdata <= X"52FF9739";
    when 16#01488# => romdata <= X"FC135372";
    when 16#01489# => romdata <= X"802EB138";
    when 16#0148A# => romdata <= X"74087009";
    when 16#0148B# => romdata <= X"F7FBFDFF";
    when 16#0148C# => romdata <= X"120670F8";
    when 16#0148D# => romdata <= X"84828180";
    when 16#0148E# => romdata <= X"06515151";
    when 16#0148F# => romdata <= X"709A3884";
    when 16#01490# => romdata <= X"15841757";
    when 16#01491# => romdata <= X"55837327";
    when 16#01492# => romdata <= X"D0387408";
    when 16#01493# => romdata <= X"76082ED0";
    when 16#01494# => romdata <= X"38747655";
    when 16#01495# => romdata <= X"52FEDF39";
    when 16#01496# => romdata <= X"800BB00C";
    when 16#01497# => romdata <= X"883D0D04";
    when 16#01498# => romdata <= X"F33D0D60";
    when 16#01499# => romdata <= X"6264725A";
    when 16#0149A# => romdata <= X"5A5E5E80";
    when 16#0149B# => romdata <= X"5C767081";
    when 16#0149C# => romdata <= X"05583381";
    when 16#0149D# => romdata <= X"F3BD1133";
    when 16#0149E# => romdata <= X"70832A70";
    when 16#0149F# => romdata <= X"81065155";
    when 16#014A0# => romdata <= X"555672E9";
    when 16#014A1# => romdata <= X"3875AD2E";
    when 16#014A2# => romdata <= X"82883875";
    when 16#014A3# => romdata <= X"AB2E8284";
    when 16#014A4# => romdata <= X"38773070";
    when 16#014A5# => romdata <= X"79078025";
    when 16#014A6# => romdata <= X"79903270";
    when 16#014A7# => romdata <= X"30707207";
    when 16#014A8# => romdata <= X"80257307";
    when 16#014A9# => romdata <= X"53575751";
    when 16#014AA# => romdata <= X"5372802E";
    when 16#014AB# => romdata <= X"873875B0";
    when 16#014AC# => romdata <= X"2E81EB38";
    when 16#014AD# => romdata <= X"778A3888";
    when 16#014AE# => romdata <= X"5875B02E";
    when 16#014AF# => romdata <= X"83388A58";
    when 16#014B0# => romdata <= X"810A5A7B";
    when 16#014B1# => romdata <= X"8438FE0A";
    when 16#014B2# => romdata <= X"5A775279";
    when 16#014B3# => romdata <= X"51F6BE3F";
    when 16#014B4# => romdata <= X"B0087853";
    when 16#014B5# => romdata <= X"7A525BF6";
    when 16#014B6# => romdata <= X"8F3FB008";
    when 16#014B7# => romdata <= X"5A807081";
    when 16#014B8# => romdata <= X"F3BD1833";
    when 16#014B9# => romdata <= X"70822A70";
    when 16#014BA# => romdata <= X"81065156";
    when 16#014BB# => romdata <= X"565A5572";
    when 16#014BC# => romdata <= X"802E80C1";
    when 16#014BD# => romdata <= X"38D01656";
    when 16#014BE# => romdata <= X"75782580";
    when 16#014BF# => romdata <= X"D7388079";
    when 16#014C0# => romdata <= X"24757B26";
    when 16#014C1# => romdata <= X"07537293";
    when 16#014C2# => romdata <= X"38747A2E";
    when 16#014C3# => romdata <= X"80EB387A";
    when 16#014C4# => romdata <= X"762580ED";
    when 16#014C5# => romdata <= X"3872802E";
    when 16#014C6# => romdata <= X"80E738FF";
    when 16#014C7# => romdata <= X"77708105";
    when 16#014C8# => romdata <= X"59335759";
    when 16#014C9# => romdata <= X"81F3BD16";
    when 16#014CA# => romdata <= X"3370822A";
    when 16#014CB# => romdata <= X"70810651";
    when 16#014CC# => romdata <= X"545472C1";
    when 16#014CD# => romdata <= X"38738306";
    when 16#014CE# => romdata <= X"5372802E";
    when 16#014CF# => romdata <= X"97387381";
    when 16#014D0# => romdata <= X"06C91755";
    when 16#014D1# => romdata <= X"53728538";
    when 16#014D2# => romdata <= X"FFA91654";
    when 16#014D3# => romdata <= X"73567776";
    when 16#014D4# => romdata <= X"24FFAB38";
    when 16#014D5# => romdata <= X"80792480";
    when 16#014D6# => romdata <= X"F0387B80";
    when 16#014D7# => romdata <= X"2E843874";
    when 16#014D8# => romdata <= X"30557C80";
    when 16#014D9# => romdata <= X"2E8C38FF";
    when 16#014DA# => romdata <= X"17537883";
    when 16#014DB# => romdata <= X"387D5372";
    when 16#014DC# => romdata <= X"7D0C74B0";
    when 16#014DD# => romdata <= X"0C8F3D0D";
    when 16#014DE# => romdata <= X"04815375";
    when 16#014DF# => romdata <= X"7B24FF95";
    when 16#014E0# => romdata <= X"38817579";
    when 16#014E1# => romdata <= X"29177870";
    when 16#014E2# => romdata <= X"81055A33";
    when 16#014E3# => romdata <= X"585659FF";
    when 16#014E4# => romdata <= X"9339815C";
    when 16#014E5# => romdata <= X"76708105";
    when 16#014E6# => romdata <= X"583356FD";
    when 16#014E7# => romdata <= X"F4398077";
    when 16#014E8# => romdata <= X"33545472";
    when 16#014E9# => romdata <= X"80F82EB2";
    when 16#014EA# => romdata <= X"387280D8";
    when 16#014EB# => romdata <= X"32703070";
    when 16#014EC# => romdata <= X"80257607";
    when 16#014ED# => romdata <= X"51515372";
    when 16#014EE# => romdata <= X"802EFDF8";
    when 16#014EF# => romdata <= X"38811733";
    when 16#014F0# => romdata <= X"82185856";
    when 16#014F1# => romdata <= X"9058FDF8";
    when 16#014F2# => romdata <= X"39810A55";
    when 16#014F3# => romdata <= X"7B8438FE";
    when 16#014F4# => romdata <= X"0A557F53";
    when 16#014F5# => romdata <= X"A2730CFF";
    when 16#014F6# => romdata <= X"89398154";
    when 16#014F7# => romdata <= X"CC39FD3D";
    when 16#014F8# => romdata <= X"0D775476";
    when 16#014F9# => romdata <= X"53755281";
    when 16#014FA# => romdata <= X"F6A00851";
    when 16#014FB# => romdata <= X"FCF23F85";
    when 16#014FC# => romdata <= X"3D0D04F3";
    when 16#014FD# => romdata <= X"3D0D6062";
    when 16#014FE# => romdata <= X"64725A5A";
    when 16#014FF# => romdata <= X"5D5D805E";
    when 16#01500# => romdata <= X"76708105";
    when 16#01501# => romdata <= X"583381F3";
    when 16#01502# => romdata <= X"BD113370";
    when 16#01503# => romdata <= X"832A7081";
    when 16#01504# => romdata <= X"06515555";
    when 16#01505# => romdata <= X"5672E938";
    when 16#01506# => romdata <= X"75AD2E81";
    when 16#01507# => romdata <= X"FF3875AB";
    when 16#01508# => romdata <= X"2E81FB38";
    when 16#01509# => romdata <= X"77307079";
    when 16#0150A# => romdata <= X"07802579";
    when 16#0150B# => romdata <= X"90327030";
    when 16#0150C# => romdata <= X"70720780";
    when 16#0150D# => romdata <= X"25730753";
    when 16#0150E# => romdata <= X"57575153";
    when 16#0150F# => romdata <= X"72802E87";
    when 16#01510# => romdata <= X"3875B02E";
    when 16#01511# => romdata <= X"81E23877";
    when 16#01512# => romdata <= X"8A388858";
    when 16#01513# => romdata <= X"75B02E83";
    when 16#01514# => romdata <= X"388A5877";
    when 16#01515# => romdata <= X"52FF51F3";
    when 16#01516# => romdata <= X"8F3FB008";
    when 16#01517# => romdata <= X"78535AFF";
    when 16#01518# => romdata <= X"51F3AA3F";
    when 16#01519# => romdata <= X"B0085B80";
    when 16#0151A# => romdata <= X"705A5581";
    when 16#0151B# => romdata <= X"F3BD1633";
    when 16#0151C# => romdata <= X"70822A70";
    when 16#0151D# => romdata <= X"81065154";
    when 16#0151E# => romdata <= X"5472802E";
    when 16#0151F# => romdata <= X"80C138D0";
    when 16#01520# => romdata <= X"16567578";
    when 16#01521# => romdata <= X"2580D738";
    when 16#01522# => romdata <= X"80792475";
    when 16#01523# => romdata <= X"7B260753";
    when 16#01524# => romdata <= X"72933874";
    when 16#01525# => romdata <= X"7A2E80EB";
    when 16#01526# => romdata <= X"387A7625";
    when 16#01527# => romdata <= X"80ED3872";
    when 16#01528# => romdata <= X"802E80E7";
    when 16#01529# => romdata <= X"38FF7770";
    when 16#0152A# => romdata <= X"81055933";
    when 16#0152B# => romdata <= X"575981F3";
    when 16#0152C# => romdata <= X"BD163370";
    when 16#0152D# => romdata <= X"822A7081";
    when 16#0152E# => romdata <= X"06515454";
    when 16#0152F# => romdata <= X"72C13873";
    when 16#01530# => romdata <= X"83065372";
    when 16#01531# => romdata <= X"802E9738";
    when 16#01532# => romdata <= X"738106C9";
    when 16#01533# => romdata <= X"17555372";
    when 16#01534# => romdata <= X"8538FFA9";
    when 16#01535# => romdata <= X"16547356";
    when 16#01536# => romdata <= X"777624FF";
    when 16#01537# => romdata <= X"AB388079";
    when 16#01538# => romdata <= X"24818938";
    when 16#01539# => romdata <= X"7D802E84";
    when 16#0153A# => romdata <= X"38743055";
    when 16#0153B# => romdata <= X"7B802E8C";
    when 16#0153C# => romdata <= X"38FF1753";
    when 16#0153D# => romdata <= X"7883387C";
    when 16#0153E# => romdata <= X"53727C0C";
    when 16#0153F# => romdata <= X"74B00C8F";
    when 16#01540# => romdata <= X"3D0D0481";
    when 16#01541# => romdata <= X"53757B24";
    when 16#01542# => romdata <= X"FF953881";
    when 16#01543# => romdata <= X"75792917";
    when 16#01544# => romdata <= X"78708105";
    when 16#01545# => romdata <= X"5A335856";
    when 16#01546# => romdata <= X"59FF9339";
    when 16#01547# => romdata <= X"815E7670";
    when 16#01548# => romdata <= X"81055833";
    when 16#01549# => romdata <= X"56FDFD39";
    when 16#0154A# => romdata <= X"80773354";
    when 16#0154B# => romdata <= X"547280F8";
    when 16#0154C# => romdata <= X"2E80C338";
    when 16#0154D# => romdata <= X"7280D832";
    when 16#0154E# => romdata <= X"70307080";
    when 16#0154F# => romdata <= X"25760751";
    when 16#01550# => romdata <= X"51537280";
    when 16#01551# => romdata <= X"2EFE8038";
    when 16#01552# => romdata <= X"81173382";
    when 16#01553# => romdata <= X"18585690";
    when 16#01554# => romdata <= X"705358FF";
    when 16#01555# => romdata <= X"51F1913F";
    when 16#01556# => romdata <= X"B0087853";
    when 16#01557# => romdata <= X"5AFF51F1";
    when 16#01558# => romdata <= X"AC3FB008";
    when 16#01559# => romdata <= X"5B80705A";
    when 16#0155A# => romdata <= X"55FE8039";
    when 16#0155B# => romdata <= X"FF605455";
    when 16#0155C# => romdata <= X"A2730CFE";
    when 16#0155D# => romdata <= X"F7398154";
    when 16#0155E# => romdata <= X"FFBA39FD";
    when 16#0155F# => romdata <= X"3D0D7754";
    when 16#01560# => romdata <= X"76537552";
    when 16#01561# => romdata <= X"81F6A008";
    when 16#01562# => romdata <= X"51FCE83F";
    when 16#01563# => romdata <= X"853D0D04";
    when 16#01564# => romdata <= X"F33D0D7F";
    when 16#01565# => romdata <= X"618B1170";
    when 16#01566# => romdata <= X"F8065C55";
    when 16#01567# => romdata <= X"555E7296";
    when 16#01568# => romdata <= X"26833890";
    when 16#01569# => romdata <= X"59807924";
    when 16#0156A# => romdata <= X"747A2607";
    when 16#0156B# => romdata <= X"53805472";
    when 16#0156C# => romdata <= X"742E0981";
    when 16#0156D# => romdata <= X"0680CB38";
    when 16#0156E# => romdata <= X"7D518BCA";
    when 16#0156F# => romdata <= X"3F7883F7";
    when 16#01570# => romdata <= X"2680C638";
    when 16#01571# => romdata <= X"78832A70";
    when 16#01572# => romdata <= X"10101081";
    when 16#01573# => romdata <= X"FDDC058C";
    when 16#01574# => romdata <= X"11085959";
    when 16#01575# => romdata <= X"5A76782E";
    when 16#01576# => romdata <= X"83B03884";
    when 16#01577# => romdata <= X"1708FC06";
    when 16#01578# => romdata <= X"568C1708";
    when 16#01579# => romdata <= X"88180871";
    when 16#0157A# => romdata <= X"8C120C88";
    when 16#0157B# => romdata <= X"120C5875";
    when 16#0157C# => romdata <= X"17841108";
    when 16#0157D# => romdata <= X"81078412";
    when 16#0157E# => romdata <= X"0C537D51";
    when 16#0157F# => romdata <= X"8B893F88";
    when 16#01580# => romdata <= X"175473B0";
    when 16#01581# => romdata <= X"0C8F3D0D";
    when 16#01582# => romdata <= X"0478892A";
    when 16#01583# => romdata <= X"79832A5B";
    when 16#01584# => romdata <= X"5372802E";
    when 16#01585# => romdata <= X"BF387886";
    when 16#01586# => romdata <= X"2AB8055A";
    when 16#01587# => romdata <= X"847327B4";
    when 16#01588# => romdata <= X"3880DB13";
    when 16#01589# => romdata <= X"5A947327";
    when 16#0158A# => romdata <= X"AB38788C";
    when 16#0158B# => romdata <= X"2A80EE05";
    when 16#0158C# => romdata <= X"5A80D473";
    when 16#0158D# => romdata <= X"279E3878";
    when 16#0158E# => romdata <= X"8F2A80F7";
    when 16#0158F# => romdata <= X"055A82D4";
    when 16#01590# => romdata <= X"73279138";
    when 16#01591# => romdata <= X"78922A80";
    when 16#01592# => romdata <= X"FC055A8A";
    when 16#01593# => romdata <= X"D4732784";
    when 16#01594# => romdata <= X"3880FE5A";
    when 16#01595# => romdata <= X"79101010";
    when 16#01596# => romdata <= X"81FDDC05";
    when 16#01597# => romdata <= X"8C110858";
    when 16#01598# => romdata <= X"5576752E";
    when 16#01599# => romdata <= X"A3388417";
    when 16#0159A# => romdata <= X"08FC0670";
    when 16#0159B# => romdata <= X"7A315556";
    when 16#0159C# => romdata <= X"738F2488";
    when 16#0159D# => romdata <= X"D5387380";
    when 16#0159E# => romdata <= X"25FEE638";
    when 16#0159F# => romdata <= X"8C170857";
    when 16#015A0# => romdata <= X"76752E09";
    when 16#015A1# => romdata <= X"8106DF38";
    when 16#015A2# => romdata <= X"811A5A81";
    when 16#015A3# => romdata <= X"FDEC0857";
    when 16#015A4# => romdata <= X"7681FDE4";
    when 16#015A5# => romdata <= X"2E82C038";
    when 16#015A6# => romdata <= X"841708FC";
    when 16#015A7# => romdata <= X"06707A31";
    when 16#015A8# => romdata <= X"5556738F";
    when 16#015A9# => romdata <= X"2481F938";
    when 16#015AA# => romdata <= X"81FDE40B";
    when 16#015AB# => romdata <= X"81FDF00C";
    when 16#015AC# => romdata <= X"81FDE40B";
    when 16#015AD# => romdata <= X"81FDEC0C";
    when 16#015AE# => romdata <= X"738025FE";
    when 16#015AF# => romdata <= X"B23883FF";
    when 16#015B0# => romdata <= X"762783DF";
    when 16#015B1# => romdata <= X"3875892A";
    when 16#015B2# => romdata <= X"76832A55";
    when 16#015B3# => romdata <= X"5372802E";
    when 16#015B4# => romdata <= X"BF387586";
    when 16#015B5# => romdata <= X"2AB80554";
    when 16#015B6# => romdata <= X"847327B4";
    when 16#015B7# => romdata <= X"3880DB13";
    when 16#015B8# => romdata <= X"54947327";
    when 16#015B9# => romdata <= X"AB38758C";
    when 16#015BA# => romdata <= X"2A80EE05";
    when 16#015BB# => romdata <= X"5480D473";
    when 16#015BC# => romdata <= X"279E3875";
    when 16#015BD# => romdata <= X"8F2A80F7";
    when 16#015BE# => romdata <= X"055482D4";
    when 16#015BF# => romdata <= X"73279138";
    when 16#015C0# => romdata <= X"75922A80";
    when 16#015C1# => romdata <= X"FC05548A";
    when 16#015C2# => romdata <= X"D4732784";
    when 16#015C3# => romdata <= X"3880FE54";
    when 16#015C4# => romdata <= X"73101010";
    when 16#015C5# => romdata <= X"81FDDC05";
    when 16#015C6# => romdata <= X"88110856";
    when 16#015C7# => romdata <= X"5874782E";
    when 16#015C8# => romdata <= X"86CF3884";
    when 16#015C9# => romdata <= X"1508FC06";
    when 16#015CA# => romdata <= X"53757327";
    when 16#015CB# => romdata <= X"8D388815";
    when 16#015CC# => romdata <= X"08557478";
    when 16#015CD# => romdata <= X"2E098106";
    when 16#015CE# => romdata <= X"EA388C15";
    when 16#015CF# => romdata <= X"0881FDDC";
    when 16#015D0# => romdata <= X"0B840508";
    when 16#015D1# => romdata <= X"718C1A0C";
    when 16#015D2# => romdata <= X"76881A0C";
    when 16#015D3# => romdata <= X"7888130C";
    when 16#015D4# => romdata <= X"788C180C";
    when 16#015D5# => romdata <= X"5D587953";
    when 16#015D6# => romdata <= X"807A2483";
    when 16#015D7# => romdata <= X"E6387282";
    when 16#015D8# => romdata <= X"2C81712B";
    when 16#015D9# => romdata <= X"5C537A7C";
    when 16#015DA# => romdata <= X"26819838";
    when 16#015DB# => romdata <= X"7B7B0653";
    when 16#015DC# => romdata <= X"7282F138";
    when 16#015DD# => romdata <= X"79FC0684";
    when 16#015DE# => romdata <= X"055A7A10";
    when 16#015DF# => romdata <= X"707D0654";
    when 16#015E0# => romdata <= X"5B7282E0";
    when 16#015E1# => romdata <= X"38841A5A";
    when 16#015E2# => romdata <= X"F1398817";
    when 16#015E3# => romdata <= X"8C110858";
    when 16#015E4# => romdata <= X"5876782E";
    when 16#015E5# => romdata <= X"098106FC";
    when 16#015E6# => romdata <= X"C238821A";
    when 16#015E7# => romdata <= X"5AFDEC39";
    when 16#015E8# => romdata <= X"78177981";
    when 16#015E9# => romdata <= X"0784190C";
    when 16#015EA# => romdata <= X"7081FDF0";
    when 16#015EB# => romdata <= X"0C7081FD";
    when 16#015EC# => romdata <= X"EC0C81FD";
    when 16#015ED# => romdata <= X"E40B8C12";
    when 16#015EE# => romdata <= X"0C8C1108";
    when 16#015EF# => romdata <= X"88120C74";
    when 16#015F0# => romdata <= X"81078412";
    when 16#015F1# => romdata <= X"0C741175";
    when 16#015F2# => romdata <= X"710C5153";
    when 16#015F3# => romdata <= X"7D5187B7";
    when 16#015F4# => romdata <= X"3F881754";
    when 16#015F5# => romdata <= X"FCAC3981";
    when 16#015F6# => romdata <= X"FDDC0B84";
    when 16#015F7# => romdata <= X"05087A54";
    when 16#015F8# => romdata <= X"5C798025";
    when 16#015F9# => romdata <= X"FEF83882";
    when 16#015FA# => romdata <= X"DA397A09";
    when 16#015FB# => romdata <= X"7C067081";
    when 16#015FC# => romdata <= X"FDDC0B84";
    when 16#015FD# => romdata <= X"050C5C7A";
    when 16#015FE# => romdata <= X"105B7A7C";
    when 16#015FF# => romdata <= X"2685387A";
    when 16#01600# => romdata <= X"85B83881";
    when 16#01601# => romdata <= X"FDDC0B88";
    when 16#01602# => romdata <= X"05087084";
    when 16#01603# => romdata <= X"1208FC06";
    when 16#01604# => romdata <= X"707C317C";
    when 16#01605# => romdata <= X"72268F72";
    when 16#01606# => romdata <= X"25075757";
    when 16#01607# => romdata <= X"5C5D5572";
    when 16#01608# => romdata <= X"802E80DB";
    when 16#01609# => romdata <= X"38797A16";
    when 16#0160A# => romdata <= X"81FDD408";
    when 16#0160B# => romdata <= X"1B90115A";
    when 16#0160C# => romdata <= X"55575B81";
    when 16#0160D# => romdata <= X"FDD008FF";
    when 16#0160E# => romdata <= X"2E8838A0";
    when 16#0160F# => romdata <= X"8F13E080";
    when 16#01610# => romdata <= X"06577652";
    when 16#01611# => romdata <= X"7D5186C0";
    when 16#01612# => romdata <= X"3FB00854";
    when 16#01613# => romdata <= X"B008FF2E";
    when 16#01614# => romdata <= X"9038B008";
    when 16#01615# => romdata <= X"76278299";
    when 16#01616# => romdata <= X"387481FD";
    when 16#01617# => romdata <= X"DC2E8291";
    when 16#01618# => romdata <= X"3881FDDC";
    when 16#01619# => romdata <= X"0B880508";
    when 16#0161A# => romdata <= X"55841508";
    when 16#0161B# => romdata <= X"FC06707A";
    when 16#0161C# => romdata <= X"317A7226";
    when 16#0161D# => romdata <= X"8F722507";
    when 16#0161E# => romdata <= X"52555372";
    when 16#0161F# => romdata <= X"83E63874";
    when 16#01620# => romdata <= X"79810784";
    when 16#01621# => romdata <= X"170C7916";
    when 16#01622# => romdata <= X"7081FDDC";
    when 16#01623# => romdata <= X"0B88050C";
    when 16#01624# => romdata <= X"75810784";
    when 16#01625# => romdata <= X"120C547E";
    when 16#01626# => romdata <= X"525785EB";
    when 16#01627# => romdata <= X"3F881754";
    when 16#01628# => romdata <= X"FAE03975";
    when 16#01629# => romdata <= X"832A7054";
    when 16#0162A# => romdata <= X"54807424";
    when 16#0162B# => romdata <= X"819B3872";
    when 16#0162C# => romdata <= X"822C8171";
    when 16#0162D# => romdata <= X"2B81FDE0";
    when 16#0162E# => romdata <= X"08077081";
    when 16#0162F# => romdata <= X"FDDC0B84";
    when 16#01630# => romdata <= X"050C7510";
    when 16#01631# => romdata <= X"101081FD";
    when 16#01632# => romdata <= X"DC058811";
    when 16#01633# => romdata <= X"08585A5D";
    when 16#01634# => romdata <= X"53778C18";
    when 16#01635# => romdata <= X"0C748818";
    when 16#01636# => romdata <= X"0C768819";
    when 16#01637# => romdata <= X"0C768C16";
    when 16#01638# => romdata <= X"0CFCF339";
    when 16#01639# => romdata <= X"797A1010";
    when 16#0163A# => romdata <= X"1081FDDC";
    when 16#0163B# => romdata <= X"05705759";
    when 16#0163C# => romdata <= X"5D8C1508";
    when 16#0163D# => romdata <= X"5776752E";
    when 16#0163E# => romdata <= X"A3388417";
    when 16#0163F# => romdata <= X"08FC0670";
    when 16#01640# => romdata <= X"7A315556";
    when 16#01641# => romdata <= X"738F2483";
    when 16#01642# => romdata <= X"CA387380";
    when 16#01643# => romdata <= X"25848138";
    when 16#01644# => romdata <= X"8C170857";
    when 16#01645# => romdata <= X"76752E09";
    when 16#01646# => romdata <= X"8106DF38";
    when 16#01647# => romdata <= X"8815811B";
    when 16#01648# => romdata <= X"70830655";
    when 16#01649# => romdata <= X"5B5572C9";
    when 16#0164A# => romdata <= X"387C8306";
    when 16#0164B# => romdata <= X"5372802E";
    when 16#0164C# => romdata <= X"FDB838FF";
    when 16#0164D# => romdata <= X"1DF81959";
    when 16#0164E# => romdata <= X"5D881808";
    when 16#0164F# => romdata <= X"782EEA38";
    when 16#01650# => romdata <= X"FDB53983";
    when 16#01651# => romdata <= X"1A53FC96";
    when 16#01652# => romdata <= X"39831470";
    when 16#01653# => romdata <= X"822C8171";
    when 16#01654# => romdata <= X"2B81FDE0";
    when 16#01655# => romdata <= X"08077081";
    when 16#01656# => romdata <= X"FDDC0B84";
    when 16#01657# => romdata <= X"050C7610";
    when 16#01658# => romdata <= X"101081FD";
    when 16#01659# => romdata <= X"DC058811";
    when 16#0165A# => romdata <= X"08595B5E";
    when 16#0165B# => romdata <= X"5153FEE1";
    when 16#0165C# => romdata <= X"3981FDA0";
    when 16#0165D# => romdata <= X"081758B0";
    when 16#0165E# => romdata <= X"08762E81";
    when 16#0165F# => romdata <= X"8D3881FD";
    when 16#01660# => romdata <= X"D008FF2E";
    when 16#01661# => romdata <= X"83EC3873";
    when 16#01662# => romdata <= X"76311881";
    when 16#01663# => romdata <= X"FDA00C73";
    when 16#01664# => romdata <= X"87067057";
    when 16#01665# => romdata <= X"5372802E";
    when 16#01666# => romdata <= X"88388873";
    when 16#01667# => romdata <= X"31701555";
    when 16#01668# => romdata <= X"5676149F";
    when 16#01669# => romdata <= X"FF06A080";
    when 16#0166A# => romdata <= X"71311770";
    when 16#0166B# => romdata <= X"547F5357";
    when 16#0166C# => romdata <= X"5383D53F";
    when 16#0166D# => romdata <= X"B00853B0";
    when 16#0166E# => romdata <= X"08FF2E81";
    when 16#0166F# => romdata <= X"A03881FD";
    when 16#01670# => romdata <= X"A0081670";
    when 16#01671# => romdata <= X"81FDA00C";
    when 16#01672# => romdata <= X"747581FD";
    when 16#01673# => romdata <= X"DC0B8805";
    when 16#01674# => romdata <= X"0C747631";
    when 16#01675# => romdata <= X"18708107";
    when 16#01676# => romdata <= X"51555658";
    when 16#01677# => romdata <= X"7B81FDDC";
    when 16#01678# => romdata <= X"2E839C38";
    when 16#01679# => romdata <= X"798F2682";
    when 16#0167A# => romdata <= X"CB38810B";
    when 16#0167B# => romdata <= X"84150C84";
    when 16#0167C# => romdata <= X"1508FC06";
    when 16#0167D# => romdata <= X"707A317A";
    when 16#0167E# => romdata <= X"72268F72";
    when 16#0167F# => romdata <= X"25075255";
    when 16#01680# => romdata <= X"5372802E";
    when 16#01681# => romdata <= X"FCF93880";
    when 16#01682# => romdata <= X"DB39B008";
    when 16#01683# => romdata <= X"9FFF0653";
    when 16#01684# => romdata <= X"72FEEB38";
    when 16#01685# => romdata <= X"7781FDA0";
    when 16#01686# => romdata <= X"0C81FDDC";
    when 16#01687# => romdata <= X"0B880508";
    when 16#01688# => romdata <= X"7B188107";
    when 16#01689# => romdata <= X"84120C55";
    when 16#0168A# => romdata <= X"81FDCC08";
    when 16#0168B# => romdata <= X"78278638";
    when 16#0168C# => romdata <= X"7781FDCC";
    when 16#0168D# => romdata <= X"0C81FDC8";
    when 16#0168E# => romdata <= X"087827FC";
    when 16#0168F# => romdata <= X"AC387781";
    when 16#01690# => romdata <= X"FDC80C84";
    when 16#01691# => romdata <= X"1508FC06";
    when 16#01692# => romdata <= X"707A317A";
    when 16#01693# => romdata <= X"72268F72";
    when 16#01694# => romdata <= X"25075255";
    when 16#01695# => romdata <= X"5372802E";
    when 16#01696# => romdata <= X"FCA53888";
    when 16#01697# => romdata <= X"39807454";
    when 16#01698# => romdata <= X"56FEDB39";
    when 16#01699# => romdata <= X"7D51829F";
    when 16#0169A# => romdata <= X"3F800BB0";
    when 16#0169B# => romdata <= X"0C8F3D0D";
    when 16#0169C# => romdata <= X"04735380";
    when 16#0169D# => romdata <= X"7424A938";
    when 16#0169E# => romdata <= X"72822C81";
    when 16#0169F# => romdata <= X"712B81FD";
    when 16#016A0# => romdata <= X"E0080770";
    when 16#016A1# => romdata <= X"81FDDC0B";
    when 16#016A2# => romdata <= X"84050C5D";
    when 16#016A3# => romdata <= X"53778C18";
    when 16#016A4# => romdata <= X"0C748818";
    when 16#016A5# => romdata <= X"0C768819";
    when 16#016A6# => romdata <= X"0C768C16";
    when 16#016A7# => romdata <= X"0CF9B739";
    when 16#016A8# => romdata <= X"83147082";
    when 16#016A9# => romdata <= X"2C81712B";
    when 16#016AA# => romdata <= X"81FDE008";
    when 16#016AB# => romdata <= X"077081FD";
    when 16#016AC# => romdata <= X"DC0B8405";
    when 16#016AD# => romdata <= X"0C5E5153";
    when 16#016AE# => romdata <= X"D4397B7B";
    when 16#016AF# => romdata <= X"065372FC";
    when 16#016B0# => romdata <= X"A338841A";
    when 16#016B1# => romdata <= X"7B105C5A";
    when 16#016B2# => romdata <= X"F139FF1A";
    when 16#016B3# => romdata <= X"8111515A";
    when 16#016B4# => romdata <= X"F7B93978";
    when 16#016B5# => romdata <= X"17798107";
    when 16#016B6# => romdata <= X"84190C8C";
    when 16#016B7# => romdata <= X"18088819";
    when 16#016B8# => romdata <= X"08718C12";
    when 16#016B9# => romdata <= X"0C88120C";
    when 16#016BA# => romdata <= X"597081FD";
    when 16#016BB# => romdata <= X"F00C7081";
    when 16#016BC# => romdata <= X"FDEC0C81";
    when 16#016BD# => romdata <= X"FDE40B8C";
    when 16#016BE# => romdata <= X"120C8C11";
    when 16#016BF# => romdata <= X"0888120C";
    when 16#016C0# => romdata <= X"74810784";
    when 16#016C1# => romdata <= X"120C7411";
    when 16#016C2# => romdata <= X"75710C51";
    when 16#016C3# => romdata <= X"53F9BD39";
    when 16#016C4# => romdata <= X"75178411";
    when 16#016C5# => romdata <= X"08810784";
    when 16#016C6# => romdata <= X"120C538C";
    when 16#016C7# => romdata <= X"17088818";
    when 16#016C8# => romdata <= X"08718C12";
    when 16#016C9# => romdata <= X"0C88120C";
    when 16#016CA# => romdata <= X"587D5180";
    when 16#016CB# => romdata <= X"DA3F8817";
    when 16#016CC# => romdata <= X"54F5CF39";
    when 16#016CD# => romdata <= X"7284150C";
    when 16#016CE# => romdata <= X"F41AF806";
    when 16#016CF# => romdata <= X"70841E08";
    when 16#016D0# => romdata <= X"81060784";
    when 16#016D1# => romdata <= X"1E0C701D";
    when 16#016D2# => romdata <= X"545B850B";
    when 16#016D3# => romdata <= X"84140C85";
    when 16#016D4# => romdata <= X"0B88140C";
    when 16#016D5# => romdata <= X"8F7B27FD";
    when 16#016D6# => romdata <= X"CF38881C";
    when 16#016D7# => romdata <= X"527D5182";
    when 16#016D8# => romdata <= X"903F81FD";
    when 16#016D9# => romdata <= X"DC0B8805";
    when 16#016DA# => romdata <= X"0881FDA0";
    when 16#016DB# => romdata <= X"085955FD";
    when 16#016DC# => romdata <= X"B7397781";
    when 16#016DD# => romdata <= X"FDA00C73";
    when 16#016DE# => romdata <= X"81FDD00C";
    when 16#016DF# => romdata <= X"FC913972";
    when 16#016E0# => romdata <= X"84150CFD";
    when 16#016E1# => romdata <= X"A3390404";
    when 16#016E2# => romdata <= X"FD3D0D80";
    when 16#016E3# => romdata <= X"0B829ECC";
    when 16#016E4# => romdata <= X"0C765186";
    when 16#016E5# => romdata <= X"CB3FB008";
    when 16#016E6# => romdata <= X"53B008FF";
    when 16#016E7# => romdata <= X"2E883872";
    when 16#016E8# => romdata <= X"B00C853D";
    when 16#016E9# => romdata <= X"0D04829E";
    when 16#016EA# => romdata <= X"CC085473";
    when 16#016EB# => romdata <= X"802EF038";
    when 16#016EC# => romdata <= X"7574710C";
    when 16#016ED# => romdata <= X"5272B00C";
    when 16#016EE# => romdata <= X"853D0D04";
    when 16#016EF# => romdata <= X"FB3D0D77";
    when 16#016F0# => romdata <= X"705256C2";
    when 16#016F1# => romdata <= X"3F81FDDC";
    when 16#016F2# => romdata <= X"0B880508";
    when 16#016F3# => romdata <= X"841108FC";
    when 16#016F4# => romdata <= X"06707B31";
    when 16#016F5# => romdata <= X"9FEF05E0";
    when 16#016F6# => romdata <= X"8006E080";
    when 16#016F7# => romdata <= X"05565653";
    when 16#016F8# => romdata <= X"A0807424";
    when 16#016F9# => romdata <= X"94388052";
    when 16#016FA# => romdata <= X"7551FF9C";
    when 16#016FB# => romdata <= X"3F81FDE4";
    when 16#016FC# => romdata <= X"08155372";
    when 16#016FD# => romdata <= X"B0082E8F";
    when 16#016FE# => romdata <= X"387551FF";
    when 16#016FF# => romdata <= X"8A3F8053";
    when 16#01700# => romdata <= X"72B00C87";
    when 16#01701# => romdata <= X"3D0D0473";
    when 16#01702# => romdata <= X"30527551";
    when 16#01703# => romdata <= X"FEFA3FB0";
    when 16#01704# => romdata <= X"08FF2EA8";
    when 16#01705# => romdata <= X"3881FDDC";
    when 16#01706# => romdata <= X"0B880508";
    when 16#01707# => romdata <= X"75753181";
    when 16#01708# => romdata <= X"0784120C";
    when 16#01709# => romdata <= X"5381FDA0";
    when 16#0170A# => romdata <= X"08743181";
    when 16#0170B# => romdata <= X"FDA00C75";
    when 16#0170C# => romdata <= X"51FED43F";
    when 16#0170D# => romdata <= X"810BB00C";
    when 16#0170E# => romdata <= X"873D0D04";
    when 16#0170F# => romdata <= X"80527551";
    when 16#01710# => romdata <= X"FEC63F81";
    when 16#01711# => romdata <= X"FDDC0B88";
    when 16#01712# => romdata <= X"0508B008";
    when 16#01713# => romdata <= X"71315653";
    when 16#01714# => romdata <= X"8F7525FF";
    when 16#01715# => romdata <= X"A438B008";
    when 16#01716# => romdata <= X"81FDD008";
    when 16#01717# => romdata <= X"3181FDA0";
    when 16#01718# => romdata <= X"0C748107";
    when 16#01719# => romdata <= X"84140C75";
    when 16#0171A# => romdata <= X"51FE9C3F";
    when 16#0171B# => romdata <= X"8053FF90";
    when 16#0171C# => romdata <= X"39F63D0D";
    when 16#0171D# => romdata <= X"7C7E545B";
    when 16#0171E# => romdata <= X"72802E82";
    when 16#0171F# => romdata <= X"83387A51";
    when 16#01720# => romdata <= X"FE843FF8";
    when 16#01721# => romdata <= X"13841108";
    when 16#01722# => romdata <= X"70FE0670";
    when 16#01723# => romdata <= X"13841108";
    when 16#01724# => romdata <= X"FC065D58";
    when 16#01725# => romdata <= X"59545881";
    when 16#01726# => romdata <= X"FDE40875";
    when 16#01727# => romdata <= X"2E82DE38";
    when 16#01728# => romdata <= X"7884160C";
    when 16#01729# => romdata <= X"80738106";
    when 16#0172A# => romdata <= X"545A727A";
    when 16#0172B# => romdata <= X"2E81D538";
    when 16#0172C# => romdata <= X"78158411";
    when 16#0172D# => romdata <= X"08810651";
    when 16#0172E# => romdata <= X"5372A038";
    when 16#0172F# => romdata <= X"78175779";
    when 16#01730# => romdata <= X"81E63888";
    when 16#01731# => romdata <= X"15085372";
    when 16#01732# => romdata <= X"81FDE42E";
    when 16#01733# => romdata <= X"82F9388C";
    when 16#01734# => romdata <= X"1508708C";
    when 16#01735# => romdata <= X"150C7388";
    when 16#01736# => romdata <= X"120C5676";
    when 16#01737# => romdata <= X"81078419";
    when 16#01738# => romdata <= X"0C761877";
    when 16#01739# => romdata <= X"710C5379";
    when 16#0173A# => romdata <= X"81913883";
    when 16#0173B# => romdata <= X"FF772781";
    when 16#0173C# => romdata <= X"C8387689";
    when 16#0173D# => romdata <= X"2A77832A";
    when 16#0173E# => romdata <= X"56537280";
    when 16#0173F# => romdata <= X"2EBF3876";
    when 16#01740# => romdata <= X"862AB805";
    when 16#01741# => romdata <= X"55847327";
    when 16#01742# => romdata <= X"B43880DB";
    when 16#01743# => romdata <= X"13559473";
    when 16#01744# => romdata <= X"27AB3876";
    when 16#01745# => romdata <= X"8C2A80EE";
    when 16#01746# => romdata <= X"055580D4";
    when 16#01747# => romdata <= X"73279E38";
    when 16#01748# => romdata <= X"768F2A80";
    when 16#01749# => romdata <= X"F7055582";
    when 16#0174A# => romdata <= X"D4732791";
    when 16#0174B# => romdata <= X"3876922A";
    when 16#0174C# => romdata <= X"80FC0555";
    when 16#0174D# => romdata <= X"8AD47327";
    when 16#0174E# => romdata <= X"843880FE";
    when 16#0174F# => romdata <= X"55741010";
    when 16#01750# => romdata <= X"1081FDDC";
    when 16#01751# => romdata <= X"05881108";
    when 16#01752# => romdata <= X"55567376";
    when 16#01753# => romdata <= X"2E82B338";
    when 16#01754# => romdata <= X"841408FC";
    when 16#01755# => romdata <= X"06537673";
    when 16#01756# => romdata <= X"278D3888";
    when 16#01757# => romdata <= X"14085473";
    when 16#01758# => romdata <= X"762E0981";
    when 16#01759# => romdata <= X"06EA388C";
    when 16#0175A# => romdata <= X"1408708C";
    when 16#0175B# => romdata <= X"1A0C7488";
    when 16#0175C# => romdata <= X"1A0C7888";
    when 16#0175D# => romdata <= X"120C5677";
    when 16#0175E# => romdata <= X"8C150C7A";
    when 16#0175F# => romdata <= X"51FC883F";
    when 16#01760# => romdata <= X"8C3D0D04";
    when 16#01761# => romdata <= X"77087871";
    when 16#01762# => romdata <= X"31597705";
    when 16#01763# => romdata <= X"88190854";
    when 16#01764# => romdata <= X"577281FD";
    when 16#01765# => romdata <= X"E42E80E0";
    when 16#01766# => romdata <= X"388C1808";
    when 16#01767# => romdata <= X"708C150C";
    when 16#01768# => romdata <= X"7388120C";
    when 16#01769# => romdata <= X"56FE8939";
    when 16#0176A# => romdata <= X"8815088C";
    when 16#0176B# => romdata <= X"1608708C";
    when 16#0176C# => romdata <= X"130C5788";
    when 16#0176D# => romdata <= X"170CFEA3";
    when 16#0176E# => romdata <= X"3976832A";
    when 16#0176F# => romdata <= X"70545580";
    when 16#01770# => romdata <= X"75248198";
    when 16#01771# => romdata <= X"3872822C";
    when 16#01772# => romdata <= X"81712B81";
    when 16#01773# => romdata <= X"FDE00807";
    when 16#01774# => romdata <= X"81FDDC0B";
    when 16#01775# => romdata <= X"84050C53";
    when 16#01776# => romdata <= X"74101010";
    when 16#01777# => romdata <= X"81FDDC05";
    when 16#01778# => romdata <= X"88110855";
    when 16#01779# => romdata <= X"56758C19";
    when 16#0177A# => romdata <= X"0C738819";
    when 16#0177B# => romdata <= X"0C778817";
    when 16#0177C# => romdata <= X"0C778C15";
    when 16#0177D# => romdata <= X"0CFF8439";
    when 16#0177E# => romdata <= X"815AFDB4";
    when 16#0177F# => romdata <= X"39781773";
    when 16#01780# => romdata <= X"81065457";
    when 16#01781# => romdata <= X"72983877";
    when 16#01782# => romdata <= X"08787131";
    when 16#01783# => romdata <= X"5977058C";
    when 16#01784# => romdata <= X"1908881A";
    when 16#01785# => romdata <= X"08718C12";
    when 16#01786# => romdata <= X"0C88120C";
    when 16#01787# => romdata <= X"57577681";
    when 16#01788# => romdata <= X"0784190C";
    when 16#01789# => romdata <= X"7781FDDC";
    when 16#0178A# => romdata <= X"0B88050C";
    when 16#0178B# => romdata <= X"81FDD808";
    when 16#0178C# => romdata <= X"7726FEC7";
    when 16#0178D# => romdata <= X"3881FDD4";
    when 16#0178E# => romdata <= X"08527A51";
    when 16#0178F# => romdata <= X"FAFE3F7A";
    when 16#01790# => romdata <= X"51FAC43F";
    when 16#01791# => romdata <= X"FEBA3981";
    when 16#01792# => romdata <= X"788C150C";
    when 16#01793# => romdata <= X"7888150C";
    when 16#01794# => romdata <= X"738C1A0C";
    when 16#01795# => romdata <= X"73881A0C";
    when 16#01796# => romdata <= X"5AFD8039";
    when 16#01797# => romdata <= X"83157082";
    when 16#01798# => romdata <= X"2C81712B";
    when 16#01799# => romdata <= X"81FDE008";
    when 16#0179A# => romdata <= X"0781FDDC";
    when 16#0179B# => romdata <= X"0B84050C";
    when 16#0179C# => romdata <= X"51537410";
    when 16#0179D# => romdata <= X"101081FD";
    when 16#0179E# => romdata <= X"DC058811";
    when 16#0179F# => romdata <= X"085556FE";
    when 16#017A0# => romdata <= X"E4397453";
    when 16#017A1# => romdata <= X"807524A7";
    when 16#017A2# => romdata <= X"3872822C";
    when 16#017A3# => romdata <= X"81712B81";
    when 16#017A4# => romdata <= X"FDE00807";
    when 16#017A5# => romdata <= X"81FDDC0B";
    when 16#017A6# => romdata <= X"84050C53";
    when 16#017A7# => romdata <= X"758C190C";
    when 16#017A8# => romdata <= X"7388190C";
    when 16#017A9# => romdata <= X"7788170C";
    when 16#017AA# => romdata <= X"778C150C";
    when 16#017AB# => romdata <= X"FDCD3983";
    when 16#017AC# => romdata <= X"1570822C";
    when 16#017AD# => romdata <= X"81712B81";
    when 16#017AE# => romdata <= X"FDE00807";
    when 16#017AF# => romdata <= X"81FDDC0B";
    when 16#017B0# => romdata <= X"84050C51";
    when 16#017B1# => romdata <= X"53D63981";
    when 16#017B2# => romdata <= X"0BB00C04";
    when 16#017B3# => romdata <= X"803D0D72";
    when 16#017B4# => romdata <= X"812E8938";
    when 16#017B5# => romdata <= X"800BB00C";
    when 16#017B6# => romdata <= X"823D0D04";
    when 16#017B7# => romdata <= X"7351B23F";
    when 16#017B8# => romdata <= X"FE3D0D82";
    when 16#017B9# => romdata <= X"9EC80851";
    when 16#017BA# => romdata <= X"708A3882";
    when 16#017BB# => romdata <= X"9ED07082";
    when 16#017BC# => romdata <= X"9EC80C51";
    when 16#017BD# => romdata <= X"70751252";
    when 16#017BE# => romdata <= X"52FF5370";
    when 16#017BF# => romdata <= X"87FB8080";
    when 16#017C0# => romdata <= X"26883870";
    when 16#017C1# => romdata <= X"829EC80C";
    when 16#017C2# => romdata <= X"715372B0";
    when 16#017C3# => romdata <= X"0C843D0D";
    when 16#017C4# => romdata <= X"0400FF39";
    when 16#017C5# => romdata <= X"00000000";
    when 16#017C6# => romdata <= X"00000000";
    when 16#017C7# => romdata <= X"00000000";
    when 16#017C8# => romdata <= X"00000000";
    when 16#017C9# => romdata <= X"00CAC5CA";
    when 16#017CA# => romdata <= X"C5C0C0C0";
    when 16#017CB# => romdata <= X"C0C0C0C0";
    when 16#017CC# => romdata <= X"C0C0C0CF";
    when 16#017CD# => romdata <= X"CFCFCF00";
    when 16#017CE# => romdata <= X"00000F0F";
    when 16#017CF# => romdata <= X"0F0F8F8F";
    when 16#017D0# => romdata <= X"CFCFCFCF";
    when 16#017D1# => romdata <= X"CFCF4F0F";
    when 16#017D2# => romdata <= X"0F0F0000";
    when 16#017D3# => romdata <= X"CFCFCFCF";
    when 16#017D4# => romdata <= X"0F0F0F0F";
    when 16#017D5# => romdata <= X"0F0F0F0F";
    when 16#017D6# => romdata <= X"0F0FFEFE";
    when 16#017D7# => romdata <= X"FEFC0000";
    when 16#017D8# => romdata <= X"CFCFCFCF";
    when 16#017D9# => romdata <= X"CFCFCFCF";
    when 16#017DA# => romdata <= X"CFCFCFCF";
    when 16#017DB# => romdata <= X"CFFFFF7E";
    when 16#017DC# => romdata <= X"7E000000";
    when 16#017DD# => romdata <= X"00000000";
    when 16#017DE# => romdata <= X"00000000";
    when 16#017DF# => romdata <= X"00000000";
    when 16#017E0# => romdata <= X"00003F3F";
    when 16#017E1# => romdata <= X"3F3F0101";
    when 16#017E2# => romdata <= X"01010101";
    when 16#017E3# => romdata <= X"01010101";
    when 16#017E4# => romdata <= X"3F3F3F3F";
    when 16#017E5# => romdata <= X"0000383C";
    when 16#017E6# => romdata <= X"3E3E3F3F";
    when 16#017E7# => romdata <= X"3F3B3B39";
    when 16#017E8# => romdata <= X"39383838";
    when 16#017E9# => romdata <= X"38383800";
    when 16#017EA# => romdata <= X"003F3F3F";
    when 16#017EB# => romdata <= X"3F383838";
    when 16#017EC# => romdata <= X"38383838";
    when 16#017ED# => romdata <= X"38383C3F";
    when 16#017EE# => romdata <= X"3F1F0F00";
    when 16#017EF# => romdata <= X"003F3F3F";
    when 16#017F0# => romdata <= X"3F030303";
    when 16#017F1# => romdata <= X"03030303";
    when 16#017F2# => romdata <= X"03033F3F";
    when 16#017F3# => romdata <= X"3F3E0000";
    when 16#017F4# => romdata <= X"00000000";
    when 16#017F5# => romdata <= X"00000000";
    when 16#017F6# => romdata <= X"00000000";
    when 16#017F7# => romdata <= X"00000000";
    when 16#017F8# => romdata <= X"00000000";
    when 16#017F9# => romdata <= X"00000000";
    when 16#017FA# => romdata <= X"00000000";
    when 16#017FB# => romdata <= X"00000000";
    when 16#017FC# => romdata <= X"00000000";
    when 16#017FD# => romdata <= X"00000000";
    when 16#017FE# => romdata <= X"00000000";
    when 16#017FF# => romdata <= X"00000000";
    when 16#01800# => romdata <= X"00000000";
    when 16#01801# => romdata <= X"00000000";
    when 16#01802# => romdata <= X"00000000";
    when 16#01803# => romdata <= X"00000000";
    when 16#01804# => romdata <= X"00000000";
    when 16#01805# => romdata <= X"00000000";
    when 16#01806# => romdata <= X"00000000";
    when 16#01807# => romdata <= X"00000000";
    when 16#01808# => romdata <= X"00000000";
    when 16#01809# => romdata <= X"00000000";
    when 16#0180A# => romdata <= X"00000000";
    when 16#0180B# => romdata <= X"00000000";
    when 16#0180C# => romdata <= X"8080C0C0";
    when 16#0180D# => romdata <= X"E0E06000";
    when 16#0180E# => romdata <= X"00000000";
    when 16#0180F# => romdata <= X"00000000";
    when 16#01810# => romdata <= X"00000000";
    when 16#01811# => romdata <= X"00000000";
    when 16#01812# => romdata <= X"00000000";
    when 16#01813# => romdata <= X"00000000";
    when 16#01814# => romdata <= X"00000000";
    when 16#01815# => romdata <= X"00000000";
    when 16#01816# => romdata <= X"00000000";
    when 16#01817# => romdata <= X"00000000";
    when 16#01818# => romdata <= X"00000000";
    when 16#01819# => romdata <= X"00000000";
    when 16#0181A# => romdata <= X"00000000";
    when 16#0181B# => romdata <= X"00000000";
    when 16#0181C# => romdata <= X"00000000";
    when 16#0181D# => romdata <= X"00000000";
    when 16#0181E# => romdata <= X"00000000";
    when 16#0181F# => romdata <= X"00000000";
    when 16#01820# => romdata <= X"00000000";
    when 16#01821# => romdata <= X"00000000";
    when 16#01822# => romdata <= X"806098EE";
    when 16#01823# => romdata <= X"77BBDDEC";
    when 16#01824# => romdata <= X"EE6E0200";
    when 16#01825# => romdata <= X"00000000";
    when 16#01826# => romdata <= X"00E08080";
    when 16#01827# => romdata <= X"E00000E0";
    when 16#01828# => romdata <= X"A0A00000";
    when 16#01829# => romdata <= X"E0000000";
    when 16#0182A# => romdata <= X"00E0C000";
    when 16#0182B# => romdata <= X"C0E00000";
    when 16#0182C# => romdata <= X"E08080E0";
    when 16#0182D# => romdata <= X"0000C020";
    when 16#0182E# => romdata <= X"20C00000";
    when 16#0182F# => romdata <= X"E0000000";
    when 16#01830# => romdata <= X"20E02000";
    when 16#01831# => romdata <= X"0020A060";
    when 16#01832# => romdata <= X"20000000";
    when 16#01833# => romdata <= X"00000000";
    when 16#01834# => romdata <= X"00000000";
    when 16#01835# => romdata <= X"00000000";
    when 16#01836# => romdata <= X"00000000";
    when 16#01837# => romdata <= X"00000000";
    when 16#01838# => romdata <= X"00000000";
    when 16#01839# => romdata <= X"00030007";
    when 16#0183A# => romdata <= X"00070701";
    when 16#0183B# => romdata <= X"00000000";
    when 16#0183C# => romdata <= X"00000000";
    when 16#0183D# => romdata <= X"00000300";
    when 16#0183E# => romdata <= X"C0030000";
    when 16#0183F# => romdata <= X"034242C0";
    when 16#01840# => romdata <= X"00C34242";
    when 16#01841# => romdata <= X"0000C380";
    when 16#01842# => romdata <= X"01C00340";
    when 16#01843# => romdata <= X"C04300C0";
    when 16#01844# => romdata <= X"43408001";
    when 16#01845# => romdata <= X"C20201C0";
    when 16#01846# => romdata <= X"00C38202";
    when 16#01847# => romdata <= X"80C00300";
    when 16#01848# => romdata <= X"00C04342";
    when 16#01849# => romdata <= X"8202C040";
    when 16#0184A# => romdata <= X"40800000";
    when 16#0184B# => romdata <= X"C0404000";
    when 16#0184C# => romdata <= X"80404000";
    when 16#0184D# => romdata <= X"00C04040";
    when 16#0184E# => romdata <= X"8000C040";
    when 16#0184F# => romdata <= X"4000C080";
    when 16#01850# => romdata <= X"00C00000";
    when 16#01851# => romdata <= X"00000000";
    when 16#01852# => romdata <= X"00000000";
    when 16#01853# => romdata <= X"00000000";
    when 16#01854# => romdata <= X"00000000";
    when 16#01855# => romdata <= X"00FF0000";
    when 16#01856# => romdata <= X"0000C645";
    when 16#01857# => romdata <= X"44800785";
    when 16#01858# => romdata <= X"45408007";
    when 16#01859# => romdata <= X"80424700";
    when 16#0185A# => romdata <= X"80474000";
    when 16#0185B# => romdata <= X"07C14344";
    when 16#0185C# => romdata <= X"00C38404";
    when 16#0185D# => romdata <= X"C30007C1";
    when 16#0185E# => romdata <= X"42418700";
    when 16#0185F# => romdata <= X"80404784";
    when 16#01860# => romdata <= X"04C34047";
    when 16#01861# => romdata <= X"8101C640";
    when 16#01862# => romdata <= X"40070505";
    when 16#01863# => romdata <= X"00040502";
    when 16#01864# => romdata <= X"00000704";
    when 16#01865# => romdata <= X"04030007";
    when 16#01866# => romdata <= X"05050007";
    when 16#01867# => romdata <= X"00020700";
    when 16#01868# => romdata <= X"00000000";
    when 16#01869# => romdata <= X"00000000";
    when 16#0186A# => romdata <= X"00000000";
    when 16#0186B# => romdata <= X"00000000";
    when 16#0186C# => romdata <= X"0000FF00";
    when 16#0186D# => romdata <= X"00000007";
    when 16#0186E# => romdata <= X"01030500";
    when 16#0186F# => romdata <= X"03040403";
    when 16#01870# => romdata <= X"00040502";
    when 16#01871# => romdata <= X"00040502";
    when 16#01872# => romdata <= X"00000705";
    when 16#01873# => romdata <= X"05000700";
    when 16#01874# => romdata <= X"02070000";
    when 16#01875# => romdata <= X"07040403";
    when 16#01876# => romdata <= X"00030404";
    when 16#01877# => romdata <= X"03000701";
    when 16#01878# => romdata <= X"03050007";
    when 16#01879# => romdata <= X"01010000";
    when 16#0187A# => romdata <= X"00000000";
    when 16#0187B# => romdata <= X"00000000";
    when 16#0187C# => romdata <= X"00000000";
    when 16#0187D# => romdata <= X"00000000";
    when 16#0187E# => romdata <= X"00000000";
    when 16#0187F# => romdata <= X"71756974";
    when 16#01880# => romdata <= X"00000000";
    when 16#01881# => romdata <= X"68656C70";
    when 16#01882# => romdata <= X"00000000";
    when 16#01883# => romdata <= X"73686F77";
    when 16#01884# => romdata <= X"2042504D";
    when 16#01885# => romdata <= X"20726567";
    when 16#01886# => romdata <= X"69737465";
    when 16#01887# => romdata <= X"72730000";
    when 16#01888# => romdata <= X"62706D00";
    when 16#01889# => romdata <= X"73686F77";
    when 16#0188A# => romdata <= X"2044434D";
    when 16#0188B# => romdata <= X"20726567";
    when 16#0188C# => romdata <= X"69737465";
    when 16#0188D# => romdata <= X"72730000";
    when 16#0188E# => romdata <= X"64636D00";
    when 16#0188F# => romdata <= X"64696167";
    when 16#01890# => romdata <= X"6E6F7365";
    when 16#01891# => romdata <= X"206F7574";
    when 16#01892# => romdata <= X"70757420";
    when 16#01893# => romdata <= X"2B206D6F";
    when 16#01894# => romdata <= X"64652028";
    when 16#01895# => romdata <= X"302D3320";
    when 16#01896# => romdata <= X"73756D20";
    when 16#01897# => romdata <= X"48205629";
    when 16#01898# => romdata <= X"00000000";
    when 16#01899# => romdata <= X"73656C65";
    when 16#0189A# => romdata <= X"63740000";
    when 16#0189B# => romdata <= X"73797374";
    when 16#0189C# => romdata <= X"656D2072";
    when 16#0189D# => romdata <= X"65736574";
    when 16#0189E# => romdata <= X"00000000";
    when 16#0189F# => romdata <= X"72657365";
    when 16#018A0# => romdata <= X"74000000";
    when 16#018A1# => romdata <= X"73686F77";
    when 16#018A2# => romdata <= X"20737973";
    when 16#018A3# => romdata <= X"74656D20";
    when 16#018A4# => romdata <= X"696E666F";
    when 16#018A5# => romdata <= X"203C7665";
    when 16#018A6# => romdata <= X"72626F73";
    when 16#018A7# => romdata <= X"653E0000";
    when 16#018A8# => romdata <= X"73797369";
    when 16#018A9# => romdata <= X"6E666F00";
    when 16#018AA# => romdata <= X"3C6C6F77";
    when 16#018AB# => romdata <= X"65723E20";
    when 16#018AC# => romdata <= X"3C757070";
    when 16#018AD# => romdata <= X"65723E20";
    when 16#018AE# => romdata <= X"73657220";
    when 16#018AF# => romdata <= X"44434D20";
    when 16#018B0# => romdata <= X"626F756E";
    when 16#018B1# => romdata <= X"64730000";
    when 16#018B2# => romdata <= X"73686F77";
    when 16#018B3# => romdata <= X"2F736574";
    when 16#018B4# => romdata <= X"20646562";
    when 16#018B5# => romdata <= X"75672072";
    when 16#018B6# => romdata <= X"65676973";
    when 16#018B7# => romdata <= X"74657273";
    when 16#018B8# => romdata <= X"203C7365";
    when 16#018B9# => romdata <= X"74206D6F";
    when 16#018BA# => romdata <= X"64653E00";
    when 16#018BB# => romdata <= X"64656275";
    when 16#018BC# => romdata <= X"67000000";
    when 16#018BD# => romdata <= X"736F7572";
    when 16#018BE# => romdata <= X"63653A20";
    when 16#018BF# => romdata <= X"2030203D";
    when 16#018C0# => romdata <= X"20696E74";
    when 16#018C1# => romdata <= X"2C203120";
    when 16#018C2# => romdata <= X"3D206578";
    when 16#018C3# => romdata <= X"74000000";
    when 16#018C4# => romdata <= X"636C6B00";
    when 16#018C5# => romdata <= X"70756C73";
    when 16#018C6# => romdata <= X"6520736F";
    when 16#018C7# => romdata <= X"75726365";
    when 16#018C8# => romdata <= X"3A203020";
    when 16#018C9# => romdata <= X"3D207465";
    when 16#018CA# => romdata <= X"73746765";
    when 16#018CB# => romdata <= X"6E2C2031";
    when 16#018CC# => romdata <= X"203D2065";
    when 16#018CD# => romdata <= X"78740000";
    when 16#018CE# => romdata <= X"6D696372";
    when 16#018CF# => romdata <= X"6F000000";
    when 16#018D0# => romdata <= X"74657374";
    when 16#018D1# => romdata <= X"67656E65";
    when 16#018D2# => romdata <= X"7261746F";
    when 16#018D3# => romdata <= X"72203C73";
    when 16#018D4# => romdata <= X"63616C65";
    when 16#018D5# => romdata <= X"723E203C";
    when 16#018D6# => romdata <= X"72657374";
    when 16#018D7# => romdata <= X"6172743E";
    when 16#018D8# => romdata <= X"00000000";
    when 16#018D9# => romdata <= X"74657374";
    when 16#018DA# => romdata <= X"67656E00";
    when 16#018DB# => romdata <= X"3C6D7574";
    when 16#018DC# => romdata <= X"655F6E3E";
    when 16#018DD# => romdata <= X"203C7273";
    when 16#018DE# => romdata <= X"745F6E3E";
    when 16#018DF# => romdata <= X"203C6270";
    when 16#018E0# => romdata <= X"625F6E3E";
    when 16#018E1# => romdata <= X"203C6F73";
    when 16#018E2# => romdata <= X"72313E20";
    when 16#018E3# => romdata <= X"3C6F7372";
    when 16#018E4# => romdata <= X"323E0000";
    when 16#018E5# => romdata <= X"64616363";
    when 16#018E6# => romdata <= X"6F6E6600";
    when 16#018E7# => romdata <= X"3C6D756C";
    when 16#018E8# => romdata <= X"7469706C";
    when 16#018E9# => romdata <= X"6965723E";
    when 16#018EA# => romdata <= X"20696E69";
    when 16#018EB# => romdata <= X"7469616C";
    when 16#018EC# => romdata <= X"697A6520";
    when 16#018ED# => romdata <= X"62756666";
    when 16#018EE# => romdata <= X"65720000";
    when 16#018EF# => romdata <= X"64616374";
    when 16#018F0# => romdata <= X"65737400";
    when 16#018F1# => romdata <= X"72657365";
    when 16#018F2# => romdata <= X"74204250";
    when 16#018F3# => romdata <= X"4D206361";
    when 16#018F4# => romdata <= X"6C63756C";
    when 16#018F5# => romdata <= X"6174696F";
    when 16#018F6# => romdata <= X"6E206572";
    when 16#018F7# => romdata <= X"726F7273";
    when 16#018F8# => romdata <= X"00000000";
    when 16#018F9# => romdata <= X"62706D72";
    when 16#018FA# => romdata <= X"65730000";
    when 16#018FB# => romdata <= X"72657365";
    when 16#018FC# => romdata <= X"74204443";
    when 16#018FD# => romdata <= X"4D206572";
    when 16#018FE# => romdata <= X"726F7273";
    when 16#018FF# => romdata <= X"00000000";
    when 16#01900# => romdata <= X"64636D72";
    when 16#01901# => romdata <= X"65730000";
    when 16#01902# => romdata <= X"73686F77";
    when 16#01903# => romdata <= X"20646562";
    when 16#01904# => romdata <= X"75672062";
    when 16#01905# => romdata <= X"75666665";
    when 16#01906# => romdata <= X"72203C6C";
    when 16#01907# => romdata <= X"656E6774";
    when 16#01908# => romdata <= X"683E0000";
    when 16#01909# => romdata <= X"636C6561";
    when 16#0190A# => romdata <= X"72206465";
    when 16#0190B# => romdata <= X"62756720";
    when 16#0190C# => romdata <= X"62756666";
    when 16#0190D# => romdata <= X"65720000";
    when 16#0190E# => romdata <= X"62636C65";
    when 16#0190F# => romdata <= X"61720000";
    when 16#01910# => romdata <= X"646F776E";
    when 16#01911# => romdata <= X"6C6F6164";
    when 16#01912# => romdata <= X"20646562";
    when 16#01913# => romdata <= X"75672062";
    when 16#01914# => romdata <= X"75666665";
    when 16#01915# => romdata <= X"72202878";
    when 16#01916# => romdata <= X"6D6F6465";
    when 16#01917# => romdata <= X"6D290000";
    when 16#01918# => romdata <= X"62726561";
    when 16#01919# => romdata <= X"64000000";
    when 16#0191A# => romdata <= X"75706C6F";
    when 16#0191B# => romdata <= X"61642064";
    when 16#0191C# => romdata <= X"65627567";
    when 16#0191D# => romdata <= X"20627566";
    when 16#0191E# => romdata <= X"66657220";
    when 16#0191F# => romdata <= X"28786D6F";
    when 16#01920# => romdata <= X"64656D29";
    when 16#01921# => romdata <= X"00000000";
    when 16#01922# => romdata <= X"62777269";
    when 16#01923# => romdata <= X"74650000";
    when 16#01924# => romdata <= X"62756666";
    when 16#01925# => romdata <= X"6572206F";
    when 16#01926# => romdata <= X"6E204C43";
    when 16#01927# => romdata <= X"44203C63";
    when 16#01928# => romdata <= X"683E203C";
    when 16#01929# => romdata <= X"636F6D62";
    when 16#0192A# => romdata <= X"3E000000";
    when 16#0192B# => romdata <= X"73636F70";
    when 16#0192C# => romdata <= X"65000000";
    when 16#0192D# => romdata <= X"64656275";
    when 16#0192E# => romdata <= X"67207472";
    when 16#0192F# => romdata <= X"61636520";
    when 16#01930# => romdata <= X"3C636C65";
    when 16#01931# => romdata <= X"61723E00";
    when 16#01932# => romdata <= X"74726163";
    when 16#01933# => romdata <= X"65000000";
    when 16#01934# => romdata <= X"73657475";
    when 16#01935# => romdata <= X"70206368";
    when 16#01936# => romdata <= X"616E6E65";
    when 16#01937# => romdata <= X"6C207465";
    when 16#01938# => romdata <= X"7374203C";
    when 16#01939# => romdata <= X"63683E20";
    when 16#0193A# => romdata <= X"3C76616C";
    when 16#0193B# => romdata <= X"302E2E37";
    when 16#0193C# => romdata <= X"3E000000";
    when 16#0193D# => romdata <= X"63687465";
    when 16#0193E# => romdata <= X"73740000";
    when 16#0193F# => romdata <= X"72756E6E";
    when 16#01940# => romdata <= X"696E6720";
    when 16#01941# => romdata <= X"6C696768";
    when 16#01942# => romdata <= X"74000000";
    when 16#01943# => romdata <= X"72756E00";
    when 16#01944# => romdata <= X"72756E20";
    when 16#01945# => romdata <= X"64697370";
    when 16#01946# => romdata <= X"6C617920";
    when 16#01947# => romdata <= X"74657374";
    when 16#01948# => romdata <= X"2066756E";
    when 16#01949# => romdata <= X"6374696F";
    when 16#0194A# => romdata <= X"6E000000";
    when 16#0194B# => romdata <= X"64697370";
    when 16#0194C# => romdata <= X"6C617900";
    when 16#0194D# => romdata <= X"73657420";
    when 16#0194E# => romdata <= X"6261636B";
    when 16#0194F# => romdata <= X"6C696768";
    when 16#01950# => romdata <= X"74203C30";
    when 16#01951# => romdata <= X"2E2E3331";
    when 16#01952# => romdata <= X"3E000000";
    when 16#01953# => romdata <= X"6261636B";
    when 16#01954# => romdata <= X"00000000";
    when 16#01955# => romdata <= X"73686F77";
    when 16#01956# => romdata <= X"206C6F67";
    when 16#01957# => romdata <= X"6F206F6E";
    when 16#01958# => romdata <= X"20676C63";
    when 16#01959# => romdata <= X"64000000";
    when 16#0195A# => romdata <= X"6C6F676F";
    when 16#0195B# => romdata <= X"00000000";
    when 16#0195C# => romdata <= X"63686563";
    when 16#0195D# => romdata <= X"6B204932";
    when 16#0195E# => romdata <= X"43206164";
    when 16#0195F# => romdata <= X"64726573";
    when 16#01960# => romdata <= X"73000000";
    when 16#01961# => romdata <= X"69326300";
    when 16#01962# => romdata <= X"72656164";
    when 16#01963# => romdata <= X"20454550";
    when 16#01964# => romdata <= X"524F4D20";
    when 16#01965# => romdata <= X"3C627573";
    when 16#01966# => romdata <= X"3E203C69";
    when 16#01967# => romdata <= X"32635F61";
    when 16#01968# => romdata <= X"6464723E";
    when 16#01969# => romdata <= X"203C6C65";
    when 16#0196A# => romdata <= X"6E677468";
    when 16#0196B# => romdata <= X"3E000000";
    when 16#0196C# => romdata <= X"65657072";
    when 16#0196D# => romdata <= X"6F6D0000";
    when 16#0196E# => romdata <= X"41444320";
    when 16#0196F# => romdata <= X"72656769";
    when 16#01970# => romdata <= X"73746572";
    when 16#01971# => romdata <= X"20747261";
    when 16#01972# => romdata <= X"6E736665";
    when 16#01973# => romdata <= X"72203C76";
    when 16#01974# => romdata <= X"616C7565";
    when 16#01975# => romdata <= X"3E000000";
    when 16#01976# => romdata <= X"61747261";
    when 16#01977# => romdata <= X"6E730000";
    when 16#01978# => romdata <= X"696E6974";
    when 16#01979# => romdata <= X"20414443";
    when 16#0197A# => romdata <= X"20726567";
    when 16#0197B# => romdata <= X"69737465";
    when 16#0197C# => romdata <= X"72730000";
    when 16#0197D# => romdata <= X"61696E69";
    when 16#0197E# => romdata <= X"74000000";
    when 16#0197F# => romdata <= X"72656164";
    when 16#01980# => romdata <= X"20636872";
    when 16#01981# => romdata <= X"6F6E7465";
    when 16#01982# => romdata <= X"6C207265";
    when 16#01983# => romdata <= X"67697374";
    when 16#01984# => romdata <= X"65727300";
    when 16#01985# => romdata <= X"63726561";
    when 16#01986# => romdata <= X"64000000";
    when 16#01987# => romdata <= X"696E6974";
    when 16#01988# => romdata <= X"20636872";
    when 16#01989# => romdata <= X"6F6E7465";
    when 16#0198A# => romdata <= X"6C207265";
    when 16#0198B# => romdata <= X"67697374";
    when 16#0198C# => romdata <= X"65727300";
    when 16#0198D# => romdata <= X"63696E69";
    when 16#0198E# => romdata <= X"74000000";
    when 16#0198F# => romdata <= X"77726974";
    when 16#01990# => romdata <= X"65206368";
    when 16#01991# => romdata <= X"726F6E74";
    when 16#01992# => romdata <= X"656C2072";
    when 16#01993# => romdata <= X"65676973";
    when 16#01994# => romdata <= X"74657220";
    when 16#01995# => romdata <= X"3C726567";
    when 16#01996# => romdata <= X"3E203C76";
    when 16#01997# => romdata <= X"616C7565";
    when 16#01998# => romdata <= X"3E000000";
    when 16#01999# => romdata <= X"63777269";
    when 16#0199A# => romdata <= X"74650000";
    when 16#0199B# => romdata <= X"616C6961";
    when 16#0199C# => romdata <= X"7320666F";
    when 16#0199D# => romdata <= X"72207800";
    when 16#0199E# => romdata <= X"6D656D00";
    when 16#0199F# => romdata <= X"77726974";
    when 16#019A0# => romdata <= X"6520776F";
    when 16#019A1# => romdata <= X"7264203C";
    when 16#019A2# => romdata <= X"61646472";
    when 16#019A3# => romdata <= X"3E203C6C";
    when 16#019A4# => romdata <= X"656E6774";
    when 16#019A5# => romdata <= X"683E203C";
    when 16#019A6# => romdata <= X"76616C75";
    when 16#019A7# => romdata <= X"65287329";
    when 16#019A8# => romdata <= X"3E000000";
    when 16#019A9# => romdata <= X"776D656D";
    when 16#019AA# => romdata <= X"00000000";
    when 16#019AB# => romdata <= X"6558616D";
    when 16#019AC# => romdata <= X"696E6520";
    when 16#019AD# => romdata <= X"6D656D6F";
    when 16#019AE# => romdata <= X"7279203C";
    when 16#019AF# => romdata <= X"61646472";
    when 16#019B0# => romdata <= X"3E203C6C";
    when 16#019B1# => romdata <= X"656E6774";
    when 16#019B2# => romdata <= X"683E0000";
    when 16#019B3# => romdata <= X"636C6561";
    when 16#019B4# => romdata <= X"72207363";
    when 16#019B5# => romdata <= X"7265656E";
    when 16#019B6# => romdata <= X"00000000";
    when 16#019B7# => romdata <= X"636C6561";
    when 16#019B8# => romdata <= X"72000000";
    when 16#019B9# => romdata <= X"65787465";
    when 16#019BA# => romdata <= X"726E616C";
    when 16#019BB# => romdata <= X"20636C6F";
    when 16#019BC# => romdata <= X"636B2000";
    when 16#019BD# => romdata <= X"61637469";
    when 16#019BE# => romdata <= X"76650A00";
    when 16#019BF# => romdata <= X"73656C65";
    when 16#019C0# => romdata <= X"63746564";
    when 16#019C1# => romdata <= X"0A000000";
    when 16#019C2# => romdata <= X"4E4F5420";
    when 16#019C3# => romdata <= X"00000000";
    when 16#019C4# => romdata <= X"6D696372";
    when 16#019C5# => romdata <= X"6F70756C";
    when 16#019C6# => romdata <= X"73652073";
    when 16#019C7# => romdata <= X"6F757263";
    when 16#019C8# => romdata <= X"653A2000";
    when 16#019C9# => romdata <= X"65787465";
    when 16#019CA# => romdata <= X"726E616C";
    when 16#019CB# => romdata <= X"00000000";
    when 16#019CC# => romdata <= X"6265616D";
    when 16#019CD# => romdata <= X"20706F73";
    when 16#019CE# => romdata <= X"6974696F";
    when 16#019CF# => romdata <= X"6E206D6F";
    when 16#019D0# => romdata <= X"6E69746F";
    when 16#019D1# => romdata <= X"72000000";
    when 16#019D2# => romdata <= X"0A0A0000";
    when 16#019D3# => romdata <= X"20286F6E";
    when 16#019D4# => romdata <= X"2073696D";
    when 16#019D5# => romdata <= X"290A0000";
    when 16#019D6# => romdata <= X"0A485720";
    when 16#019D7# => romdata <= X"73796E74";
    when 16#019D8# => romdata <= X"68657369";
    when 16#019D9# => romdata <= X"7A65643A";
    when 16#019DA# => romdata <= X"20000000";
    when 16#019DB# => romdata <= X"0A535720";
    when 16#019DC# => romdata <= X"636F6D70";
    when 16#019DD# => romdata <= X"696C6564";
    when 16#019DE# => romdata <= X"2020203A";
    when 16#019DF# => romdata <= X"20536570";
    when 16#019E0# => romdata <= X"20203920";
    when 16#019E1# => romdata <= X"32303131";
    when 16#019E2# => romdata <= X"20203134";
    when 16#019E3# => romdata <= X"3A31363A";
    when 16#019E4# => romdata <= X"34340000";
    when 16#019E5# => romdata <= X"0A737973";
    when 16#019E6# => romdata <= X"74656D20";
    when 16#019E7# => romdata <= X"636C6F63";
    when 16#019E8# => romdata <= X"6B20203A";
    when 16#019E9# => romdata <= X"20000000";
    when 16#019EA# => romdata <= X"204D487A";
    when 16#019EB# => romdata <= X"0A000000";
    when 16#019EC# => romdata <= X"44454255";
    when 16#019ED# => romdata <= X"47204D4F";
    when 16#019EE# => romdata <= X"44450000";
    when 16#019EF# => romdata <= X"20282B44";
    when 16#019F0# => romdata <= X"56492900";
    when 16#019F1# => romdata <= X"20282B64";
    when 16#019F2# => romdata <= X"65627567";
    when 16#019F3# => romdata <= X"20627566";
    when 16#019F4# => romdata <= X"66657220";
    when 16#019F5# => romdata <= X"7472616E";
    when 16#019F6# => romdata <= X"73666572";
    when 16#019F7# => romdata <= X"29000000";
    when 16#019F8# => romdata <= X"204F4E0A";
    when 16#019F9# => romdata <= X"00000000";
    when 16#019FA# => romdata <= X"6265616D";
    when 16#019FB# => romdata <= X"20706F73";
    when 16#019FC# => romdata <= X"6974696F";
    when 16#019FD# => romdata <= X"6E206D6F";
    when 16#019FE# => romdata <= X"6E69746F";
    when 16#019FF# => romdata <= X"720A0000";
    when 16#01A00# => romdata <= X"0A536570";
    when 16#01A01# => romdata <= X"20203920";
    when 16#01A02# => romdata <= X"32303131";
    when 16#01A03# => romdata <= X"20203134";
    when 16#01A04# => romdata <= X"3A31363A";
    when 16#01A05# => romdata <= X"34340000";
    when 16#01A06# => romdata <= X"0A696E69";
    when 16#01A07# => romdata <= X"74204144";
    when 16#01A08# => romdata <= X"43000000";
    when 16#01A09# => romdata <= X"0A696E69";
    when 16#01A0A# => romdata <= X"7420434C";
    when 16#01A0B# => romdata <= X"4B000000";
    when 16#01A0C# => romdata <= X"0A696E69";
    when 16#01A0D# => romdata <= X"74204441";
    when 16#01A0E# => romdata <= X"43000000";
    when 16#01A0F# => romdata <= X"0A696E69";
    when 16#01A10# => romdata <= X"74204250";
    when 16#01A11# => romdata <= X"4D000000";
    when 16#01A12# => romdata <= X"202D2D3E";
    when 16#01A13# => romdata <= X"20455252";
    when 16#01A14# => romdata <= X"4F520000";
    when 16#01A15# => romdata <= X"4552524F";
    when 16#01A16# => romdata <= X"523A2074";
    when 16#01A17# => romdata <= X"6F6F206D";
    when 16#01A18# => romdata <= X"75636820";
    when 16#01A19# => romdata <= X"636F6D6D";
    when 16#01A1A# => romdata <= X"616E6473";
    when 16#01A1B# => romdata <= X"2E0A0000";
    when 16#01A1C# => romdata <= X"3E200000";
    when 16#01A1D# => romdata <= X"636F6D6D";
    when 16#01A1E# => romdata <= X"616E6420";
    when 16#01A1F# => romdata <= X"6E6F7420";
    when 16#01A20# => romdata <= X"666F756E";
    when 16#01A21# => romdata <= X"642E0A00";
    when 16#01A22# => romdata <= X"73757070";
    when 16#01A23# => romdata <= X"6F727465";
    when 16#01A24# => romdata <= X"6420636F";
    when 16#01A25# => romdata <= X"6D6D616E";
    when 16#01A26# => romdata <= X"64733A0A";
    when 16#01A27# => romdata <= X"0A000000";
    when 16#01A28# => romdata <= X"202D2000";
    when 16#01A29# => romdata <= X"76656E64";
    when 16#01A2A# => romdata <= X"6F723F20";
    when 16#01A2B# => romdata <= X"20000000";
    when 16#01A2C# => romdata <= X"485A4452";
    when 16#01A2D# => romdata <= X"20202020";
    when 16#01A2E# => romdata <= X"20000000";
    when 16#01A2F# => romdata <= X"67616973";
    when 16#01A30# => romdata <= X"6C657220";
    when 16#01A31# => romdata <= X"20000000";
    when 16#01A32# => romdata <= X"4148422F";
    when 16#01A33# => romdata <= X"41504220";
    when 16#01A34# => romdata <= X"42726964";
    when 16#01A35# => romdata <= X"67650000";
    when 16#01A36# => romdata <= X"45534120";
    when 16#01A37# => romdata <= X"20202020";
    when 16#01A38# => romdata <= X"20000000";
    when 16#01A39# => romdata <= X"756E6B6E";
    when 16#01A3A# => romdata <= X"6F776E20";
    when 16#01A3B# => romdata <= X"64657669";
    when 16#01A3C# => romdata <= X"63650000";
    when 16#01A3D# => romdata <= X"4C656F6E";
    when 16#01A3E# => romdata <= X"32204D65";
    when 16#01A3F# => romdata <= X"6D6F7279";
    when 16#01A40# => romdata <= X"20436F6E";
    when 16#01A41# => romdata <= X"74726F6C";
    when 16#01A42# => romdata <= X"6C657200";
    when 16#01A43# => romdata <= X"47522031";
    when 16#01A44# => romdata <= X"302F3130";
    when 16#01A45# => romdata <= X"30204D62";
    when 16#01A46# => romdata <= X"69742045";
    when 16#01A47# => romdata <= X"74686572";
    when 16#01A48# => romdata <= X"6E657420";
    when 16#01A49# => romdata <= X"4D414300";
    when 16#01A4A# => romdata <= X"64696666";
    when 16#01A4B# => romdata <= X"6572656E";
    when 16#01A4C# => romdata <= X"7469616C";
    when 16#01A4D# => romdata <= X"20637572";
    when 16#01A4E# => romdata <= X"72656E74";
    when 16#01A4F# => romdata <= X"206D6F6E";
    when 16#01A50# => romdata <= X"69746F72";
    when 16#01A51# => romdata <= X"00000000";
    when 16#01A52# => romdata <= X"64656275";
    when 16#01A53# => romdata <= X"67207472";
    when 16#01A54# => romdata <= X"61636572";
    when 16#01A55# => romdata <= X"206D656D";
    when 16#01A56# => romdata <= X"6F727900";
    when 16#01A57# => romdata <= X"4541444F";
    when 16#01A58# => romdata <= X"47533130";
    when 16#01A59# => romdata <= X"32206469";
    when 16#01A5A# => romdata <= X"73706C61";
    when 16#01A5B# => romdata <= X"79206472";
    when 16#01A5C# => romdata <= X"69766572";
    when 16#01A5D# => romdata <= X"00000000";
    when 16#01A5E# => romdata <= X"64656275";
    when 16#01A5F# => romdata <= X"67206275";
    when 16#01A60# => romdata <= X"66666572";
    when 16#01A61# => romdata <= X"20636F6E";
    when 16#01A62# => romdata <= X"74726F6C";
    when 16#01A63# => romdata <= X"00000000";
    when 16#01A64# => romdata <= X"74726967";
    when 16#01A65# => romdata <= X"67657220";
    when 16#01A66# => romdata <= X"67656E65";
    when 16#01A67# => romdata <= X"7261746F";
    when 16#01A68# => romdata <= X"72000000";
    when 16#01A69# => romdata <= X"64656275";
    when 16#01A6A# => romdata <= X"6720636F";
    when 16#01A6B# => romdata <= X"6E736F6C";
    when 16#01A6C# => romdata <= X"65000000";
    when 16#01A6D# => romdata <= X"44434D20";
    when 16#01A6E# => romdata <= X"70686173";
    when 16#01A6F# => romdata <= X"65207368";
    when 16#01A70# => romdata <= X"69667420";
    when 16#01A71# => romdata <= X"636F6E74";
    when 16#01A72# => romdata <= X"726F6C00";
    when 16#01A73# => romdata <= X"5A505520";
    when 16#01A74# => romdata <= X"4D656D6F";
    when 16#01A75# => romdata <= X"72792077";
    when 16#01A76# => romdata <= X"72617070";
    when 16#01A77# => romdata <= X"65720000";
    when 16#01A78# => romdata <= X"5A505520";
    when 16#01A79# => romdata <= X"41484220";
    when 16#01A7A# => romdata <= X"57726170";
    when 16#01A7B# => romdata <= X"70657200";
    when 16#01A7C# => romdata <= X"56474120";
    when 16#01A7D# => romdata <= X"636F6E74";
    when 16#01A7E# => romdata <= X"726F6C6C";
    when 16#01A7F# => romdata <= X"65720000";
    when 16#01A80# => romdata <= X"4D6F6475";
    when 16#01A81# => romdata <= X"6C617220";
    when 16#01A82# => romdata <= X"54696D65";
    when 16#01A83# => romdata <= X"7220556E";
    when 16#01A84# => romdata <= X"69740000";
    when 16#01A85# => romdata <= X"47656E65";
    when 16#01A86# => romdata <= X"72616C20";
    when 16#01A87# => romdata <= X"50757270";
    when 16#01A88# => romdata <= X"6F736520";
    when 16#01A89# => romdata <= X"492F4F20";
    when 16#01A8A# => romdata <= X"706F7274";
    when 16#01A8B# => romdata <= X"00000000";
    when 16#01A8C# => romdata <= X"47656E65";
    when 16#01A8D# => romdata <= X"72696320";
    when 16#01A8E# => romdata <= X"55415254";
    when 16#01A8F# => romdata <= X"00000000";
    when 16#01A90# => romdata <= X"414D4241";
    when 16#01A91# => romdata <= X"20577261";
    when 16#01A92# => romdata <= X"70706572";
    when 16#01A93# => romdata <= X"20666F72";
    when 16#01A94# => romdata <= X"204F4320";
    when 16#01A95# => romdata <= X"4932432D";
    when 16#01A96# => romdata <= X"6D617374";
    when 16#01A97# => romdata <= X"65720000";
    when 16#01A98# => romdata <= X"53504920";
    when 16#01A99# => romdata <= X"4D656D6F";
    when 16#01A9A# => romdata <= X"72792043";
    when 16#01A9B# => romdata <= X"6F6E7472";
    when 16#01A9C# => romdata <= X"6F6C6C65";
    when 16#01A9D# => romdata <= X"72000000";
    when 16#01A9E# => romdata <= X"4475616C";
    when 16#01A9F# => romdata <= X"2D706F72";
    when 16#01AA0# => romdata <= X"74204148";
    when 16#01AA1# => romdata <= X"42205352";
    when 16#01AA2# => romdata <= X"414D206D";
    when 16#01AA3# => romdata <= X"6F64756C";
    when 16#01AA4# => romdata <= X"65000000";
    when 16#01AA5# => romdata <= X"20206170";
    when 16#01AA6# => romdata <= X"62736C76";
    when 16#01AA7# => romdata <= X"00000000";
    when 16#01AA8# => romdata <= X"76656E64";
    when 16#01AA9# => romdata <= X"20307800";
    when 16#01AAA# => romdata <= X"64657620";
    when 16#01AAB# => romdata <= X"30780000";
    when 16#01AAC# => romdata <= X"76657220";
    when 16#01AAD# => romdata <= X"00000000";
    when 16#01AAE# => romdata <= X"69727120";
    when 16#01AAF# => romdata <= X"00000000";
    when 16#01AB0# => romdata <= X"61646472";
    when 16#01AB1# => romdata <= X"20307800";
    when 16#01AB2# => romdata <= X"6168626D";
    when 16#01AB3# => romdata <= X"73740000";
    when 16#01AB4# => romdata <= X"61686273";
    when 16#01AB5# => romdata <= X"6C760000";
    when 16#01AB6# => romdata <= X"000018DB";
    when 16#01AB7# => romdata <= X"0000197F";
    when 16#01AB8# => romdata <= X"00001973";
    when 16#01AB9# => romdata <= X"00001967";
    when 16#01ABA# => romdata <= X"0000195B";
    when 16#01ABB# => romdata <= X"0000194F";
    when 16#01ABC# => romdata <= X"00001943";
    when 16#01ABD# => romdata <= X"00001937";
    when 16#01ABE# => romdata <= X"0000192B";
    when 16#01ABF# => romdata <= X"0000191F";
    when 16#01AC0# => romdata <= X"00001913";
    when 16#01AC1# => romdata <= X"04580808";
    when 16#01AC2# => romdata <= X"20FF0000";
    when 16#01AC3# => romdata <= X"00006B14";
    when 16#01AC4# => romdata <= X"00006BF4";
    when 16#01AC5# => romdata <= X"02010305";
    when 16#01AC6# => romdata <= X"05070501";
    when 16#01AC7# => romdata <= X"03030505";
    when 16#01AC8# => romdata <= X"02030104";
    when 16#01AC9# => romdata <= X"05050505";
    when 16#01ACA# => romdata <= X"05050505";
    when 16#01ACB# => romdata <= X"05050101";
    when 16#01ACC# => romdata <= X"04050404";
    when 16#01ACD# => romdata <= X"07050505";
    when 16#01ACE# => romdata <= X"05050505";
    when 16#01ACF# => romdata <= X"05030405";
    when 16#01AD0# => romdata <= X"05050505";
    when 16#01AD1# => romdata <= X"05050505";
    when 16#01AD2# => romdata <= X"05050505";
    when 16#01AD3# => romdata <= X"05050503";
    when 16#01AD4# => romdata <= X"04030505";
    when 16#01AD5# => romdata <= X"02050504";
    when 16#01AD6# => romdata <= X"05050405";
    when 16#01AD7# => romdata <= X"04010204";
    when 16#01AD8# => romdata <= X"02050404";
    when 16#01AD9# => romdata <= X"05050404";
    when 16#01ADA# => romdata <= X"04040507";
    when 16#01ADB# => romdata <= X"05040404";
    when 16#01ADC# => romdata <= X"02040500";
    when 16#01ADD# => romdata <= X"04050200";
    when 16#01ADE# => romdata <= X"04080303";
    when 16#01ADF# => romdata <= X"04090003";
    when 16#01AE0# => romdata <= X"06000000";
    when 16#01AE1# => romdata <= X"00020204";
    when 16#01AE2# => romdata <= X"04040400";
    when 16#01AE3# => romdata <= X"04060003";
    when 16#01AE4# => romdata <= X"05000000";
    when 16#01AE5# => romdata <= X"00000404";
    when 16#01AE6# => romdata <= X"05050204";
    when 16#01AE7# => romdata <= X"05060305";
    when 16#01AE8# => romdata <= X"04030705";
    when 16#01AE9# => romdata <= X"04050303";
    when 16#01AEA# => romdata <= X"02040502";
    when 16#01AEB# => romdata <= X"03020405";
    when 16#01AEC# => romdata <= X"06060604";
    when 16#01AED# => romdata <= X"05050505";
    when 16#01AEE# => romdata <= X"05050504";
    when 16#01AEF# => romdata <= X"04040404";
    when 16#01AF0# => romdata <= X"03030303";
    when 16#01AF1# => romdata <= X"05050505";
    when 16#01AF2# => romdata <= X"05050505";
    when 16#01AF3# => romdata <= X"05040404";
    when 16#01AF4# => romdata <= X"04050404";
    when 16#01AF5# => romdata <= X"04040404";
    when 16#01AF6# => romdata <= X"04040503";
    when 16#01AF7# => romdata <= X"04040404";
    when 16#01AF8# => romdata <= X"02020303";
    when 16#01AF9# => romdata <= X"04040404";
    when 16#01AFA# => romdata <= X"04040405";
    when 16#01AFB# => romdata <= X"04040404";
    when 16#01AFC# => romdata <= X"04030303";
    when 16#01AFD# => romdata <= X"00005F07";
    when 16#01AFE# => romdata <= X"0007741C";
    when 16#01AFF# => romdata <= X"771C172E";
    when 16#01B00# => romdata <= X"6A3E2B3A";
    when 16#01B01# => romdata <= X"06493608";
    when 16#01B02# => romdata <= X"36493036";
    when 16#01B03# => romdata <= X"49597648";
    when 16#01B04# => romdata <= X"073C4281";
    when 16#01B05# => romdata <= X"81423C0A";
    when 16#01B06# => romdata <= X"041F040A";
    when 16#01B07# => romdata <= X"08083E08";
    when 16#01B08# => romdata <= X"08806008";
    when 16#01B09# => romdata <= X"080840C0";
    when 16#01B0A# => romdata <= X"300C033E";
    when 16#01B0B# => romdata <= X"4141413E";
    when 16#01B0C# => romdata <= X"44427F40";
    when 16#01B0D# => romdata <= X"40466151";
    when 16#01B0E# => romdata <= X"49462241";
    when 16#01B0F# => romdata <= X"49493618";
    when 16#01B10# => romdata <= X"14127F10";
    when 16#01B11# => romdata <= X"27454545";
    when 16#01B12# => romdata <= X"393E4949";
    when 16#01B13# => romdata <= X"49300101";
    when 16#01B14# => romdata <= X"710D0336";
    when 16#01B15# => romdata <= X"49494936";
    when 16#01B16# => romdata <= X"06494929";
    when 16#01B17# => romdata <= X"1E36D008";
    when 16#01B18# => romdata <= X"14224114";
    when 16#01B19# => romdata <= X"14141414";
    when 16#01B1A# => romdata <= X"41221408";
    when 16#01B1B# => romdata <= X"02510906";
    when 16#01B1C# => romdata <= X"3C4299A5";
    when 16#01B1D# => romdata <= X"BD421C7C";
    when 16#01B1E# => romdata <= X"1211127C";
    when 16#01B1F# => romdata <= X"7F494949";
    when 16#01B20# => romdata <= X"363E4141";
    when 16#01B21# => romdata <= X"41227F41";
    when 16#01B22# => romdata <= X"41413E7F";
    when 16#01B23# => romdata <= X"49494941";
    when 16#01B24# => romdata <= X"7F090909";
    when 16#01B25# => romdata <= X"013E4149";
    when 16#01B26# => romdata <= X"497A7F08";
    when 16#01B27# => romdata <= X"08087F41";
    when 16#01B28# => romdata <= X"7F414041";
    when 16#01B29# => romdata <= X"413F7F08";
    when 16#01B2A# => romdata <= X"1422417F";
    when 16#01B2B# => romdata <= X"40404040";
    when 16#01B2C# => romdata <= X"7F060C06";
    when 16#01B2D# => romdata <= X"7F7F0608";
    when 16#01B2E# => romdata <= X"307F3E41";
    when 16#01B2F# => romdata <= X"41413E7F";
    when 16#01B30# => romdata <= X"09090906";
    when 16#01B31# => romdata <= X"3E4161C1";
    when 16#01B32# => romdata <= X"BE7F0919";
    when 16#01B33# => romdata <= X"29462649";
    when 16#01B34# => romdata <= X"49493201";
    when 16#01B35# => romdata <= X"017F0101";
    when 16#01B36# => romdata <= X"3F404040";
    when 16#01B37# => romdata <= X"3F073840";
    when 16#01B38# => romdata <= X"38071F60";
    when 16#01B39# => romdata <= X"1F601F63";
    when 16#01B3A# => romdata <= X"14081463";
    when 16#01B3B# => romdata <= X"01067806";
    when 16#01B3C# => romdata <= X"01615149";
    when 16#01B3D# => romdata <= X"45437F41";
    when 16#01B3E# => romdata <= X"41030C30";
    when 16#01B3F# => romdata <= X"C041417F";
    when 16#01B40# => romdata <= X"04020102";
    when 16#01B41# => romdata <= X"04808080";
    when 16#01B42# => romdata <= X"80800102";
    when 16#01B43# => romdata <= X"20545454";
    when 16#01B44# => romdata <= X"787F4444";
    when 16#01B45# => romdata <= X"44383844";
    when 16#01B46# => romdata <= X"44443844";
    when 16#01B47# => romdata <= X"44447F38";
    when 16#01B48# => romdata <= X"54545458";
    when 16#01B49# => romdata <= X"087E0901";
    when 16#01B4A# => romdata <= X"18A4A4A4";
    when 16#01B4B# => romdata <= X"787F0404";
    when 16#01B4C# => romdata <= X"787D807D";
    when 16#01B4D# => romdata <= X"7F102844";
    when 16#01B4E# => romdata <= X"3F407C04";
    when 16#01B4F# => romdata <= X"7804787C";
    when 16#01B50# => romdata <= X"04047838";
    when 16#01B51# => romdata <= X"444438FC";
    when 16#01B52# => romdata <= X"24242418";
    when 16#01B53# => romdata <= X"18242424";
    when 16#01B54# => romdata <= X"FC7C0804";
    when 16#01B55# => romdata <= X"04485454";
    when 16#01B56# => romdata <= X"24043F44";
    when 16#01B57# => romdata <= X"403C4040";
    when 16#01B58# => romdata <= X"7C1C2040";
    when 16#01B59# => romdata <= X"201C1C60";
    when 16#01B5A# => romdata <= X"601C6060";
    when 16#01B5B# => romdata <= X"1C442810";
    when 16#01B5C# => romdata <= X"28449CA0";
    when 16#01B5D# => romdata <= X"601C6454";
    when 16#01B5E# => romdata <= X"544C187E";
    when 16#01B5F# => romdata <= X"8181FFFF";
    when 16#01B60# => romdata <= X"81817E18";
    when 16#01B61# => romdata <= X"18040810";
    when 16#01B62# => romdata <= X"0C143E55";
    when 16#01B63# => romdata <= X"55FF8181";
    when 16#01B64# => romdata <= X"81FF8060";
    when 16#01B65# => romdata <= X"80608060";
    when 16#01B66# => romdata <= X"60600060";
    when 16#01B67# => romdata <= X"60006060";
    when 16#01B68# => romdata <= X"047F0414";
    when 16#01B69# => romdata <= X"7F140201";
    when 16#01B6A# => romdata <= X"01024629";
    when 16#01B6B# => romdata <= X"1608344A";
    when 16#01B6C# => romdata <= X"31483000";
    when 16#01B6D# => romdata <= X"18243E41";
    when 16#01B6E# => romdata <= X"227F4941";
    when 16#01B6F# => romdata <= X"03040403";
    when 16#01B70# => romdata <= X"03040304";
    when 16#01B71# => romdata <= X"04030403";
    when 16#01B72# => romdata <= X"183C3C18";
    when 16#01B73# => romdata <= X"08080808";
    when 16#01B74# => romdata <= X"03010203";
    when 16#01B75# => romdata <= X"020E020E";
    when 16#01B76# => romdata <= X"060E0048";
    when 16#01B77# => romdata <= X"30384438";
    when 16#01B78# => romdata <= X"54483844";
    when 16#01B79# => romdata <= X"FE44487E";
    when 16#01B7A# => romdata <= X"49014438";
    when 16#01B7B# => romdata <= X"28384403";
    when 16#01B7C# => romdata <= X"147C1403";
    when 16#01B7D# => romdata <= X"E7E74E55";
    when 16#01B7E# => romdata <= X"55390101";
    when 16#01B7F# => romdata <= X"0001011C";
    when 16#01B80# => romdata <= X"2A555522";
    when 16#01B81# => romdata <= X"1C1D151E";
    when 16#01B82# => romdata <= X"18240018";
    when 16#01B83# => romdata <= X"24080808";
    when 16#01B84# => romdata <= X"18080808";
    when 16#01B85# => romdata <= X"3C42BD95";
    when 16#01B86# => romdata <= X"A9423C01";
    when 16#01B87# => romdata <= X"01010101";
    when 16#01B88# => romdata <= X"06090906";
    when 16#01B89# => romdata <= X"44445F44";
    when 16#01B8A# => romdata <= X"44191512";
    when 16#01B8B# => romdata <= X"15150A02";
    when 16#01B8C# => romdata <= X"01FC2020";
    when 16#01B8D# => romdata <= X"1C0E7F01";
    when 16#01B8E# => romdata <= X"7F011818";
    when 16#01B8F# => romdata <= X"00804002";
    when 16#01B90# => romdata <= X"1F060909";
    when 16#01B91# => romdata <= X"06241800";
    when 16#01B92# => romdata <= X"2418824F";
    when 16#01B93# => romdata <= X"304C62F1";
    when 16#01B94# => romdata <= X"824F300C";
    when 16#01B95# => romdata <= X"D2B1955F";
    when 16#01B96# => romdata <= X"304C62F1";
    when 16#01B97# => romdata <= X"30484520";
    when 16#01B98# => romdata <= X"60392E38";
    when 16#01B99# => romdata <= X"6060382E";
    when 16#01B9A# => romdata <= X"3960701D";
    when 16#01B9B# => romdata <= X"131D7072";
    when 16#01B9C# => romdata <= X"1D121E71";
    when 16#01B9D# => romdata <= X"701D121D";
    when 16#01B9E# => romdata <= X"70603B25";
    when 16#01B9F# => romdata <= X"3B607E11";
    when 16#01BA0# => romdata <= X"7F49411E";
    when 16#01BA1# => romdata <= X"2161927C";
    when 16#01BA2# => romdata <= X"5556447C";
    when 16#01BA3# => romdata <= X"5655447C";
    when 16#01BA4# => romdata <= X"5655467D";
    when 16#01BA5# => romdata <= X"54544545";
    when 16#01BA6# => romdata <= X"7E44447E";
    when 16#01BA7# => romdata <= X"45467D46";
    when 16#01BA8# => romdata <= X"457C4508";
    when 16#01BA9# => romdata <= X"7F49413E";
    when 16#01BAA# => romdata <= X"7E091222";
    when 16#01BAB# => romdata <= X"7D384546";
    when 16#01BAC# => romdata <= X"44383844";
    when 16#01BAD# => romdata <= X"46453838";
    when 16#01BAE# => romdata <= X"46454638";
    when 16#01BAF# => romdata <= X"3A454546";
    when 16#01BB0# => romdata <= X"39384544";
    when 16#01BB1# => romdata <= X"45382214";
    when 16#01BB2# => romdata <= X"081422BC";
    when 16#01BB3# => romdata <= X"625A463D";
    when 16#01BB4# => romdata <= X"3C41423C";
    when 16#01BB5# => romdata <= X"3C42413C";
    when 16#01BB6# => romdata <= X"3C42413E";
    when 16#01BB7# => romdata <= X"3D40403D";
    when 16#01BB8# => romdata <= X"0608F209";
    when 16#01BB9# => romdata <= X"067F2222";
    when 16#01BBA# => romdata <= X"1CFE0989";
    when 16#01BBB# => romdata <= X"76205556";
    when 16#01BBC# => romdata <= X"78205655";
    when 16#01BBD# => romdata <= X"78225555";
    when 16#01BBE# => romdata <= X"7A235556";
    when 16#01BBF# => romdata <= X"7B205554";
    when 16#01BC0# => romdata <= X"79275557";
    when 16#01BC1# => romdata <= X"78205438";
    when 16#01BC2# => romdata <= X"54483844";
    when 16#01BC3# => romdata <= X"C4385556";
    when 16#01BC4# => romdata <= X"58385655";
    when 16#01BC5# => romdata <= X"583A5555";
    when 16#01BC6# => romdata <= X"5A395454";
    when 16#01BC7# => romdata <= X"59017A7A";
    when 16#01BC8# => romdata <= X"01027902";
    when 16#01BC9# => romdata <= X"02780260";
    when 16#01BCA# => romdata <= X"91927C7B";
    when 16#01BCB# => romdata <= X"090A7338";
    when 16#01BCC# => romdata <= X"45463838";
    when 16#01BCD# => romdata <= X"4645383A";
    when 16#01BCE# => romdata <= X"45453A3B";
    when 16#01BCF# => romdata <= X"45463B39";
    when 16#01BD0# => romdata <= X"44443908";
    when 16#01BD1# => romdata <= X"082A0808";
    when 16#01BD2# => romdata <= X"B8644C3A";
    when 16#01BD3# => romdata <= X"3C41427C";
    when 16#01BD4# => romdata <= X"3C42417C";
    when 16#01BD5# => romdata <= X"3A41417A";
    when 16#01BD6# => romdata <= X"3D40407D";
    when 16#01BD7# => romdata <= X"986219FF";
    when 16#01BD8# => romdata <= X"423C9A60";
    when 16#01BD9# => romdata <= X"1A000000";
    when 16#01BDA# => romdata <= X"69326320";
    when 16#01BDB# => romdata <= X"4456490A";
    when 16#01BDC# => romdata <= X"00000000";
    when 16#01BDD# => romdata <= X"69326320";
    when 16#01BDE# => romdata <= X"464D430A";
    when 16#01BDF# => romdata <= X"00000000";
    when 16#01BE0# => romdata <= X"61646472";
    when 16#01BE1# => romdata <= X"6573733A";
    when 16#01BE2# => romdata <= X"20307800";
    when 16#01BE3# => romdata <= X"2020202D";
    when 16#01BE4# => romdata <= X"2D3E2020";
    when 16#01BE5# => romdata <= X"2041434B";
    when 16#01BE6# => romdata <= X"0A000000";
    when 16#01BE7# => romdata <= X"72656164";
    when 16#01BE8# => romdata <= X"20646174";
    when 16#01BE9# => romdata <= X"61202800";
    when 16#01BEA# => romdata <= X"20627974";
    when 16#01BEB# => romdata <= X"65732920";
    when 16#01BEC# => romdata <= X"66726F6D";
    when 16#01BED# => romdata <= X"20493243";
    when 16#01BEE# => romdata <= X"2D616464";
    when 16#01BEF# => romdata <= X"72657373";
    when 16#01BF0# => romdata <= X"20307800";
    when 16#01BF1# => romdata <= X"6E6F6163";
    when 16#01BF2# => romdata <= X"6B200000";
    when 16#01BF3# => romdata <= X"6368726F";
    when 16#01BF4# => romdata <= X"6E74656C";
    when 16#01BF5# => romdata <= X"20726567";
    when 16#01BF6# => romdata <= X"20307800";
    when 16#01BF7# => romdata <= X"3A203078";
    when 16#01BF8# => romdata <= X"00000000";
    when 16#01BF9# => romdata <= X"206E6163";
    when 16#01BFA# => romdata <= X"6B000000";
    when 16#01BFB# => romdata <= X"6572726F";
    when 16#01BFC# => romdata <= X"7220286E";
    when 16#01BFD# => romdata <= X"61636B29";
    when 16#01BFE# => romdata <= X"0A000000";
    when 16#01BFF# => romdata <= X"0A202063";
    when 16#01C00# => romdata <= X"68616E6E";
    when 16#01C01# => romdata <= X"656C2033";
    when 16#01C02# => romdata <= X"20696E70";
    when 16#01C03# => romdata <= X"7574206F";
    when 16#01C04# => romdata <= X"76657266";
    when 16#01C05# => romdata <= X"6C6F7700";
    when 16#01C06# => romdata <= X"0A202063";
    when 16#01C07# => romdata <= X"68616E6E";
    when 16#01C08# => romdata <= X"656C2032";
    when 16#01C09# => romdata <= X"20696E70";
    when 16#01C0A# => romdata <= X"7574206F";
    when 16#01C0B# => romdata <= X"76657266";
    when 16#01C0C# => romdata <= X"6C6F7700";
    when 16#01C0D# => romdata <= X"0A202063";
    when 16#01C0E# => romdata <= X"68616E6E";
    when 16#01C0F# => romdata <= X"656C2031";
    when 16#01C10# => romdata <= X"20696E70";
    when 16#01C11# => romdata <= X"7574206F";
    when 16#01C12# => romdata <= X"76657266";
    when 16#01C13# => romdata <= X"6C6F7700";
    when 16#01C14# => romdata <= X"0A202063";
    when 16#01C15# => romdata <= X"68616E6E";
    when 16#01C16# => romdata <= X"656C2030";
    when 16#01C17# => romdata <= X"20696E70";
    when 16#01C18# => romdata <= X"7574206F";
    when 16#01C19# => romdata <= X"76657266";
    when 16#01C1A# => romdata <= X"6C6F7700";
    when 16#01C1B# => romdata <= X"0A202063";
    when 16#01C1C# => romdata <= X"68616E6E";
    when 16#01C1D# => romdata <= X"656C2033";
    when 16#01C1E# => romdata <= X"20717561";
    when 16#01C1F# => romdata <= X"6473756D";
    when 16#01C20# => romdata <= X"206F7665";
    when 16#01C21# => romdata <= X"72666C6F";
    when 16#01C22# => romdata <= X"77000000";
    when 16#01C23# => romdata <= X"0A202063";
    when 16#01C24# => romdata <= X"68616E6E";
    when 16#01C25# => romdata <= X"656C2032";
    when 16#01C26# => romdata <= X"20717561";
    when 16#01C27# => romdata <= X"6473756D";
    when 16#01C28# => romdata <= X"206F7665";
    when 16#01C29# => romdata <= X"72666C6F";
    when 16#01C2A# => romdata <= X"77000000";
    when 16#01C2B# => romdata <= X"0A202063";
    when 16#01C2C# => romdata <= X"68616E6E";
    when 16#01C2D# => romdata <= X"656C2031";
    when 16#01C2E# => romdata <= X"20717561";
    when 16#01C2F# => romdata <= X"6473756D";
    when 16#01C30# => romdata <= X"206F7665";
    when 16#01C31# => romdata <= X"72666C6F";
    when 16#01C32# => romdata <= X"77000000";
    when 16#01C33# => romdata <= X"0A202063";
    when 16#01C34# => romdata <= X"68616E6E";
    when 16#01C35# => romdata <= X"656C2030";
    when 16#01C36# => romdata <= X"20717561";
    when 16#01C37# => romdata <= X"6473756D";
    when 16#01C38# => romdata <= X"206F7665";
    when 16#01C39# => romdata <= X"72666C6F";
    when 16#01C3A# => romdata <= X"77000000";
    when 16#01C3B# => romdata <= X"0A202073";
    when 16#01C3C# => romdata <= X"756D2073";
    when 16#01C3D# => romdata <= X"63616C65";
    when 16#01C3E# => romdata <= X"72206F76";
    when 16#01C3F# => romdata <= X"6572666C";
    when 16#01C40# => romdata <= X"6F770000";
    when 16#01C41# => romdata <= X"0A202073";
    when 16#01C42# => romdata <= X"756D2076";
    when 16#01C43# => romdata <= X"616C7565";
    when 16#01C44# => romdata <= X"20637574";
    when 16#01C45# => romdata <= X"74656400";
    when 16#01C46# => romdata <= X"0A202063";
    when 16#01C47# => romdata <= X"68616E6E";
    when 16#01C48# => romdata <= X"656C2033";
    when 16#01C49# => romdata <= X"20646976";
    when 16#01C4A# => romdata <= X"6964656E";
    when 16#01C4B# => romdata <= X"64206375";
    when 16#01C4C# => romdata <= X"74746564";
    when 16#01C4D# => romdata <= X"00000000";
    when 16#01C4E# => romdata <= X"0A202063";
    when 16#01C4F# => romdata <= X"68616E6E";
    when 16#01C50# => romdata <= X"656C2033";
    when 16#01C51# => romdata <= X"206E6F69";
    when 16#01C52# => romdata <= X"73652063";
    when 16#01C53# => romdata <= X"6F6D7065";
    when 16#01C54# => romdata <= X"6E736174";
    when 16#01C55# => romdata <= X"696F6E20";
    when 16#01C56# => romdata <= X"746F2062";
    when 16#01C57# => romdata <= X"69670000";
    when 16#01C58# => romdata <= X"0A202063";
    when 16#01C59# => romdata <= X"68616E6E";
    when 16#01C5A# => romdata <= X"656C2033";
    when 16#01C5B# => romdata <= X"206E6F69";
    when 16#01C5C# => romdata <= X"73652076";
    when 16#01C5D# => romdata <= X"616C7565";
    when 16#01C5E# => romdata <= X"20637574";
    when 16#01C5F# => romdata <= X"74656400";
    when 16#01C60# => romdata <= X"0A202063";
    when 16#01C61# => romdata <= X"68616E6E";
    when 16#01C62# => romdata <= X"656C2032";
    when 16#01C63# => romdata <= X"20646976";
    when 16#01C64# => romdata <= X"6964656E";
    when 16#01C65# => romdata <= X"64206375";
    when 16#01C66# => romdata <= X"74746564";
    when 16#01C67# => romdata <= X"00000000";
    when 16#01C68# => romdata <= X"0A202063";
    when 16#01C69# => romdata <= X"68616E6E";
    when 16#01C6A# => romdata <= X"656C2032";
    when 16#01C6B# => romdata <= X"206E6F69";
    when 16#01C6C# => romdata <= X"73652063";
    when 16#01C6D# => romdata <= X"6F6D7065";
    when 16#01C6E# => romdata <= X"6E736174";
    when 16#01C6F# => romdata <= X"696F6E20";
    when 16#01C70# => romdata <= X"746F2062";
    when 16#01C71# => romdata <= X"69670000";
    when 16#01C72# => romdata <= X"0A202063";
    when 16#01C73# => romdata <= X"68616E6E";
    when 16#01C74# => romdata <= X"656C2032";
    when 16#01C75# => romdata <= X"206E6F69";
    when 16#01C76# => romdata <= X"73652076";
    when 16#01C77# => romdata <= X"616C7565";
    when 16#01C78# => romdata <= X"20637574";
    when 16#01C79# => romdata <= X"74656400";
    when 16#01C7A# => romdata <= X"0A202063";
    when 16#01C7B# => romdata <= X"68616E6E";
    when 16#01C7C# => romdata <= X"656C2031";
    when 16#01C7D# => romdata <= X"20646976";
    when 16#01C7E# => romdata <= X"6964656E";
    when 16#01C7F# => romdata <= X"64206375";
    when 16#01C80# => romdata <= X"74746564";
    when 16#01C81# => romdata <= X"00000000";
    when 16#01C82# => romdata <= X"0A202063";
    when 16#01C83# => romdata <= X"68616E6E";
    when 16#01C84# => romdata <= X"656C2031";
    when 16#01C85# => romdata <= X"206E6F69";
    when 16#01C86# => romdata <= X"73652063";
    when 16#01C87# => romdata <= X"6F6D7065";
    when 16#01C88# => romdata <= X"6E736174";
    when 16#01C89# => romdata <= X"696F6E20";
    when 16#01C8A# => romdata <= X"746F2062";
    when 16#01C8B# => romdata <= X"69670000";
    when 16#01C8C# => romdata <= X"0A202063";
    when 16#01C8D# => romdata <= X"68616E6E";
    when 16#01C8E# => romdata <= X"656C2031";
    when 16#01C8F# => romdata <= X"206E6F69";
    when 16#01C90# => romdata <= X"73652076";
    when 16#01C91# => romdata <= X"616C7565";
    when 16#01C92# => romdata <= X"20637574";
    when 16#01C93# => romdata <= X"74656400";
    when 16#01C94# => romdata <= X"0A202063";
    when 16#01C95# => romdata <= X"68616E6E";
    when 16#01C96# => romdata <= X"656C2030";
    when 16#01C97# => romdata <= X"20646976";
    when 16#01C98# => romdata <= X"6964656E";
    when 16#01C99# => romdata <= X"64206375";
    when 16#01C9A# => romdata <= X"74746564";
    when 16#01C9B# => romdata <= X"00000000";
    when 16#01C9C# => romdata <= X"0A202063";
    when 16#01C9D# => romdata <= X"68616E6E";
    when 16#01C9E# => romdata <= X"656C2030";
    when 16#01C9F# => romdata <= X"206E6F69";
    when 16#01CA0# => romdata <= X"73652063";
    when 16#01CA1# => romdata <= X"6F6D7065";
    when 16#01CA2# => romdata <= X"6E736174";
    when 16#01CA3# => romdata <= X"696F6E20";
    when 16#01CA4# => romdata <= X"746F2062";
    when 16#01CA5# => romdata <= X"69670000";
    when 16#01CA6# => romdata <= X"0A202063";
    when 16#01CA7# => romdata <= X"68616E6E";
    when 16#01CA8# => romdata <= X"656C2030";
    when 16#01CA9# => romdata <= X"206E6F69";
    when 16#01CAA# => romdata <= X"73652076";
    when 16#01CAB# => romdata <= X"616C7565";
    when 16#01CAC# => romdata <= X"20637574";
    when 16#01CAD# => romdata <= X"74656400";
    when 16#01CAE# => romdata <= X"0A202073";
    when 16#01CAF# => romdata <= X"6F667477";
    when 16#01CB0# => romdata <= X"61726520";
    when 16#01CB1# => romdata <= X"6572726F";
    when 16#01CB2# => romdata <= X"72000000";
    when 16#01CB3# => romdata <= X"0A657874";
    when 16#01CB4# => romdata <= X"65726E61";
    when 16#01CB5# => romdata <= X"6C20636C";
    when 16#01CB6# => romdata <= X"6F636B20";
    when 16#01CB7# => romdata <= X"20202020";
    when 16#01CB8# => romdata <= X"2020203A";
    when 16#01CB9# => romdata <= X"20000000";
    when 16#01CBA# => romdata <= X"61637469";
    when 16#01CBB# => romdata <= X"76650000";
    when 16#01CBC# => romdata <= X"0A6D6963";
    when 16#01CBD# => romdata <= X"726F7075";
    when 16#01CBE# => romdata <= X"6C736520";
    when 16#01CBF# => romdata <= X"736F7572";
    when 16#01CC0# => romdata <= X"63652020";
    when 16#01CC1# => romdata <= X"2020203A";
    when 16#01CC2# => romdata <= X"20000000";
    when 16#01CC3# => romdata <= X"0A6D6963";
    when 16#01CC4# => romdata <= X"726F7075";
    when 16#01CC5# => romdata <= X"6C736520";
    when 16#01CC6# => romdata <= X"6576656E";
    when 16#01CC7# => romdata <= X"74206C69";
    when 16#01CC8# => romdata <= X"6D69743A";
    when 16#01CC9# => romdata <= X"20000000";
    when 16#01CCA# => romdata <= X"0A6D6561";
    when 16#01CCB# => romdata <= X"73757265";
    when 16#01CCC# => romdata <= X"6D656E74";
    when 16#01CCD# => romdata <= X"206C656E";
    when 16#01CCE# => romdata <= X"67746820";
    when 16#01CCF# => romdata <= X"2020203A";
    when 16#01CD0# => romdata <= X"20000000";
    when 16#01CD1# => romdata <= X"0A626561";
    when 16#01CD2# => romdata <= X"6D20706F";
    when 16#01CD3# => romdata <= X"73697469";
    when 16#01CD4# => romdata <= X"6F6E206D";
    when 16#01CD5# => romdata <= X"6F6E6974";
    when 16#01CD6# => romdata <= X"6F722072";
    when 16#01CD7# => romdata <= X"65676973";
    when 16#01CD8# => romdata <= X"74657273";
    when 16#01CD9# => romdata <= X"00000000";
    when 16#01CDA# => romdata <= X"0A202020";
    when 16#01CDB# => romdata <= X"20202020";
    when 16#01CDC# => romdata <= X"20202020";
    when 16#01CDD# => romdata <= X"20202020";
    when 16#01CDE# => romdata <= X"20202020";
    when 16#01CDF# => romdata <= X"20202020";
    when 16#01CE0# => romdata <= X"20636861";
    when 16#01CE1# => romdata <= X"6E6E656C";
    when 16#01CE2# => romdata <= X"20302020";
    when 16#01CE3# => romdata <= X"20636861";
    when 16#01CE4# => romdata <= X"6E6E656C";
    when 16#01CE5# => romdata <= X"20312020";
    when 16#01CE6# => romdata <= X"20636861";
    when 16#01CE7# => romdata <= X"6E6E656C";
    when 16#01CE8# => romdata <= X"20322020";
    when 16#01CE9# => romdata <= X"20636861";
    when 16#01CEA# => romdata <= X"6E6E656C";
    when 16#01CEB# => romdata <= X"20330000";
    when 16#01CEC# => romdata <= X"0A202020";
    when 16#01CED# => romdata <= X"20202020";
    when 16#01CEE# => romdata <= X"20202020";
    when 16#01CEF# => romdata <= X"20202020";
    when 16#01CF0# => romdata <= X"20202020";
    when 16#01CF1# => romdata <= X"20202020";
    when 16#01CF2# => romdata <= X"202D2D2D";
    when 16#01CF3# => romdata <= X"2D20686F";
    when 16#01CF4# => romdata <= X"72697A6F";
    when 16#01CF5# => romdata <= X"6E74616C";
    when 16#01CF6# => romdata <= X"202D2D2D";
    when 16#01CF7# => romdata <= X"2D2D2020";
    when 16#01CF8# => romdata <= X"202D2D2D";
    when 16#01CF9# => romdata <= X"2D2D2D20";
    when 16#01CFA# => romdata <= X"76657274";
    when 16#01CFB# => romdata <= X"6963616C";
    when 16#01CFC# => romdata <= X"202D2D2D";
    when 16#01CFD# => romdata <= X"2D2D0000";
    when 16#01CFE# => romdata <= X"0A736361";
    when 16#01CFF# => romdata <= X"6C657220";
    when 16#01D00# => romdata <= X"76616C75";
    when 16#01D01# => romdata <= X"65732020";
    when 16#01D02# => romdata <= X"20202020";
    when 16#01D03# => romdata <= X"20202020";
    when 16#01D04# => romdata <= X"20000000";
    when 16#01D05# => romdata <= X"0A6E6F69";
    when 16#01D06# => romdata <= X"73652063";
    when 16#01D07# => romdata <= X"6F6D7065";
    when 16#01D08# => romdata <= X"6E736174";
    when 16#01D09# => romdata <= X"696F6E20";
    when 16#01D0A# => romdata <= X"20202020";
    when 16#01D0B# => romdata <= X"20000000";
    when 16#01D0C# => romdata <= X"0A6D6561";
    when 16#01D0D# => romdata <= X"73757265";
    when 16#01D0E# => romdata <= X"6D656E74";
    when 16#01D0F# => romdata <= X"20202020";
    when 16#01D10# => romdata <= X"20202020";
    when 16#01D11# => romdata <= X"20202020";
    when 16#01D12# => romdata <= X"20000000";
    when 16#01D13# => romdata <= X"0A73616D";
    when 16#01D14# => romdata <= X"706C6573";
    when 16#01D15# => romdata <= X"20286469";
    when 16#01D16# => romdata <= X"76292020";
    when 16#01D17# => romdata <= X"20202020";
    when 16#01D18# => romdata <= X"3A200000";
    when 16#01D19# => romdata <= X"0A73756D";
    when 16#01D1A# => romdata <= X"20636861";
    when 16#01D1B# => romdata <= X"6E6E656C";
    when 16#01D1C# => romdata <= X"20736361";
    when 16#01D1D# => romdata <= X"6C657220";
    when 16#01D1E# => romdata <= X"3A200000";
    when 16#01D1F# => romdata <= X"0A73756D";
    when 16#01D20# => romdata <= X"20636861";
    when 16#01D21# => romdata <= X"6E6E656C";
    when 16#01D22# => romdata <= X"20202020";
    when 16#01D23# => romdata <= X"20202020";
    when 16#01D24# => romdata <= X"3A200000";
    when 16#01D25# => romdata <= X"0A0A706F";
    when 16#01D26# => romdata <= X"73697469";
    when 16#01D27# => romdata <= X"6F6E2063";
    when 16#01D28# => romdata <= X"6F6D7075";
    when 16#01D29# => romdata <= X"74617469";
    when 16#01D2A# => romdata <= X"6F6E0000";
    when 16#01D2B# => romdata <= X"0A202073";
    when 16#01D2C# => romdata <= X"63616C65";
    when 16#01D2D# => romdata <= X"72207661";
    when 16#01D2E# => romdata <= X"6C756573";
    when 16#01D2F# => romdata <= X"20202020";
    when 16#01D30# => romdata <= X"20202020";
    when 16#01D31# => romdata <= X"20000000";
    when 16#01D32# => romdata <= X"0A20206F";
    when 16#01D33# => romdata <= X"66667365";
    when 16#01D34# => romdata <= X"74202020";
    when 16#01D35# => romdata <= X"20202020";
    when 16#01D36# => romdata <= X"20202020";
    when 16#01D37# => romdata <= X"20202020";
    when 16#01D38# => romdata <= X"20000000";
    when 16#01D39# => romdata <= X"0A6F7574";
    when 16#01D3A# => romdata <= X"70757420";
    when 16#01D3B# => romdata <= X"73656C65";
    when 16#01D3C# => romdata <= X"6374203A";
    when 16#01D3D# => romdata <= X"20000000";
    when 16#01D3E# => romdata <= X"64697265";
    when 16#01D3F# => romdata <= X"6374206D";
    when 16#01D40# => romdata <= X"6F646500";
    when 16#01D41# => romdata <= X"0A63616C";
    when 16#01D42# => romdata <= X"63207374";
    when 16#01D43# => romdata <= X"61746520";
    when 16#01D44# => romdata <= X"2020203A";
    when 16#01D45# => romdata <= X"20307800";
    when 16#01D46# => romdata <= X"76657274";
    when 16#01D47# => romdata <= X"6963616C";
    when 16#01D48# => romdata <= X"00000000";
    when 16#01D49# => romdata <= X"686F7269";
    when 16#01D4A# => romdata <= X"7A6F6E74";
    when 16#01D4B# => romdata <= X"616C0000";
    when 16#01D4C# => romdata <= X"73756D00";
    when 16#01D4D# => romdata <= X"6368616E";
    when 16#01D4E# => romdata <= X"6E656C20";
    when 16#01D4F# => romdata <= X"33000000";
    when 16#01D50# => romdata <= X"6368616E";
    when 16#01D51# => romdata <= X"6E656C20";
    when 16#01D52# => romdata <= X"32000000";
    when 16#01D53# => romdata <= X"6368616E";
    when 16#01D54# => romdata <= X"6E656C20";
    when 16#01D55# => romdata <= X"31000000";
    when 16#01D56# => romdata <= X"6368616E";
    when 16#01D57# => romdata <= X"6E656C20";
    when 16#01D58# => romdata <= X"30000000";
    when 16#01D59# => romdata <= X"636C6B3A";
    when 16#01D5A# => romdata <= X"20000000";
    when 16#01D5B# => romdata <= X"494E5400";
    when 16#01D5C# => romdata <= X"6D70756C";
    when 16#01D5D# => romdata <= X"733A2000";
    when 16#01D5E# => romdata <= X"65787400";
    when 16#01D5F# => romdata <= X"0A6D6561";
    when 16#01D60# => romdata <= X"732E206C";
    when 16#01D61# => romdata <= X"656E6774";
    when 16#01D62# => romdata <= X"683A2000";
    when 16#01D63# => romdata <= X"0A636830";
    when 16#01D64# => romdata <= X"3A200000";
    when 16#01D65# => romdata <= X"6368313A";
    when 16#01D66# => romdata <= X"20000000";
    when 16#01D67# => romdata <= X"0A636832";
    when 16#01D68# => romdata <= X"3A200000";
    when 16#01D69# => romdata <= X"6368333A";
    when 16#01D6A# => romdata <= X"20000000";
    when 16#01D6B# => romdata <= X"0A73706C";
    when 16#01D6C# => romdata <= X"3A200000";
    when 16#01D6D# => romdata <= X"73756D3A";
    when 16#01D6E# => romdata <= X"20000000";
    when 16#01D6F# => romdata <= X"0A6F7574";
    when 16#01D70# => romdata <= X"7075743A";
    when 16#01D71# => romdata <= X"20000000";
    when 16#01D72# => romdata <= X"7467656E";
    when 16#01D73# => romdata <= X"00000000";
    when 16#01D74# => romdata <= X"0A63616C";
    when 16#01D75# => romdata <= X"63207374";
    when 16#01D76# => romdata <= X"6174653A";
    when 16#01D77# => romdata <= X"20000000";
    when 16#01D78# => romdata <= X"63683320";
    when 16#01D79# => romdata <= X"696E7020";
    when 16#01D7A# => romdata <= X"6F762020";
    when 16#01D7B# => romdata <= X"00000000";
    when 16#01D7C# => romdata <= X"63683220";
    when 16#01D7D# => romdata <= X"696E7020";
    when 16#01D7E# => romdata <= X"6F762020";
    when 16#01D7F# => romdata <= X"00000000";
    when 16#01D80# => romdata <= X"63683120";
    when 16#01D81# => romdata <= X"696E7020";
    when 16#01D82# => romdata <= X"6F762020";
    when 16#01D83# => romdata <= X"00000000";
    when 16#01D84# => romdata <= X"63683020";
    when 16#01D85# => romdata <= X"696E7020";
    when 16#01D86# => romdata <= X"6F762020";
    when 16#01D87# => romdata <= X"00000000";
    when 16#01D88# => romdata <= X"63683320";
    when 16#01D89# => romdata <= X"73756D20";
    when 16#01D8A# => romdata <= X"6F762020";
    when 16#01D8B# => romdata <= X"00000000";
    when 16#01D8C# => romdata <= X"63683220";
    when 16#01D8D# => romdata <= X"73756D20";
    when 16#01D8E# => romdata <= X"6F762020";
    when 16#01D8F# => romdata <= X"00000000";
    when 16#01D90# => romdata <= X"63683120";
    when 16#01D91# => romdata <= X"73756D20";
    when 16#01D92# => romdata <= X"6F762020";
    when 16#01D93# => romdata <= X"00000000";
    when 16#01D94# => romdata <= X"63683020";
    when 16#01D95# => romdata <= X"73756D20";
    when 16#01D96# => romdata <= X"6F762020";
    when 16#01D97# => romdata <= X"00000000";
    when 16#01D98# => romdata <= X"73756D20";
    when 16#01D99# => romdata <= X"73636C20";
    when 16#01D9A# => romdata <= X"6F762020";
    when 16#01D9B# => romdata <= X"00000000";
    when 16#01D9C# => romdata <= X"73756D20";
    when 16#01D9D# => romdata <= X"63757420";
    when 16#01D9E# => romdata <= X"20000000";
    when 16#01D9F# => romdata <= X"63683320";
    when 16#01DA0# => romdata <= X"64697620";
    when 16#01DA1# => romdata <= X"63757420";
    when 16#01DA2# => romdata <= X"20000000";
    when 16#01DA3# => romdata <= X"63683320";
    when 16#01DA4# => romdata <= X"6E736520";
    when 16#01DA5# => romdata <= X"636D7020";
    when 16#01DA6# => romdata <= X"20000000";
    when 16#01DA7# => romdata <= X"63683320";
    when 16#01DA8# => romdata <= X"6E736520";
    when 16#01DA9# => romdata <= X"63757420";
    when 16#01DAA# => romdata <= X"20000000";
    when 16#01DAB# => romdata <= X"63683220";
    when 16#01DAC# => romdata <= X"64697620";
    when 16#01DAD# => romdata <= X"63757420";
    when 16#01DAE# => romdata <= X"20000000";
    when 16#01DAF# => romdata <= X"63683220";
    when 16#01DB0# => romdata <= X"6E736520";
    when 16#01DB1# => romdata <= X"636D7020";
    when 16#01DB2# => romdata <= X"20000000";
    when 16#01DB3# => romdata <= X"63683220";
    when 16#01DB4# => romdata <= X"6E736520";
    when 16#01DB5# => romdata <= X"63757420";
    when 16#01DB6# => romdata <= X"20000000";
    when 16#01DB7# => romdata <= X"63683120";
    when 16#01DB8# => romdata <= X"64697620";
    when 16#01DB9# => romdata <= X"63757420";
    when 16#01DBA# => romdata <= X"20000000";
    when 16#01DBB# => romdata <= X"63683120";
    when 16#01DBC# => romdata <= X"6E736520";
    when 16#01DBD# => romdata <= X"636D7020";
    when 16#01DBE# => romdata <= X"20000000";
    when 16#01DBF# => romdata <= X"63683120";
    when 16#01DC0# => romdata <= X"6E736520";
    when 16#01DC1# => romdata <= X"63757420";
    when 16#01DC2# => romdata <= X"20000000";
    when 16#01DC3# => romdata <= X"63683020";
    when 16#01DC4# => romdata <= X"64697620";
    when 16#01DC5# => romdata <= X"63757420";
    when 16#01DC6# => romdata <= X"20000000";
    when 16#01DC7# => romdata <= X"63683020";
    when 16#01DC8# => romdata <= X"6E736520";
    when 16#01DC9# => romdata <= X"636D7020";
    when 16#01DCA# => romdata <= X"20000000";
    when 16#01DCB# => romdata <= X"63683020";
    when 16#01DCC# => romdata <= X"6E736520";
    when 16#01DCD# => romdata <= X"63757420";
    when 16#01DCE# => romdata <= X"20000000";
    when 16#01DCF# => romdata <= X"736F6674";
    when 16#01DD0# => romdata <= X"20657272";
    when 16#01DD1# => romdata <= X"20200000";
    when 16#01DD2# => romdata <= X"0000350D";
    when 16#01DD3# => romdata <= X"00003503";
    when 16#01DD4# => romdata <= X"000034F9";
    when 16#01DD5# => romdata <= X"000034EF";
    when 16#01DD6# => romdata <= X"000034E5";
    when 16#01DD7# => romdata <= X"000034DC";
    when 16#01DD8# => romdata <= X"000034D3";
    when 16#01DD9# => romdata <= X"00003676";
    when 16#01DDA# => romdata <= X"000039D3";
    when 16#01DDB# => romdata <= X"000039C9";
    when 16#01DDC# => romdata <= X"000039BF";
    when 16#01DDD# => romdata <= X"000039B5";
    when 16#01DDE# => romdata <= X"000039AB";
    when 16#01DDF# => romdata <= X"000039A1";
    when 16#01DE0# => romdata <= X"0A202044";
    when 16#01DE1# => romdata <= X"434D2061";
    when 16#01DE2# => romdata <= X"63746976";
    when 16#01DE3# => romdata <= X"65000000";
    when 16#01DE4# => romdata <= X"0A202044";
    when 16#01DE5# => romdata <= X"434D204E";
    when 16#01DE6# => romdata <= X"4F542061";
    when 16#01DE7# => romdata <= X"63746976";
    when 16#01DE8# => romdata <= X"65000000";
    when 16#01DE9# => romdata <= X"0A202075";
    when 16#01DEA# => romdata <= X"70706572";
    when 16#01DEB# => romdata <= X"20626F75";
    when 16#01DEC# => romdata <= X"6E64206F";
    when 16#01DED# => romdata <= X"76657266";
    when 16#01DEE# => romdata <= X"6C6F7700";
    when 16#01DEF# => romdata <= X"0A20206C";
    when 16#01DF0# => romdata <= X"6F776572";
    when 16#01DF1# => romdata <= X"20626F75";
    when 16#01DF2# => romdata <= X"6E642075";
    when 16#01DF3# => romdata <= X"6E646572";
    when 16#01DF4# => romdata <= X"666C6F77";
    when 16#01DF5# => romdata <= X"00000000";
    when 16#01DF6# => romdata <= X"0A202063";
    when 16#01DF7# => romdata <= X"6F6E6E65";
    when 16#01DF8# => romdata <= X"6374696F";
    when 16#01DF9# => romdata <= X"6E206C6F";
    when 16#01DFA# => romdata <= X"73740000";
    when 16#01DFB# => romdata <= X"0A202074";
    when 16#01DFC# => romdata <= X"696D656F";
    when 16#01DFD# => romdata <= X"75740000";
    when 16#01DFE# => romdata <= X"0A646174";
    when 16#01DFF# => romdata <= X"6120696E";
    when 16#01E00# => romdata <= X"20202020";
    when 16#01E01# => romdata <= X"203A2000";
    when 16#01E02# => romdata <= X"0A73756D";
    when 16#01E03# => romdata <= X"20696E20";
    when 16#01E04# => romdata <= X"20202020";
    when 16#01E05# => romdata <= X"203A2000";
    when 16#01E06# => romdata <= X"0A617665";
    when 16#01E07# => romdata <= X"72616765";
    when 16#01E08# => romdata <= X"20202020";
    when 16#01E09# => romdata <= X"203A2000";
    when 16#01E0A# => romdata <= X"0A6C6F77";
    when 16#01E0B# => romdata <= X"65722062";
    when 16#01E0C# => romdata <= X"6F756E64";
    when 16#01E0D# => romdata <= X"203A2000";
    when 16#01E0E# => romdata <= X"0A757070";
    when 16#01E0F# => romdata <= X"65722062";
    when 16#01E10# => romdata <= X"6F756E64";
    when 16#01E11# => romdata <= X"203A2000";
    when 16#01E12# => romdata <= X"0A737461";
    when 16#01E13# => romdata <= X"74652020";
    when 16#01E14# => romdata <= X"20202020";
    when 16#01E15# => romdata <= X"203A2030";
    when 16#01E16# => romdata <= X"78000000";
    when 16#01E17# => romdata <= X"0A307800";
    when 16#01E18# => romdata <= X"786D6F64";
    when 16#01E19# => romdata <= X"656D2074";
    when 16#01E1A# => romdata <= X"72616E73";
    when 16#01E1B# => romdata <= X"6D69742E";
    when 16#01E1C# => romdata <= X"2E2E0A00";
    when 16#01E1D# => romdata <= X"20627974";
    when 16#01E1E# => romdata <= X"65732074";
    when 16#01E1F# => romdata <= X"72616E73";
    when 16#01E20# => romdata <= X"6D697474";
    when 16#01E21# => romdata <= X"65640A00";
    when 16#01E22# => romdata <= X"63616E63";
    when 16#01E23# => romdata <= X"656C0A00";
    when 16#01E24# => romdata <= X"72657472";
    when 16#01E25# => romdata <= X"79206F75";
    when 16#01E26# => romdata <= X"740A0000";
    when 16#01E27# => romdata <= X"786D6F64";
    when 16#01E28# => romdata <= X"656D2072";
    when 16#01E29# => romdata <= X"65636569";
    when 16#01E2A# => romdata <= X"76652E2E";
    when 16#01E2B# => romdata <= X"2E0A0000";
    when 16#01E2C# => romdata <= X"20627974";
    when 16#01E2D# => romdata <= X"65732072";
    when 16#01E2E# => romdata <= X"65636569";
    when 16#01E2F# => romdata <= X"7665640A";
    when 16#01E30# => romdata <= X"00000000";
    when 16#01E31# => romdata <= X"72782062";
    when 16#01E32# => romdata <= X"75666665";
    when 16#01E33# => romdata <= X"72206675";
    when 16#01E34# => romdata <= X"6C6C0A00";
    when 16#01E35# => romdata <= X"74696D65";
    when 16#01E36# => romdata <= X"206F7574";
    when 16#01E37# => romdata <= X"0A000000";
    when 16#01E38# => romdata <= X"64656275";
    when 16#01E39# => romdata <= X"67207265";
    when 16#01E3A# => romdata <= X"67697374";
    when 16#01E3B# => romdata <= X"65727300";
    when 16#01E3C# => romdata <= X"0A6D6F64";
    when 16#01E3D# => romdata <= X"65202020";
    when 16#01E3E# => romdata <= X"20202020";
    when 16#01E3F# => romdata <= X"203A2000";
    when 16#01E40# => romdata <= X"0A616464";
    when 16#01E41# => romdata <= X"72657373";
    when 16#01E42# => romdata <= X"20302020";
    when 16#01E43# => romdata <= X"203A2030";
    when 16#01E44# => romdata <= X"78000000";
    when 16#01E45# => romdata <= X"0A616464";
    when 16#01E46# => romdata <= X"72657373";
    when 16#01E47# => romdata <= X"20312020";
    when 16#01E48# => romdata <= X"203A2030";
    when 16#01E49# => romdata <= X"78000000";
    when 16#01E4A# => romdata <= X"0A627566";
    when 16#01E4B# => romdata <= X"66657220";
    when 16#01E4C# => romdata <= X"73697A65";
    when 16#01E4D# => romdata <= X"203A2000";
    when 16#01E4E# => romdata <= X"0A646562";
    when 16#01E4F# => romdata <= X"75672074";
    when 16#01E50# => romdata <= X"72616365";
    when 16#01E51# => romdata <= X"206D656D";
    when 16#01E52# => romdata <= X"6F727900";
    when 16#01E53# => romdata <= X"0A74696D";
    when 16#01E54# => romdata <= X"65207374";
    when 16#01E55# => romdata <= X"616D7020";
    when 16#01E56# => romdata <= X"20202073";
    when 16#01E57# => romdata <= X"74617465";
    when 16#01E58# => romdata <= X"00000000";
    when 16#01E59# => romdata <= X"20203078";
    when 16#01E5A# => romdata <= X"00000000";
    when 16#01E5B# => romdata <= X"6D61783A";
    when 16#01E5C# => romdata <= X"20000000";
    when 16#01E5D# => romdata <= X"6D696E3A";
    when 16#01E5E# => romdata <= X"20000000";
    when 16#01E5F# => romdata <= X"63683A20";
    when 16#01E60# => romdata <= X"00000000";
    when 16#01E61# => romdata <= X"73706C3A";
    when 16#01E62# => romdata <= X"20000000";
    when 16#01E63# => romdata <= X"30622020";
    when 16#01E64# => romdata <= X"20202020";
    when 16#01E65# => romdata <= X"20202020";
    when 16#01E66# => romdata <= X"20202020";
    when 16#01E67# => romdata <= X"20202020";
    when 16#01E68# => romdata <= X"20202020";
    when 16#01E69# => romdata <= X"20202020";
    when 16#01E6A# => romdata <= X"20202020";
    when 16#01E6B# => romdata <= X"20200000";
    when 16#01E6C# => romdata <= X"20202020";
    when 16#01E6D# => romdata <= X"20202020";
    when 16#01E6E# => romdata <= X"00000000";
    when 16#01E6F# => romdata <= X"00202020";
    when 16#01E70# => romdata <= X"20202020";
    when 16#01E71# => romdata <= X"20202828";
    when 16#01E72# => romdata <= X"28282820";
    when 16#01E73# => romdata <= X"20202020";
    when 16#01E74# => romdata <= X"20202020";
    when 16#01E75# => romdata <= X"20202020";
    when 16#01E76# => romdata <= X"20202020";
    when 16#01E77# => romdata <= X"20881010";
    when 16#01E78# => romdata <= X"10101010";
    when 16#01E79# => romdata <= X"10101010";
    when 16#01E7A# => romdata <= X"10101010";
    when 16#01E7B# => romdata <= X"10040404";
    when 16#01E7C# => romdata <= X"04040404";
    when 16#01E7D# => romdata <= X"04040410";
    when 16#01E7E# => romdata <= X"10101010";
    when 16#01E7F# => romdata <= X"10104141";
    when 16#01E80# => romdata <= X"41414141";
    when 16#01E81# => romdata <= X"01010101";
    when 16#01E82# => romdata <= X"01010101";
    when 16#01E83# => romdata <= X"01010101";
    when 16#01E84# => romdata <= X"01010101";
    when 16#01E85# => romdata <= X"01010101";
    when 16#01E86# => romdata <= X"10101010";
    when 16#01E87# => romdata <= X"10104242";
    when 16#01E88# => romdata <= X"42424242";
    when 16#01E89# => romdata <= X"02020202";
    when 16#01E8A# => romdata <= X"02020202";
    when 16#01E8B# => romdata <= X"02020202";
    when 16#01E8C# => romdata <= X"02020202";
    when 16#01E8D# => romdata <= X"02020202";
    when 16#01E8E# => romdata <= X"10101010";
    when 16#01E8F# => romdata <= X"20000000";
    when 16#01E90# => romdata <= X"00000000";
    when 16#01E91# => romdata <= X"00000000";
    when 16#01E92# => romdata <= X"00000000";
    when 16#01E93# => romdata <= X"00000000";
    when 16#01E94# => romdata <= X"00000000";
    when 16#01E95# => romdata <= X"00000000";
    when 16#01E96# => romdata <= X"00000000";
    when 16#01E97# => romdata <= X"00000000";
    when 16#01E98# => romdata <= X"00000000";
    when 16#01E99# => romdata <= X"00000000";
    when 16#01E9A# => romdata <= X"00000000";
    when 16#01E9B# => romdata <= X"00000000";
    when 16#01E9C# => romdata <= X"00000000";
    when 16#01E9D# => romdata <= X"00000000";
    when 16#01E9E# => romdata <= X"00000000";
    when 16#01E9F# => romdata <= X"00000000";
    when 16#01EA0# => romdata <= X"00000000";
    when 16#01EA1# => romdata <= X"00000000";
    when 16#01EA2# => romdata <= X"00000000";
    when 16#01EA3# => romdata <= X"00000000";
    when 16#01EA4# => romdata <= X"00000000";
    when 16#01EA5# => romdata <= X"00000000";
    when 16#01EA6# => romdata <= X"00000000";
    when 16#01EA7# => romdata <= X"00000000";
    when 16#01EA8# => romdata <= X"00000000";
    when 16#01EA9# => romdata <= X"00000000";
    when 16#01EAA# => romdata <= X"00000000";
    when 16#01EAB# => romdata <= X"00000000";
    when 16#01EAC# => romdata <= X"00000000";
    when 16#01EAD# => romdata <= X"00000000";
    when 16#01EAE# => romdata <= X"00000000";
    when 16#01EAF# => romdata <= X"00000000";
    when 16#01EB0# => romdata <= X"80000C00";
    when 16#01EB1# => romdata <= X"00000000";
    when 16#01EB2# => romdata <= X"80000900";
    when 16#01EB3# => romdata <= X"80000800";
    when 16#01EB4# => romdata <= X"00000000";
    when 16#01EB5# => romdata <= X"00000000";
    when 16#01EB6# => romdata <= X"FF000000";
    when 16#01EB7# => romdata <= X"00000000";
    when 16#01EB8# => romdata <= X"80000B00";
    when 16#01EB9# => romdata <= X"00FFFFFF";
    when 16#01EBA# => romdata <= X"FF00FFFF";
    when 16#01EBB# => romdata <= X"FFFF00FF";
    when 16#01EBC# => romdata <= X"FFFFFF00";
    when 16#01EBD# => romdata <= X"00000000";
    when 16#01EBE# => romdata <= X"00000000";
    when 16#01EBF# => romdata <= X"80000F00";
    when 16#01EC0# => romdata <= X"80000A00";
    when 16#01EC1# => romdata <= X"80000700";
    when 16#01EC2# => romdata <= X"80000600";
    when 16#01EC3# => romdata <= X"80000400";
    when 16#01EC4# => romdata <= X"80000200";
    when 16#01EC5# => romdata <= X"80000100";
    when 16#01EC6# => romdata <= X"80000004";
    when 16#01EC7# => romdata <= X"80000000";
    when 16#01EC8# => romdata <= X"00007B24";
    when 16#01EC9# => romdata <= X"00000000";
    when 16#01ECA# => romdata <= X"00007D8C";
    when 16#01ECB# => romdata <= X"00007DE8";
    when 16#01ECC# => romdata <= X"00007E44";
    when 16#01ECD# => romdata <= X"00000000";
    when 16#01ECE# => romdata <= X"00000000";
    when 16#01ECF# => romdata <= X"00000000";
    when 16#01ED0# => romdata <= X"00000000";
    when 16#01ED1# => romdata <= X"00000000";
    when 16#01ED2# => romdata <= X"00000000";
    when 16#01ED3# => romdata <= X"00000000";
    when 16#01ED4# => romdata <= X"00000000";
    when 16#01ED5# => romdata <= X"00000000";
    when 16#01ED6# => romdata <= X"00006838";
    when 16#01ED7# => romdata <= X"00000000";
    when 16#01ED8# => romdata <= X"00000000";
    when 16#01ED9# => romdata <= X"00000000";
    when 16#01EDA# => romdata <= X"00000000";
    when 16#01EDB# => romdata <= X"00000000";
    when 16#01EDC# => romdata <= X"00000000";
    when 16#01EDD# => romdata <= X"00000000";
    when 16#01EDE# => romdata <= X"00000000";
    when 16#01EDF# => romdata <= X"00000000";
    when 16#01EE0# => romdata <= X"00000000";
    when 16#01EE1# => romdata <= X"00000000";
    when 16#01EE2# => romdata <= X"00000000";
    when 16#01EE3# => romdata <= X"00000000";
    when 16#01EE4# => romdata <= X"00000000";
    when 16#01EE5# => romdata <= X"00000000";
    when 16#01EE6# => romdata <= X"00000000";
    when 16#01EE7# => romdata <= X"00000000";
    when 16#01EE8# => romdata <= X"00000000";
    when 16#01EE9# => romdata <= X"00000000";
    when 16#01EEA# => romdata <= X"00000000";
    when 16#01EEB# => romdata <= X"00000000";
    when 16#01EEC# => romdata <= X"00000000";
    when 16#01EED# => romdata <= X"00000000";
    when 16#01EEE# => romdata <= X"00000000";
    when 16#01EEF# => romdata <= X"00000000";
    when 16#01EF0# => romdata <= X"00000000";
    when 16#01EF1# => romdata <= X"00000000";
    when 16#01EF2# => romdata <= X"00000000";
    when 16#01EF3# => romdata <= X"00000001";
    when 16#01EF4# => romdata <= X"330EABCD";
    when 16#01EF5# => romdata <= X"1234E66D";
    when 16#01EF6# => romdata <= X"DEEC0005";
    when 16#01EF7# => romdata <= X"000B0000";
    when 16#01EF8# => romdata <= X"00000000";
    when 16#01EF9# => romdata <= X"00000000";
    when 16#01EFA# => romdata <= X"00000000";
    when 16#01EFB# => romdata <= X"00000000";
    when 16#01EFC# => romdata <= X"00000000";
    when 16#01EFD# => romdata <= X"00000000";
    when 16#01EFE# => romdata <= X"00000000";
    when 16#01EFF# => romdata <= X"00000000";
    when 16#01F00# => romdata <= X"00000000";
    when 16#01F01# => romdata <= X"00000000";
    when 16#01F02# => romdata <= X"00000000";
    when 16#01F03# => romdata <= X"00000000";
    when 16#01F04# => romdata <= X"00000000";
    when 16#01F05# => romdata <= X"00000000";
    when 16#01F06# => romdata <= X"00000000";
    when 16#01F07# => romdata <= X"00000000";
    when 16#01F08# => romdata <= X"00000000";
    when 16#01F09# => romdata <= X"00000000";
    when 16#01F0A# => romdata <= X"00000000";
    when 16#01F0B# => romdata <= X"00000000";
    when 16#01F0C# => romdata <= X"00000000";
    when 16#01F0D# => romdata <= X"00000000";
    when 16#01F0E# => romdata <= X"00000000";
    when 16#01F0F# => romdata <= X"00000000";
    when 16#01F10# => romdata <= X"00000000";
    when 16#01F11# => romdata <= X"00000000";
    when 16#01F12# => romdata <= X"00000000";
    when 16#01F13# => romdata <= X"00000000";
    when 16#01F14# => romdata <= X"00000000";
    when 16#01F15# => romdata <= X"00000000";
    when 16#01F16# => romdata <= X"00000000";
    when 16#01F17# => romdata <= X"00000000";
    when 16#01F18# => romdata <= X"00000000";
    when 16#01F19# => romdata <= X"00000000";
    when 16#01F1A# => romdata <= X"00000000";
    when 16#01F1B# => romdata <= X"00000000";
    when 16#01F1C# => romdata <= X"00000000";
    when 16#01F1D# => romdata <= X"00000000";
    when 16#01F1E# => romdata <= X"00000000";
    when 16#01F1F# => romdata <= X"00000000";
    when 16#01F20# => romdata <= X"00000000";
    when 16#01F21# => romdata <= X"00000000";
    when 16#01F22# => romdata <= X"00000000";
    when 16#01F23# => romdata <= X"00000000";
    when 16#01F24# => romdata <= X"00000000";
    when 16#01F25# => romdata <= X"00000000";
    when 16#01F26# => romdata <= X"00000000";
    when 16#01F27# => romdata <= X"00000000";
    when 16#01F28# => romdata <= X"00000000";
    when 16#01F29# => romdata <= X"00000000";
    when 16#01F2A# => romdata <= X"00000000";
    when 16#01F2B# => romdata <= X"00000000";
    when 16#01F2C# => romdata <= X"00000000";
    when 16#01F2D# => romdata <= X"00000000";
    when 16#01F2E# => romdata <= X"00000000";
    when 16#01F2F# => romdata <= X"00000000";
    when 16#01F30# => romdata <= X"00000000";
    when 16#01F31# => romdata <= X"00000000";
    when 16#01F32# => romdata <= X"00000000";
    when 16#01F33# => romdata <= X"00000000";
    when 16#01F34# => romdata <= X"00000000";
    when 16#01F35# => romdata <= X"00000000";
    when 16#01F36# => romdata <= X"00000000";
    when 16#01F37# => romdata <= X"00000000";
    when 16#01F38# => romdata <= X"00000000";
    when 16#01F39# => romdata <= X"00000000";
    when 16#01F3A# => romdata <= X"00000000";
    when 16#01F3B# => romdata <= X"00000000";
    when 16#01F3C# => romdata <= X"00000000";
    when 16#01F3D# => romdata <= X"00000000";
    when 16#01F3E# => romdata <= X"00000000";
    when 16#01F3F# => romdata <= X"00000000";
    when 16#01F40# => romdata <= X"00000000";
    when 16#01F41# => romdata <= X"00000000";
    when 16#01F42# => romdata <= X"00000000";
    when 16#01F43# => romdata <= X"00000000";
    when 16#01F44# => romdata <= X"00000000";
    when 16#01F45# => romdata <= X"00000000";
    when 16#01F46# => romdata <= X"00000000";
    when 16#01F47# => romdata <= X"00000000";
    when 16#01F48# => romdata <= X"00000000";
    when 16#01F49# => romdata <= X"00000000";
    when 16#01F4A# => romdata <= X"00000000";
    when 16#01F4B# => romdata <= X"00000000";
    when 16#01F4C# => romdata <= X"00000000";
    when 16#01F4D# => romdata <= X"00000000";
    when 16#01F4E# => romdata <= X"00000000";
    when 16#01F4F# => romdata <= X"00000000";
    when 16#01F50# => romdata <= X"00000000";
    when 16#01F51# => romdata <= X"00000000";
    when 16#01F52# => romdata <= X"00000000";
    when 16#01F53# => romdata <= X"00000000";
    when 16#01F54# => romdata <= X"00000000";
    when 16#01F55# => romdata <= X"00000000";
    when 16#01F56# => romdata <= X"00000000";
    when 16#01F57# => romdata <= X"00000000";
    when 16#01F58# => romdata <= X"00000000";
    when 16#01F59# => romdata <= X"00000000";
    when 16#01F5A# => romdata <= X"00000000";
    when 16#01F5B# => romdata <= X"00000000";
    when 16#01F5C# => romdata <= X"00000000";
    when 16#01F5D# => romdata <= X"00000000";
    when 16#01F5E# => romdata <= X"00000000";
    when 16#01F5F# => romdata <= X"00000000";
    when 16#01F60# => romdata <= X"00000000";
    when 16#01F61# => romdata <= X"00000000";
    when 16#01F62# => romdata <= X"00000000";
    when 16#01F63# => romdata <= X"00000000";
    when 16#01F64# => romdata <= X"00000000";
    when 16#01F65# => romdata <= X"00000000";
    when 16#01F66# => romdata <= X"00000000";
    when 16#01F67# => romdata <= X"00000000";
    when 16#01F68# => romdata <= X"00000000";
    when 16#01F69# => romdata <= X"00000000";
    when 16#01F6A# => romdata <= X"00000000";
    when 16#01F6B# => romdata <= X"00000000";
    when 16#01F6C# => romdata <= X"00000000";
    when 16#01F6D# => romdata <= X"00000000";
    when 16#01F6E# => romdata <= X"00000000";
    when 16#01F6F# => romdata <= X"00000000";
    when 16#01F70# => romdata <= X"00000000";
    when 16#01F71# => romdata <= X"00000000";
    when 16#01F72# => romdata <= X"00000000";
    when 16#01F73# => romdata <= X"00000000";
    when 16#01F74# => romdata <= X"00000000";
    when 16#01F75# => romdata <= X"00000000";
    when 16#01F76# => romdata <= X"00000000";
    when 16#01F77# => romdata <= X"00000000";
    when 16#01F78# => romdata <= X"00000000";
    when 16#01F79# => romdata <= X"00000000";
    when 16#01F7A# => romdata <= X"00000000";
    when 16#01F7B# => romdata <= X"00000000";
    when 16#01F7C# => romdata <= X"00000000";
    when 16#01F7D# => romdata <= X"00000000";
    when 16#01F7E# => romdata <= X"00000000";
    when 16#01F7F# => romdata <= X"00000000";
    when 16#01F80# => romdata <= X"00000000";
    when 16#01F81# => romdata <= X"00000000";
    when 16#01F82# => romdata <= X"00000000";
    when 16#01F83# => romdata <= X"00000000";
    when 16#01F84# => romdata <= X"00000000";
    when 16#01F85# => romdata <= X"00000000";
    when 16#01F86# => romdata <= X"00000000";
    when 16#01F87# => romdata <= X"00000000";
    when 16#01F88# => romdata <= X"00000000";
    when 16#01F89# => romdata <= X"00000000";
    when 16#01F8A# => romdata <= X"00000000";
    when 16#01F8B# => romdata <= X"00000000";
    when 16#01F8C# => romdata <= X"00000000";
    when 16#01F8D# => romdata <= X"00000000";
    when 16#01F8E# => romdata <= X"00000000";
    when 16#01F8F# => romdata <= X"00000000";
    when 16#01F90# => romdata <= X"00000000";
    when 16#01F91# => romdata <= X"00000000";
    when 16#01F92# => romdata <= X"00000000";
    when 16#01F93# => romdata <= X"00000000";
    when 16#01F94# => romdata <= X"00000000";
    when 16#01F95# => romdata <= X"00000000";
    when 16#01F96# => romdata <= X"00000000";
    when 16#01F97# => romdata <= X"00000000";
    when 16#01F98# => romdata <= X"00000000";
    when 16#01F99# => romdata <= X"00000000";
    when 16#01F9A# => romdata <= X"00000000";
    when 16#01F9B# => romdata <= X"00000000";
    when 16#01F9C# => romdata <= X"00000000";
    when 16#01F9D# => romdata <= X"00000000";
    when 16#01F9E# => romdata <= X"00000000";
    when 16#01F9F# => romdata <= X"00000000";
    when 16#01FA0# => romdata <= X"00000000";
    when 16#01FA1# => romdata <= X"00000000";
    when 16#01FA2# => romdata <= X"00000000";
    when 16#01FA3# => romdata <= X"00000000";
    when 16#01FA4# => romdata <= X"00000000";
    when 16#01FA5# => romdata <= X"00000000";
    when 16#01FA6# => romdata <= X"00000000";
    when 16#01FA7# => romdata <= X"00000000";
    when 16#01FA8# => romdata <= X"00000000";
    when 16#01FA9# => romdata <= X"00000000";
    when 16#01FAA# => romdata <= X"00000000";
    when 16#01FAB# => romdata <= X"00000000";
    when 16#01FAC# => romdata <= X"00000000";
    when 16#01FAD# => romdata <= X"00000000";
    when 16#01FAE# => romdata <= X"00000000";
    when 16#01FAF# => romdata <= X"00000000";
    when 16#01FB0# => romdata <= X"00000000";
    when 16#01FB1# => romdata <= X"00000000";
    when 16#01FB2# => romdata <= X"00000000";
    when 16#01FB3# => romdata <= X"00000000";
    when 16#01FB4# => romdata <= X"FFFFFFFF";
    when 16#01FB5# => romdata <= X"00000000";
    when 16#01FB6# => romdata <= X"00020000";
    when 16#01FB7# => romdata <= X"00000000";
    when 16#01FB8# => romdata <= X"00000000";
    when 16#01FB9# => romdata <= X"00007EDC";
    when 16#01FBA# => romdata <= X"00007EDC";
    when 16#01FBB# => romdata <= X"00007EE4";
    when 16#01FBC# => romdata <= X"00007EE4";
    when 16#01FBD# => romdata <= X"00007EEC";
    when 16#01FBE# => romdata <= X"00007EEC";
    when 16#01FBF# => romdata <= X"00007EF4";
    when 16#01FC0# => romdata <= X"00007EF4";
    when 16#01FC1# => romdata <= X"00007EFC";
    when 16#01FC2# => romdata <= X"00007EFC";
    when 16#01FC3# => romdata <= X"00007F04";
    when 16#01FC4# => romdata <= X"00007F04";
    when 16#01FC5# => romdata <= X"00007F0C";
    when 16#01FC6# => romdata <= X"00007F0C";
    when 16#01FC7# => romdata <= X"00007F14";
    when 16#01FC8# => romdata <= X"00007F14";
    when 16#01FC9# => romdata <= X"00007F1C";
    when 16#01FCA# => romdata <= X"00007F1C";
    when 16#01FCB# => romdata <= X"00007F24";
    when 16#01FCC# => romdata <= X"00007F24";
    when 16#01FCD# => romdata <= X"00007F2C";
    when 16#01FCE# => romdata <= X"00007F2C";
    when 16#01FCF# => romdata <= X"00007F34";
    when 16#01FD0# => romdata <= X"00007F34";
    when 16#01FD1# => romdata <= X"00007F3C";
    when 16#01FD2# => romdata <= X"00007F3C";
    when 16#01FD3# => romdata <= X"00007F44";
    when 16#01FD4# => romdata <= X"00007F44";
    when 16#01FD5# => romdata <= X"00007F4C";
    when 16#01FD6# => romdata <= X"00007F4C";
    when 16#01FD7# => romdata <= X"00007F54";
    when 16#01FD8# => romdata <= X"00007F54";
    when 16#01FD9# => romdata <= X"00007F5C";
    when 16#01FDA# => romdata <= X"00007F5C";
    when 16#01FDB# => romdata <= X"00007F64";
    when 16#01FDC# => romdata <= X"00007F64";
    when 16#01FDD# => romdata <= X"00007F6C";
    when 16#01FDE# => romdata <= X"00007F6C";
    when 16#01FDF# => romdata <= X"00007F74";
    when 16#01FE0# => romdata <= X"00007F74";
    when 16#01FE1# => romdata <= X"00007F7C";
    when 16#01FE2# => romdata <= X"00007F7C";
    when 16#01FE3# => romdata <= X"00007F84";
    when 16#01FE4# => romdata <= X"00007F84";
    when 16#01FE5# => romdata <= X"00007F8C";
    when 16#01FE6# => romdata <= X"00007F8C";
    when 16#01FE7# => romdata <= X"00007F94";
    when 16#01FE8# => romdata <= X"00007F94";
    when 16#01FE9# => romdata <= X"00007F9C";
    when 16#01FEA# => romdata <= X"00007F9C";
    when 16#01FEB# => romdata <= X"00007FA4";
    when 16#01FEC# => romdata <= X"00007FA4";
    when 16#01FED# => romdata <= X"00007FAC";
    when 16#01FEE# => romdata <= X"00007FAC";
    when 16#01FEF# => romdata <= X"00007FB4";
    when 16#01FF0# => romdata <= X"00007FB4";
    when 16#01FF1# => romdata <= X"00007FBC";
    when 16#01FF2# => romdata <= X"00007FBC";
    when 16#01FF3# => romdata <= X"00007FC4";
    when 16#01FF4# => romdata <= X"00007FC4";
    when 16#01FF5# => romdata <= X"00007FCC";
    when 16#01FF6# => romdata <= X"00007FCC";
    when 16#01FF7# => romdata <= X"00007FD4";
    when 16#01FF8# => romdata <= X"00007FD4";
    when 16#01FF9# => romdata <= X"00007FDC";
    when 16#01FFA# => romdata <= X"00007FDC";
    when 16#01FFB# => romdata <= X"00007FE4";
    when 16#01FFC# => romdata <= X"00007FE4";
    when 16#01FFD# => romdata <= X"00007FEC";
    when 16#01FFE# => romdata <= X"00007FEC";
    when 16#01FFF# => romdata <= X"00007FF4";
    when 16#02000# => romdata <= X"00007FF4";
    when 16#02001# => romdata <= X"00007FFC";
    when 16#02002# => romdata <= X"00007FFC";
    when 16#02003# => romdata <= X"00008004";
    when 16#02004# => romdata <= X"00008004";
    when 16#02005# => romdata <= X"0000800C";
    when 16#02006# => romdata <= X"0000800C";
    when 16#02007# => romdata <= X"00008014";
    when 16#02008# => romdata <= X"00008014";
    when 16#02009# => romdata <= X"0000801C";
    when 16#0200A# => romdata <= X"0000801C";
    when 16#0200B# => romdata <= X"00008024";
    when 16#0200C# => romdata <= X"00008024";
    when 16#0200D# => romdata <= X"0000802C";
    when 16#0200E# => romdata <= X"0000802C";
    when 16#0200F# => romdata <= X"00008034";
    when 16#02010# => romdata <= X"00008034";
    when 16#02011# => romdata <= X"0000803C";
    when 16#02012# => romdata <= X"0000803C";
    when 16#02013# => romdata <= X"00008044";
    when 16#02014# => romdata <= X"00008044";
    when 16#02015# => romdata <= X"0000804C";
    when 16#02016# => romdata <= X"0000804C";
    when 16#02017# => romdata <= X"00008054";
    when 16#02018# => romdata <= X"00008054";
    when 16#02019# => romdata <= X"0000805C";
    when 16#0201A# => romdata <= X"0000805C";
    when 16#0201B# => romdata <= X"00008064";
    when 16#0201C# => romdata <= X"00008064";
    when 16#0201D# => romdata <= X"0000806C";
    when 16#0201E# => romdata <= X"0000806C";
    when 16#0201F# => romdata <= X"00008074";
    when 16#02020# => romdata <= X"00008074";
    when 16#02021# => romdata <= X"0000807C";
    when 16#02022# => romdata <= X"0000807C";
    when 16#02023# => romdata <= X"00008084";
    when 16#02024# => romdata <= X"00008084";
    when 16#02025# => romdata <= X"0000808C";
    when 16#02026# => romdata <= X"0000808C";
    when 16#02027# => romdata <= X"00008094";
    when 16#02028# => romdata <= X"00008094";
    when 16#02029# => romdata <= X"0000809C";
    when 16#0202A# => romdata <= X"0000809C";
    when 16#0202B# => romdata <= X"000080A4";
    when 16#0202C# => romdata <= X"000080A4";
    when 16#0202D# => romdata <= X"000080AC";
    when 16#0202E# => romdata <= X"000080AC";
    when 16#0202F# => romdata <= X"000080B4";
    when 16#02030# => romdata <= X"000080B4";
    when 16#02031# => romdata <= X"000080BC";
    when 16#02032# => romdata <= X"000080BC";
    when 16#02033# => romdata <= X"000080C4";
    when 16#02034# => romdata <= X"000080C4";
    when 16#02035# => romdata <= X"000080CC";
    when 16#02036# => romdata <= X"000080CC";
    when 16#02037# => romdata <= X"000080D4";
    when 16#02038# => romdata <= X"000080D4";
    when 16#02039# => romdata <= X"000080DC";
    when 16#0203A# => romdata <= X"000080DC";
    when 16#0203B# => romdata <= X"000080E4";
    when 16#0203C# => romdata <= X"000080E4";
    when 16#0203D# => romdata <= X"000080EC";
    when 16#0203E# => romdata <= X"000080EC";
    when 16#0203F# => romdata <= X"000080F4";
    when 16#02040# => romdata <= X"000080F4";
    when 16#02041# => romdata <= X"000080FC";
    when 16#02042# => romdata <= X"000080FC";
    when 16#02043# => romdata <= X"00008104";
    when 16#02044# => romdata <= X"00008104";
    when 16#02045# => romdata <= X"0000810C";
    when 16#02046# => romdata <= X"0000810C";
    when 16#02047# => romdata <= X"00008114";
    when 16#02048# => romdata <= X"00008114";
    when 16#02049# => romdata <= X"0000811C";
    when 16#0204A# => romdata <= X"0000811C";
    when 16#0204B# => romdata <= X"00008124";
    when 16#0204C# => romdata <= X"00008124";
    when 16#0204D# => romdata <= X"0000812C";
    when 16#0204E# => romdata <= X"0000812C";
    when 16#0204F# => romdata <= X"00008134";
    when 16#02050# => romdata <= X"00008134";
    when 16#02051# => romdata <= X"0000813C";
    when 16#02052# => romdata <= X"0000813C";
    when 16#02053# => romdata <= X"00008144";
    when 16#02054# => romdata <= X"00008144";
    when 16#02055# => romdata <= X"0000814C";
    when 16#02056# => romdata <= X"0000814C";
    when 16#02057# => romdata <= X"00008154";
    when 16#02058# => romdata <= X"00008154";
    when 16#02059# => romdata <= X"0000815C";
    when 16#0205A# => romdata <= X"0000815C";
    when 16#0205B# => romdata <= X"00008164";
    when 16#0205C# => romdata <= X"00008164";
    when 16#0205D# => romdata <= X"0000816C";
    when 16#0205E# => romdata <= X"0000816C";
    when 16#0205F# => romdata <= X"00008174";
    when 16#02060# => romdata <= X"00008174";
    when 16#02061# => romdata <= X"0000817C";
    when 16#02062# => romdata <= X"0000817C";
    when 16#02063# => romdata <= X"00008184";
    when 16#02064# => romdata <= X"00008184";
    when 16#02065# => romdata <= X"0000818C";
    when 16#02066# => romdata <= X"0000818C";
    when 16#02067# => romdata <= X"00008194";
    when 16#02068# => romdata <= X"00008194";
    when 16#02069# => romdata <= X"0000819C";
    when 16#0206A# => romdata <= X"0000819C";
    when 16#0206B# => romdata <= X"000081A4";
    when 16#0206C# => romdata <= X"000081A4";
    when 16#0206D# => romdata <= X"000081AC";
    when 16#0206E# => romdata <= X"000081AC";
    when 16#0206F# => romdata <= X"000081B4";
    when 16#02070# => romdata <= X"000081B4";
    when 16#02071# => romdata <= X"000081BC";
    when 16#02072# => romdata <= X"000081BC";
    when 16#02073# => romdata <= X"000081C4";
    when 16#02074# => romdata <= X"000081C4";
    when 16#02075# => romdata <= X"000081CC";
    when 16#02076# => romdata <= X"000081CC";
    when 16#02077# => romdata <= X"000081D4";
    when 16#02078# => romdata <= X"000081D4";
    when 16#02079# => romdata <= X"000081DC";
    when 16#0207A# => romdata <= X"000081DC";
    when 16#0207B# => romdata <= X"000081E4";
    when 16#0207C# => romdata <= X"000081E4";
    when 16#0207D# => romdata <= X"000081EC";
    when 16#0207E# => romdata <= X"000081EC";
    when 16#0207F# => romdata <= X"000081F4";
    when 16#02080# => romdata <= X"000081F4";
    when 16#02081# => romdata <= X"000081FC";
    when 16#02082# => romdata <= X"000081FC";
    when 16#02083# => romdata <= X"00008204";
    when 16#02084# => romdata <= X"00008204";
    when 16#02085# => romdata <= X"0000820C";
    when 16#02086# => romdata <= X"0000820C";
    when 16#02087# => romdata <= X"00008214";
    when 16#02088# => romdata <= X"00008214";
    when 16#02089# => romdata <= X"0000821C";
    when 16#0208A# => romdata <= X"0000821C";
    when 16#0208B# => romdata <= X"00008224";
    when 16#0208C# => romdata <= X"00008224";
    when 16#0208D# => romdata <= X"0000822C";
    when 16#0208E# => romdata <= X"0000822C";
    when 16#0208F# => romdata <= X"00008234";
    when 16#02090# => romdata <= X"00008234";
    when 16#02091# => romdata <= X"0000823C";
    when 16#02092# => romdata <= X"0000823C";
    when 16#02093# => romdata <= X"00008244";
    when 16#02094# => romdata <= X"00008244";
    when 16#02095# => romdata <= X"0000824C";
    when 16#02096# => romdata <= X"0000824C";
    when 16#02097# => romdata <= X"00008254";
    when 16#02098# => romdata <= X"00008254";
    when 16#02099# => romdata <= X"0000825C";
    when 16#0209A# => romdata <= X"0000825C";
    when 16#0209B# => romdata <= X"00008264";
    when 16#0209C# => romdata <= X"00008264";
    when 16#0209D# => romdata <= X"0000826C";
    when 16#0209E# => romdata <= X"0000826C";
    when 16#0209F# => romdata <= X"00008274";
    when 16#020A0# => romdata <= X"00008274";
    when 16#020A1# => romdata <= X"0000827C";
    when 16#020A2# => romdata <= X"0000827C";
    when 16#020A3# => romdata <= X"00008284";
    when 16#020A4# => romdata <= X"00008284";
    when 16#020A5# => romdata <= X"0000828C";
    when 16#020A6# => romdata <= X"0000828C";
    when 16#020A7# => romdata <= X"00008294";
    when 16#020A8# => romdata <= X"00008294";
    when 16#020A9# => romdata <= X"0000829C";
    when 16#020AA# => romdata <= X"0000829C";
    when 16#020AB# => romdata <= X"000082A4";
    when 16#020AC# => romdata <= X"000082A4";
    when 16#020AD# => romdata <= X"000082AC";
    when 16#020AE# => romdata <= X"000082AC";
    when 16#020AF# => romdata <= X"000082B4";
    when 16#020B0# => romdata <= X"000082B4";
    when 16#020B1# => romdata <= X"000082BC";
    when 16#020B2# => romdata <= X"000082BC";
    when 16#020B3# => romdata <= X"000082C4";
    when 16#020B4# => romdata <= X"000082C4";
    when 16#020B5# => romdata <= X"000082CC";
    when 16#020B6# => romdata <= X"000082CC";
    when 16#020B7# => romdata <= X"000082D4";
    when 16#020B8# => romdata <= X"000082D4";
    when 16#020B9# => romdata <= X"000082D4";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
