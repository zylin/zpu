library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;


library zylin;
use zylin.zpu_config.all;
use zylin.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBit downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(0 to ((2**(maxAddrBit+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
0 => x"800b0b0b",
1 => x"0b0b8070",
2 => x"0b0b80e5",
3 => x"d00c3a0b",
4 => x"0b0bbed7",
5 => x"04000000",
6 => x"00000000",
7 => x"00000000",
8 => x"80088408",
9 => x"88080b0b",
10 => x"0bbfa72d",
11 => x"880c840c",
12 => x"800c0400",
13 => x"00000000",
14 => x"00000000",
15 => x"00000000",
16 => x"71fd0608",
17 => x"72830609",
18 => x"81058205",
19 => x"832b2a83",
20 => x"ffff0652",
21 => x"0b0b0400",
22 => x"00000000",
23 => x"00000000",
24 => x"71fd0608",
25 => x"83ffff73",
26 => x"83060981",
27 => x"05820583",
28 => x"2b2b0906",
29 => x"7383ffff",
30 => x"0b0b0b0b",
31 => x"83a70400",
32 => x"72098105",
33 => x"72057373",
34 => x"09060906",
35 => x"73097306",
36 => x"070a8106",
37 => x"530b0b51",
38 => x"04000000",
39 => x"00000000",
40 => x"72722473",
41 => x"732e0753",
42 => x"0b0b5104",
43 => x"00000000",
44 => x"00000000",
45 => x"00000000",
46 => x"00000000",
47 => x"00000000",
48 => x"71737109",
49 => x"71068106",
50 => x"30720a10",
51 => x"0a720a10",
52 => x"0a31050a",
53 => x"81065151",
54 => x"530b0b51",
55 => x"04000000",
56 => x"72722673",
57 => x"732e0753",
58 => x"0b0b5104",
59 => x"00000000",
60 => x"00000000",
61 => x"00000000",
62 => x"00000000",
63 => x"00000000",
64 => x"00000000",
65 => x"00000000",
66 => x"00000000",
67 => x"00000000",
68 => x"00000000",
69 => x"00000000",
70 => x"00000000",
71 => x"00000000",
72 => x"0b0b0b88",
73 => x"c6040000",
74 => x"00000000",
75 => x"00000000",
76 => x"00000000",
77 => x"00000000",
78 => x"00000000",
79 => x"00000000",
80 => x"720a722b",
81 => x"0a530b0b",
82 => x"51040000",
83 => x"00000000",
84 => x"00000000",
85 => x"00000000",
86 => x"00000000",
87 => x"00000000",
88 => x"72729f06",
89 => x"0981050b",
90 => x"0b0b88a7",
91 => x"05040000",
92 => x"00000000",
93 => x"00000000",
94 => x"00000000",
95 => x"00000000",
96 => x"72722aff",
97 => x"739f062a",
98 => x"0974090a",
99 => x"8106ff05",
100 => x"0607530b",
101 => x"0b510400",
102 => x"00000000",
103 => x"00000000",
104 => x"7171530b",
105 => x"0b510406",
106 => x"73830609",
107 => x"81058205",
108 => x"832b0b2b",
109 => x"0772fc06",
110 => x"0c515104",
111 => x"00000000",
112 => x"72098105",
113 => x"72050970",
114 => x"81050906",
115 => x"0a810653",
116 => x"0b0b5104",
117 => x"00000000",
118 => x"00000000",
119 => x"00000000",
120 => x"72098105",
121 => x"72050970",
122 => x"81050906",
123 => x"0a098106",
124 => x"530b0b51",
125 => x"04000000",
126 => x"00000000",
127 => x"00000000",
128 => x"71098105",
129 => x"520b0b04",
130 => x"00000000",
131 => x"00000000",
132 => x"00000000",
133 => x"00000000",
134 => x"00000000",
135 => x"00000000",
136 => x"72720981",
137 => x"0505530b",
138 => x"0b510400",
139 => x"00000000",
140 => x"00000000",
141 => x"00000000",
142 => x"00000000",
143 => x"00000000",
144 => x"72097206",
145 => x"73730906",
146 => x"07530b0b",
147 => x"51040000",
148 => x"00000000",
149 => x"00000000",
150 => x"00000000",
151 => x"00000000",
152 => x"71fc0608",
153 => x"72830609",
154 => x"81058305",
155 => x"1010102a",
156 => x"81ff0652",
157 => x"0b0b0400",
158 => x"00000000",
159 => x"00000000",
160 => x"71fc0608",
161 => x"0b0b80e5",
162 => x"bc738306",
163 => x"10100508",
164 => x"060b0b0b",
165 => x"88ac0400",
166 => x"00000000",
167 => x"00000000",
168 => x"80088408",
169 => x"88087575",
170 => x"0b0b0ba3",
171 => x"fa2d5050",
172 => x"80085688",
173 => x"0c840c80",
174 => x"0c510400",
175 => x"00000000",
176 => x"80088408",
177 => x"88087575",
178 => x"0b0b0ba4",
179 => x"ca2d5050",
180 => x"80085688",
181 => x"0c840c80",
182 => x"0c510400",
183 => x"00000000",
184 => x"72097081",
185 => x"0509060a",
186 => x"8106ff05",
187 => x"70540b0b",
188 => x"71067309",
189 => x"727405ff",
190 => x"05060751",
191 => x"51510400",
192 => x"72097081",
193 => x"0509060a",
194 => x"098106ff",
195 => x"0570540b",
196 => x"0b710673",
197 => x"09727405",
198 => x"ff050607",
199 => x"51515104",
200 => x"05ff0504",
201 => x"00000000",
202 => x"00000000",
203 => x"00000000",
204 => x"00000000",
205 => x"00000000",
206 => x"00000000",
207 => x"00000000",
208 => x"810b0b0b",
209 => x"80e5cc0c",
210 => x"51040000",
211 => x"00000000",
212 => x"00000000",
213 => x"00000000",
214 => x"00000000",
215 => x"00000000",
216 => x"71810552",
217 => x"0b0b0400",
218 => x"00000000",
219 => x"00000000",
220 => x"00000000",
221 => x"00000000",
222 => x"00000000",
223 => x"00000000",
224 => x"00000000",
225 => x"00000000",
226 => x"00000000",
227 => x"00000000",
228 => x"00000000",
229 => x"00000000",
230 => x"00000000",
231 => x"00000000",
232 => x"02840572",
233 => x"10100552",
234 => x"0b0b0400",
235 => x"00000000",
236 => x"00000000",
237 => x"00000000",
238 => x"00000000",
239 => x"00000000",
240 => x"00000000",
241 => x"00000000",
242 => x"00000000",
243 => x"00000000",
244 => x"00000000",
245 => x"00000000",
246 => x"00000000",
247 => x"00000000",
248 => x"717105ff",
249 => x"0571530b",
250 => x"0b510400",
251 => x"00000000",
252 => x"00000000",
253 => x"00000000",
254 => x"00000000",
255 => x"00000000",
256 => x"84803f80",
257 => x"cef23f04",
258 => x"10101010",
259 => x"10101010",
260 => x"10101010",
261 => x"10101010",
262 => x"10101010",
263 => x"10101010",
264 => x"10101010",
265 => x"10101053",
266 => x"0b0b5104",
267 => x"7381ff06",
268 => x"73830609",
269 => x"81058305",
270 => x"1010102b",
271 => x"0772fc06",
272 => x"0c515104",
273 => x"3c047272",
274 => x"80728106",
275 => x"ff050972",
276 => x"06057110",
277 => x"520b0b72",
278 => x"0a100a53",
279 => x"0b0b72e9",
280 => x"38515153",
281 => x"0b0b5104",
282 => x"70700b0b",
283 => x"80f5c008",
284 => x"520b0b84",
285 => x"0b720508",
286 => x"70810651",
287 => x"510b0b70",
288 => x"f2387108",
289 => x"81ff0680",
290 => x"0c505004",
291 => x"70700b0b",
292 => x"80f5c008",
293 => x"520b0b84",
294 => x"0b720508",
295 => x"700a100a",
296 => x"70810651",
297 => x"51510b0b",
298 => x"70ed3873",
299 => x"720c5050",
300 => x"0480e5cc",
301 => x"08802ea8",
302 => x"38838080",
303 => x"0b0b0b80",
304 => x"f5c00c82",
305 => x"a0800b0b",
306 => x"0b80f5c4",
307 => x"0c829080",
308 => x"0b80f5d4",
309 => x"0c0b0b80",
310 => x"f5c80b80",
311 => x"f5d80c04",
312 => x"f8808080",
313 => x"a40b0b0b",
314 => x"80f5c00c",
315 => x"f8808082",
316 => x"800b0b0b",
317 => x"80f5c40c",
318 => x"f8808084",
319 => x"800b80f5",
320 => x"d40cf880",
321 => x"8080940b",
322 => x"80f5d80c",
323 => x"f8808080",
324 => x"9c0b80f5",
325 => x"d00cf880",
326 => x"8080a00b",
327 => x"80f5dc0c",
328 => x"04f23d0d",
329 => x"600b0b80",
330 => x"f5c40856",
331 => x"5d82750c",
332 => x"8059805a",
333 => x"800b8f3d",
334 => x"71101017",
335 => x"70085957",
336 => x"5d5b8076",
337 => x"81ff067c",
338 => x"832b5658",
339 => x"520b0b0b",
340 => x"76530b0b",
341 => x"7b5198c6",
342 => x"3f7d7f7a",
343 => x"72077c72",
344 => x"07717160",
345 => x"8105415f",
346 => x"5d5b5957",
347 => x"557a8724",
348 => x"80c1380b",
349 => x"0b80f5c4",
350 => x"087b1010",
351 => x"71057008",
352 => x"58515580",
353 => x"7681ff06",
354 => x"7c832b56",
355 => x"58520b0b",
356 => x"0b76530b",
357 => x"0b7b5198",
358 => x"853f7d7f",
359 => x"7a72077c",
360 => x"72077171",
361 => x"60810541",
362 => x"5f5d5b59",
363 => x"5755877b",
364 => x"25c13876",
365 => x"7d0c7784",
366 => x"1e0c7c80",
367 => x"0c903d0d",
368 => x"04707080",
369 => x"f5cc3351",
370 => x"0b0b70b2",
371 => x"3880e5d8",
372 => x"08700852",
373 => x"0b0b520b",
374 => x"0b0b7080",
375 => x"2e9a3884",
376 => x"720580e5",
377 => x"d80c702d",
378 => x"80e5d808",
379 => x"7008520b",
380 => x"0b520b0b",
381 => x"0b70e838",
382 => x"810b80f5",
383 => x"cc345050",
384 => x"0404700b",
385 => x"0b80f5bc",
386 => x"08802e8e",
387 => x"380b0b0b",
388 => x"0b800b80",
389 => x"2e098106",
390 => x"83385004",
391 => x"0b0b80f5",
392 => x"bc510b0b",
393 => x"0bf3d93f",
394 => x"50040470",
395 => x"70028f05",
396 => x"33520b0b",
397 => x"0b0b718a",
398 => x"2e893871",
399 => x"51fccd3f",
400 => x"5050048d",
401 => x"51fcc53f",
402 => x"7151fcc0",
403 => x"3f505004",
404 => x"cd3d0db6",
405 => x"3d707084",
406 => x"05520b0b",
407 => x"088cab5d",
408 => x"56a63d5f",
409 => x"5d807570",
410 => x"81055733",
411 => x"765c5559",
412 => x"0b730b79",
413 => x"2e80ca38",
414 => x"8f3d5c73",
415 => x"a52e0981",
416 => x"0680cf38",
417 => x"79708105",
418 => x"5b33540b",
419 => x"0b7380e4",
420 => x"2e81c838",
421 => x"7380e424",
422 => x"80d13873",
423 => x"80e32ea8",
424 => x"3880520b",
425 => x"0ba5517a",
426 => x"2d80520b",
427 => x"0b73517a",
428 => x"2d821959",
429 => x"79708105",
430 => x"5b33540b",
431 => x"0b73ffbb",
432 => x"3878800c",
433 => x"b53d0d04",
434 => x"7c841e83",
435 => x"72053356",
436 => x"5e578052",
437 => x"0b0b7351",
438 => x"7a2d8119",
439 => x"7a708105",
440 => x"5c335559",
441 => x"0b73ff93",
442 => x"38d73973",
443 => x"80f32e09",
444 => x"8106ffad",
445 => x"387c841e",
446 => x"7108595e",
447 => x"56807733",
448 => x"56560b74",
449 => x"0b762e8d",
450 => x"38811670",
451 => x"1870335a",
452 => x"555677f5",
453 => x"38ff1655",
454 => x"807625ff",
455 => x"97387670",
456 => x"81055833",
457 => x"5880520b",
458 => x"0b77517a",
459 => x"2d811975",
460 => x"ff175757",
461 => x"59807625",
462 => x"fefa3876",
463 => x"70810558",
464 => x"33588052",
465 => x"0b0b7751",
466 => x"7a2d8119",
467 => x"75ff1757",
468 => x"57590b75",
469 => x"8024c738",
470 => x"feda397c",
471 => x"841e7108",
472 => x"70719f2c",
473 => x"59530b0b",
474 => x"595e5680",
475 => x"7524818d",
476 => x"38757e7d",
477 => x"58595580",
478 => x"57740b77",
479 => x"2e098106",
480 => x"bc38b07c",
481 => x"3402b905",
482 => x"567b0b76",
483 => x"2e9938ff",
484 => x"16560b0b",
485 => x"75337870",
486 => x"81055a34",
487 => x"8117577b",
488 => x"762e0981",
489 => x"06e93880",
490 => x"7834767e",
491 => x"ff720557",
492 => x"58560b0b",
493 => x"758024fe",
494 => x"e538fdf8",
495 => x"398a7536",
496 => x"0b0b80d7",
497 => x"b005540b",
498 => x"0b733376",
499 => x"70810558",
500 => x"348a7535",
501 => x"550b0b74",
502 => x"802effad",
503 => x"388a7536",
504 => x"0b0b80d7",
505 => x"b005540b",
506 => x"0b733376",
507 => x"70810558",
508 => x"348a7535",
509 => x"550b0b74",
510 => x"c438ff8d",
511 => x"3974520b",
512 => x"0b76530b",
513 => x"0bb53dff",
514 => x"b8055192",
515 => x"dc3fa43d",
516 => x"0856fedd",
517 => x"397080c1",
518 => x"0b81c48c",
519 => x"34800b81",
520 => x"c5e40c70",
521 => x"800c5004",
522 => x"7070800b",
523 => x"81c48c33",
524 => x"520b0b52",
525 => x"0b0b0b70",
526 => x"80c12e98",
527 => x"387181c5",
528 => x"e4080781",
529 => x"c5e40c80",
530 => x"c20b81c4",
531 => x"90347080",
532 => x"0c505004",
533 => x"810b81c5",
534 => x"e4080781",
535 => x"c5e40c80",
536 => x"c20b81c4",
537 => x"90347080",
538 => x"0c505004",
539 => x"70707070",
540 => x"7570088a",
541 => x"05530b0b",
542 => x"530b0b81",
543 => x"c48c3351",
544 => x"0b0b7080",
545 => x"c12e8c38",
546 => x"73f13870",
547 => x"800c5050",
548 => x"505004ff",
549 => x"72057081",
550 => x"c4880831",
551 => x"740c800c",
552 => x"50505050",
553 => x"04fc3d0d",
554 => x"81c49408",
555 => x"550b0b74",
556 => x"802e8e38",
557 => x"76750871",
558 => x"0c81c494",
559 => x"0856540b",
560 => x"0b8c1553",
561 => x"0b0b81c4",
562 => x"8808520b",
563 => x"0b8a518e",
564 => x"e93f7380",
565 => x"0c863d0d",
566 => x"04fb3d0d",
567 => x"77700856",
568 => x"56b0530b",
569 => x"0b81c494",
570 => x"08520b0b",
571 => x"7451a1ff",
572 => x"3f850b8c",
573 => x"170c850b",
574 => x"8c160c75",
575 => x"08750c81",
576 => x"c4940854",
577 => x"0b0b7380",
578 => x"2e8c3873",
579 => x"08750c81",
580 => x"c4940854",
581 => x"0b0b8c14",
582 => x"530b0b81",
583 => x"c4880852",
584 => x"0b0b8a51",
585 => x"8e943f84",
586 => x"1508b738",
587 => x"860b8c16",
588 => x"0c881552",
589 => x"0b0b8816",
590 => x"08518d96",
591 => x"3f81c494",
592 => x"08700876",
593 => x"0c540b0b",
594 => x"8c157054",
595 => x"0b0b540b",
596 => x"0b8a520b",
597 => x"0b730851",
598 => x"8de03f73",
599 => x"800c873d",
600 => x"0d047508",
601 => x"540b0bb0",
602 => x"530b0b73",
603 => x"520b0b75",
604 => x"51a0fc3f",
605 => x"73800c87",
606 => x"3d0d04e1",
607 => x"3d0db051",
608 => x"93833f80",
609 => x"0881c484",
610 => x"0cb05192",
611 => x"f83f8008",
612 => x"81c4940c",
613 => x"81c48408",
614 => x"80080c80",
615 => x"0b800884",
616 => x"050c820b",
617 => x"80088805",
618 => x"0ca80b80",
619 => x"088c050c",
620 => x"9f530b0b",
621 => x"0b0b80d7",
622 => x"bc520b0b",
623 => x"80089005",
624 => x"51a0ac3f",
625 => x"993d5c9f",
626 => x"530b0b0b",
627 => x"0b80d7dc",
628 => x"520b0b7b",
629 => x"51a0983f",
630 => x"8a0b8182",
631 => x"cc0c0b0b",
632 => x"80e28051",
633 => x"f8ea3f0b",
634 => x"0b80d7fc",
635 => x"51f8e13f",
636 => x"0b0b80e2",
637 => x"8051f8d8",
638 => x"3f80e5e0",
639 => x"08802e8a",
640 => x"a1380b0b",
641 => x"80d8ac51",
642 => x"f8c63f0b",
643 => x"0b80e280",
644 => x"51f8bd3f",
645 => x"80e5dc08",
646 => x"520b0b0b",
647 => x"0b80d8d8",
648 => x"51f8ad3f",
649 => x"8051b488",
650 => x"3f800880",
651 => x"f5ec0c81",
652 => x"0b923d5c",
653 => x"58800b80",
654 => x"e5dc0825",
655 => x"8383388e",
656 => x"3d5d80c1",
657 => x"0b81c48c",
658 => x"34810b81",
659 => x"c5e40c80",
660 => x"c20b81c4",
661 => x"9034825e",
662 => x"835a9f53",
663 => x"0b0b0b0b",
664 => x"80d98852",
665 => x"0b0b7a51",
666 => x"9f853f81",
667 => x"5f807b53",
668 => x"0b0b7c52",
669 => x"0b0b558c",
670 => x"f43f8008",
671 => x"752e0981",
672 => x"06833881",
673 => x"550b0b74",
674 => x"81c5e40c",
675 => x"7d705755",
676 => x"0b0b7483",
677 => x"25a63874",
678 => x"101015fd",
679 => x"0540a13d",
680 => x"ffbc0553",
681 => x"0b0b8352",
682 => x"0b0b7551",
683 => x"8b8c3f81",
684 => x"1e705f70",
685 => x"5755830b",
686 => x"7524dc38",
687 => x"7f540b0b",
688 => x"74530b0b",
689 => x"80f5f052",
690 => x"0b0b81c4",
691 => x"9c518af6",
692 => x"3f81c494",
693 => x"08700857",
694 => x"57b0530b",
695 => x"0b76520b",
696 => x"0b75519e",
697 => x"8a3f850b",
698 => x"8c180c85",
699 => x"0b8c170c",
700 => x"7608760c",
701 => x"81c49408",
702 => x"550b0b74",
703 => x"802e8a38",
704 => x"7408760c",
705 => x"81c49408",
706 => x"558c1553",
707 => x"0b0b81c4",
708 => x"8808520b",
709 => x"0b8a518a",
710 => x"a13f8416",
711 => x"08888c38",
712 => x"860b8c17",
713 => x"0c881652",
714 => x"0b0b8817",
715 => x"085189a2",
716 => x"3f81c494",
717 => x"08700877",
718 => x"0c578c16",
719 => x"70540b0b",
720 => x"558a520b",
721 => x"0b740851",
722 => x"89f03f80",
723 => x"c10b81c4",
724 => x"90335656",
725 => x"0b0b7575",
726 => x"26a83880",
727 => x"c3520b0b",
728 => x"75518adb",
729 => x"3f80087f",
730 => x"2e87ff38",
731 => x"81167081",
732 => x"ff0681c4",
733 => x"9033520b",
734 => x"0b57550b",
735 => x"0b747627",
736 => x"da38797e",
737 => x"29607072",
738 => x"35704172",
739 => x"72317087",
740 => x"2972315e",
741 => x"530b0b8a",
742 => x"0581c48c",
743 => x"3381c488",
744 => x"085a520b",
745 => x"0b520b0b",
746 => x"58550b76",
747 => x"80c12e87",
748 => x"f03878f6",
749 => x"38811858",
750 => x"80e5dc08",
751 => x"7825fd82",
752 => x"388051b0",
753 => x"eb3f8008",
754 => x"81c4800c",
755 => x"0b0b80d9",
756 => x"a851f4fc",
757 => x"3f0b0b80",
758 => x"e28051f4",
759 => x"f33f0b0b",
760 => x"80d9b851",
761 => x"f4ea3f0b",
762 => x"0b80e280",
763 => x"51f4e13f",
764 => x"81c48808",
765 => x"520b0b0b",
766 => x"0b80d9f0",
767 => x"51f4d13f",
768 => x"85520b0b",
769 => x"0b0b80da",
770 => x"8c51f4c4",
771 => x"3f81c5e4",
772 => x"08520b0b",
773 => x"0b0b80da",
774 => x"a851f4b4",
775 => x"3f81520b",
776 => x"0b0b0b80",
777 => x"da8c51f4",
778 => x"a73f81c4",
779 => x"8c33520b",
780 => x"0b0b0b80",
781 => x"dac451f4",
782 => x"973f80c1",
783 => x"520b0b0b",
784 => x"0b80dae0",
785 => x"51f4893f",
786 => x"81c49033",
787 => x"520b0b0b",
788 => x"0b80dafc",
789 => x"51f3f93f",
790 => x"80c2520b",
791 => x"0b0b0b80",
792 => x"dae051f3",
793 => x"eb3f81c4",
794 => x"bc08520b",
795 => x"0b0b0b80",
796 => x"db9851f3",
797 => x"db3f8752",
798 => x"0b0b0b0b",
799 => x"80da8c51",
800 => x"f3ce3f81",
801 => x"82cc0852",
802 => x"0b0b0b0b",
803 => x"80dbb451",
804 => x"f3be3f0b",
805 => x"0b80dbd0",
806 => x"51f3b53f",
807 => x"0b0b80db",
808 => x"fc51f3ac",
809 => x"3f81c494",
810 => x"08700853",
811 => x"0b0b560b",
812 => x"0b80dc88",
813 => x"51f3993f",
814 => x"0b0b80dc",
815 => x"a451f390",
816 => x"3f81c494",
817 => x"08847105",
818 => x"08530b0b",
819 => x"5d0b0b80",
820 => x"dcd851f2",
821 => x"fb3f8052",
822 => x"0b0b0b0b",
823 => x"80da8c51",
824 => x"f2ee3f81",
825 => x"c4940888",
826 => x"71050853",
827 => x"0b0b580b",
828 => x"0b80dcf4",
829 => x"51f2d93f",
830 => x"82520b0b",
831 => x"0b0b80da",
832 => x"8c51f2cc",
833 => x"3f81c494",
834 => x"088c7105",
835 => x"08530b0b",
836 => x"590b0b80",
837 => x"dd9051f2",
838 => x"b73f9152",
839 => x"0b0b0b0b",
840 => x"80da8c51",
841 => x"f2aa3f81",
842 => x"c4940890",
843 => x"05520b0b",
844 => x"0b0b80dd",
845 => x"ac51f298",
846 => x"3f0b0b80",
847 => x"ddc851f2",
848 => x"8f3f0b0b",
849 => x"80de8051",
850 => x"f2863f81",
851 => x"c4840870",
852 => x"08530b0b",
853 => x"570b0b80",
854 => x"dc8851f1",
855 => x"f33f0b0b",
856 => x"80de9451",
857 => x"f1ea3f81",
858 => x"c4840884",
859 => x"71050853",
860 => x"0b0b550b",
861 => x"0b80dcd8",
862 => x"51f1d53f",
863 => x"80520b0b",
864 => x"0b0b80da",
865 => x"8c51f1c8",
866 => x"3f81c484",
867 => x"08887105",
868 => x"08530b0b",
869 => x"560b0b80",
870 => x"dcf451f1",
871 => x"b33f8152",
872 => x"0b0b0b0b",
873 => x"80da8c51",
874 => x"f1a63f81",
875 => x"c484088c",
876 => x"71050853",
877 => x"0b0b5d0b",
878 => x"0b80dd90",
879 => x"51f1913f",
880 => x"92520b0b",
881 => x"0b0b80da",
882 => x"8c51f184",
883 => x"3f81c484",
884 => x"08900552",
885 => x"0b0b0b0b",
886 => x"80ddac51",
887 => x"f0f23f0b",
888 => x"0b80ddc8",
889 => x"51f0e93f",
890 => x"7d520b0b",
891 => x"0b0b80de",
892 => x"d451f0dc",
893 => x"3f85520b",
894 => x"0b0b0b80",
895 => x"da8c51f0",
896 => x"cf3f7952",
897 => x"0b0b0b0b",
898 => x"80def051",
899 => x"f0c23f8d",
900 => x"520b0b0b",
901 => x"0b80da8c",
902 => x"51f0b53f",
903 => x"7f520b0b",
904 => x"0b0b80df",
905 => x"8c51f0a8",
906 => x"3f87520b",
907 => x"0b0b0b80",
908 => x"da8c51f0",
909 => x"9b3f7e52",
910 => x"0b0b0b0b",
911 => x"80dfa851",
912 => x"f08e3f81",
913 => x"520b0b0b",
914 => x"0b80da8c",
915 => x"51f0813f",
916 => x"7b520b0b",
917 => x"0b0b80df",
918 => x"c451eff4",
919 => x"3f0b0b80",
920 => x"dfe051ef",
921 => x"eb3f7a52",
922 => x"0b0b0b0b",
923 => x"80e09851",
924 => x"efde3f0b",
925 => x"0b80e0b4",
926 => x"51efd53f",
927 => x"0b0b80e2",
928 => x"8051efcc",
929 => x"3f81c480",
930 => x"0880f5ec",
931 => x"08317080",
932 => x"f5e80c52",
933 => x"0b0b0b0b",
934 => x"80e0ec51",
935 => x"efb23f80",
936 => x"f5e80856",
937 => x"810b7625",
938 => x"819d3880",
939 => x"e5dc0870",
940 => x"77bd84c0",
941 => x"293580f5",
942 => x"e00c7671",
943 => x"3580f5e4",
944 => x"0c768ddd",
945 => x"297187e8",
946 => x"293581c4",
947 => x"980c5b0b",
948 => x"0b80e0fc",
949 => x"51eef93f",
950 => x"80f5e008",
951 => x"520b0b0b",
952 => x"0b80e1ac",
953 => x"51eee93f",
954 => x"0b0b80e1",
955 => x"b451eee0",
956 => x"3f80f5e4",
957 => x"08520b0b",
958 => x"0b0b80e1",
959 => x"ac51eed0",
960 => x"3f81c498",
961 => x"08520b0b",
962 => x"0b0b80e1",
963 => x"e451eec0",
964 => x"3f0b0b80",
965 => x"e28051ee",
966 => x"b73f800b",
967 => x"800ca13d",
968 => x"0d040b0b",
969 => x"80e28451",
970 => x"f5de3976",
971 => x"0856b053",
972 => x"0b0b7552",
973 => x"0b0b7651",
974 => x"95b53f80",
975 => x"c10b81c4",
976 => x"90335656",
977 => x"f88e390b",
978 => x"0b80e2b4",
979 => x"51ee813f",
980 => x"0b0b80e2",
981 => x"ec51edf8",
982 => x"3f0b0b80",
983 => x"e28051ed",
984 => x"ef3f800b",
985 => x"800ca13d",
986 => x"0d04a13d",
987 => x"ffb80552",
988 => x"0b0b8051",
989 => x"80dc3f9f",
990 => x"530b0b0b",
991 => x"0b80e38c",
992 => x"520b0b7a",
993 => x"5194e83f",
994 => x"777881c4",
995 => x"880c8117",
996 => x"7081ff06",
997 => x"81c49033",
998 => x"520b0b58",
999 => x"565af7db",
1000 => x"39ff1570",
1001 => x"77317e0c",
1002 => x"59800b81",
1003 => x"19595980",
1004 => x"e5dc0878",
1005 => x"25f58b38",
1006 => x"f8873970",
1007 => x"70738232",
1008 => x"70307072",
1009 => x"07802580",
1010 => x"0c520b0b",
1011 => x"520b0b50",
1012 => x"50047070",
1013 => x"70747671",
1014 => x"530b0b54",
1015 => x"0b0b520b",
1016 => x"0b0b0b71",
1017 => x"822e8338",
1018 => x"83517181",
1019 => x"2e9a3881",
1020 => x"72269f38",
1021 => x"71822eb8",
1022 => x"3871842e",
1023 => x"a9387073",
1024 => x"0c70800c",
1025 => x"50505004",
1026 => x"80e40b81",
1027 => x"c4880825",
1028 => x"8b388073",
1029 => x"0c70800c",
1030 => x"50505004",
1031 => x"83730c70",
1032 => x"800c5050",
1033 => x"50048273",
1034 => x"0c70800c",
1035 => x"50505004",
1036 => x"81730c70",
1037 => x"800c5050",
1038 => x"50047074",
1039 => x"74148205",
1040 => x"710c800c",
1041 => x"5004f73d",
1042 => x"0d7b7d7f",
1043 => x"61857205",
1044 => x"70822b75",
1045 => x"71057074",
1046 => x"71708405",
1047 => x"530b0b0c",
1048 => x"5a5a5d5b",
1049 => x"760c7980",
1050 => x"f8180c79",
1051 => x"86720552",
1052 => x"0b0b5758",
1053 => x"5a5a7676",
1054 => x"249e3876",
1055 => x"b329822b",
1056 => x"79710551",
1057 => x"530b0b76",
1058 => x"73708405",
1059 => x"550c8114",
1060 => x"540b0b75",
1061 => x"7425f038",
1062 => x"7681cc29",
1063 => x"19fc7105",
1064 => x"088105fc",
1065 => x"72050c7a",
1066 => x"1970089f",
1067 => x"a073050c",
1068 => x"5856850b",
1069 => x"81c4880c",
1070 => x"75800c8b",
1071 => x"3d0d0470",
1072 => x"70700293",
1073 => x"05335180",
1074 => x"02840597",
1075 => x"0533540b",
1076 => x"0b520b0b",
1077 => x"70732e88",
1078 => x"3871800c",
1079 => x"50505004",
1080 => x"7081c48c",
1081 => x"34810b80",
1082 => x"0c505050",
1083 => x"04f83d0d",
1084 => x"7a7c5956",
1085 => x"820b8319",
1086 => x"55550b0b",
1087 => x"74167033",
1088 => x"75335b51",
1089 => x"530b0b72",
1090 => x"792e80cf",
1091 => x"3880c10b",
1092 => x"81168116",
1093 => x"56565782",
1094 => x"7525df38",
1095 => x"ffa91770",
1096 => x"81ff0655",
1097 => x"590b7382",
1098 => x"26833887",
1099 => x"5581530b",
1100 => x"0b7680d2",
1101 => x"2e9e3877",
1102 => x"520b0b75",
1103 => x"5193b53f",
1104 => x"80530b0b",
1105 => x"72800825",
1106 => x"8b388715",
1107 => x"81c4880c",
1108 => x"81530b0b",
1109 => x"72800c8a",
1110 => x"3d0d0472",
1111 => x"81c48c34",
1112 => x"827525ff",
1113 => x"9538ffb4",
1114 => x"39f93d0d",
1115 => x"797b7d54",
1116 => x"0b0b5872",
1117 => x"59773079",
1118 => x"70307072",
1119 => x"079f2a73",
1120 => x"71315a52",
1121 => x"0b0b5977",
1122 => x"0b795673",
1123 => x"0c530b0b",
1124 => x"73847305",
1125 => x"0c540b0b",
1126 => x"800c893d",
1127 => x"0d04f93d",
1128 => x"0d797b7d",
1129 => x"7f56540b",
1130 => x"0b520b0b",
1131 => x"540b0b72",
1132 => x"802ea638",
1133 => x"70577158",
1134 => x"a0733152",
1135 => x"0b0b800b",
1136 => x"7225a638",
1137 => x"7770742b",
1138 => x"5770732a",
1139 => x"78752b07",
1140 => x"56510b74",
1141 => x"76530b0b",
1142 => x"510b0b70",
1143 => x"740c7184",
1144 => x"150c7380",
1145 => x"0c893d0d",
1146 => x"04805677",
1147 => x"72302b55",
1148 => x"0b0b7476",
1149 => x"530b0b51",
1150 => x"e039fb3d",
1151 => x"0d777955",
1152 => x"5580560b",
1153 => x"0b757524",
1154 => x"b5388074",
1155 => x"24a53880",
1156 => x"530b0b73",
1157 => x"520b0b74",
1158 => x"5180f33f",
1159 => x"8008540b",
1160 => x"0b75802e",
1161 => x"87388008",
1162 => x"30540b0b",
1163 => x"73800c87",
1164 => x"3d0d0473",
1165 => x"30768132",
1166 => x"57540b0b",
1167 => x"d2397430",
1168 => x"55815673",
1169 => x"8025c838",
1170 => x"ea39fa3d",
1171 => x"0d787a57",
1172 => x"5580570b",
1173 => x"0b767524",
1174 => x"ae38759f",
1175 => x"2c540b0b",
1176 => x"81530b0b",
1177 => x"75743274",
1178 => x"31520b0b",
1179 => x"74519f3f",
1180 => x"8008540b",
1181 => x"0b76802e",
1182 => x"87388008",
1183 => x"30540b0b",
1184 => x"73800c88",
1185 => x"3d0d0474",
1186 => x"30558157",
1187 => x"cd39fc3d",
1188 => x"0d767853",
1189 => x"0b0b540b",
1190 => x"0b81530b",
1191 => x"0b807473",
1192 => x"26520b0b",
1193 => x"5572802e",
1194 => x"9e387080",
1195 => x"2eb73880",
1196 => x"7224b238",
1197 => x"71107310",
1198 => x"75722653",
1199 => x"0b0b540b",
1200 => x"0b520b0b",
1201 => x"72e43873",
1202 => x"51788338",
1203 => x"74510b0b",
1204 => x"70800c86",
1205 => x"3d0d0472",
1206 => x"0a100a72",
1207 => x"0a100a53",
1208 => x"0b0b530b",
1209 => x"0b72802e",
1210 => x"de387174",
1211 => x"26e93873",
1212 => x"72317574",
1213 => x"07740a10",
1214 => x"0a740a10",
1215 => x"0a555556",
1216 => x"540b0be1",
1217 => x"39707073",
1218 => x"520b0b80",
1219 => x"eea80851",
1220 => x"953f5050",
1221 => x"04707073",
1222 => x"520b0b80",
1223 => x"eea80851",
1224 => x"92dc3f50",
1225 => x"5004f43d",
1226 => x"0d7e608b",
1227 => x"710570f8",
1228 => x"065b5555",
1229 => x"5d729626",
1230 => x"83389058",
1231 => x"800b7824",
1232 => x"74792607",
1233 => x"5580540b",
1234 => x"0b74742e",
1235 => x"09810680",
1236 => x"d5387c51",
1237 => x"8edf3f77",
1238 => x"83f72680",
1239 => x"d0387783",
1240 => x"2a701010",
1241 => x"1080e6a0",
1242 => x"058c7105",
1243 => x"08585854",
1244 => x"0b0b7577",
1245 => x"2e828a38",
1246 => x"841608fc",
1247 => x"068c1708",
1248 => x"88180871",
1249 => x"8c72050c",
1250 => x"8872050c",
1251 => x"5b760584",
1252 => x"71050881",
1253 => x"07847205",
1254 => x"0c530b0b",
1255 => x"7c518e96",
1256 => x"3f881654",
1257 => x"0b0b7380",
1258 => x"0c8e3d0d",
1259 => x"0477892a",
1260 => x"78832a58",
1261 => x"540b0b73",
1262 => x"802ebf38",
1263 => x"77862ab8",
1264 => x"05578474",
1265 => x"27b43880",
1266 => x"db145794",
1267 => x"7427ab38",
1268 => x"778c2a80",
1269 => x"ee055780",
1270 => x"d474279e",
1271 => x"38778f2a",
1272 => x"80f70557",
1273 => x"82d47427",
1274 => x"91387792",
1275 => x"2a80fc05",
1276 => x"578ad474",
1277 => x"27843880",
1278 => x"fe570b0b",
1279 => x"76101010",
1280 => x"80e6a005",
1281 => x"8c710508",
1282 => x"56530b0b",
1283 => x"74732ea6",
1284 => x"38841508",
1285 => x"fc067079",
1286 => x"3155560b",
1287 => x"738f2489",
1288 => x"d2387380",
1289 => x"2589d438",
1290 => x"8c150855",
1291 => x"0b0b7473",
1292 => x"2e098106",
1293 => x"dc388117",
1294 => x"5980e6b0",
1295 => x"08560b0b",
1296 => x"7580e6a8",
1297 => x"2e82f938",
1298 => x"841608fc",
1299 => x"06707931",
1300 => x"55550b73",
1301 => x"8f2480c2",
1302 => x"3880e6a8",
1303 => x"0b80e6b4",
1304 => x"0c80e6a8",
1305 => x"0b80e6b0",
1306 => x"0c807424",
1307 => x"80e83874",
1308 => x"16847105",
1309 => x"08810784",
1310 => x"72050c53",
1311 => x"0b0bfe9c",
1312 => x"3988168c",
1313 => x"71050857",
1314 => x"590b750b",
1315 => x"792e0981",
1316 => x"06fde538",
1317 => x"821459ff",
1318 => x"a0397716",
1319 => x"78810784",
1320 => x"180c7080",
1321 => x"e6b40c70",
1322 => x"80e6b00c",
1323 => x"80e6a80b",
1324 => x"8c72050c",
1325 => x"8c710508",
1326 => x"8872050c",
1327 => x"74810784",
1328 => x"72050c74",
1329 => x"0574710c",
1330 => x"5b7c518b",
1331 => x"e93f8816",
1332 => x"540b0bfd",
1333 => x"d13983ff",
1334 => x"752783c1",
1335 => x"3874892a",
1336 => x"75832a54",
1337 => x"0b0b540b",
1338 => x"0b73802e",
1339 => x"80cb3874",
1340 => x"862ab805",
1341 => x"530b0b84",
1342 => x"7427be38",
1343 => x"80db1453",
1344 => x"0b0b9474",
1345 => x"27b33874",
1346 => x"8c2a80ee",
1347 => x"05530b0b",
1348 => x"80d47427",
1349 => x"a438748f",
1350 => x"2a80f705",
1351 => x"530b0b82",
1352 => x"d4742795",
1353 => x"3874922a",
1354 => x"80fc0553",
1355 => x"0b0b8ad4",
1356 => x"74278638",
1357 => x"80fe530b",
1358 => x"0b721010",
1359 => x"1080e6a0",
1360 => x"05887105",
1361 => x"0855570b",
1362 => x"730b772e",
1363 => x"86cd3884",
1364 => x"1408fc06",
1365 => x"5b740b7b",
1366 => x"278f3888",
1367 => x"1408540b",
1368 => x"0b73772e",
1369 => x"098106e7",
1370 => x"388c1408",
1371 => x"80e6a00b",
1372 => x"84050871",
1373 => x"8c190c75",
1374 => x"88190c77",
1375 => x"8873050c",
1376 => x"5c57758c",
1377 => x"150c7853",
1378 => x"0b0b8079",
1379 => x"2483be38",
1380 => x"72822c81",
1381 => x"712b5656",
1382 => x"0b747b26",
1383 => x"80d1387a",
1384 => x"7506570b",
1385 => x"0b7682bc",
1386 => x"3878fc06",
1387 => x"84055974",
1388 => x"10707c06",
1389 => x"55550b73",
1390 => x"82aa3884",
1391 => x"1959f039",
1392 => x"80e6a00b",
1393 => x"84050879",
1394 => x"540b0b5b",
1395 => x"788025c0",
1396 => x"3882fa39",
1397 => x"74097b06",
1398 => x"7080e6a0",
1399 => x"0b84050c",
1400 => x"5b741055",
1401 => x"0b0b747b",
1402 => x"26853874",
1403 => x"85f33880",
1404 => x"e6a00b88",
1405 => x"05087084",
1406 => x"720508fc",
1407 => x"06707b31",
1408 => x"7b72268f",
1409 => x"7225075d",
1410 => x"575c5c55",
1411 => x"78802e80",
1412 => x"e3387915",
1413 => x"80e69808",
1414 => x"19907105",
1415 => x"59540b0b",
1416 => x"5680e694",
1417 => x"08ff2e89",
1418 => x"38a08f73",
1419 => x"05e08006",
1420 => x"570b0b76",
1421 => x"520b0b7c",
1422 => x"5188fc3f",
1423 => x"8008540b",
1424 => x"0b8008ff",
1425 => x"2e903880",
1426 => x"08762782",
1427 => x"c2387480",
1428 => x"e6a02e82",
1429 => x"ba3880e6",
1430 => x"a00b8805",
1431 => x"08558415",
1432 => x"08fc0670",
1433 => x"79317972",
1434 => x"268f7225",
1435 => x"075d555a",
1436 => x"7a849b38",
1437 => x"77810784",
1438 => x"160c7715",
1439 => x"7080e6a0",
1440 => x"0b88050c",
1441 => x"74810784",
1442 => x"72050c56",
1443 => x"7c5188a6",
1444 => x"3f881554",
1445 => x"0b0b7380",
1446 => x"0c8e3d0d",
1447 => x"0474832a",
1448 => x"70540b0b",
1449 => x"540b0b80",
1450 => x"742481a9",
1451 => x"3872822c",
1452 => x"81712b80",
1453 => x"e6a40807",
1454 => x"7080e6a0",
1455 => x"0b84050c",
1456 => x"75101010",
1457 => x"80e6a005",
1458 => x"88710508",
1459 => x"718c1b0c",
1460 => x"70881b0c",
1461 => x"79887305",
1462 => x"0c57555c",
1463 => x"55758c15",
1464 => x"0cfda339",
1465 => x"78791010",
1466 => x"1080e6a0",
1467 => x"0570565b",
1468 => x"5c8c1408",
1469 => x"560b0b75",
1470 => x"742ea738",
1471 => x"841608fc",
1472 => x"06707931",
1473 => x"58530b0b",
1474 => x"768f2484",
1475 => x"98387680",
1476 => x"2584de38",
1477 => x"8c160856",
1478 => x"0b0b7574",
1479 => x"2e098106",
1480 => x"db388814",
1481 => x"811a7083",
1482 => x"06555a54",
1483 => x"0b0b72c1",
1484 => x"387b8306",
1485 => x"560b0b75",
1486 => x"802efd98",
1487 => x"38ff1cf8",
1488 => x"1b5b5c88",
1489 => x"1a087a2e",
1490 => x"e838fd95",
1491 => x"39831953",
1492 => x"0b0bfcbc",
1493 => x"39831470",
1494 => x"822c8171",
1495 => x"2b80e6a4",
1496 => x"08077080",
1497 => x"e6a00b84",
1498 => x"050c7610",
1499 => x"101080e6",
1500 => x"a0058871",
1501 => x"0508718c",
1502 => x"1c0c7088",
1503 => x"1c0c7a88",
1504 => x"73050c58",
1505 => x"530b0b5d",
1506 => x"56530b0b",
1507 => x"fecf3980",
1508 => x"e5e40817",
1509 => x"59800876",
1510 => x"2e819438",
1511 => x"80e69408",
1512 => x"ff2e84b7",
1513 => x"38737631",
1514 => x"1980e5e4",
1515 => x"0c738706",
1516 => x"7056530b",
1517 => x"0b72802e",
1518 => x"88388873",
1519 => x"31701555",
1520 => x"5576149f",
1521 => x"ff06a080",
1522 => x"71311670",
1523 => x"540b0b7e",
1524 => x"530b0b51",
1525 => x"530b0b85",
1526 => x"de3f8008",
1527 => x"568008ff",
1528 => x"2e81a238",
1529 => x"80e5e408",
1530 => x"73057080",
1531 => x"e5e40c74",
1532 => x"7580e6a0",
1533 => x"0b88050c",
1534 => x"77763115",
1535 => x"81075556",
1536 => x"597a80e6",
1537 => x"a02e83e0",
1538 => x"38798f26",
1539 => x"838d3881",
1540 => x"0b84150c",
1541 => x"841508fc",
1542 => x"06707931",
1543 => x"7972268f",
1544 => x"7225075d",
1545 => x"555a7a80",
1546 => x"2efcc938",
1547 => x"80e03980",
1548 => x"089fff06",
1549 => x"550b0b74",
1550 => x"fee23878",
1551 => x"80e5e40c",
1552 => x"80e6a00b",
1553 => x"8805087a",
1554 => x"18810784",
1555 => x"72050c55",
1556 => x"80e69008",
1557 => x"79278638",
1558 => x"7880e690",
1559 => x"0c80e68c",
1560 => x"087927fb",
1561 => x"f9387880",
1562 => x"e68c0c84",
1563 => x"1508fc06",
1564 => x"70793179",
1565 => x"72268f72",
1566 => x"25075d55",
1567 => x"5a7a802e",
1568 => x"fbf2388a",
1569 => x"39807457",
1570 => x"530b0bfe",
1571 => x"d7397c51",
1572 => x"84a43f80",
1573 => x"0b800c8e",
1574 => x"3d0d0480",
1575 => x"7324a538",
1576 => x"72822c81",
1577 => x"712b80e6",
1578 => x"a4080770",
1579 => x"80e6a00b",
1580 => x"84050c5c",
1581 => x"5a768c17",
1582 => x"0c738817",
1583 => x"0c758818",
1584 => x"0cf9bf39",
1585 => x"83730570",
1586 => x"822c8171",
1587 => x"2b80e6a4",
1588 => x"08077080",
1589 => x"e6a00b84",
1590 => x"050c5d5b",
1591 => x"530b0bd5",
1592 => x"397a7506",
1593 => x"5c0b0b7b",
1594 => x"fbfa3884",
1595 => x"19751056",
1596 => x"59ef39ff",
1597 => x"17810559",
1598 => x"f6bf398c",
1599 => x"15088816",
1600 => x"08718c72",
1601 => x"050c8872",
1602 => x"050c5975",
1603 => x"15847105",
1604 => x"08810784",
1605 => x"72050c58",
1606 => x"7c51839a",
1607 => x"3f881554",
1608 => x"0b0bfaf2",
1609 => x"39771678",
1610 => x"81078418",
1611 => x"0c8c1708",
1612 => x"88180871",
1613 => x"8c72050c",
1614 => x"8872050c",
1615 => x"5c7080e6",
1616 => x"b40c7080",
1617 => x"e6b00c80",
1618 => x"e6a80b8c",
1619 => x"72050c8c",
1620 => x"71050888",
1621 => x"72050c77",
1622 => x"81078472",
1623 => x"050c7705",
1624 => x"77710c55",
1625 => x"7c5182ce",
1626 => x"3f881654",
1627 => x"0b0bf4b6",
1628 => x"39721684",
1629 => x"71050881",
1630 => x"07847205",
1631 => x"0c588c16",
1632 => x"08881708",
1633 => x"718c7205",
1634 => x"0c887205",
1635 => x"0c577c51",
1636 => x"82a43f88",
1637 => x"16540b0b",
1638 => x"f48c3972",
1639 => x"84150cf4",
1640 => x"1af80670",
1641 => x"841d0881",
1642 => x"0607841d",
1643 => x"0c701c55",
1644 => x"56850b84",
1645 => x"150c850b",
1646 => x"88150c8f",
1647 => x"7627fd90",
1648 => x"38881b52",
1649 => x"0b0b7c51",
1650 => x"85b43f80",
1651 => x"e6a00b88",
1652 => x"050880e5",
1653 => x"e4085a55",
1654 => x"fcf63978",
1655 => x"80e5e40c",
1656 => x"7380e694",
1657 => x"0cfbc639",
1658 => x"7284150c",
1659 => x"fce239fb",
1660 => x"3d0d7770",
1661 => x"7a7c5855",
1662 => x"530b0b56",
1663 => x"8f752781",
1664 => x"85387276",
1665 => x"07830651",
1666 => x"0b0b7080",
1667 => x"f9387573",
1668 => x"520b0b54",
1669 => x"0b0b7070",
1670 => x"8405520b",
1671 => x"0b087470",
1672 => x"8405560c",
1673 => x"73717084",
1674 => x"05530b0b",
1675 => x"08717084",
1676 => x"05530b0b",
1677 => x"0c717084",
1678 => x"05530b0b",
1679 => x"08717084",
1680 => x"05530b0b",
1681 => x"0c717084",
1682 => x"05530b0b",
1683 => x"08717084",
1684 => x"05530b0b",
1685 => x"0cf01656",
1686 => x"540b0b74",
1687 => x"8f26ffb6",
1688 => x"38837527",
1689 => x"99387070",
1690 => x"8405520b",
1691 => x"0b087470",
1692 => x"8405560c",
1693 => x"fc15550b",
1694 => x"0b748326",
1695 => x"e9387371",
1696 => x"540b0b52",
1697 => x"0b0bff15",
1698 => x"510b0b70",
1699 => x"ff2e9f38",
1700 => x"72708105",
1701 => x"540b0b33",
1702 => x"72708105",
1703 => x"540b0b34",
1704 => x"ff710551",
1705 => x"0b0b70ff",
1706 => x"2e098106",
1707 => x"e3387580",
1708 => x"0c873d0d",
1709 => x"04040470",
1710 => x"70707080",
1711 => x"0b81c5e8",
1712 => x"0c765188",
1713 => x"d93f8008",
1714 => x"530b0b80",
1715 => x"08ff2e89",
1716 => x"3872800c",
1717 => x"50505050",
1718 => x"0481c5e8",
1719 => x"08540b0b",
1720 => x"73802eed",
1721 => x"38757471",
1722 => x"0c520b0b",
1723 => x"72800c50",
1724 => x"50505004",
1725 => x"fb3d0d77",
1726 => x"79707207",
1727 => x"8306530b",
1728 => x"0b540b0b",
1729 => x"520b0b70",
1730 => x"9b387173",
1731 => x"7308540b",
1732 => x"0b56540b",
1733 => x"0b717308",
1734 => x"2e80d838",
1735 => x"7375540b",
1736 => x"0b520b0b",
1737 => x"0b0b7133",
1738 => x"7081ff06",
1739 => x"520b0b54",
1740 => x"0b0b7080",
1741 => x"2ea53872",
1742 => x"3355700b",
1743 => x"752e0981",
1744 => x"069c3881",
1745 => x"72058114",
1746 => x"71337081",
1747 => x"ff06540b",
1748 => x"0b56540b",
1749 => x"0b520b0b",
1750 => x"70dd3872",
1751 => x"33557381",
1752 => x"ff067581",
1753 => x"ff067171",
1754 => x"31800c55",
1755 => x"520b0b87",
1756 => x"3d0d0471",
1757 => x"09f7fbfd",
1758 => x"ff730506",
1759 => x"f8848281",
1760 => x"8006520b",
1761 => x"0b0b0b71",
1762 => x"9f388414",
1763 => x"84167108",
1764 => x"540b0b56",
1765 => x"540b0b71",
1766 => x"75082ed7",
1767 => x"38737554",
1768 => x"0b0b520b",
1769 => x"0bfefd39",
1770 => x"800b800c",
1771 => x"873d0d04",
1772 => x"fb3d0d77",
1773 => x"70520b0b",
1774 => x"56fdfa3f",
1775 => x"80e6a00b",
1776 => x"88050884",
1777 => x"710508fc",
1778 => x"06707b31",
1779 => x"9fef05e0",
1780 => x"8006e080",
1781 => x"05520b0b",
1782 => x"5555a080",
1783 => x"75249838",
1784 => x"80520b0b",
1785 => x"7551fdcf",
1786 => x"3f80e6a8",
1787 => x"0814530b",
1788 => x"0b728008",
1789 => x"2e913875",
1790 => x"51fdbb3f",
1791 => x"80530b0b",
1792 => x"72800c87",
1793 => x"3d0d0474",
1794 => x"30520b0b",
1795 => x"7551fda7",
1796 => x"3f8008ff",
1797 => x"2eab3880",
1798 => x"e6a00b88",
1799 => x"05087476",
1800 => x"31810784",
1801 => x"72050c53",
1802 => x"0b0b80e5",
1803 => x"e4087531",
1804 => x"80e5e40c",
1805 => x"7551fcfe",
1806 => x"3f810b80",
1807 => x"0c873d0d",
1808 => x"0480520b",
1809 => x"0b7551fc",
1810 => x"ee3f80e6",
1811 => x"a00b8805",
1812 => x"08800871",
1813 => x"31540b0b",
1814 => x"540b0b8f",
1815 => x"7325ff97",
1816 => x"38800880",
1817 => x"e6940831",
1818 => x"80e5e40c",
1819 => x"72810784",
1820 => x"150c7551",
1821 => x"fcc03f80",
1822 => x"530b0bff",
1823 => x"8339f73d",
1824 => x"0d7b7d54",
1825 => x"0b0b5a72",
1826 => x"802e82ab",
1827 => x"387951fc",
1828 => x"a43ff873",
1829 => x"05847105",
1830 => x"0870fe06",
1831 => x"70730584",
1832 => x"710508fc",
1833 => x"065c5758",
1834 => x"540b0b57",
1835 => x"80e6a808",
1836 => x"742e838b",
1837 => x"38778415",
1838 => x"0c807381",
1839 => x"0656590b",
1840 => x"740b792e",
1841 => x"81f53877",
1842 => x"14847105",
1843 => x"08810656",
1844 => x"530b0b74",
1845 => x"a3387716",
1846 => x"56788287",
1847 => x"38881408",
1848 => x"550b0b74",
1849 => x"80e6a82e",
1850 => x"83a7388c",
1851 => x"1408708c",
1852 => x"170c7588",
1853 => x"72050c58",
1854 => x"75810784",
1855 => x"180c7517",
1856 => x"76710c54",
1857 => x"0b0b7881",
1858 => x"a93883ff",
1859 => x"762781e5",
1860 => x"3875892a",
1861 => x"76832a54",
1862 => x"0b0b540b",
1863 => x"0b73802e",
1864 => x"80cb3875",
1865 => x"862ab805",
1866 => x"530b0b84",
1867 => x"7427be38",
1868 => x"80db1453",
1869 => x"0b0b9474",
1870 => x"27b33875",
1871 => x"8c2a80ee",
1872 => x"05530b0b",
1873 => x"80d47427",
1874 => x"a438758f",
1875 => x"2a80f705",
1876 => x"530b0b82",
1877 => x"d4742795",
1878 => x"3875922a",
1879 => x"80fc0553",
1880 => x"0b0b8ad4",
1881 => x"74278638",
1882 => x"80fe530b",
1883 => x"0b721010",
1884 => x"1080e6a0",
1885 => x"05887105",
1886 => x"0855550b",
1887 => x"730b752e",
1888 => x"82da3884",
1889 => x"1408fc06",
1890 => x"59750b79",
1891 => x"278f3888",
1892 => x"1408540b",
1893 => x"0b73752e",
1894 => x"098106e7",
1895 => x"388c1408",
1896 => x"708c190c",
1897 => x"7488190c",
1898 => x"77887205",
1899 => x"0c55768c",
1900 => x"150c7951",
1901 => x"fa803f8b",
1902 => x"3d0d0476",
1903 => x"08777131",
1904 => x"58760588",
1905 => x"18085656",
1906 => x"0b7480e6",
1907 => x"a82e80ea",
1908 => x"388c1708",
1909 => x"708c170c",
1910 => x"75887205",
1911 => x"0c530b0b",
1912 => x"fde53988",
1913 => x"14088c15",
1914 => x"08708c73",
1915 => x"050c5988",
1916 => x"190cfe84",
1917 => x"3975832a",
1918 => x"70540b0b",
1919 => x"540b0b80",
1920 => x"742481a2",
1921 => x"3872822c",
1922 => x"81712b80",
1923 => x"e6a40807",
1924 => x"80e6a00b",
1925 => x"84050c74",
1926 => x"10101080",
1927 => x"e6a00588",
1928 => x"71050871",
1929 => x"8c1b0c70",
1930 => x"881b0c79",
1931 => x"8873050c",
1932 => x"565a5576",
1933 => x"8c150cfe",
1934 => x"f9398159",
1935 => x"fd893977",
1936 => x"16738106",
1937 => x"540b0b55",
1938 => x"729a3876",
1939 => x"08777131",
1940 => x"5875058c",
1941 => x"18088819",
1942 => x"08718c72",
1943 => x"050c8872",
1944 => x"050c5555",
1945 => x"0b0b7481",
1946 => x"0784180c",
1947 => x"7680e6a0",
1948 => x"0b88050c",
1949 => x"80e69c08",
1950 => x"7526feb6",
1951 => x"3880e698",
1952 => x"08520b0b",
1953 => x"7951faa8",
1954 => x"3f7951f8",
1955 => x"a93ffea7",
1956 => x"3981778c",
1957 => x"170c7788",
1958 => x"170c758c",
1959 => x"190c7588",
1960 => x"190c59fc",
1961 => x"d3398314",
1962 => x"70822c81",
1963 => x"712b80e6",
1964 => x"a4080780",
1965 => x"e6a00b84",
1966 => x"050c7510",
1967 => x"101080e6",
1968 => x"a0058871",
1969 => x"0508718c",
1970 => x"1c0c7088",
1971 => x"1c0c7a88",
1972 => x"73050c57",
1973 => x"5b56530b",
1974 => x"0bfed839",
1975 => x"807324a3",
1976 => x"3872822c",
1977 => x"81712b80",
1978 => x"e6a40807",
1979 => x"80e6a00b",
1980 => x"84050c58",
1981 => x"748c180c",
1982 => x"7388180c",
1983 => x"7688160c",
1984 => x"fdac3983",
1985 => x"73057082",
1986 => x"2c81712b",
1987 => x"80e6a408",
1988 => x"0780e6a0",
1989 => x"0b84050c",
1990 => x"59530b0b",
1991 => x"d7397070",
1992 => x"7081c5ec",
1993 => x"08510b0b",
1994 => x"708a3881",
1995 => x"c5f47081",
1996 => x"c5ec0c51",
1997 => x"740b7105",
1998 => x"520b0bff",
1999 => x"530b0b71",
2000 => x"87fb8080",
2001 => x"268a3871",
2002 => x"81c5ec0c",
2003 => x"70530b0b",
2004 => x"72800c50",
2005 => x"50500470",
2006 => x"70707080",
2007 => x"0b80e5d0",
2008 => x"08540b0b",
2009 => x"540b0b72",
2010 => x"812e9d38",
2011 => x"7381c5f0",
2012 => x"0ccabe3f",
2013 => x"c98a3f80",
2014 => x"f5a8520b",
2015 => x"0b8151d3",
2016 => x"fa3f8008",
2017 => x"518a8f3f",
2018 => x"7281c5f0",
2019 => x"0ccaa23f",
2020 => x"c8ee3f80",
2021 => x"f5a8520b",
2022 => x"0b8151d3",
2023 => x"de3f8008",
2024 => x"5189f33f",
2025 => x"00ff3900",
2026 => x"ff39f53d",
2027 => x"0d7e6081",
2028 => x"c5f00870",
2029 => x"5b585b5b",
2030 => x"7580c538",
2031 => x"777a25a2",
2032 => x"38771b70",
2033 => x"337081ff",
2034 => x"06585859",
2035 => x"758a2e99",
2036 => x"387681ff",
2037 => x"0651c9b4",
2038 => x"3f811858",
2039 => x"790b7824",
2040 => x"e0387980",
2041 => x"0c8d3d0d",
2042 => x"048d51c9",
2043 => x"9f3f7833",
2044 => x"7081ff06",
2045 => x"520b0b57",
2046 => x"c9923f81",
2047 => x"1858dd39",
2048 => x"79557a54",
2049 => x"0b0b7d53",
2050 => x"0b0b8552",
2051 => x"0b0b8d3d",
2052 => x"fc0551c8",
2053 => x"af3f8008",
2054 => x"5688f43f",
2055 => x"7b80080c",
2056 => x"75800c8d",
2057 => x"3d0d04f6",
2058 => x"3d0d7d7f",
2059 => x"81c5f008",
2060 => x"705a585a",
2061 => x"5a7580ca",
2062 => x"38767925",
2063 => x"b638761a",
2064 => x"58c8a53f",
2065 => x"80087834",
2066 => x"800b8008",
2067 => x"81ff0657",
2068 => x"580b758a",
2069 => x"2ea83875",
2070 => x"8d327030",
2071 => x"7080257a",
2072 => x"07515156",
2073 => x"0b0b7580",
2074 => x"c0388117",
2075 => x"57780b77",
2076 => x"24cc3876",
2077 => x"560b0b75",
2078 => x"800c8c3d",
2079 => x"0d048158",
2080 => x"d6397855",
2081 => x"79540b0b",
2082 => x"7c530b0b",
2083 => x"84520b0b",
2084 => x"8c3dfc05",
2085 => x"51c7ad3f",
2086 => x"80085687",
2087 => x"f23f7a80",
2088 => x"080c7580",
2089 => x"0c8c3d0d",
2090 => x"04811756",
2091 => x"c839f93d",
2092 => x"0d795781",
2093 => x"c5f00880",
2094 => x"2eb23876",
2095 => x"518ac03f",
2096 => x"7b567a55",
2097 => x"80088105",
2098 => x"540b0b76",
2099 => x"530b0b82",
2100 => x"520b0b89",
2101 => x"3dfc0551",
2102 => x"c6ea3f80",
2103 => x"085787af",
2104 => x"3f778008",
2105 => x"0c76800c",
2106 => x"893d0d04",
2107 => x"87a13f85",
2108 => x"0b80080c",
2109 => x"ff0b800c",
2110 => x"893d0d04",
2111 => x"fb3d0d81",
2112 => x"c5f00870",
2113 => x"56540b0b",
2114 => x"73883874",
2115 => x"800c873d",
2116 => x"0d047753",
2117 => x"0b0b8352",
2118 => x"0b0b873d",
2119 => x"fc0551c6",
2120 => x"a33f8008",
2121 => x"540b0b86",
2122 => x"e63f7580",
2123 => x"080c7380",
2124 => x"0c873d0d",
2125 => x"04ff0b80",
2126 => x"0c04fb3d",
2127 => x"0d775581",
2128 => x"c5f00880",
2129 => x"2eae3874",
2130 => x"5189b43f",
2131 => x"80088105",
2132 => x"540b0b74",
2133 => x"530b0b87",
2134 => x"520b0b87",
2135 => x"3dfc0551",
2136 => x"c5e23f80",
2137 => x"085586a7",
2138 => x"3f758008",
2139 => x"0c74800c",
2140 => x"873d0d04",
2141 => x"86993f85",
2142 => x"0b80080c",
2143 => x"ff0b800c",
2144 => x"873d0d04",
2145 => x"fa3d0d81",
2146 => x"c5f00880",
2147 => x"2ea8387a",
2148 => x"5579540b",
2149 => x"0b78530b",
2150 => x"0b86520b",
2151 => x"0b883dfc",
2152 => x"0551c5a0",
2153 => x"3f800856",
2154 => x"85e53f76",
2155 => x"80080c75",
2156 => x"800c883d",
2157 => x"0d0485d7",
2158 => x"3f9d0b80",
2159 => x"080cff0b",
2160 => x"800c883d",
2161 => x"0d04f73d",
2162 => x"0d7b7d5b",
2163 => x"59bc530b",
2164 => x"0b80520b",
2165 => x"0b795186",
2166 => x"fd3f8070",
2167 => x"56579856",
2168 => x"74197033",
2169 => x"70782b79",
2170 => x"078118f8",
2171 => x"1a5a5859",
2172 => x"55588475",
2173 => x"24ea3876",
2174 => x"7a238419",
2175 => x"58807056",
2176 => x"57985674",
2177 => x"18703370",
2178 => x"782b7907",
2179 => x"8118f81a",
2180 => x"5a585951",
2181 => x"540b0b84",
2182 => x"7524e838",
2183 => x"76821b23",
2184 => x"88195880",
2185 => x"70565798",
2186 => x"56741870",
2187 => x"3370782b",
2188 => x"79078118",
2189 => x"f81a5a58",
2190 => x"5951540b",
2191 => x"0b847524",
2192 => x"e8387684",
2193 => x"1b0c8c19",
2194 => x"58807056",
2195 => x"57985674",
2196 => x"18703370",
2197 => x"782b7907",
2198 => x"8118f81a",
2199 => x"5a585951",
2200 => x"540b0b84",
2201 => x"7524e838",
2202 => x"76881b23",
2203 => x"90195880",
2204 => x"70565798",
2205 => x"56741870",
2206 => x"3370782b",
2207 => x"79078118",
2208 => x"f81a5a58",
2209 => x"5951540b",
2210 => x"0b847524",
2211 => x"e838768a",
2212 => x"1b239419",
2213 => x"58807056",
2214 => x"57985674",
2215 => x"18703370",
2216 => x"782b7907",
2217 => x"8118f81a",
2218 => x"5a585951",
2219 => x"540b0b84",
2220 => x"7524e838",
2221 => x"768c1b23",
2222 => x"98195880",
2223 => x"70565798",
2224 => x"56741870",
2225 => x"3370782b",
2226 => x"79078118",
2227 => x"f81a5a58",
2228 => x"5951540b",
2229 => x"0b847524",
2230 => x"e838768e",
2231 => x"1b239c19",
2232 => x"58807056",
2233 => x"57b85674",
2234 => x"18703370",
2235 => x"782b7907",
2236 => x"8118f81a",
2237 => x"5a58595a",
2238 => x"540b0b88",
2239 => x"7524e838",
2240 => x"76901b0c",
2241 => x"8b3d0d04",
2242 => x"e93d0d6a",
2243 => x"81c5f008",
2244 => x"57570b75",
2245 => x"933880c0",
2246 => x"800b8418",
2247 => x"0c75ac18",
2248 => x"0c75800c",
2249 => x"993d0d04",
2250 => x"893d7055",
2251 => x"6a540b0b",
2252 => x"558a520b",
2253 => x"0b993dff",
2254 => x"bc0551c2",
2255 => x"873f8008",
2256 => x"77530b0b",
2257 => x"75520b0b",
2258 => x"56fcfb3f",
2259 => x"82c13f77",
2260 => x"80080c75",
2261 => x"800c993d",
2262 => x"0d04e93d",
2263 => x"0d695781",
2264 => x"c5f00880",
2265 => x"2ebd3876",
2266 => x"5185943f",
2267 => x"893d7056",
2268 => x"80088105",
2269 => x"5577540b",
2270 => x"0b568f52",
2271 => x"0b0b993d",
2272 => x"ffbc0551",
2273 => x"c1be3f80",
2274 => x"086b530b",
2275 => x"0b76520b",
2276 => x"0b57fcb2",
2277 => x"3f81f83f",
2278 => x"7780080c",
2279 => x"76800c99",
2280 => x"3d0d0481",
2281 => x"ea3f850b",
2282 => x"80080cff",
2283 => x"0b800c99",
2284 => x"3d0d04fc",
2285 => x"3d0d8154",
2286 => x"0b0b81c5",
2287 => x"f0088838",
2288 => x"73800c86",
2289 => x"3d0d0476",
2290 => x"530b0b97",
2291 => x"b9520b0b",
2292 => x"863dfc05",
2293 => x"51c0ed3f",
2294 => x"8008540b",
2295 => x"0b81b03f",
2296 => x"7480080c",
2297 => x"73800c86",
2298 => x"3d0d04f4",
2299 => x"3d0d7e80",
2300 => x"f5d40870",
2301 => x"0881ff06",
2302 => x"913df805",
2303 => x"540b0b51",
2304 => x"5959c29d",
2305 => x"3f775780",
2306 => x"540b0b76",
2307 => x"557b7d58",
2308 => x"520b0b0b",
2309 => x"76530b0b",
2310 => x"8e3df005",
2311 => x"5184dc3f",
2312 => x"797b5879",
2313 => x"0c76841a",
2314 => x"0c78800c",
2315 => x"8e3d0d04",
2316 => x"f43d0d7e",
2317 => x"80f5d408",
2318 => x"70087081",
2319 => x"ff06923d",
2320 => x"f8055551",
2321 => x"5a5759c1",
2322 => x"d83f7757",
2323 => x"800b8b3d",
2324 => x"59540b0b",
2325 => x"76557b7d",
2326 => x"58520b0b",
2327 => x"0b76530b",
2328 => x"0b775184",
2329 => x"963f8056",
2330 => x"bd84c076",
2331 => x"5555797b",
2332 => x"58520b0b",
2333 => x"0b76530b",
2334 => x"0b775183",
2335 => x"fe3f7a57",
2336 => x"78802e84",
2337 => x"3876790c",
2338 => x"76800c8e",
2339 => x"3d0d0480",
2340 => x"eea80880",
2341 => x"0c04f73d",
2342 => x"0d7b80ee",
2343 => x"a80882c8",
2344 => x"7105085a",
2345 => x"540b0b5a",
2346 => x"77802e80",
2347 => x"eb388188",
2348 => x"18841908",
2349 => x"ff058171",
2350 => x"2b595559",
2351 => x"80742481",
2352 => x"80388074",
2353 => x"2480c138",
2354 => x"73822b78",
2355 => x"71058805",
2356 => x"56568180",
2357 => x"19087706",
2358 => x"530b0b72",
2359 => x"802e80c3",
2360 => x"38781670",
2361 => x"08530b0b",
2362 => x"530b0b79",
2363 => x"51740853",
2364 => x"0b0b722d",
2365 => x"ff14fc17",
2366 => x"fc177981",
2367 => x"2c5a5757",
2368 => x"540b0b73",
2369 => x"8025cb38",
2370 => x"7708580b",
2371 => x"0b77ff9e",
2372 => x"3880eea8",
2373 => x"08530b0b",
2374 => x"bc730508",
2375 => x"a9387951",
2376 => x"f5823f74",
2377 => x"08530b0b",
2378 => x"722dff14",
2379 => x"fc17fc17",
2380 => x"79812c5a",
2381 => x"5757540b",
2382 => x"0b738025",
2383 => x"ff9438c8",
2384 => x"398057fe",
2385 => x"fd397251",
2386 => x"bc730508",
2387 => x"540b0b73",
2388 => x"2d7951f4",
2389 => x"cf3ffb3d",
2390 => x"0d777a71",
2391 => x"028c05a3",
2392 => x"05335854",
2393 => x"0b0b540b",
2394 => x"0b568373",
2395 => x"2780e738",
2396 => x"75830651",
2397 => x"0b0b7080",
2398 => x"dd387488",
2399 => x"2b750770",
2400 => x"71902b07",
2401 => x"55518f73",
2402 => x"27b33873",
2403 => x"72708405",
2404 => x"540b0b0c",
2405 => x"71747170",
2406 => x"8405530b",
2407 => x"0b0c7471",
2408 => x"70840553",
2409 => x"0b0b0c74",
2410 => x"71708405",
2411 => x"530b0b0c",
2412 => x"f014540b",
2413 => x"0b520b0b",
2414 => x"728f26cf",
2415 => x"38837327",
2416 => x"95387372",
2417 => x"70840554",
2418 => x"0b0b0cfc",
2419 => x"7305530b",
2420 => x"0b728326",
2421 => x"ed38ff73",
2422 => x"05510b0b",
2423 => x"70ff2e98",
2424 => x"38747270",
2425 => x"8105540b",
2426 => x"0b34ff71",
2427 => x"05510b0b",
2428 => x"70ff2e09",
2429 => x"8106ea38",
2430 => x"75800c87",
2431 => x"3d0d0470",
2432 => x"70707075",
2433 => x"70718306",
2434 => x"530b0b55",
2435 => x"520b0b70",
2436 => x"80c53871",
2437 => x"70087009",
2438 => x"f7fbfdff",
2439 => x"720506f8",
2440 => x"84828180",
2441 => x"06540b0b",
2442 => x"520b0b53",
2443 => x"0b0b71a3",
2444 => x"38847305",
2445 => x"70087009",
2446 => x"f7fbfdff",
2447 => x"720506f8",
2448 => x"84828180",
2449 => x"06540b0b",
2450 => x"520b0b53",
2451 => x"0b0b7180",
2452 => x"2edf3872",
2453 => x"520b0b0b",
2454 => x"0b713353",
2455 => x"0b0b7280",
2456 => x"2e8f3881",
2457 => x"72057033",
2458 => x"540b0b52",
2459 => x"0b0b72f3",
2460 => x"38717431",
2461 => x"800c5050",
2462 => x"505004e4",
2463 => x"3d0d6ea1",
2464 => x"3d08a33d",
2465 => x"0859575f",
2466 => x"80764d77",
2467 => x"4ea33d08",
2468 => x"a53d0857",
2469 => x"4b0b754c",
2470 => x"5e0b0b7d",
2471 => x"6c2487b2",
2472 => x"38806a24",
2473 => x"87cd3869",
2474 => x"6b58566b",
2475 => x"6d5d460b",
2476 => x"7b477544",
2477 => x"76450b0b",
2478 => x"64646868",
2479 => x"5c5c5656",
2480 => x"0b7481f5",
2481 => x"38787627",
2482 => x"82dd3875",
2483 => x"81ff2683",
2484 => x"2b5583ff",
2485 => x"ff76278c",
2486 => x"389055fe",
2487 => x"800a7627",
2488 => x"83389855",
2489 => x"750b752a",
2490 => x"80e3bc05",
2491 => x"7033a077",
2492 => x"31713157",
2493 => x"55577480",
2494 => x"2e953875",
2495 => x"752ba076",
2496 => x"317a772b",
2497 => x"7c722a07",
2498 => x"7c782b5d",
2499 => x"5b59560b",
2500 => x"0b75902a",
2501 => x"7683ffff",
2502 => x"0671540b",
2503 => x"0b7a530b",
2504 => x"0b595788",
2505 => x"bf3f8008",
2506 => x"5b88a53f",
2507 => x"80088008",
2508 => x"79297c90",
2509 => x"2b7c902a",
2510 => x"07565659",
2511 => x"73752794",
2512 => x"388008ff",
2513 => x"05761555",
2514 => x"59757426",
2515 => x"87387474",
2516 => x"2687f438",
2517 => x"76520b0b",
2518 => x"73753151",
2519 => x"88863f80",
2520 => x"085587ec",
2521 => x"3f800880",
2522 => x"0879297b",
2523 => x"83ffff06",
2524 => x"77902b07",
2525 => x"56595773",
2526 => x"78279638",
2527 => x"8008ff05",
2528 => x"76155557",
2529 => x"75742689",
2530 => x"38777426",
2531 => x"77713158",
2532 => x"5678902b",
2533 => x"77075880",
2534 => x"5b0b0b7a",
2535 => x"4077417f",
2536 => x"0b615654",
2537 => x"0b0b7d80",
2538 => x"dd38737f",
2539 => x"0c747f84",
2540 => x"050c7e80",
2541 => x"0c9e3d0d",
2542 => x"0480705c",
2543 => x"58747926",
2544 => x"d8387481",
2545 => x"ff26832b",
2546 => x"577483ff",
2547 => x"ff2682bd",
2548 => x"3874772a",
2549 => x"80e3bc05",
2550 => x"7033a079",
2551 => x"31713159",
2552 => x"5c5d7682",
2553 => x"cf387654",
2554 => x"0b0b7479",
2555 => x"27853881",
2556 => x"540b0b79",
2557 => x"76277407",
2558 => x"59815878",
2559 => x"ff993876",
2560 => x"58805bff",
2561 => x"94397352",
2562 => x"0b0b7453",
2563 => x"0b0b9e3d",
2564 => x"e80551d2",
2565 => x"d43f6769",
2566 => x"567f0c74",
2567 => x"7f84050c",
2568 => x"7e800c9e",
2569 => x"3d0d0475",
2570 => x"802e81d2",
2571 => x"387581ff",
2572 => x"26832b55",
2573 => x"83ffff76",
2574 => x"278c3890",
2575 => x"55fe800a",
2576 => x"76278338",
2577 => x"9855750b",
2578 => x"752a80e3",
2579 => x"bc057033",
2580 => x"a0773171",
2581 => x"31575e54",
2582 => x"0b0b7484",
2583 => x"b8387876",
2584 => x"31540b0b",
2585 => x"8176902a",
2586 => x"7783ffff",
2587 => x"065f5d5b",
2588 => x"0b7b520b",
2589 => x"0b735185",
2590 => x"eb3f8008",
2591 => x"5785d13f",
2592 => x"80088008",
2593 => x"7e297890",
2594 => x"2b7c902a",
2595 => x"07565659",
2596 => x"73752794",
2597 => x"388008ff",
2598 => x"05761555",
2599 => x"59757426",
2600 => x"87387474",
2601 => x"26859738",
2602 => x"7b520b0b",
2603 => x"73753151",
2604 => x"85b23f80",
2605 => x"08558598",
2606 => x"3f800880",
2607 => x"087e297b",
2608 => x"83ffff06",
2609 => x"77902b07",
2610 => x"56595773",
2611 => x"78279638",
2612 => x"8008ff05",
2613 => x"76155557",
2614 => x"75742689",
2615 => x"38777426",
2616 => x"77713158",
2617 => x"5a78902b",
2618 => x"77077b41",
2619 => x"410b7f0b",
2620 => x"6156540b",
2621 => x"0b7d802e",
2622 => x"fdb038fe",
2623 => x"89397552",
2624 => x"0b0b8151",
2625 => x"84ca3f80",
2626 => x"0856fea1",
2627 => x"399057fe",
2628 => x"800a7527",
2629 => x"fdbb3898",
2630 => x"75712a80",
2631 => x"e3bc0570",
2632 => x"33a07331",
2633 => x"7131530b",
2634 => x"0b5d5e57",
2635 => x"0b0b7680",
2636 => x"2efdb338",
2637 => x"a0773175",
2638 => x"782b7772",
2639 => x"2a077779",
2640 => x"2b7b7a2b",
2641 => x"7d742a07",
2642 => x"7d7b2b73",
2643 => x"902a7483",
2644 => x"ffff0671",
2645 => x"597f772a",
2646 => x"585e5c41",
2647 => x"5f585c54",
2648 => x"0b0b8480",
2649 => x"3f800854",
2650 => x"0b0b83e4",
2651 => x"3f800880",
2652 => x"08792975",
2653 => x"902b7e90",
2654 => x"2a075656",
2655 => x"59737527",
2656 => x"99388008",
2657 => x"ff057b15",
2658 => x"55597a74",
2659 => x"268c3873",
2660 => x"75278738",
2661 => x"ff197b15",
2662 => x"55597652",
2663 => x"0b0b7375",
2664 => x"315183c0",
2665 => x"3f800855",
2666 => x"83a63f80",
2667 => x"08800879",
2668 => x"297d83ff",
2669 => x"ff067790",
2670 => x"2b075659",
2671 => x"57737827",
2672 => x"99388008",
2673 => x"ff057b15",
2674 => x"55577a74",
2675 => x"268c3873",
2676 => x"78278738",
2677 => x"ff177b15",
2678 => x"55570b73",
2679 => x"78317990",
2680 => x"2b780770",
2681 => x"83ffff06",
2682 => x"71902a79",
2683 => x"83ffff06",
2684 => x"7a902a73",
2685 => x"72297373",
2686 => x"29747329",
2687 => x"76742973",
2688 => x"902a0572",
2689 => x"05575543",
2690 => x"5f5b585a",
2691 => x"57595a74",
2692 => x"7c278638",
2693 => x"84808017",
2694 => x"5774902a",
2695 => x"177983ff",
2696 => x"ff067684",
2697 => x"80802905",
2698 => x"57570b0b",
2699 => x"767a269a",
2700 => x"38767a32",
2701 => x"70307072",
2702 => x"07802556",
2703 => x"5a5b7c76",
2704 => x"27fad438",
2705 => x"73802efa",
2706 => x"ce38ff18",
2707 => x"58805bfa",
2708 => x"c839ff76",
2709 => x"530b0b77",
2710 => x"540b0b9f",
2711 => x"3de80552",
2712 => x"0b0b5ece",
2713 => x"843f6769",
2714 => x"574c0b75",
2715 => x"4d698025",
2716 => x"f8b5387d",
2717 => x"096a6c5c",
2718 => x"530b0b7a",
2719 => x"540b0b9f",
2720 => x"3de80552",
2721 => x"0b0b5ecd",
2722 => x"e03f6769",
2723 => x"714c704d",
2724 => x"5856f897",
2725 => x"39a07531",
2726 => x"76762b7a",
2727 => x"772b7c73",
2728 => x"2a077c78",
2729 => x"2b72902a",
2730 => x"7383ffff",
2731 => x"0671587e",
2732 => x"762a5742",
2733 => x"405d5d57",
2734 => x"5881a93f",
2735 => x"80085781",
2736 => x"8f3f8008",
2737 => x"80087e29",
2738 => x"78902b7d",
2739 => x"902a0756",
2740 => x"56597375",
2741 => x"27993880",
2742 => x"08ff0576",
2743 => x"15555975",
2744 => x"74268c38",
2745 => x"73752787",
2746 => x"38ff1976",
2747 => x"1555597b",
2748 => x"520b0b73",
2749 => x"75315180",
2750 => x"eb3f8008",
2751 => x"5580d13f",
2752 => x"80088008",
2753 => x"7e297c83",
2754 => x"ffff0670",
2755 => x"78902b07",
2756 => x"51565858",
2757 => x"73772799",
2758 => x"388008ff",
2759 => x"05761555",
2760 => x"58757426",
2761 => x"8c387377",
2762 => x"278738ff",
2763 => x"18761555",
2764 => x"5878902b",
2765 => x"78077478",
2766 => x"31555bfa",
2767 => x"b339ff19",
2768 => x"76155559",
2769 => x"fae239ff",
2770 => x"19761555",
2771 => x"59f88539",
2772 => x"70707080",
2773 => x"530b0b75",
2774 => x"520b0b74",
2775 => x"51ceaf3f",
2776 => x"50505004",
2777 => x"70707081",
2778 => x"530b0b75",
2779 => x"520b0b74",
2780 => x"51ce9b3f",
2781 => x"50505004",
2782 => x"707080f5",
2783 => x"b00bfc05",
2784 => x"7008520b",
2785 => x"0b520b0b",
2786 => x"0b70ff2e",
2787 => x"9738702d",
2788 => x"fc720570",
2789 => x"08520b0b",
2790 => x"520b0b0b",
2791 => x"70ff2e09",
2792 => x"8106eb38",
2793 => x"50500404",
2794 => x"ffb4963f",
2795 => x"04000000",
2796 => x"30313233",
2797 => x"34353637",
2798 => x"38390000",
2799 => x"44485259",
2800 => x"53544f4e",
2801 => x"45205052",
2802 => x"4f475241",
2803 => x"4d2c2053",
2804 => x"4f4d4520",
2805 => x"53545249",
2806 => x"4e470000",
2807 => x"44485259",
2808 => x"53544f4e",
2809 => x"45205052",
2810 => x"4f475241",
2811 => x"4d2c2031",
2812 => x"27535420",
2813 => x"53545249",
2814 => x"4e470000",
2815 => x"44687279",
2816 => x"73746f6e",
2817 => x"65204265",
2818 => x"6e63686d",
2819 => x"61726b2c",
2820 => x"20566572",
2821 => x"73696f6e",
2822 => x"20322e31",
2823 => x"20284c61",
2824 => x"6e677561",
2825 => x"67653a20",
2826 => x"43290a00",
2827 => x"50726f67",
2828 => x"72616d20",
2829 => x"636f6d70",
2830 => x"696c6564",
2831 => x"20776974",
2832 => x"68202772",
2833 => x"65676973",
2834 => x"74657227",
2835 => x"20617474",
2836 => x"72696275",
2837 => x"74650a00",
2838 => x"45786563",
2839 => x"7574696f",
2840 => x"6e207374",
2841 => x"61727473",
2842 => x"2c202564",
2843 => x"2072756e",
2844 => x"73207468",
2845 => x"726f7567",
2846 => x"68204468",
2847 => x"72797374",
2848 => x"6f6e650a",
2849 => x"00000000",
2850 => x"44485259",
2851 => x"53544f4e",
2852 => x"45205052",
2853 => x"4f475241",
2854 => x"4d2c2032",
2855 => x"274e4420",
2856 => x"53545249",
2857 => x"4e470000",
2858 => x"45786563",
2859 => x"7574696f",
2860 => x"6e20656e",
2861 => x"64730a00",
2862 => x"46696e61",
2863 => x"6c207661",
2864 => x"6c756573",
2865 => x"206f6620",
2866 => x"74686520",
2867 => x"76617269",
2868 => x"61626c65",
2869 => x"73207573",
2870 => x"65642069",
2871 => x"6e207468",
2872 => x"65206265",
2873 => x"6e63686d",
2874 => x"61726b3a",
2875 => x"0a000000",
2876 => x"496e745f",
2877 => x"476c6f62",
2878 => x"3a202020",
2879 => x"20202020",
2880 => x"20202020",
2881 => x"2025640a",
2882 => x"00000000",
2883 => x"20202020",
2884 => x"20202020",
2885 => x"73686f75",
2886 => x"6c642062",
2887 => x"653a2020",
2888 => x"2025640a",
2889 => x"00000000",
2890 => x"426f6f6c",
2891 => x"5f476c6f",
2892 => x"623a2020",
2893 => x"20202020",
2894 => x"20202020",
2895 => x"2025640a",
2896 => x"00000000",
2897 => x"43685f31",
2898 => x"5f476c6f",
2899 => x"623a2020",
2900 => x"20202020",
2901 => x"20202020",
2902 => x"2025630a",
2903 => x"00000000",
2904 => x"20202020",
2905 => x"20202020",
2906 => x"73686f75",
2907 => x"6c642062",
2908 => x"653a2020",
2909 => x"2025630a",
2910 => x"00000000",
2911 => x"43685f32",
2912 => x"5f476c6f",
2913 => x"623a2020",
2914 => x"20202020",
2915 => x"20202020",
2916 => x"2025630a",
2917 => x"00000000",
2918 => x"4172725f",
2919 => x"315f476c",
2920 => x"6f625b38",
2921 => x"5d3a2020",
2922 => x"20202020",
2923 => x"2025640a",
2924 => x"00000000",
2925 => x"4172725f",
2926 => x"325f476c",
2927 => x"6f625b38",
2928 => x"5d5b375d",
2929 => x"3a202020",
2930 => x"2025640a",
2931 => x"00000000",
2932 => x"20202020",
2933 => x"20202020",
2934 => x"73686f75",
2935 => x"6c642062",
2936 => x"653a2020",
2937 => x"204e756d",
2938 => x"6265725f",
2939 => x"4f665f52",
2940 => x"756e7320",
2941 => x"2b203130",
2942 => x"0a000000",
2943 => x"5074725f",
2944 => x"476c6f62",
2945 => x"2d3e0a00",
2946 => x"20205074",
2947 => x"725f436f",
2948 => x"6d703a20",
2949 => x"20202020",
2950 => x"20202020",
2951 => x"2025640a",
2952 => x"00000000",
2953 => x"20202020",
2954 => x"20202020",
2955 => x"73686f75",
2956 => x"6c642062",
2957 => x"653a2020",
2958 => x"2028696d",
2959 => x"706c656d",
2960 => x"656e7461",
2961 => x"74696f6e",
2962 => x"2d646570",
2963 => x"656e6465",
2964 => x"6e74290a",
2965 => x"00000000",
2966 => x"20204469",
2967 => x"7363723a",
2968 => x"20202020",
2969 => x"20202020",
2970 => x"20202020",
2971 => x"2025640a",
2972 => x"00000000",
2973 => x"2020456e",
2974 => x"756d5f43",
2975 => x"6f6d703a",
2976 => x"20202020",
2977 => x"20202020",
2978 => x"2025640a",
2979 => x"00000000",
2980 => x"2020496e",
2981 => x"745f436f",
2982 => x"6d703a20",
2983 => x"20202020",
2984 => x"20202020",
2985 => x"2025640a",
2986 => x"00000000",
2987 => x"20205374",
2988 => x"725f436f",
2989 => x"6d703a20",
2990 => x"20202020",
2991 => x"20202020",
2992 => x"2025730a",
2993 => x"00000000",
2994 => x"20202020",
2995 => x"20202020",
2996 => x"73686f75",
2997 => x"6c642062",
2998 => x"653a2020",
2999 => x"20444852",
3000 => x"5953544f",
3001 => x"4e452050",
3002 => x"524f4752",
3003 => x"414d2c20",
3004 => x"534f4d45",
3005 => x"20535452",
3006 => x"494e470a",
3007 => x"00000000",
3008 => x"4e657874",
3009 => x"5f507472",
3010 => x"5f476c6f",
3011 => x"622d3e0a",
3012 => x"00000000",
3013 => x"20202020",
3014 => x"20202020",
3015 => x"73686f75",
3016 => x"6c642062",
3017 => x"653a2020",
3018 => x"2028696d",
3019 => x"706c656d",
3020 => x"656e7461",
3021 => x"74696f6e",
3022 => x"2d646570",
3023 => x"656e6465",
3024 => x"6e74292c",
3025 => x"2073616d",
3026 => x"65206173",
3027 => x"2061626f",
3028 => x"76650a00",
3029 => x"496e745f",
3030 => x"315f4c6f",
3031 => x"633a2020",
3032 => x"20202020",
3033 => x"20202020",
3034 => x"2025640a",
3035 => x"00000000",
3036 => x"496e745f",
3037 => x"325f4c6f",
3038 => x"633a2020",
3039 => x"20202020",
3040 => x"20202020",
3041 => x"2025640a",
3042 => x"00000000",
3043 => x"496e745f",
3044 => x"335f4c6f",
3045 => x"633a2020",
3046 => x"20202020",
3047 => x"20202020",
3048 => x"2025640a",
3049 => x"00000000",
3050 => x"456e756d",
3051 => x"5f4c6f63",
3052 => x"3a202020",
3053 => x"20202020",
3054 => x"20202020",
3055 => x"2025640a",
3056 => x"00000000",
3057 => x"5374725f",
3058 => x"315f4c6f",
3059 => x"633a2020",
3060 => x"20202020",
3061 => x"20202020",
3062 => x"2025730a",
3063 => x"00000000",
3064 => x"20202020",
3065 => x"20202020",
3066 => x"73686f75",
3067 => x"6c642062",
3068 => x"653a2020",
3069 => x"20444852",
3070 => x"5953544f",
3071 => x"4e452050",
3072 => x"524f4752",
3073 => x"414d2c20",
3074 => x"31275354",
3075 => x"20535452",
3076 => x"494e470a",
3077 => x"00000000",
3078 => x"5374725f",
3079 => x"325f4c6f",
3080 => x"633a2020",
3081 => x"20202020",
3082 => x"20202020",
3083 => x"2025730a",
3084 => x"00000000",
3085 => x"20202020",
3086 => x"20202020",
3087 => x"73686f75",
3088 => x"6c642062",
3089 => x"653a2020",
3090 => x"20444852",
3091 => x"5953544f",
3092 => x"4e452050",
3093 => x"524f4752",
3094 => x"414d2c20",
3095 => x"32274e44",
3096 => x"20535452",
3097 => x"494e470a",
3098 => x"00000000",
3099 => x"55736572",
3100 => x"2074696d",
3101 => x"653a2025",
3102 => x"640a0000",
3103 => x"4d696372",
3104 => x"6f736563",
3105 => x"6f6e6473",
3106 => x"20666f72",
3107 => x"206f6e65",
3108 => x"2072756e",
3109 => x"20746872",
3110 => x"6f756768",
3111 => x"20446872",
3112 => x"7973746f",
3113 => x"6e653a20",
3114 => x"00000000",
3115 => x"2564200a",
3116 => x"00000000",
3117 => x"44687279",
3118 => x"73746f6e",
3119 => x"65732070",
3120 => x"65722053",
3121 => x"65636f6e",
3122 => x"643a2020",
3123 => x"20202020",
3124 => x"20202020",
3125 => x"20202020",
3126 => x"20202020",
3127 => x"20202020",
3128 => x"00000000",
3129 => x"56415820",
3130 => x"4d495053",
3131 => x"20726174",
3132 => x"696e6720",
3133 => x"2a203130",
3134 => x"3030203d",
3135 => x"20256420",
3136 => x"0a000000",
3137 => x"50726f67",
3138 => x"72616d20",
3139 => x"636f6d70",
3140 => x"696c6564",
3141 => x"20776974",
3142 => x"686f7574",
3143 => x"20277265",
3144 => x"67697374",
3145 => x"65722720",
3146 => x"61747472",
3147 => x"69627574",
3148 => x"650a0000",
3149 => x"4d656173",
3150 => x"75726564",
3151 => x"2074696d",
3152 => x"6520746f",
3153 => x"6f20736d",
3154 => x"616c6c20",
3155 => x"746f206f",
3156 => x"62746169",
3157 => x"6e206d65",
3158 => x"616e696e",
3159 => x"6766756c",
3160 => x"20726573",
3161 => x"756c7473",
3162 => x"0a000000",
3163 => x"506c6561",
3164 => x"73652069",
3165 => x"6e637265",
3166 => x"61736520",
3167 => x"6e756d62",
3168 => x"6572206f",
3169 => x"66207275",
3170 => x"6e730a00",
3171 => x"44485259",
3172 => x"53544f4e",
3173 => x"45205052",
3174 => x"4f475241",
3175 => x"4d2c2033",
3176 => x"27524420",
3177 => x"53545249",
3178 => x"4e470000",
3179 => x"43000000",
3180 => x"64756d6d",
3181 => x"792e6578",
3182 => x"65000000",
3183 => x"00010202",
3184 => x"03030303",
3185 => x"04040404",
3186 => x"04040404",
3187 => x"05050505",
3188 => x"05050505",
3189 => x"05050505",
3190 => x"05050505",
3191 => x"06060606",
3192 => x"06060606",
3193 => x"06060606",
3194 => x"06060606",
3195 => x"06060606",
3196 => x"06060606",
3197 => x"06060606",
3198 => x"06060606",
3199 => x"07070707",
3200 => x"07070707",
3201 => x"07070707",
3202 => x"07070707",
3203 => x"07070707",
3204 => x"07070707",
3205 => x"07070707",
3206 => x"07070707",
3207 => x"07070707",
3208 => x"07070707",
3209 => x"07070707",
3210 => x"07070707",
3211 => x"07070707",
3212 => x"07070707",
3213 => x"07070707",
3214 => x"07070707",
3215 => x"08080808",
3216 => x"08080808",
3217 => x"08080808",
3218 => x"08080808",
3219 => x"08080808",
3220 => x"08080808",
3221 => x"08080808",
3222 => x"08080808",
3223 => x"08080808",
3224 => x"08080808",
3225 => x"08080808",
3226 => x"08080808",
3227 => x"08080808",
3228 => x"08080808",
3229 => x"08080808",
3230 => x"08080808",
3231 => x"08080808",
3232 => x"08080808",
3233 => x"08080808",
3234 => x"08080808",
3235 => x"08080808",
3236 => x"08080808",
3237 => x"08080808",
3238 => x"08080808",
3239 => x"08080808",
3240 => x"08080808",
3241 => x"08080808",
3242 => x"08080808",
3243 => x"08080808",
3244 => x"08080808",
3245 => x"08080808",
3246 => x"08080808",
3247 => x"00ffffff",
3248 => x"ff00ffff",
3249 => x"ffff00ff",
3250 => x"ffffff00",
3251 => x"00000000",
3252 => x"00000000",
3253 => x"00000000",
3254 => x"00003ab8",
3255 => x"000186a0", -- iterations
3256 => x"00000000",
3257 => x"00000000",
3258 => x"00000000",
3259 => x"00000000",
3260 => x"00000000",
3261 => x"00000000",
3262 => x"00000000",
3263 => x"00000000",
3264 => x"00000000",
3265 => x"00000000",
3266 => x"00000000",
3267 => x"00000000",
3268 => x"00000000",
3269 => x"ffffffff",
3270 => x"00000000",
3271 => x"00020000",
3272 => x"00000000",
3273 => x"00000000",
3274 => x"00003320",
3275 => x"00003320",
3276 => x"00003328",
3277 => x"00003328",
3278 => x"00003330",
3279 => x"00003330",
3280 => x"00003338",
3281 => x"00003338",
3282 => x"00003340",
3283 => x"00003340",
3284 => x"00003348",
3285 => x"00003348",
3286 => x"00003350",
3287 => x"00003350",
3288 => x"00003358",
3289 => x"00003358",
3290 => x"00003360",
3291 => x"00003360",
3292 => x"00003368",
3293 => x"00003368",
3294 => x"00003370",
3295 => x"00003370",
3296 => x"00003378",
3297 => x"00003378",
3298 => x"00003380",
3299 => x"00003380",
3300 => x"00003388",
3301 => x"00003388",
3302 => x"00003390",
3303 => x"00003390",
3304 => x"00003398",
3305 => x"00003398",
3306 => x"000033a0",
3307 => x"000033a0",
3308 => x"000033a8",
3309 => x"000033a8",
3310 => x"000033b0",
3311 => x"000033b0",
3312 => x"000033b8",
3313 => x"000033b8",
3314 => x"000033c0",
3315 => x"000033c0",
3316 => x"000033c8",
3317 => x"000033c8",
3318 => x"000033d0",
3319 => x"000033d0",
3320 => x"000033d8",
3321 => x"000033d8",
3322 => x"000033e0",
3323 => x"000033e0",
3324 => x"000033e8",
3325 => x"000033e8",
3326 => x"000033f0",
3327 => x"000033f0",
3328 => x"000033f8",
3329 => x"000033f8",
3330 => x"00003400",
3331 => x"00003400",
3332 => x"00003408",
3333 => x"00003408",
3334 => x"00003410",
3335 => x"00003410",
3336 => x"00003418",
3337 => x"00003418",
3338 => x"00003420",
3339 => x"00003420",
3340 => x"00003428",
3341 => x"00003428",
3342 => x"00003430",
3343 => x"00003430",
3344 => x"00003438",
3345 => x"00003438",
3346 => x"00003440",
3347 => x"00003440",
3348 => x"00003448",
3349 => x"00003448",
3350 => x"00003450",
3351 => x"00003450",
3352 => x"00003458",
3353 => x"00003458",
3354 => x"00003460",
3355 => x"00003460",
3356 => x"00003468",
3357 => x"00003468",
3358 => x"00003470",
3359 => x"00003470",
3360 => x"00003478",
3361 => x"00003478",
3362 => x"00003480",
3363 => x"00003480",
3364 => x"00003488",
3365 => x"00003488",
3366 => x"00003490",
3367 => x"00003490",
3368 => x"00003498",
3369 => x"00003498",
3370 => x"000034a0",
3371 => x"000034a0",
3372 => x"000034a8",
3373 => x"000034a8",
3374 => x"000034b0",
3375 => x"000034b0",
3376 => x"000034b8",
3377 => x"000034b8",
3378 => x"000034c0",
3379 => x"000034c0",
3380 => x"000034c8",
3381 => x"000034c8",
3382 => x"000034d0",
3383 => x"000034d0",
3384 => x"000034d8",
3385 => x"000034d8",
3386 => x"000034e0",
3387 => x"000034e0",
3388 => x"000034e8",
3389 => x"000034e8",
3390 => x"000034f0",
3391 => x"000034f0",
3392 => x"000034f8",
3393 => x"000034f8",
3394 => x"00003500",
3395 => x"00003500",
3396 => x"00003508",
3397 => x"00003508",
3398 => x"00003510",
3399 => x"00003510",
3400 => x"00003518",
3401 => x"00003518",
3402 => x"00003520",
3403 => x"00003520",
3404 => x"00003528",
3405 => x"00003528",
3406 => x"00003530",
3407 => x"00003530",
3408 => x"00003538",
3409 => x"00003538",
3410 => x"00003540",
3411 => x"00003540",
3412 => x"00003548",
3413 => x"00003548",
3414 => x"00003550",
3415 => x"00003550",
3416 => x"00003558",
3417 => x"00003558",
3418 => x"00003560",
3419 => x"00003560",
3420 => x"00003568",
3421 => x"00003568",
3422 => x"00003570",
3423 => x"00003570",
3424 => x"00003578",
3425 => x"00003578",
3426 => x"00003580",
3427 => x"00003580",
3428 => x"00003588",
3429 => x"00003588",
3430 => x"00003590",
3431 => x"00003590",
3432 => x"00003598",
3433 => x"00003598",
3434 => x"000035a0",
3435 => x"000035a0",
3436 => x"000035a8",
3437 => x"000035a8",
3438 => x"000035b0",
3439 => x"000035b0",
3440 => x"000035b8",
3441 => x"000035b8",
3442 => x"000035c0",
3443 => x"000035c0",
3444 => x"000035c8",
3445 => x"000035c8",
3446 => x"000035d0",
3447 => x"000035d0",
3448 => x"000035d8",
3449 => x"000035d8",
3450 => x"000035e0",
3451 => x"000035e0",
3452 => x"000035e8",
3453 => x"000035e8",
3454 => x"000035f0",
3455 => x"000035f0",
3456 => x"000035f8",
3457 => x"000035f8",
3458 => x"00003600",
3459 => x"00003600",
3460 => x"00003608",
3461 => x"00003608",
3462 => x"00003610",
3463 => x"00003610",
3464 => x"00003618",
3465 => x"00003618",
3466 => x"00003620",
3467 => x"00003620",
3468 => x"00003628",
3469 => x"00003628",
3470 => x"00003630",
3471 => x"00003630",
3472 => x"00003638",
3473 => x"00003638",
3474 => x"00003640",
3475 => x"00003640",
3476 => x"00003648",
3477 => x"00003648",
3478 => x"00003650",
3479 => x"00003650",
3480 => x"00003658",
3481 => x"00003658",
3482 => x"00003660",
3483 => x"00003660",
3484 => x"00003668",
3485 => x"00003668",
3486 => x"00003670",
3487 => x"00003670",
3488 => x"00003678",
3489 => x"00003678",
3490 => x"00003680",
3491 => x"00003680",
3492 => x"00003688",
3493 => x"00003688",
3494 => x"00003690",
3495 => x"00003690",
3496 => x"00003698",
3497 => x"00003698",
3498 => x"000036a0",
3499 => x"000036a0",
3500 => x"000036a8",
3501 => x"000036a8",
3502 => x"000036b0",
3503 => x"000036b0",
3504 => x"000036b8",
3505 => x"000036b8",
3506 => x"000036c0",
3507 => x"000036c0",
3508 => x"000036c8",
3509 => x"000036c8",
3510 => x"000036d0",
3511 => x"000036d0",
3512 => x"000036d8",
3513 => x"000036d8",
3514 => x"000036e0",
3515 => x"000036e0",
3516 => x"000036e8",
3517 => x"000036e8",
3518 => x"000036f0",
3519 => x"000036f0",
3520 => x"000036f8",
3521 => x"000036f8",
3522 => x"00003700",
3523 => x"00003700",
3524 => x"00003708",
3525 => x"00003708",
3526 => x"00003710",
3527 => x"00003710",
3528 => x"00003718",
3529 => x"00003718",
3530 => x"0000372c",
3531 => x"00000000",
3532 => x"00003994",
3533 => x"000039f0",
3534 => x"00003a4c",
3535 => x"00000000",
3536 => x"00000000",
3537 => x"00000000",
3538 => x"00000000",
3539 => x"00000000",
3540 => x"00000000",
3541 => x"00000000",
3542 => x"00000000",
3543 => x"00000000",
3544 => x"000031ac",
3545 => x"00000000",
3546 => x"00000000",
3547 => x"00000000",
3548 => x"00000000",
3549 => x"00000000",
3550 => x"00000000",
3551 => x"00000000",
3552 => x"00000000",
3553 => x"00000000",
3554 => x"00000000",
3555 => x"00000000",
3556 => x"00000000",
3557 => x"00000000",
3558 => x"00000000",
3559 => x"00000000",
3560 => x"00000000",
3561 => x"00000000",
3562 => x"00000000",
3563 => x"00000000",
3564 => x"00000000",
3565 => x"00000000",
3566 => x"00000000",
3567 => x"00000000",
3568 => x"00000000",
3569 => x"00000000",
3570 => x"00000000",
3571 => x"00000000",
3572 => x"00000000",
3573 => x"00000001",
3574 => x"330eabcd",
3575 => x"1234e66d",
3576 => x"deec0005",
3577 => x"000b0000",
3578 => x"00000000",
3579 => x"00000000",
3580 => x"00000000",
3581 => x"00000000",
3582 => x"00000000",
3583 => x"00000000",
3584 => x"00000000",
3585 => x"00000000",
3586 => x"00000000",
3587 => x"00000000",
3588 => x"00000000",
3589 => x"00000000",
3590 => x"00000000",
3591 => x"00000000",
3592 => x"00000000",
3593 => x"00000000",
3594 => x"00000000",
3595 => x"00000000",
3596 => x"00000000",
3597 => x"00000000",
3598 => x"00000000",
3599 => x"00000000",
3600 => x"00000000",
3601 => x"00000000",
3602 => x"00000000",
3603 => x"00000000",
3604 => x"00000000",
3605 => x"00000000",
3606 => x"00000000",
3607 => x"00000000",
3608 => x"00000000",
3609 => x"00000000",
3610 => x"00000000",
3611 => x"00000000",
3612 => x"00000000",
3613 => x"00000000",
3614 => x"00000000",
3615 => x"00000000",
3616 => x"00000000",
3617 => x"00000000",
3618 => x"00000000",
3619 => x"00000000",
3620 => x"00000000",
3621 => x"00000000",
3622 => x"00000000",
3623 => x"00000000",
3624 => x"00000000",
3625 => x"00000000",
3626 => x"00000000",
3627 => x"00000000",
3628 => x"00000000",
3629 => x"00000000",
3630 => x"00000000",
3631 => x"00000000",
3632 => x"00000000",
3633 => x"00000000",
3634 => x"00000000",
3635 => x"00000000",
3636 => x"00000000",
3637 => x"00000000",
3638 => x"00000000",
3639 => x"00000000",
3640 => x"00000000",
3641 => x"00000000",
3642 => x"00000000",
3643 => x"00000000",
3644 => x"00000000",
3645 => x"00000000",
3646 => x"00000000",
3647 => x"00000000",
3648 => x"00000000",
3649 => x"00000000",
3650 => x"00000000",
3651 => x"00000000",
3652 => x"00000000",
3653 => x"00000000",
3654 => x"00000000",
3655 => x"00000000",
3656 => x"00000000",
3657 => x"00000000",
3658 => x"00000000",
3659 => x"00000000",
3660 => x"00000000",
3661 => x"00000000",
3662 => x"00000000",
3663 => x"00000000",
3664 => x"00000000",
3665 => x"00000000",
3666 => x"00000000",
3667 => x"00000000",
3668 => x"00000000",
3669 => x"00000000",
3670 => x"00000000",
3671 => x"00000000",
3672 => x"00000000",
3673 => x"00000000",
3674 => x"00000000",
3675 => x"00000000",
3676 => x"00000000",
3677 => x"00000000",
3678 => x"00000000",
3679 => x"00000000",
3680 => x"00000000",
3681 => x"00000000",
3682 => x"00000000",
3683 => x"00000000",
3684 => x"00000000",
3685 => x"00000000",
3686 => x"00000000",
3687 => x"00000000",
3688 => x"00000000",
3689 => x"00000000",
3690 => x"00000000",
3691 => x"00000000",
3692 => x"00000000",
3693 => x"00000000",
3694 => x"00000000",
3695 => x"00000000",
3696 => x"00000000",
3697 => x"00000000",
3698 => x"00000000",
3699 => x"00000000",
3700 => x"00000000",
3701 => x"00000000",
3702 => x"00000000",
3703 => x"00000000",
3704 => x"00000000",
3705 => x"00000000",
3706 => x"00000000",
3707 => x"00000000",
3708 => x"00000000",
3709 => x"00000000",
3710 => x"00000000",
3711 => x"00000000",
3712 => x"00000000",
3713 => x"00000000",
3714 => x"00000000",
3715 => x"00000000",
3716 => x"00000000",
3717 => x"00000000",
3718 => x"00000000",
3719 => x"00000000",
3720 => x"00000000",
3721 => x"00000000",
3722 => x"00000000",
3723 => x"00000000",
3724 => x"00000000",
3725 => x"00000000",
3726 => x"00000000",
3727 => x"00000000",
3728 => x"00000000",
3729 => x"00000000",
3730 => x"00000000",
3731 => x"00000000",
3732 => x"00000000",
3733 => x"00000000",
3734 => x"00000000",
3735 => x"00000000",
3736 => x"00000000",
3737 => x"00000000",
3738 => x"00000000",
3739 => x"00000000",
3740 => x"00000000",
3741 => x"00000000",
3742 => x"00000000",
3743 => x"00000000",
3744 => x"00000000",
3745 => x"00000000",
3746 => x"00000000",
3747 => x"00000000",
3748 => x"00000000",
3749 => x"00000000",
3750 => x"00000000",
3751 => x"00000000",
3752 => x"00000000",
3753 => x"00000000",
3754 => x"000031b0",
3755 => x"ffffffff",
3756 => x"00000000",
3757 => x"ffffffff",
3758 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(conv_integer(memAAddr)) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(conv_integer(memAAddr));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(conv_integer(memBAddr)) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(conv_integer(memBAddr));
		end if;
	end if;
end process;




end dualport_ram_arch;
