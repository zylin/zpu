
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 15;
constant bytes : integer := 28492;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B80F5";
    when 16#00001# => romdata <= X"E4040000";
    when 16#00002# => romdata <= X"00000000";
    when 16#00003# => romdata <= X"00000000";
    when 16#00004# => romdata <= X"00000000";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"0B0B80F8";
    when 16#00009# => romdata <= X"CB040000";
    when 16#0000A# => romdata <= X"00000000";
    when 16#0000B# => romdata <= X"00000000";
    when 16#0000C# => romdata <= X"00000000";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B80F7";
    when 16#00049# => romdata <= X"FD040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B80F7E0";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B81CE";
    when 16#000A2# => romdata <= X"D0738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B80";
    when 16#000A5# => romdata <= X"F7E30400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"0B0B80F8";
    when 16#000A9# => romdata <= X"B2040000";
    when 16#000AA# => romdata <= X"00000000";
    when 16#000AB# => romdata <= X"00000000";
    when 16#000AC# => romdata <= X"00000000";
    when 16#000AD# => romdata <= X"00000000";
    when 16#000AE# => romdata <= X"00000000";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"0B0B80F8";
    when 16#000B1# => romdata <= X"99040000";
    when 16#000B2# => romdata <= X"00000000";
    when 16#000B3# => romdata <= X"00000000";
    when 16#000B4# => romdata <= X"00000000";
    when 16#000B5# => romdata <= X"00000000";
    when 16#000B6# => romdata <= X"00000000";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"81CEE00C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"FF3D0D02";
    when 16#00101# => romdata <= X"8F053370";
    when 16#00102# => romdata <= X"525280F5";
    when 16#00103# => romdata <= X"A63F7151";
    when 16#00104# => romdata <= X"80F6943F";
    when 16#00105# => romdata <= X"71B00C83";
    when 16#00106# => romdata <= X"3D0D04FF";
    when 16#00107# => romdata <= X"3D0D81CE";
    when 16#00108# => romdata <= X"BC08B811";
    when 16#00109# => romdata <= X"08535180";
    when 16#0010A# => romdata <= X"0BB8120C";
    when 16#0010B# => romdata <= X"71B00C83";
    when 16#0010C# => romdata <= X"3D0D0480";
    when 16#0010D# => romdata <= X"0B81F1F0";
    when 16#0010E# => romdata <= X"34800BB0";
    when 16#0010F# => romdata <= X"0C04FB3D";
    when 16#00110# => romdata <= X"0D815180";
    when 16#00111# => romdata <= X"C7CE3FB0";
    when 16#00112# => romdata <= X"08538251";
    when 16#00113# => romdata <= X"80C7C53F";
    when 16#00114# => romdata <= X"B00856B0";
    when 16#00115# => romdata <= X"08833890";
    when 16#00116# => romdata <= X"5672FC06";
    when 16#00117# => romdata <= X"5575812E";
    when 16#00118# => romdata <= X"80FB3880";
    when 16#00119# => romdata <= X"54737627";
    when 16#0011A# => romdata <= X"AD387383";
    when 16#0011B# => romdata <= X"06537280";
    when 16#0011C# => romdata <= X"2EB23881";
    when 16#0011D# => romdata <= X"C2C05180";
    when 16#0011E# => romdata <= X"F0923F74";
    when 16#0011F# => romdata <= X"70840556";
    when 16#00120# => romdata <= X"0852A051";
    when 16#00121# => romdata <= X"80F0A83F";
    when 16#00122# => romdata <= X"A05180EF";
    when 16#00123# => romdata <= X"E53F8114";
    when 16#00124# => romdata <= X"54757426";
    when 16#00125# => romdata <= X"D5388A51";
    when 16#00126# => romdata <= X"80EFD73F";
    when 16#00127# => romdata <= X"800BB00C";
    when 16#00128# => romdata <= X"873D0D04";
    when 16#00129# => romdata <= X"81A7D051";
    when 16#0012A# => romdata <= X"80EFE13F";
    when 16#0012B# => romdata <= X"7452A051";
    when 16#0012C# => romdata <= X"80EFFC3F";
    when 16#0012D# => romdata <= X"81B4BC51";
    when 16#0012E# => romdata <= X"80EFD13F";
    when 16#0012F# => romdata <= X"81C2C051";
    when 16#00130# => romdata <= X"80EFC93F";
    when 16#00131# => romdata <= X"74708405";
    when 16#00132# => romdata <= X"560852A0";
    when 16#00133# => romdata <= X"5180EFDF";
    when 16#00134# => romdata <= X"3FA05180";
    when 16#00135# => romdata <= X"EF9C3F81";
    when 16#00136# => romdata <= X"1454FFB5";
    when 16#00137# => romdata <= X"3981C2C0";
    when 16#00138# => romdata <= X"5180EFA8";
    when 16#00139# => romdata <= X"3F740852";
    when 16#0013A# => romdata <= X"A05180EF";
    when 16#0013B# => romdata <= X"C23F8A51";
    when 16#0013C# => romdata <= X"80EEFF3F";
    when 16#0013D# => romdata <= X"800BB00C";
    when 16#0013E# => romdata <= X"873D0D04";
    when 16#0013F# => romdata <= X"FC3D0D81";
    when 16#00140# => romdata <= X"5180C690";
    when 16#00141# => romdata <= X"3FB00852";
    when 16#00142# => romdata <= X"825180C4";
    when 16#00143# => romdata <= X"D53FB008";
    when 16#00144# => romdata <= X"81FF0672";
    when 16#00145# => romdata <= X"56538354";
    when 16#00146# => romdata <= X"72802EA2";
    when 16#00147# => romdata <= X"38735180";
    when 16#00148# => romdata <= X"C5F23F81";
    when 16#00149# => romdata <= X"147081FF";
    when 16#0014A# => romdata <= X"06FF1570";
    when 16#0014B# => romdata <= X"81FF06B0";
    when 16#0014C# => romdata <= X"08797084";
    when 16#0014D# => romdata <= X"055B0C56";
    when 16#0014E# => romdata <= X"52555272";
    when 16#0014F# => romdata <= X"E03872B0";
    when 16#00150# => romdata <= X"0C863D0D";
    when 16#00151# => romdata <= X"04803D0D";
    when 16#00152# => romdata <= X"8C5180EE";
    when 16#00153# => romdata <= X"A53F800B";
    when 16#00154# => romdata <= X"B00C823D";
    when 16#00155# => romdata <= X"0D04FB3D";
    when 16#00156# => romdata <= X"0D800B81";
    when 16#00157# => romdata <= X"A7D45256";
    when 16#00158# => romdata <= X"80EEA93F";
    when 16#00159# => romdata <= X"75557410";
    when 16#0015A# => romdata <= X"81FE0653";
    when 16#0015B# => romdata <= X"81D05281";
    when 16#0015C# => romdata <= X"CEE80851";
    when 16#0015D# => romdata <= X"80D2D33F";
    when 16#0015E# => romdata <= X"B008982B";
    when 16#0015F# => romdata <= X"54807424";
    when 16#00160# => romdata <= X"A23881A7";
    when 16#00161# => romdata <= X"E05180EE";
    when 16#00162# => romdata <= X"833F7452";
    when 16#00163# => romdata <= X"885180EE";
    when 16#00164# => romdata <= X"9E3F81A7";
    when 16#00165# => romdata <= X"EC5180ED";
    when 16#00166# => romdata <= X"F33F8116";
    when 16#00167# => romdata <= X"7083FFFF";
    when 16#00168# => romdata <= X"06575481";
    when 16#00169# => romdata <= X"157081FF";
    when 16#0016A# => romdata <= X"0670982B";
    when 16#0016B# => romdata <= X"52565473";
    when 16#0016C# => romdata <= X"8025FFB2";
    when 16#0016D# => romdata <= X"3875B00C";
    when 16#0016E# => romdata <= X"873D0D04";
    when 16#0016F# => romdata <= X"F33D0D7F";
    when 16#00170# => romdata <= X"02840580";
    when 16#00171# => romdata <= X"C3053302";
    when 16#00172# => romdata <= X"880580C6";
    when 16#00173# => romdata <= X"052281A7";
    when 16#00174# => romdata <= X"FC545B55";
    when 16#00175# => romdata <= X"5880EDB4";
    when 16#00176# => romdata <= X"3F785180";
    when 16#00177# => romdata <= X"EEF83F81";
    when 16#00178# => romdata <= X"A8885180";
    when 16#00179# => romdata <= X"EDA63F73";
    when 16#0017A# => romdata <= X"52885180";
    when 16#0017B# => romdata <= X"EDC13F81";
    when 16#0017C# => romdata <= X"A8A45180";
    when 16#0017D# => romdata <= X"ED963F80";
    when 16#0017E# => romdata <= X"57767927";
    when 16#0017F# => romdata <= X"81A13873";
    when 16#00180# => romdata <= X"108E3D5D";
    when 16#00181# => romdata <= X"5A7981FF";
    when 16#00182# => romdata <= X"06538190";
    when 16#00183# => romdata <= X"52775180";
    when 16#00184# => romdata <= X"D1B83F76";
    when 16#00185# => romdata <= X"882A5390";
    when 16#00186# => romdata <= X"52775180";
    when 16#00187# => romdata <= X"D1AC3F76";
    when 16#00188# => romdata <= X"81FF0653";
    when 16#00189# => romdata <= X"90527751";
    when 16#0018A# => romdata <= X"80D19F3F";
    when 16#0018B# => romdata <= X"811A7081";
    when 16#0018C# => romdata <= X"FF065455";
    when 16#0018D# => romdata <= X"81905277";
    when 16#0018E# => romdata <= X"5180D18E";
    when 16#0018F# => romdata <= X"3F805380";
    when 16#00190# => romdata <= X"E0527751";
    when 16#00191# => romdata <= X"80D1833F";
    when 16#00192# => romdata <= X"B008982B";
    when 16#00193# => romdata <= X"54807424";
    when 16#00194# => romdata <= X"8A388818";
    when 16#00195# => romdata <= X"087081FF";
    when 16#00196# => romdata <= X"065C567A";
    when 16#00197# => romdata <= X"81FF0681";
    when 16#00198# => romdata <= X"C2C05256";
    when 16#00199# => romdata <= X"80ECA53F";
    when 16#0019A# => romdata <= X"75528851";
    when 16#0019B# => romdata <= X"80ECC03F";
    when 16#0019C# => romdata <= X"81B29851";
    when 16#0019D# => romdata <= X"80EC953F";
    when 16#0019E# => romdata <= X"E0165480";
    when 16#0019F# => romdata <= X"DF7427B6";
    when 16#001A0# => romdata <= X"38768706";
    when 16#001A1# => romdata <= X"701D5755";
    when 16#001A2# => romdata <= X"A0763474";
    when 16#001A3# => romdata <= X"872EB938";
    when 16#001A4# => romdata <= X"81177083";
    when 16#001A5# => romdata <= X"FFFF0658";
    when 16#001A6# => romdata <= X"55787726";
    when 16#001A7# => romdata <= X"FEE73880";
    when 16#001A8# => romdata <= X"E00B8C19";
    when 16#001A9# => romdata <= X"0C8C1808";
    when 16#001AA# => romdata <= X"70812A81";
    when 16#001AB# => romdata <= X"06585A76";
    when 16#001AC# => romdata <= X"F4388F3D";
    when 16#001AD# => romdata <= X"0D047687";
    when 16#001AE# => romdata <= X"06701D55";
    when 16#001AF# => romdata <= X"55757434";
    when 16#001B0# => romdata <= X"74872E09";
    when 16#001B1# => romdata <= X"8106C938";
    when 16#001B2# => romdata <= X"7B5180EB";
    when 16#001B3# => romdata <= X"BF3F8A51";
    when 16#001B4# => romdata <= X"80EB9F3F";
    when 16#001B5# => romdata <= X"81177083";
    when 16#001B6# => romdata <= X"FFFF0658";
    when 16#001B7# => romdata <= X"55787726";
    when 16#001B8# => romdata <= X"FEA338FF";
    when 16#001B9# => romdata <= X"BA39FB3D";
    when 16#001BA# => romdata <= X"0D815180";
    when 16#001BB# => romdata <= X"C0F43FB0";
    when 16#001BC# => romdata <= X"0881FF06";
    when 16#001BD# => romdata <= X"54825180";
    when 16#001BE# => romdata <= X"C29A3FB0";
    when 16#001BF# => romdata <= X"0881FF06";
    when 16#001C0# => romdata <= X"56835180";
    when 16#001C1# => romdata <= X"C0DC3FB0";
    when 16#001C2# => romdata <= X"0883FFFF";
    when 16#001C3# => romdata <= X"0655739C";
    when 16#001C4# => romdata <= X"3881CEE8";
    when 16#001C5# => romdata <= X"08547484";
    when 16#001C6# => romdata <= X"38818055";
    when 16#001C7# => romdata <= X"74537552";
    when 16#001C8# => romdata <= X"7351FD98";
    when 16#001C9# => romdata <= X"3F74B00C";
    when 16#001CA# => romdata <= X"873D0D04";
    when 16#001CB# => romdata <= X"81CEEC08";
    when 16#001CC# => romdata <= X"54E439F8";
    when 16#001CD# => romdata <= X"3D0D02AA";
    when 16#001CE# => romdata <= X"052281CE";
    when 16#001CF# => romdata <= X"C43381F7";
    when 16#001D0# => romdata <= X"06585876";
    when 16#001D1# => romdata <= X"81CEC434";
    when 16#001D2# => romdata <= X"81CEE808";
    when 16#001D3# => romdata <= X"5580C053";
    when 16#001D4# => romdata <= X"81905274";
    when 16#001D5# => romdata <= X"5180CEF2";
    when 16#001D6# => romdata <= X"3F745180";
    when 16#001D7# => romdata <= X"CF9E3FB0";
    when 16#001D8# => romdata <= X"0881FF06";
    when 16#001D9# => romdata <= X"5473802E";
    when 16#001DA# => romdata <= X"84903876";
    when 16#001DB# => romdata <= X"5380D052";
    when 16#001DC# => romdata <= X"745180CE";
    when 16#001DD# => romdata <= X"D53F8059";
    when 16#001DE# => romdata <= X"8F5781CE";
    when 16#001DF# => romdata <= X"C43381FE";
    when 16#001E0# => romdata <= X"06547381";
    when 16#001E1# => romdata <= X"CEC43481";
    when 16#001E2# => romdata <= X"CEE80874";
    when 16#001E3# => romdata <= X"575580C0";
    when 16#001E4# => romdata <= X"53819052";
    when 16#001E5# => romdata <= X"745180CE";
    when 16#001E6# => romdata <= X"B13F7451";
    when 16#001E7# => romdata <= X"80CEDD3F";
    when 16#001E8# => romdata <= X"B00881FF";
    when 16#001E9# => romdata <= X"06547380";
    when 16#001EA# => romdata <= X"2E83C438";
    when 16#001EB# => romdata <= X"755380D0";
    when 16#001EC# => romdata <= X"52745180";
    when 16#001ED# => romdata <= X"CE943F77";
    when 16#001EE# => romdata <= X"772C8106";
    when 16#001EF# => romdata <= X"5574802E";
    when 16#001F0# => romdata <= X"83A23881";
    when 16#001F1# => romdata <= X"CEC43382";
    when 16#001F2# => romdata <= X"07547381";
    when 16#001F3# => romdata <= X"CEC43481";
    when 16#001F4# => romdata <= X"CEE80874";
    when 16#001F5# => romdata <= X"575580C0";
    when 16#001F6# => romdata <= X"53819052";
    when 16#001F7# => romdata <= X"745180CD";
    when 16#001F8# => romdata <= X"E93F7451";
    when 16#001F9# => romdata <= X"80CE953F";
    when 16#001FA# => romdata <= X"B00881FF";
    when 16#001FB# => romdata <= X"06547380";
    when 16#001FC# => romdata <= X"2E82E638";
    when 16#001FD# => romdata <= X"755380D0";
    when 16#001FE# => romdata <= X"52745180";
    when 16#001FF# => romdata <= X"CDCC3F81";
    when 16#00200# => romdata <= X"CEE80855";
    when 16#00201# => romdata <= X"80C15381";
    when 16#00202# => romdata <= X"90527451";
    when 16#00203# => romdata <= X"80CDBB3F";
    when 16#00204# => romdata <= X"745180CD";
    when 16#00205# => romdata <= X"E73FB008";
    when 16#00206# => romdata <= X"81FF0656";
    when 16#00207# => romdata <= X"75802E82";
    when 16#00208# => romdata <= X"8C388053";
    when 16#00209# => romdata <= X"80E05274";
    when 16#0020A# => romdata <= X"5180CD9E";
    when 16#0020B# => romdata <= X"3F745180";
    when 16#0020C# => romdata <= X"CDCA3FB0";
    when 16#0020D# => romdata <= X"0881FF06";
    when 16#0020E# => romdata <= X"5473802E";
    when 16#0020F# => romdata <= X"81EF3888";
    when 16#00210# => romdata <= X"15087090";
    when 16#00211# => romdata <= X"2B70902C";
    when 16#00212# => romdata <= X"56565673";
    when 16#00213# => romdata <= X"822A8106";
    when 16#00214# => romdata <= X"5473802E";
    when 16#00215# => romdata <= X"8D388177";
    when 16#00216# => romdata <= X"2B790770";
    when 16#00217# => romdata <= X"83FFFF06";
    when 16#00218# => romdata <= X"5A5681CE";
    when 16#00219# => romdata <= X"C4338107";
    when 16#0021A# => romdata <= X"547381CE";
    when 16#0021B# => romdata <= X"C43481CE";
    when 16#0021C# => romdata <= X"E8087457";
    when 16#0021D# => romdata <= X"5580C053";
    when 16#0021E# => romdata <= X"81905274";
    when 16#0021F# => romdata <= X"5180CCCA";
    when 16#00220# => romdata <= X"3F745180";
    when 16#00221# => romdata <= X"CCF63FB0";
    when 16#00222# => romdata <= X"0881FF06";
    when 16#00223# => romdata <= X"5473802E";
    when 16#00224# => romdata <= X"81A83875";
    when 16#00225# => romdata <= X"5380D052";
    when 16#00226# => romdata <= X"745180CC";
    when 16#00227# => romdata <= X"AD3F7681";
    when 16#00228# => romdata <= X"800A2981";
    when 16#00229# => romdata <= X"FF0A0570";
    when 16#0022A# => romdata <= X"982C5856";
    when 16#0022B# => romdata <= X"768025FD";
    when 16#0022C# => romdata <= X"C93881CE";
    when 16#0022D# => romdata <= X"C4338207";
    when 16#0022E# => romdata <= X"577681CE";
    when 16#0022F# => romdata <= X"C43481CE";
    when 16#00230# => romdata <= X"E8085580";
    when 16#00231# => romdata <= X"C0538190";
    when 16#00232# => romdata <= X"52745180";
    when 16#00233# => romdata <= X"CBFC3F74";
    when 16#00234# => romdata <= X"5180CCA8";
    when 16#00235# => romdata <= X"3FB00881";
    when 16#00236# => romdata <= X"FF065877";
    when 16#00237# => romdata <= X"802E81B8";
    when 16#00238# => romdata <= X"38765380";
    when 16#00239# => romdata <= X"D0527451";
    when 16#0023A# => romdata <= X"80CBDF3F";
    when 16#0023B# => romdata <= X"81CEC433";
    when 16#0023C# => romdata <= X"88075776";
    when 16#0023D# => romdata <= X"81CEC434";
    when 16#0023E# => romdata <= X"81CEE808";
    when 16#0023F# => romdata <= X"5580C053";
    when 16#00240# => romdata <= X"81905274";
    when 16#00241# => romdata <= X"5180CBC2";
    when 16#00242# => romdata <= X"3F745180";
    when 16#00243# => romdata <= X"CBEE3FB0";
    when 16#00244# => romdata <= X"0881FF06";
    when 16#00245# => romdata <= X"5877802E";
    when 16#00246# => romdata <= X"80EF3876";
    when 16#00247# => romdata <= X"5380D052";
    when 16#00248# => romdata <= X"745180CB";
    when 16#00249# => romdata <= X"A53F78B0";
    when 16#0024A# => romdata <= X"0C8A3D0D";
    when 16#0024B# => romdata <= X"0481A8A8";
    when 16#0024C# => romdata <= X"5180E6D8";
    when 16#0024D# => romdata <= X"3FFF54FE";
    when 16#0024E# => romdata <= X"923981A8";
    when 16#0024F# => romdata <= X"A85180E6";
    when 16#00250# => romdata <= X"CB3F7681";
    when 16#00251# => romdata <= X"800A2981";
    when 16#00252# => romdata <= X"FF0A0570";
    when 16#00253# => romdata <= X"982C5856";
    when 16#00254# => romdata <= X"768025FC";
    when 16#00255# => romdata <= X"A538FEDA";
    when 16#00256# => romdata <= X"3981A8A8";
    when 16#00257# => romdata <= X"5180E6AC";
    when 16#00258# => romdata <= X"3FFD9C39";
    when 16#00259# => romdata <= X"81CEC433";
    when 16#0025A# => romdata <= X"81FD0654";
    when 16#0025B# => romdata <= X"FCDC3981";
    when 16#0025C# => romdata <= X"A8A85180";
    when 16#0025D# => romdata <= X"E6963FFC";
    when 16#0025E# => romdata <= X"BE3981A8";
    when 16#0025F# => romdata <= X"A85180E6";
    when 16#00260# => romdata <= X"8B3F8059";
    when 16#00261# => romdata <= X"8F57FBF2";
    when 16#00262# => romdata <= X"3981A8A8";
    when 16#00263# => romdata <= X"5180E5FC";
    when 16#00264# => romdata <= X"3F78B00C";
    when 16#00265# => romdata <= X"8A3D0D04";
    when 16#00266# => romdata <= X"81A8A851";
    when 16#00267# => romdata <= X"80E5ED3F";
    when 16#00268# => romdata <= X"FECA39FF";
    when 16#00269# => romdata <= X"3D0D8151";
    when 16#0026A# => romdata <= X"BBB83FB0";
    when 16#0026B# => romdata <= X"0881FF06";
    when 16#0026C# => romdata <= X"52818051";
    when 16#0026D# => romdata <= X"FAFD3F82";
    when 16#0026E# => romdata <= X"8051FAF7";
    when 16#0026F# => romdata <= X"3F848351";
    when 16#00270# => romdata <= X"FAF13F86";
    when 16#00271# => romdata <= X"F151FAEB";
    when 16#00272# => romdata <= X"3F71832B";
    when 16#00273# => romdata <= X"88830751";
    when 16#00274# => romdata <= X"FAE13F71";
    when 16#00275# => romdata <= X"B00C833D";
    when 16#00276# => romdata <= X"0D04FE3D";
    when 16#00277# => romdata <= X"0D029305";
    when 16#00278# => romdata <= X"33028405";
    when 16#00279# => romdata <= X"97053354";
    when 16#0027A# => romdata <= X"52717327";
    when 16#0027B# => romdata <= X"9438A051";
    when 16#0027C# => romdata <= X"80E4FF3F";
    when 16#0027D# => romdata <= X"81127081";
    when 16#0027E# => romdata <= X"FF065152";
    when 16#0027F# => romdata <= X"727226EE";
    when 16#00280# => romdata <= X"38843D0D";
    when 16#00281# => romdata <= X"04FE3D0D";
    when 16#00282# => romdata <= X"74708106";
    when 16#00283# => romdata <= X"53537185";
    when 16#00284# => romdata <= X"D0387281";
    when 16#00285# => romdata <= X"2A708106";
    when 16#00286# => romdata <= X"51527185";
    when 16#00287# => romdata <= X"AC387282";
    when 16#00288# => romdata <= X"2A708106";
    when 16#00289# => romdata <= X"51527185";
    when 16#0028A# => romdata <= X"88387283";
    when 16#0028B# => romdata <= X"2A708106";
    when 16#0028C# => romdata <= X"51527184";
    when 16#0028D# => romdata <= X"E4387284";
    when 16#0028E# => romdata <= X"2A708106";
    when 16#0028F# => romdata <= X"51527184";
    when 16#00290# => romdata <= X"C0387285";
    when 16#00291# => romdata <= X"2A708106";
    when 16#00292# => romdata <= X"51527184";
    when 16#00293# => romdata <= X"9C387286";
    when 16#00294# => romdata <= X"2A708106";
    when 16#00295# => romdata <= X"51527183";
    when 16#00296# => romdata <= X"F8387287";
    when 16#00297# => romdata <= X"2A708106";
    when 16#00298# => romdata <= X"51527183";
    when 16#00299# => romdata <= X"D4387288";
    when 16#0029A# => romdata <= X"2A708106";
    when 16#0029B# => romdata <= X"51527183";
    when 16#0029C# => romdata <= X"B0387289";
    when 16#0029D# => romdata <= X"2A708106";
    when 16#0029E# => romdata <= X"51527183";
    when 16#0029F# => romdata <= X"8C38728A";
    when 16#002A0# => romdata <= X"2A708106";
    when 16#002A1# => romdata <= X"51527182";
    when 16#002A2# => romdata <= X"E838728B";
    when 16#002A3# => romdata <= X"2A708106";
    when 16#002A4# => romdata <= X"51527182";
    when 16#002A5# => romdata <= X"C438728C";
    when 16#002A6# => romdata <= X"2A708106";
    when 16#002A7# => romdata <= X"51527182";
    when 16#002A8# => romdata <= X"A038728D";
    when 16#002A9# => romdata <= X"2A708106";
    when 16#002AA# => romdata <= X"51527181";
    when 16#002AB# => romdata <= X"FC38728E";
    when 16#002AC# => romdata <= X"2A708106";
    when 16#002AD# => romdata <= X"51527181";
    when 16#002AE# => romdata <= X"D838728F";
    when 16#002AF# => romdata <= X"2A708106";
    when 16#002B0# => romdata <= X"51527181";
    when 16#002B1# => romdata <= X"B4387290";
    when 16#002B2# => romdata <= X"2A708106";
    when 16#002B3# => romdata <= X"51527181";
    when 16#002B4# => romdata <= X"90387291";
    when 16#002B5# => romdata <= X"2A708106";
    when 16#002B6# => romdata <= X"51527180";
    when 16#002B7# => romdata <= X"EC387292";
    when 16#002B8# => romdata <= X"2A708106";
    when 16#002B9# => romdata <= X"51527180";
    when 16#002BA# => romdata <= X"C8387293";
    when 16#002BB# => romdata <= X"2A708106";
    when 16#002BC# => romdata <= X"515271A6";
    when 16#002BD# => romdata <= X"3872942A";
    when 16#002BE# => romdata <= X"70810651";
    when 16#002BF# => romdata <= X"52718B38";
    when 16#002C0# => romdata <= X"80732483";
    when 16#002C1# => romdata <= X"F438843D";
    when 16#002C2# => romdata <= X"0D0481A8";
    when 16#002C3# => romdata <= X"E05180E2";
    when 16#002C4# => romdata <= X"FB3F7280";
    when 16#002C5# => romdata <= X"25F03883";
    when 16#002C6# => romdata <= X"E03981A8";
    when 16#002C7# => romdata <= X"FC5180E2";
    when 16#002C8# => romdata <= X"EB3F7294";
    when 16#002C9# => romdata <= X"2A708106";
    when 16#002CA# => romdata <= X"51527180";
    when 16#002CB# => romdata <= X"2ED238DA";
    when 16#002CC# => romdata <= X"3981A998";
    when 16#002CD# => romdata <= X"5180E2D4";
    when 16#002CE# => romdata <= X"3F72932A";
    when 16#002CF# => romdata <= X"70810651";
    when 16#002D0# => romdata <= X"5271802E";
    when 16#002D1# => romdata <= X"FFAF38D2";
    when 16#002D2# => romdata <= X"3981A9B4";
    when 16#002D3# => romdata <= X"5180E2BC";
    when 16#002D4# => romdata <= X"3F72922A";
    when 16#002D5# => romdata <= X"70810651";
    when 16#002D6# => romdata <= X"5271802E";
    when 16#002D7# => romdata <= X"FF8C38D1";
    when 16#002D8# => romdata <= X"3981A9D0";
    when 16#002D9# => romdata <= X"5180E2A4";
    when 16#002DA# => romdata <= X"3F72912A";
    when 16#002DB# => romdata <= X"70810651";
    when 16#002DC# => romdata <= X"5271802E";
    when 16#002DD# => romdata <= X"FEE838D1";
    when 16#002DE# => romdata <= X"3981A9F0";
    when 16#002DF# => romdata <= X"5180E28C";
    when 16#002E0# => romdata <= X"3F72902A";
    when 16#002E1# => romdata <= X"70810651";
    when 16#002E2# => romdata <= X"5271802E";
    when 16#002E3# => romdata <= X"FEC438D1";
    when 16#002E4# => romdata <= X"3981AA90";
    when 16#002E5# => romdata <= X"5180E1F4";
    when 16#002E6# => romdata <= X"3F728F2A";
    when 16#002E7# => romdata <= X"70810651";
    when 16#002E8# => romdata <= X"5271802E";
    when 16#002E9# => romdata <= X"FEA038D1";
    when 16#002EA# => romdata <= X"3981AAB0";
    when 16#002EB# => romdata <= X"5180E1DC";
    when 16#002EC# => romdata <= X"3F728E2A";
    when 16#002ED# => romdata <= X"70810651";
    when 16#002EE# => romdata <= X"5271802E";
    when 16#002EF# => romdata <= X"FDFC38D1";
    when 16#002F0# => romdata <= X"3981AAD0";
    when 16#002F1# => romdata <= X"5180E1C4";
    when 16#002F2# => romdata <= X"3F728D2A";
    when 16#002F3# => romdata <= X"70810651";
    when 16#002F4# => romdata <= X"5271802E";
    when 16#002F5# => romdata <= X"FDD838D1";
    when 16#002F6# => romdata <= X"3981AAE4";
    when 16#002F7# => romdata <= X"5180E1AC";
    when 16#002F8# => romdata <= X"3F728C2A";
    when 16#002F9# => romdata <= X"70810651";
    when 16#002FA# => romdata <= X"5271802E";
    when 16#002FB# => romdata <= X"FDB438D1";
    when 16#002FC# => romdata <= X"3981AB84";
    when 16#002FD# => romdata <= X"5180E194";
    when 16#002FE# => romdata <= X"3F728B2A";
    when 16#002FF# => romdata <= X"70810651";
    when 16#00300# => romdata <= X"5271802E";
    when 16#00301# => romdata <= X"FD9038D1";
    when 16#00302# => romdata <= X"3981ABAC";
    when 16#00303# => romdata <= X"5180E0FC";
    when 16#00304# => romdata <= X"3F728A2A";
    when 16#00305# => romdata <= X"70810651";
    when 16#00306# => romdata <= X"5271802E";
    when 16#00307# => romdata <= X"FCEC38D1";
    when 16#00308# => romdata <= X"3981ABCC";
    when 16#00309# => romdata <= X"5180E0E4";
    when 16#0030A# => romdata <= X"3F72892A";
    when 16#0030B# => romdata <= X"70810651";
    when 16#0030C# => romdata <= X"5271802E";
    when 16#0030D# => romdata <= X"FCC838D1";
    when 16#0030E# => romdata <= X"3981ABEC";
    when 16#0030F# => romdata <= X"5180E0CC";
    when 16#00310# => romdata <= X"3F72882A";
    when 16#00311# => romdata <= X"70810651";
    when 16#00312# => romdata <= X"5271802E";
    when 16#00313# => romdata <= X"FCA438D1";
    when 16#00314# => romdata <= X"3981AC94";
    when 16#00315# => romdata <= X"5180E0B4";
    when 16#00316# => romdata <= X"3F72872A";
    when 16#00317# => romdata <= X"70810651";
    when 16#00318# => romdata <= X"5271802E";
    when 16#00319# => romdata <= X"FC8038D1";
    when 16#0031A# => romdata <= X"3981ACB4";
    when 16#0031B# => romdata <= X"5180E09C";
    when 16#0031C# => romdata <= X"3F72862A";
    when 16#0031D# => romdata <= X"70810651";
    when 16#0031E# => romdata <= X"5271802E";
    when 16#0031F# => romdata <= X"FBDC38D1";
    when 16#00320# => romdata <= X"3981ACD4";
    when 16#00321# => romdata <= X"5180E084";
    when 16#00322# => romdata <= X"3F72852A";
    when 16#00323# => romdata <= X"70810651";
    when 16#00324# => romdata <= X"5271802E";
    when 16#00325# => romdata <= X"FBB838D1";
    when 16#00326# => romdata <= X"3981ACFC";
    when 16#00327# => romdata <= X"5180DFEC";
    when 16#00328# => romdata <= X"3F72842A";
    when 16#00329# => romdata <= X"70810651";
    when 16#0032A# => romdata <= X"5271802E";
    when 16#0032B# => romdata <= X"FB9438D1";
    when 16#0032C# => romdata <= X"3981AD9C";
    when 16#0032D# => romdata <= X"5180DFD4";
    when 16#0032E# => romdata <= X"3F72832A";
    when 16#0032F# => romdata <= X"70810651";
    when 16#00330# => romdata <= X"5271802E";
    when 16#00331# => romdata <= X"FAF038D1";
    when 16#00332# => romdata <= X"3981ADBC";
    when 16#00333# => romdata <= X"5180DFBC";
    when 16#00334# => romdata <= X"3F72822A";
    when 16#00335# => romdata <= X"70810651";
    when 16#00336# => romdata <= X"5271802E";
    when 16#00337# => romdata <= X"FACC38D1";
    when 16#00338# => romdata <= X"3981ADE4";
    when 16#00339# => romdata <= X"5180DFA4";
    when 16#0033A# => romdata <= X"3F72812A";
    when 16#0033B# => romdata <= X"70810651";
    when 16#0033C# => romdata <= X"5271802E";
    when 16#0033D# => romdata <= X"FAA838D1";
    when 16#0033E# => romdata <= X"3981AE84";
    when 16#0033F# => romdata <= X"5180DF8C";
    when 16#00340# => romdata <= X"3F843D0D";
    when 16#00341# => romdata <= X"04FD3D0D";
    when 16#00342# => romdata <= X"81AE9851";
    when 16#00343# => romdata <= X"80DEFD3F";
    when 16#00344# => romdata <= X"81CEF408";
    when 16#00345# => romdata <= X"7008709E";
    when 16#00346# => romdata <= X"2A708106";
    when 16#00347# => romdata <= X"51525553";
    when 16#00348# => romdata <= X"81547283";
    when 16#00349# => romdata <= X"38725473";
    when 16#0034A# => romdata <= X"802E88C4";
    when 16#0034B# => romdata <= X"3881AEB4";
    when 16#0034C# => romdata <= X"5180DED8";
    when 16#0034D# => romdata <= X"3F81AEBC";
    when 16#0034E# => romdata <= X"5180DED0";
    when 16#0034F# => romdata <= X"3F81CEF4";
    when 16#00350# => romdata <= X"08841108";
    when 16#00351# => romdata <= X"709D2A81";
    when 16#00352# => romdata <= X"06515553";
    when 16#00353# => romdata <= X"73802E87";
    when 16#00354# => romdata <= X"B03881AE";
    when 16#00355# => romdata <= X"D85180DE";
    when 16#00356# => romdata <= X"B33F81AE";
    when 16#00357# => romdata <= X"E45180DE";
    when 16#00358# => romdata <= X"AB3F81CE";
    when 16#00359# => romdata <= X"BC0880D4";
    when 16#0035A# => romdata <= X"11085254";
    when 16#0035B# => romdata <= X"80DFE73F";
    when 16#0035C# => romdata <= X"81AF8051";
    when 16#0035D# => romdata <= X"80DE953F";
    when 16#0035E# => romdata <= X"81CEBC08";
    when 16#0035F# => romdata <= X"80D01108";
    when 16#00360# => romdata <= X"525380DF";
    when 16#00361# => romdata <= X"D13F8A51";
    when 16#00362# => romdata <= X"80DDE73F";
    when 16#00363# => romdata <= X"81AF9C51";
    when 16#00364# => romdata <= X"80DDF93F";
    when 16#00365# => romdata <= X"81AFC051";
    when 16#00366# => romdata <= X"80DDF13F";
    when 16#00367# => romdata <= X"81B08851";
    when 16#00368# => romdata <= X"80DDE93F";
    when 16#00369# => romdata <= X"81B0D051";
    when 16#0036A# => romdata <= X"80DDE13F";
    when 16#0036B# => romdata <= X"81CEBC08";
    when 16#0036C# => romdata <= X"70085254";
    when 16#0036D# => romdata <= X"80DF9F3F";
    when 16#0036E# => romdata <= X"B00881FF";
    when 16#0036F# => romdata <= X"0653728C";
    when 16#00370# => romdata <= X"279438A0";
    when 16#00371# => romdata <= X"5180DDAA";
    when 16#00372# => romdata <= X"3F811370";
    when 16#00373# => romdata <= X"81FF0651";
    when 16#00374# => romdata <= X"538C7326";
    when 16#00375# => romdata <= X"EE3881CE";
    when 16#00376# => romdata <= X"BC088411";
    when 16#00377# => romdata <= X"08525480";
    when 16#00378# => romdata <= X"DEF43FB0";
    when 16#00379# => romdata <= X"0881FF06";
    when 16#0037A# => romdata <= X"53728C27";
    when 16#0037B# => romdata <= X"9438A051";
    when 16#0037C# => romdata <= X"80DCFF3F";
    when 16#0037D# => romdata <= X"81137081";
    when 16#0037E# => romdata <= X"FF065153";
    when 16#0037F# => romdata <= X"8C7326EE";
    when 16#00380# => romdata <= X"3881CEBC";
    when 16#00381# => romdata <= X"08881108";
    when 16#00382# => romdata <= X"525480DE";
    when 16#00383# => romdata <= X"C93FB008";
    when 16#00384# => romdata <= X"81FF0653";
    when 16#00385# => romdata <= X"728C2794";
    when 16#00386# => romdata <= X"38A05180";
    when 16#00387# => romdata <= X"DCD43F81";
    when 16#00388# => romdata <= X"137081FF";
    when 16#00389# => romdata <= X"0651538C";
    when 16#0038A# => romdata <= X"7326EE38";
    when 16#0038B# => romdata <= X"81CEBC08";
    when 16#0038C# => romdata <= X"8C110852";
    when 16#0038D# => romdata <= X"5480DE9E";
    when 16#0038E# => romdata <= X"3FB00881";
    when 16#0038F# => romdata <= X"FF065372";
    when 16#00390# => romdata <= X"8C279438";
    when 16#00391# => romdata <= X"A05180DC";
    when 16#00392# => romdata <= X"A93F8113";
    when 16#00393# => romdata <= X"7081FF06";
    when 16#00394# => romdata <= X"51538C73";
    when 16#00395# => romdata <= X"26EE3881";
    when 16#00396# => romdata <= X"B0EC5180";
    when 16#00397# => romdata <= X"DCAE3F81";
    when 16#00398# => romdata <= X"CEBC0890";
    when 16#00399# => romdata <= X"11085254";
    when 16#0039A# => romdata <= X"80DDEB3F";
    when 16#0039B# => romdata <= X"B00881FF";
    when 16#0039C# => romdata <= X"0653728C";
    when 16#0039D# => romdata <= X"279438A0";
    when 16#0039E# => romdata <= X"5180DBF6";
    when 16#0039F# => romdata <= X"3F811370";
    when 16#003A0# => romdata <= X"81FF0651";
    when 16#003A1# => romdata <= X"538C7326";
    when 16#003A2# => romdata <= X"EE3881CE";
    when 16#003A3# => romdata <= X"BC089411";
    when 16#003A4# => romdata <= X"08525480";
    when 16#003A5# => romdata <= X"DDC03FB0";
    when 16#003A6# => romdata <= X"0881FF06";
    when 16#003A7# => romdata <= X"53728C27";
    when 16#003A8# => romdata <= X"9438A051";
    when 16#003A9# => romdata <= X"80DBCB3F";
    when 16#003AA# => romdata <= X"81137081";
    when 16#003AB# => romdata <= X"FF065153";
    when 16#003AC# => romdata <= X"8C7326EE";
    when 16#003AD# => romdata <= X"3881CEBC";
    when 16#003AE# => romdata <= X"08981108";
    when 16#003AF# => romdata <= X"525480DD";
    when 16#003B0# => romdata <= X"953FB008";
    when 16#003B1# => romdata <= X"81FF0653";
    when 16#003B2# => romdata <= X"728C2794";
    when 16#003B3# => romdata <= X"38A05180";
    when 16#003B4# => romdata <= X"DBA03F81";
    when 16#003B5# => romdata <= X"137081FF";
    when 16#003B6# => romdata <= X"0651538C";
    when 16#003B7# => romdata <= X"7326EE38";
    when 16#003B8# => romdata <= X"81CEBC08";
    when 16#003B9# => romdata <= X"9C110852";
    when 16#003BA# => romdata <= X"5480DCEA";
    when 16#003BB# => romdata <= X"3FB00881";
    when 16#003BC# => romdata <= X"FF065372";
    when 16#003BD# => romdata <= X"8C279438";
    when 16#003BE# => romdata <= X"A05180DA";
    when 16#003BF# => romdata <= X"F53F8113";
    when 16#003C0# => romdata <= X"7081FF06";
    when 16#003C1# => romdata <= X"51538C73";
    when 16#003C2# => romdata <= X"26EE3881";
    when 16#003C3# => romdata <= X"B1885180";
    when 16#003C4# => romdata <= X"DAFA3F81";
    when 16#003C5# => romdata <= X"CEBC0854";
    when 16#003C6# => romdata <= X"810BB015";
    when 16#003C7# => romdata <= X"0CB01408";
    when 16#003C8# => romdata <= X"53728025";
    when 16#003C9# => romdata <= X"F838A014";
    when 16#003CA# => romdata <= X"085180DC";
    when 16#003CB# => romdata <= X"A93FB008";
    when 16#003CC# => romdata <= X"81FF0653";
    when 16#003CD# => romdata <= X"728C2794";
    when 16#003CE# => romdata <= X"38A05180";
    when 16#003CF# => romdata <= X"DAB43F81";
    when 16#003D0# => romdata <= X"137081FF";
    when 16#003D1# => romdata <= X"0654548C";
    when 16#003D2# => romdata <= X"7326EE38";
    when 16#003D3# => romdata <= X"81CEBC08";
    when 16#003D4# => romdata <= X"A4110852";
    when 16#003D5# => romdata <= X"5380DBFE";
    when 16#003D6# => romdata <= X"3FB00881";
    when 16#003D7# => romdata <= X"FF065372";
    when 16#003D8# => romdata <= X"8C279438";
    when 16#003D9# => romdata <= X"A05180DA";
    when 16#003DA# => romdata <= X"893F8113";
    when 16#003DB# => romdata <= X"7081FF06";
    when 16#003DC# => romdata <= X"54548C73";
    when 16#003DD# => romdata <= X"26EE3881";
    when 16#003DE# => romdata <= X"CEBC08A8";
    when 16#003DF# => romdata <= X"11085253";
    when 16#003E0# => romdata <= X"80DBD33F";
    when 16#003E1# => romdata <= X"B00881FF";
    when 16#003E2# => romdata <= X"0653728C";
    when 16#003E3# => romdata <= X"279438A0";
    when 16#003E4# => romdata <= X"5180D9DE";
    when 16#003E5# => romdata <= X"3F811370";
    when 16#003E6# => romdata <= X"81FF0654";
    when 16#003E7# => romdata <= X"548C7326";
    when 16#003E8# => romdata <= X"EE3881CE";
    when 16#003E9# => romdata <= X"BC08AC11";
    when 16#003EA# => romdata <= X"08525380";
    when 16#003EB# => romdata <= X"DBA83FB0";
    when 16#003EC# => romdata <= X"0881FF06";
    when 16#003ED# => romdata <= X"53728C27";
    when 16#003EE# => romdata <= X"9438A051";
    when 16#003EF# => romdata <= X"80D9B33F";
    when 16#003F0# => romdata <= X"81137081";
    when 16#003F1# => romdata <= X"FF065454";
    when 16#003F2# => romdata <= X"8C7326EE";
    when 16#003F3# => romdata <= X"3881B1A4";
    when 16#003F4# => romdata <= X"5180D9B8";
    when 16#003F5# => romdata <= X"3F81CEBC";
    when 16#003F6# => romdata <= X"0880E011";
    when 16#003F7# => romdata <= X"08525380";
    when 16#003F8# => romdata <= X"DAF43F81";
    when 16#003F9# => romdata <= X"B1B85180";
    when 16#003FA# => romdata <= X"D9A23F81";
    when 16#003FB# => romdata <= X"CEBC08B0";
    when 16#003FC# => romdata <= X"1108FE0A";
    when 16#003FD# => romdata <= X"06525480";
    when 16#003FE# => romdata <= X"DADC3F81";
    when 16#003FF# => romdata <= X"CEBC0854";
    when 16#00400# => romdata <= X"800BB015";
    when 16#00401# => romdata <= X"0C81B1CC";
    when 16#00402# => romdata <= X"5180D980";
    when 16#00403# => romdata <= X"3F81B1E4";
    when 16#00404# => romdata <= X"5180D8F8";
    when 16#00405# => romdata <= X"3F81CEBC";
    when 16#00406# => romdata <= X"0880C011";
    when 16#00407# => romdata <= X"08525380";
    when 16#00408# => romdata <= X"DAB43FB0";
    when 16#00409# => romdata <= X"0881FF06";
    when 16#0040A# => romdata <= X"53729827";
    when 16#0040B# => romdata <= X"9438A051";
    when 16#0040C# => romdata <= X"80D8BF3F";
    when 16#0040D# => romdata <= X"81137081";
    when 16#0040E# => romdata <= X"FF065454";
    when 16#0040F# => romdata <= X"987326EE";
    when 16#00410# => romdata <= X"3881CEBC";
    when 16#00411# => romdata <= X"0880C811";
    when 16#00412# => romdata <= X"08525380";
    when 16#00413# => romdata <= X"DA883FB0";
    when 16#00414# => romdata <= X"0881FF06";
    when 16#00415# => romdata <= X"53729827";
    when 16#00416# => romdata <= X"9438A051";
    when 16#00417# => romdata <= X"80D8933F";
    when 16#00418# => romdata <= X"81137081";
    when 16#00419# => romdata <= X"FF065454";
    when 16#0041A# => romdata <= X"987326EE";
    when 16#0041B# => romdata <= X"3881B280";
    when 16#0041C# => romdata <= X"5180D898";
    when 16#0041D# => romdata <= X"3F81CEBC";
    when 16#0041E# => romdata <= X"0880C411";
    when 16#0041F# => romdata <= X"08525380";
    when 16#00420# => romdata <= X"D9D43FB0";
    when 16#00421# => romdata <= X"0881FF06";
    when 16#00422# => romdata <= X"53729827";
    when 16#00423# => romdata <= X"9438A051";
    when 16#00424# => romdata <= X"80D7DF3F";
    when 16#00425# => romdata <= X"81137081";
    when 16#00426# => romdata <= X"FF065454";
    when 16#00427# => romdata <= X"987326EE";
    when 16#00428# => romdata <= X"3881CEBC";
    when 16#00429# => romdata <= X"0880CC11";
    when 16#0042A# => romdata <= X"08525380";
    when 16#0042B# => romdata <= X"D9A83FB0";
    when 16#0042C# => romdata <= X"0881FF06";
    when 16#0042D# => romdata <= X"53729827";
    when 16#0042E# => romdata <= X"9438A051";
    when 16#0042F# => romdata <= X"80D7B33F";
    when 16#00430# => romdata <= X"81137081";
    when 16#00431# => romdata <= X"FF065454";
    when 16#00432# => romdata <= X"987326EE";
    when 16#00433# => romdata <= X"388A5180";
    when 16#00434# => romdata <= X"D7A03F81";
    when 16#00435# => romdata <= X"CEBC08B4";
    when 16#00436# => romdata <= X"110881B2";
    when 16#00437# => romdata <= X"9C535153";
    when 16#00438# => romdata <= X"80D7A93F";
    when 16#00439# => romdata <= X"725180D8";
    when 16#0043A# => romdata <= X"ED3FA051";
    when 16#0043B# => romdata <= X"80D7833F";
    when 16#0043C# => romdata <= X"72862681";
    when 16#0043D# => romdata <= X"8E387210";
    when 16#0043E# => romdata <= X"1081BEC0";
    when 16#0043F# => romdata <= X"05547308";
    when 16#00440# => romdata <= X"0481B2B0";
    when 16#00441# => romdata <= X"5180D784";
    when 16#00442# => romdata <= X"3F81AEE4";
    when 16#00443# => romdata <= X"5180D6FC";
    when 16#00444# => romdata <= X"3F81CEBC";
    when 16#00445# => romdata <= X"0880D411";
    when 16#00446# => romdata <= X"08525480";
    when 16#00447# => romdata <= X"D8B83F81";
    when 16#00448# => romdata <= X"AF805180";
    when 16#00449# => romdata <= X"D6E63F81";
    when 16#0044A# => romdata <= X"CEBC0880";
    when 16#0044B# => romdata <= X"D0110852";
    when 16#0044C# => romdata <= X"5380D8A2";
    when 16#0044D# => romdata <= X"3F8A5180";
    when 16#0044E# => romdata <= X"D6B83F81";
    when 16#0044F# => romdata <= X"AF9C5180";
    when 16#00450# => romdata <= X"D6CA3F81";
    when 16#00451# => romdata <= X"AFC05180";
    when 16#00452# => romdata <= X"D6C23F81";
    when 16#00453# => romdata <= X"B0885180";
    when 16#00454# => romdata <= X"D6BA3F81";
    when 16#00455# => romdata <= X"B0D05180";
    when 16#00456# => romdata <= X"D6B23F81";
    when 16#00457# => romdata <= X"CEBC0870";
    when 16#00458# => romdata <= X"08525480";
    when 16#00459# => romdata <= X"D7F03FB0";
    when 16#0045A# => romdata <= X"0881FF06";
    when 16#0045B# => romdata <= X"53F8CF39";
    when 16#0045C# => romdata <= X"81B2B851";
    when 16#0045D# => romdata <= X"80D6953F";
    when 16#0045E# => romdata <= X"F7B33981";
    when 16#0045F# => romdata <= X"B2C05180";
    when 16#00460# => romdata <= X"D68A3F81";
    when 16#00461# => romdata <= X"CEBC08B8";
    when 16#00462# => romdata <= X"110881B2";
    when 16#00463# => romdata <= X"CC535454";
    when 16#00464# => romdata <= X"80D5F93F";
    when 16#00465# => romdata <= X"7252A051";
    when 16#00466# => romdata <= X"80D6943F";
    when 16#00467# => romdata <= X"7251F0E5";
    when 16#00468# => romdata <= X"3F8A5180";
    when 16#00469# => romdata <= X"D5CC3F80";
    when 16#0046A# => romdata <= X"0BB00C85";
    when 16#0046B# => romdata <= X"3D0D0481";
    when 16#0046C# => romdata <= X"B2E05180";
    when 16#0046D# => romdata <= X"D5D63FCB";
    when 16#0046E# => romdata <= X"3981B2EC";
    when 16#0046F# => romdata <= X"5180D5CC";
    when 16#00470# => romdata <= X"3FC13981";
    when 16#00471# => romdata <= X"B2F85180";
    when 16#00472# => romdata <= X"D5C23FFF";
    when 16#00473# => romdata <= X"B63981B2";
    when 16#00474# => romdata <= X"FC5180D5";
    when 16#00475# => romdata <= X"B73FFFAB";
    when 16#00476# => romdata <= X"3981B388";
    when 16#00477# => romdata <= X"5180D5AC";
    when 16#00478# => romdata <= X"3FFFA039";
    when 16#00479# => romdata <= X"81B39451";
    when 16#0047A# => romdata <= X"80D5A13F";
    when 16#0047B# => romdata <= X"FF9539FE";
    when 16#0047C# => romdata <= X"3D0D8151";
    when 16#0047D# => romdata <= X"AAEC3FB0";
    when 16#0047E# => romdata <= X"0881FF06";
    when 16#0047F# => romdata <= X"81CEBC08";
    when 16#00480# => romdata <= X"71B4120C";
    when 16#00481# => romdata <= X"53B00C84";
    when 16#00482# => romdata <= X"3D0D04FE";
    when 16#00483# => romdata <= X"3D0D880A";
    when 16#00484# => romdata <= X"53840A0B";
    when 16#00485# => romdata <= X"81CEB808";
    when 16#00486# => romdata <= X"8C110851";
    when 16#00487# => romdata <= X"52528071";
    when 16#00488# => romdata <= X"27953880";
    when 16#00489# => romdata <= X"73708405";
    when 16#0048A# => romdata <= X"550C8072";
    when 16#0048B# => romdata <= X"70840554";
    when 16#0048C# => romdata <= X"0CFF1151";
    when 16#0048D# => romdata <= X"70ED3880";
    when 16#0048E# => romdata <= X"0BB00C84";
    when 16#0048F# => romdata <= X"3D0D04FA";
    when 16#00490# => romdata <= X"3D0D880A";
    when 16#00491# => romdata <= X"57840A56";
    when 16#00492# => romdata <= X"8151AA96";
    when 16#00493# => romdata <= X"3FB00883";
    when 16#00494# => romdata <= X"FFFF0654";
    when 16#00495# => romdata <= X"73833890";
    when 16#00496# => romdata <= X"54805574";
    when 16#00497# => romdata <= X"742781C2";
    when 16#00498# => romdata <= X"38750870";
    when 16#00499# => romdata <= X"902C5253";
    when 16#0049A# => romdata <= X"80D5EB3F";
    when 16#0049B# => romdata <= X"B00881FF";
    when 16#0049C# => romdata <= X"0652718A";
    when 16#0049D# => romdata <= X"279438A0";
    when 16#0049E# => romdata <= X"5180D3F6";
    when 16#0049F# => romdata <= X"3F811270";
    when 16#004A0# => romdata <= X"81FF0651";
    when 16#004A1# => romdata <= X"528A7226";
    when 16#004A2# => romdata <= X"EE387290";
    when 16#004A3# => romdata <= X"2B70902C";
    when 16#004A4# => romdata <= X"525280D5";
    when 16#004A5# => romdata <= X"C13FB008";
    when 16#004A6# => romdata <= X"81FF0652";
    when 16#004A7# => romdata <= X"718A2794";
    when 16#004A8# => romdata <= X"38A05180";
    when 16#004A9# => romdata <= X"D3CC3F81";
    when 16#004AA# => romdata <= X"127081FF";
    when 16#004AB# => romdata <= X"0653538A";
    when 16#004AC# => romdata <= X"7226EE38";
    when 16#004AD# => romdata <= X"76087090";
    when 16#004AE# => romdata <= X"2C525380";
    when 16#004AF# => romdata <= X"D5983FB0";
    when 16#004B0# => romdata <= X"0881FF06";
    when 16#004B1# => romdata <= X"52718A27";
    when 16#004B2# => romdata <= X"9438A051";
    when 16#004B3# => romdata <= X"80D3A33F";
    when 16#004B4# => romdata <= X"81127081";
    when 16#004B5# => romdata <= X"FF065152";
    when 16#004B6# => romdata <= X"8A7226EE";
    when 16#004B7# => romdata <= X"3872902B";
    when 16#004B8# => romdata <= X"70902C52";
    when 16#004B9# => romdata <= X"5280D4EE";
    when 16#004BA# => romdata <= X"3FB00881";
    when 16#004BB# => romdata <= X"FF065271";
    when 16#004BC# => romdata <= X"8A279438";
    when 16#004BD# => romdata <= X"A05180D2";
    when 16#004BE# => romdata <= X"F93F8112";
    when 16#004BF# => romdata <= X"7081FF06";
    when 16#004C0# => romdata <= X"53538A72";
    when 16#004C1# => romdata <= X"26EE388A";
    when 16#004C2# => romdata <= X"5180D2E6";
    when 16#004C3# => romdata <= X"3F841784";
    when 16#004C4# => romdata <= X"17811770";
    when 16#004C5# => romdata <= X"83FFFF06";
    when 16#004C6# => romdata <= X"58545757";
    when 16#004C7# => romdata <= X"737526FE";
    when 16#004C8# => romdata <= X"C03873B0";
    when 16#004C9# => romdata <= X"0C883D0D";
    when 16#004CA# => romdata <= X"04FD3D0D";
    when 16#004CB# => romdata <= X"8151A8B2";
    when 16#004CC# => romdata <= X"3FB00881";
    when 16#004CD# => romdata <= X"FF065473";
    when 16#004CE# => romdata <= X"802EA438";
    when 16#004CF# => romdata <= X"73842690";
    when 16#004D0# => romdata <= X"3881CEB8";
    when 16#004D1# => romdata <= X"0874710C";
    when 16#004D2# => romdata <= X"5373B00C";
    when 16#004D3# => romdata <= X"853D0D04";
    when 16#004D4# => romdata <= X"81CEB808";
    when 16#004D5# => romdata <= X"5380730C";
    when 16#004D6# => romdata <= X"73B00C85";
    when 16#004D7# => romdata <= X"3D0D0481";
    when 16#004D8# => romdata <= X"B4A05180";
    when 16#004D9# => romdata <= X"D2A63F81";
    when 16#004DA# => romdata <= X"B4B05180";
    when 16#004DB# => romdata <= X"D29E3F81";
    when 16#004DC# => romdata <= X"CEB80870";
    when 16#004DD# => romdata <= X"08525380";
    when 16#004DE# => romdata <= X"D3DC3F81";
    when 16#004DF# => romdata <= X"B4C05180";
    when 16#004E0# => romdata <= X"D28A3F81";
    when 16#004E1# => romdata <= X"CEB80884";
    when 16#004E2# => romdata <= X"11085353";
    when 16#004E3# => romdata <= X"A05180D2";
    when 16#004E4# => romdata <= X"9E3F81B4";
    when 16#004E5# => romdata <= X"D45180D1";
    when 16#004E6# => romdata <= X"F33F81CE";
    when 16#004E7# => romdata <= X"B8088811";
    when 16#004E8# => romdata <= X"085353A0";
    when 16#004E9# => romdata <= X"5180D287";
    when 16#004EA# => romdata <= X"3F81B4E8";
    when 16#004EB# => romdata <= X"5180D1DC";
    when 16#004EC# => romdata <= X"3F81CEB8";
    when 16#004ED# => romdata <= X"088C1108";
    when 16#004EE# => romdata <= X"525380D3";
    when 16#004EF# => romdata <= X"993F8A51";
    when 16#004F0# => romdata <= X"80D1AF3F";
    when 16#004F1# => romdata <= X"73B00C85";
    when 16#004F2# => romdata <= X"3D0D04BC";
    when 16#004F3# => romdata <= X"0802BC0C";
    when 16#004F4# => romdata <= X"F93D0D02";
    when 16#004F5# => romdata <= X"BC08FC05";
    when 16#004F6# => romdata <= X"0C880A0B";
    when 16#004F7# => romdata <= X"BC08F405";
    when 16#004F8# => romdata <= X"0CFC3D0D";
    when 16#004F9# => romdata <= X"823DBC08";
    when 16#004FA# => romdata <= X"F0050C81";
    when 16#004FB# => romdata <= X"51A6F33F";
    when 16#004FC# => romdata <= X"B00881FF";
    when 16#004FD# => romdata <= X"06BC08F8";
    when 16#004FE# => romdata <= X"050C8251";
    when 16#004FF# => romdata <= X"A6E43FB0";
    when 16#00500# => romdata <= X"08BC08F0";
    when 16#00501# => romdata <= X"05082383";
    when 16#00502# => romdata <= X"51A6D73F";
    when 16#00503# => romdata <= X"B008BC08";
    when 16#00504# => romdata <= X"F0050882";
    when 16#00505# => romdata <= X"05238451";
    when 16#00506# => romdata <= X"A6C83FB0";
    when 16#00507# => romdata <= X"08BC08F0";
    when 16#00508# => romdata <= X"05088405";
    when 16#00509# => romdata <= X"238551A6";
    when 16#0050A# => romdata <= X"B93FB008";
    when 16#0050B# => romdata <= X"BC08F005";
    when 16#0050C# => romdata <= X"08860523";
    when 16#0050D# => romdata <= X"8651A6AA";
    when 16#0050E# => romdata <= X"3FB008BC";
    when 16#0050F# => romdata <= X"08F00508";
    when 16#00510# => romdata <= X"88052387";
    when 16#00511# => romdata <= X"51A69B3F";
    when 16#00512# => romdata <= X"B008BC08";
    when 16#00513# => romdata <= X"F005088A";
    when 16#00514# => romdata <= X"05238851";
    when 16#00515# => romdata <= X"A68C3FB0";
    when 16#00516# => romdata <= X"08BC08F0";
    when 16#00517# => romdata <= X"05088C05";
    when 16#00518# => romdata <= X"238951A5";
    when 16#00519# => romdata <= X"FD3FB008";
    when 16#0051A# => romdata <= X"BC08F005";
    when 16#0051B# => romdata <= X"088E0523";
    when 16#0051C# => romdata <= X"800B81CE";
    when 16#0051D# => romdata <= X"B808708C";
    when 16#0051E# => romdata <= X"050851BC";
    when 16#0051F# => romdata <= X"08E4050C";
    when 16#00520# => romdata <= X"BC08EC05";
    when 16#00521# => romdata <= X"0CBC08EC";
    when 16#00522# => romdata <= X"0508BC08";
    when 16#00523# => romdata <= X"E4050827";
    when 16#00524# => romdata <= X"818F38BC";
    when 16#00525# => romdata <= X"08E40508";
    when 16#00526# => romdata <= X"BC08E805";
    when 16#00527# => romdata <= X"0CBC08F8";
    when 16#00528# => romdata <= X"0508802E";
    when 16#00529# => romdata <= X"81B638BC";
    when 16#0052A# => romdata <= X"08EC0508";
    when 16#0052B# => romdata <= X"10BC08F0";
    when 16#0052C# => romdata <= X"05080570";
    when 16#0052D# => romdata <= X"22BC08F4";
    when 16#0052E# => romdata <= X"05088205";
    when 16#0052F# => romdata <= X"2271902B";
    when 16#00530# => romdata <= X"07BC08F4";
    when 16#00531# => romdata <= X"05080CBC";
    when 16#00532# => romdata <= X"08E4050C";
    when 16#00533# => romdata <= X"BC08F805";
    when 16#00534# => romdata <= X"0CBC08EC";
    when 16#00535# => romdata <= X"05088105";
    when 16#00536# => romdata <= X"7081FF06";
    when 16#00537# => romdata <= X"BC08E405";
    when 16#00538# => romdata <= X"0CBC08F8";
    when 16#00539# => romdata <= X"050C860B";
    when 16#0053A# => romdata <= X"BC08EC05";
    when 16#0053B# => romdata <= X"08278838";
    when 16#0053C# => romdata <= X"800BBC08";
    when 16#0053D# => romdata <= X"E4050CBC";
    when 16#0053E# => romdata <= X"08E40508";
    when 16#0053F# => romdata <= X"BC08F405";
    when 16#00540# => romdata <= X"088405BC";
    when 16#00541# => romdata <= X"08E80508";
    when 16#00542# => romdata <= X"FF05BC08";
    when 16#00543# => romdata <= X"E8050CBC";
    when 16#00544# => romdata <= X"08F4050C";
    when 16#00545# => romdata <= X"BC08EC05";
    when 16#00546# => romdata <= X"0CBC08E8";
    when 16#00547# => romdata <= X"0508FF87";
    when 16#00548# => romdata <= X"38BC08FC";
    when 16#00549# => romdata <= X"05080D80";
    when 16#0054A# => romdata <= X"0BB00C89";
    when 16#0054B# => romdata <= X"3D0DBC0C";
    when 16#0054C# => romdata <= X"04BC08E4";
    when 16#0054D# => romdata <= X"0508BC08";
    when 16#0054E# => romdata <= X"F4050884";
    when 16#0054F# => romdata <= X"05BC08E8";
    when 16#00550# => romdata <= X"0508FF05";
    when 16#00551# => romdata <= X"BC08E805";
    when 16#00552# => romdata <= X"0CBC08F4";
    when 16#00553# => romdata <= X"050CBC08";
    when 16#00554# => romdata <= X"EC050CBC";
    when 16#00555# => romdata <= X"08E80508";
    when 16#00556# => romdata <= X"802EC638";
    when 16#00557# => romdata <= X"BC08EC05";
    when 16#00558# => romdata <= X"0810BC08";
    when 16#00559# => romdata <= X"F0050805";
    when 16#0055A# => romdata <= X"70227090";
    when 16#0055B# => romdata <= X"2BBC08F4";
    when 16#0055C# => romdata <= X"050808FC";
    when 16#0055D# => romdata <= X"80800671";
    when 16#0055E# => romdata <= X"902C07BC";
    when 16#0055F# => romdata <= X"08F40508";
    when 16#00560# => romdata <= X"0C52BC08";
    when 16#00561# => romdata <= X"E4050CBC";
    when 16#00562# => romdata <= X"08F8050C";
    when 16#00563# => romdata <= X"800BBC08";
    when 16#00564# => romdata <= X"E4050CBC";
    when 16#00565# => romdata <= X"08EC0508";
    when 16#00566# => romdata <= X"8626FF95";
    when 16#00567# => romdata <= X"38BC08EC";
    when 16#00568# => romdata <= X"05088105";
    when 16#00569# => romdata <= X"7081FF06";
    when 16#0056A# => romdata <= X"BC08F405";
    when 16#0056B# => romdata <= X"088405BC";
    when 16#0056C# => romdata <= X"08E80508";
    when 16#0056D# => romdata <= X"FF05BC08";
    when 16#0056E# => romdata <= X"E8050CBC";
    when 16#0056F# => romdata <= X"08F4050C";
    when 16#00570# => romdata <= X"BC08EC05";
    when 16#00571# => romdata <= X"0CBC08E4";
    when 16#00572# => romdata <= X"050CBC08";
    when 16#00573# => romdata <= X"E80508FF";
    when 16#00574# => romdata <= X"8B38FECD";
    when 16#00575# => romdata <= X"39FB3D0D";
    when 16#00576# => romdata <= X"029F0533";
    when 16#00577# => romdata <= X"79982B70";
    when 16#00578# => romdata <= X"982C5154";
    when 16#00579# => romdata <= X"55810A54";
    when 16#0057A# => romdata <= X"805672E8";
    when 16#0057B# => romdata <= X"25BD38E8";
    when 16#0057C# => romdata <= X"53751081";
    when 16#0057D# => romdata <= X"07738180";
    when 16#0057E# => romdata <= X"0A298180";
    when 16#0057F# => romdata <= X"0A057098";
    when 16#00580# => romdata <= X"2C515456";
    when 16#00581# => romdata <= X"807324E9";
    when 16#00582# => romdata <= X"38807325";
    when 16#00583# => romdata <= X"80C73873";
    when 16#00584# => romdata <= X"812A810A";
    when 16#00585# => romdata <= X"07738180";
    when 16#00586# => romdata <= X"0A2981FF";
    when 16#00587# => romdata <= X"0A057098";
    when 16#00588# => romdata <= X"2C515454";
    when 16#00589# => romdata <= X"728024E7";
    when 16#0058A# => romdata <= X"38AB3997";
    when 16#0058B# => romdata <= X"73259A38";
    when 16#0058C# => romdata <= X"9774812A";
    when 16#0058D# => romdata <= X"810A0771";
    when 16#0058E# => romdata <= X"81800A29";
    when 16#0058F# => romdata <= X"81FF0A05";
    when 16#00590# => romdata <= X"70982C51";
    when 16#00591# => romdata <= X"525553DC";
    when 16#00592# => romdata <= X"39807324";
    when 16#00593# => romdata <= X"FFA33872";
    when 16#00594# => romdata <= X"8024FFBB";
    when 16#00595# => romdata <= X"38745280";
    when 16#00596# => romdata <= X"51B3AF3F";
    when 16#00597# => romdata <= X"7381FF06";
    when 16#00598# => romdata <= X"51B4AD3F";
    when 16#00599# => romdata <= X"74528151";
    when 16#0059A# => romdata <= X"B3A03F73";
    when 16#0059B# => romdata <= X"882A7081";
    when 16#0059C# => romdata <= X"FF065253";
    when 16#0059D# => romdata <= X"B49A3F74";
    when 16#0059E# => romdata <= X"528251B3";
    when 16#0059F# => romdata <= X"8D3F7390";
    when 16#005A0# => romdata <= X"2A7081FF";
    when 16#005A1# => romdata <= X"065253B4";
    when 16#005A2# => romdata <= X"873F7452";
    when 16#005A3# => romdata <= X"8351B2FA";
    when 16#005A4# => romdata <= X"3F73982A";
    when 16#005A5# => romdata <= X"51B3F93F";
    when 16#005A6# => romdata <= X"74528451";
    when 16#005A7# => romdata <= X"B2EC3F75";
    when 16#005A8# => romdata <= X"81FF0651";
    when 16#005A9# => romdata <= X"B3EA3F74";
    when 16#005AA# => romdata <= X"528551B2";
    when 16#005AB# => romdata <= X"DD3F7588";
    when 16#005AC# => romdata <= X"2A7081FF";
    when 16#005AD# => romdata <= X"065253B3";
    when 16#005AE# => romdata <= X"D73F7452";
    when 16#005AF# => romdata <= X"8651B2CA";
    when 16#005B0# => romdata <= X"3F75902A";
    when 16#005B1# => romdata <= X"7081FF06";
    when 16#005B2# => romdata <= X"5254B3C4";
    when 16#005B3# => romdata <= X"3F745287";
    when 16#005B4# => romdata <= X"51B2B73F";
    when 16#005B5# => romdata <= X"75982A51";
    when 16#005B6# => romdata <= X"B3B63F87";
    when 16#005B7# => romdata <= X"3D0D04F2";
    when 16#005B8# => romdata <= X"3D0D0280";
    when 16#005B9# => romdata <= X"C3053302";
    when 16#005BA# => romdata <= X"840580C7";
    when 16#005BB# => romdata <= X"05338180";
    when 16#005BC# => romdata <= X"0A712B98";
    when 16#005BD# => romdata <= X"2A81CEB8";
    when 16#005BE# => romdata <= X"088C1108";
    when 16#005BF# => romdata <= X"71084453";
    when 16#005C0# => romdata <= X"565C5557";
    when 16#005C1# => romdata <= X"80730C80";
    when 16#005C2# => romdata <= X"7071725C";
    when 16#005C3# => romdata <= X"5A5E5B80";
    when 16#005C4# => romdata <= X"56757A27";
    when 16#005C5# => romdata <= X"80D73881";
    when 16#005C6# => romdata <= X"772783CE";
    when 16#005C7# => romdata <= X"387783FF";
    when 16#005C8# => romdata <= X"FF068119";
    when 16#005C9# => romdata <= X"71101084";
    when 16#005CA# => romdata <= X"0A057930";
    when 16#005CB# => romdata <= X"7A823270";
    when 16#005CC# => romdata <= X"30728025";
    when 16#005CD# => romdata <= X"71802507";
    when 16#005CE# => romdata <= X"56585841";
    when 16#005CF# => romdata <= X"57595C7B";
    when 16#005D0# => romdata <= X"802E83D5";
    when 16#005D1# => romdata <= X"38821522";
    when 16#005D2# => romdata <= X"5372902B";
    when 16#005D3# => romdata <= X"70902C54";
    when 16#005D4# => romdata <= X"55727B25";
    when 16#005D5# => romdata <= X"8338725B";
    when 16#005D6# => romdata <= X"7C732583";
    when 16#005D7# => romdata <= X"38725D81";
    when 16#005D8# => romdata <= X"167081FF";
    when 16#005D9# => romdata <= X"06575E79";
    when 16#005DA# => romdata <= X"7626FFB1";
    when 16#005DB# => romdata <= X"38811970";
    when 16#005DC# => romdata <= X"81FF065A";
    when 16#005DD# => romdata <= X"5680E579";
    when 16#005DE# => romdata <= X"27FF9438";
    when 16#005DF# => romdata <= X"987D3590";
    when 16#005E0# => romdata <= X"2B70902C";
    when 16#005E1# => romdata <= X"7C309871";
    when 16#005E2# => romdata <= X"35902B70";
    when 16#005E3# => romdata <= X"902C5C5C";
    when 16#005E4# => romdata <= X"55565477";
    when 16#005E5# => romdata <= X"54777525";
    when 16#005E6# => romdata <= X"83387454";
    when 16#005E7# => romdata <= X"73902B70";
    when 16#005E8# => romdata <= X"902C5D55";
    when 16#005E9# => romdata <= X"7B54807C";
    when 16#005EA# => romdata <= X"2583D738";
    when 16#005EB# => romdata <= X"73902B70";
    when 16#005EC# => romdata <= X"902C5F56";
    when 16#005ED# => romdata <= X"80705D58";
    when 16#005EE# => romdata <= X"80705A56";
    when 16#005EF# => romdata <= X"757A2780";
    when 16#005F0# => romdata <= X"E4388177";
    when 16#005F1# => romdata <= X"27838C38";
    when 16#005F2# => romdata <= X"7783FFFF";
    when 16#005F3# => romdata <= X"06811971";
    when 16#005F4# => romdata <= X"1010840A";
    when 16#005F5# => romdata <= X"0579307A";
    when 16#005F6# => romdata <= X"82327030";
    when 16#005F7# => romdata <= X"72802571";
    when 16#005F8# => romdata <= X"80250753";
    when 16#005F9# => romdata <= X"51575357";
    when 16#005FA# => romdata <= X"59547380";
    when 16#005FB# => romdata <= X"2E83A438";
    when 16#005FC# => romdata <= X"82152254";
    when 16#005FD# => romdata <= X"73902B70";
    when 16#005FE# => romdata <= X"902C719F";
    when 16#005FF# => romdata <= X"2C707232";
    when 16#00600# => romdata <= X"7131799F";
    when 16#00601# => romdata <= X"2C707B32";
    when 16#00602# => romdata <= X"71315154";
    when 16#00603# => romdata <= X"51565653";
    when 16#00604# => romdata <= X"72742583";
    when 16#00605# => romdata <= X"38745681";
    when 16#00606# => romdata <= X"197081FF";
    when 16#00607# => romdata <= X"065A5579";
    when 16#00608# => romdata <= X"7926FFA4";
    when 16#00609# => romdata <= X"387D7635";
    when 16#0060A# => romdata <= X"982B7098";
    when 16#0060B# => romdata <= X"2C53547B";
    when 16#0060C# => romdata <= X"51FBA23F";
    when 16#0060D# => romdata <= X"811C7081";
    when 16#0060E# => romdata <= X"FF065D59";
    when 16#0060F# => romdata <= X"80E57C27";
    when 16#00610# => romdata <= X"FEF63881";
    when 16#00611# => romdata <= X"CEB8087F";
    when 16#00612# => romdata <= X"710C5880";
    when 16#00613# => romdata <= X"5281C394";
    when 16#00614# => romdata <= X"51B3AD3F";
    when 16#00615# => romdata <= X"81F2D408";
    when 16#00616# => romdata <= X"80F5C40B";
    when 16#00617# => romdata <= X"81F2D40C";
    when 16#00618# => romdata <= X"5F805280";
    when 16#00619# => romdata <= X"51AFA33F";
    when 16#0061A# => romdata <= X"81B4F851";
    when 16#0061B# => romdata <= X"80C89D3F";
    when 16#0061C# => romdata <= X"7C5180C9";
    when 16#0061D# => romdata <= X"E13F8052";
    when 16#0061E# => romdata <= X"8751AF8E";
    when 16#0061F# => romdata <= X"3F81B580";
    when 16#00620# => romdata <= X"5180C888";
    when 16#00621# => romdata <= X"3F7A5180";
    when 16#00622# => romdata <= X"C9CC3F80";
    when 16#00623# => romdata <= X"D2528051";
    when 16#00624# => romdata <= X"AEF83F81";
    when 16#00625# => romdata <= X"B5885180";
    when 16#00626# => romdata <= X"C7F23F76";
    when 16#00627# => romdata <= X"5180C9B6";
    when 16#00628# => romdata <= X"3F80C052";
    when 16#00629# => romdata <= X"8751AEE2";
    when 16#0062A# => romdata <= X"3F81B590";
    when 16#0062B# => romdata <= X"5180C7DC";
    when 16#0062C# => romdata <= X"3F7980E6";
    when 16#0062D# => romdata <= X"295180C9";
    when 16#0062E# => romdata <= X"9D3F7E81";
    when 16#0062F# => romdata <= X"F2D40C90";
    when 16#00630# => romdata <= X"3D0D0474";
    when 16#00631# => romdata <= X"22537290";
    when 16#00632# => romdata <= X"2B70902C";
    when 16#00633# => romdata <= X"545C727B";
    when 16#00634# => romdata <= X"25833872";
    when 16#00635# => romdata <= X"5B7C7325";
    when 16#00636# => romdata <= X"8338725D";
    when 16#00637# => romdata <= X"81167081";
    when 16#00638# => romdata <= X"FF06575E";
    when 16#00639# => romdata <= X"757A27FD";
    when 16#0063A# => romdata <= X"84387783";
    when 16#0063B# => romdata <= X"FFFF0681";
    when 16#0063C# => romdata <= X"19711010";
    when 16#0063D# => romdata <= X"880A0579";
    when 16#0063E# => romdata <= X"307A8232";
    when 16#0063F# => romdata <= X"70307280";
    when 16#00640# => romdata <= X"25718025";
    when 16#00641# => romdata <= X"07565840";
    when 16#00642# => romdata <= X"41575954";
    when 16#00643# => romdata <= X"73802EFF";
    when 16#00644# => romdata <= X"B2388215";
    when 16#00645# => romdata <= X"2253FFAE";
    when 16#00646# => romdata <= X"39742253";
    when 16#00647# => romdata <= X"FCAB3974";
    when 16#00648# => romdata <= X"22547390";
    when 16#00649# => romdata <= X"2B70902C";
    when 16#0064A# => romdata <= X"719F2C70";
    when 16#0064B# => romdata <= X"72327131";
    when 16#0064C# => romdata <= X"799F2C70";
    when 16#0064D# => romdata <= X"7B327131";
    when 16#0064E# => romdata <= X"51545156";
    when 16#0064F# => romdata <= X"56537274";
    when 16#00650# => romdata <= X"25833874";
    when 16#00651# => romdata <= X"56811970";
    when 16#00652# => romdata <= X"81FF065A";
    when 16#00653# => romdata <= X"55787A27";
    when 16#00654# => romdata <= X"FDD33877";
    when 16#00655# => romdata <= X"83FFFF06";
    when 16#00656# => romdata <= X"81197110";
    when 16#00657# => romdata <= X"10880A05";
    when 16#00658# => romdata <= X"79307A82";
    when 16#00659# => romdata <= X"32703072";
    when 16#0065A# => romdata <= X"80257180";
    when 16#0065B# => romdata <= X"25075351";
    when 16#0065C# => romdata <= X"57535759";
    when 16#0065D# => romdata <= X"5473802E";
    when 16#0065E# => romdata <= X"FFA53882";
    when 16#0065F# => romdata <= X"152254FF";
    when 16#00660# => romdata <= X"A1398170";
    when 16#00661# => romdata <= X"902B7090";
    when 16#00662# => romdata <= X"2C405754";
    when 16#00663# => romdata <= X"80705D58";
    when 16#00664# => romdata <= X"FCA63974";
    when 16#00665# => romdata <= X"2254FCDC";
    when 16#00666# => romdata <= X"39FA3D0D";
    when 16#00667# => romdata <= X"8A5180C5";
    when 16#00668# => romdata <= X"D13F97B9";
    when 16#00669# => romdata <= X"3F9A8553";
    when 16#0066A# => romdata <= X"81B59852";
    when 16#0066B# => romdata <= X"81B5AC51";
    when 16#0066C# => romdata <= X"97BE3FA3";
    when 16#0066D# => romdata <= X"EF5381B5";
    when 16#0066E# => romdata <= X"B05281B5";
    when 16#0066F# => romdata <= X"D85197B0";
    when 16#00670# => romdata <= X"3FBBEB53";
    when 16#00671# => romdata <= X"81B5E052";
    when 16#00672# => romdata <= X"81B5F051";
    when 16#00673# => romdata <= X"97A23FBB";
    when 16#00674# => romdata <= X"D25381B5";
    when 16#00675# => romdata <= X"F85281B6";
    when 16#00676# => romdata <= X"94519794";
    when 16#00677# => romdata <= X"3FA6A953";
    when 16#00678# => romdata <= X"81B69C52";
    when 16#00679# => romdata <= X"81B6C051";
    when 16#0067A# => romdata <= X"97863FBE";
    when 16#0067B# => romdata <= X"AE5381B6";
    when 16#0067C# => romdata <= X"C85281B6";
    when 16#0067D# => romdata <= X"E85196F8";
    when 16#0067E# => romdata <= X"3FBFCC53";
    when 16#0067F# => romdata <= X"81B6EC52";
    when 16#00680# => romdata <= X"81B79051";
    when 16#00681# => romdata <= X"96EA3FBC";
    when 16#00682# => romdata <= X"825381B7";
    when 16#00683# => romdata <= X"985281B2";
    when 16#00684# => romdata <= X"B05196DC";
    when 16#00685# => romdata <= X"3FBCC353";
    when 16#00686# => romdata <= X"81B7BC52";
    when 16#00687# => romdata <= X"81B7E451";
    when 16#00688# => romdata <= X"96CE3FBD";
    when 16#00689# => romdata <= X"EB5381B7";
    when 16#0068A# => romdata <= X"EC5281B8";
    when 16#0068B# => romdata <= X"8C5196C0";
    when 16#0068C# => romdata <= X"3F889B53";
    when 16#0068D# => romdata <= X"81B89452";
    when 16#0068E# => romdata <= X"81B8B051";
    when 16#0068F# => romdata <= X"96B23FA4";
    when 16#00690# => romdata <= X"BF5381B8";
    when 16#00691# => romdata <= X"B85281B8";
    when 16#00692# => romdata <= X"845196A4";
    when 16#00693# => romdata <= X"3FA48B53";
    when 16#00694# => romdata <= X"81B8D452";
    when 16#00695# => romdata <= X"81B8E851";
    when 16#00696# => romdata <= X"96963FB9";
    when 16#00697# => romdata <= X"905381B8";
    when 16#00698# => romdata <= X"F05281B9";
    when 16#00699# => romdata <= X"8C519688";
    when 16#0069A# => romdata <= X"3FB9B653";
    when 16#0069B# => romdata <= X"81B99452";
    when 16#0069C# => romdata <= X"81B9A851";
    when 16#0069D# => romdata <= X"95FA3FA7";
    when 16#0069E# => romdata <= X"CB5381B9";
    when 16#0069F# => romdata <= X"B05281B9";
    when 16#006A0# => romdata <= X"D45195EC";
    when 16#006A1# => romdata <= X"3F80C0AA";
    when 16#006A2# => romdata <= X"5381B9DC";
    when 16#006A3# => romdata <= X"5281B9EC";
    when 16#006A4# => romdata <= X"5195DD3F";
    when 16#006A5# => romdata <= X"80C2F553";
    when 16#006A6# => romdata <= X"81B9F052";
    when 16#006A7# => romdata <= X"81BA8C51";
    when 16#006A8# => romdata <= X"95CE3FBB";
    when 16#006A9# => romdata <= X"985381BA";
    when 16#006AA# => romdata <= X"945281BA";
    when 16#006AB# => romdata <= X"AC5195C0";
    when 16#006AC# => romdata <= X"3F80C2FD";
    when 16#006AD# => romdata <= X"5381BAB4";
    when 16#006AE# => romdata <= X"5281BAC8";
    when 16#006AF# => romdata <= X"5195B13F";
    when 16#006B0# => romdata <= X"8AD65381";
    when 16#006B1# => romdata <= X"BAD05281";
    when 16#006B2# => romdata <= X"BAE45195";
    when 16#006B3# => romdata <= X"A33F8DE6";
    when 16#006B4# => romdata <= X"5381BAE8";
    when 16#006B5# => romdata <= X"5281BB90";
    when 16#006B6# => romdata <= X"5195953F";
    when 16#006B7# => romdata <= X"BBB45381";
    when 16#006B8# => romdata <= X"BB985281";
    when 16#006B9# => romdata <= X"BBB85195";
    when 16#006BA# => romdata <= X"873F93A3";
    when 16#006BB# => romdata <= X"5381BBC0";
    when 16#006BC# => romdata <= X"5281BBD4";
    when 16#006BD# => romdata <= X"5194F93F";
    when 16#006BE# => romdata <= X"88BE5381";
    when 16#006BF# => romdata <= X"BBDC5281";
    when 16#006C0# => romdata <= X"BBE85194";
    when 16#006C1# => romdata <= X"EB3F89FC";
    when 16#006C2# => romdata <= X"5381BBEC";
    when 16#006C3# => romdata <= X"5281BC94";
    when 16#006C4# => romdata <= X"5194DD3F";
    when 16#006C5# => romdata <= X"88BE5381";
    when 16#006C6# => romdata <= X"BC9C5281";
    when 16#006C7# => romdata <= X"B4D05194";
    when 16#006C8# => romdata <= X"CF3F8AC5";
    when 16#006C9# => romdata <= X"5381BCAC";
    when 16#006CA# => romdata <= X"5281BCBC";
    when 16#006CB# => romdata <= X"5194C13F";
    when 16#006CC# => romdata <= X"88B35381";
    when 16#006CD# => romdata <= X"A7DC5281";
    when 16#006CE# => romdata <= X"A7C05194";
    when 16#006CF# => romdata <= X"B33F80D1";
    when 16#006D0# => romdata <= X"C65381A7";
    when 16#006D1# => romdata <= X"DC5281A7";
    when 16#006D2# => romdata <= X"C85194A4";
    when 16#006D3# => romdata <= X"3F9AF73F";
    when 16#006D4# => romdata <= X"94EA3F81";
    when 16#006D5# => romdata <= X"0B81F1F0";
    when 16#006D6# => romdata <= X"3481DED0";
    when 16#006D7# => romdata <= X"337081FF";
    when 16#006D8# => romdata <= X"06555573";
    when 16#006D9# => romdata <= X"B23880C6";
    when 16#006DA# => romdata <= X"953FB008";
    when 16#006DB# => romdata <= X"903894DA";
    when 16#006DC# => romdata <= X"3F81F1F0";
    when 16#006DD# => romdata <= X"335675E1";
    when 16#006DE# => romdata <= X"38883D0D";
    when 16#006DF# => romdata <= X"0480C691";
    when 16#006E0# => romdata <= X"3FB00881";
    when 16#006E1# => romdata <= X"FF065195";
    when 16#006E2# => romdata <= X"AF3F94BE";
    when 16#006E3# => romdata <= X"3F81F1F0";
    when 16#006E4# => romdata <= X"335675C5";
    when 16#006E5# => romdata <= X"38E33980";
    when 16#006E6# => romdata <= X"0B81DED0";
    when 16#006E7# => romdata <= X"349BC73F";
    when 16#006E8# => romdata <= X"81CEF408";
    when 16#006E9# => romdata <= X"70087087";
    when 16#006EA# => romdata <= X"2A810652";
    when 16#006EB# => romdata <= X"57547380";
    when 16#006EC# => romdata <= X"2E8F3876";
    when 16#006ED# => romdata <= X"802E81C5";
    when 16#006EE# => romdata <= X"38FF1770";
    when 16#006EF# => romdata <= X"81FF0658";
    when 16#006F0# => romdata <= X"5475862A";
    when 16#006F1# => romdata <= X"81065574";
    when 16#006F2# => romdata <= X"802EAA38";
    when 16#006F3# => romdata <= X"7680F738";
    when 16#006F4# => romdata <= X"81960B81";
    when 16#006F5# => romdata <= X"CEF40884";
    when 16#006F6# => romdata <= X"110870EF";
    when 16#006F7# => romdata <= X"FF0A06AE";
    when 16#006F8# => romdata <= X"800A0784";
    when 16#006F9# => romdata <= X"130C5784";
    when 16#006FA# => romdata <= X"110870BE";
    when 16#006FB# => romdata <= X"800A0784";
    when 16#006FC# => romdata <= X"130C5755";
    when 16#006FD# => romdata <= X"5775852A";
    when 16#006FE# => romdata <= X"81065574";
    when 16#006FF# => romdata <= X"802E9638";
    when 16#00700# => romdata <= X"76BA3881";
    when 16#00701# => romdata <= X"960B81CE";
    when 16#00702# => romdata <= X"BC08B811";
    when 16#00703# => romdata <= X"08575557";
    when 16#00704# => romdata <= X"800BB815";
    when 16#00705# => romdata <= X"0C75842A";
    when 16#00706# => romdata <= X"81065675";
    when 16#00707# => romdata <= X"802EFEC6";
    when 16#00708# => romdata <= X"3876802E";
    when 16#00709# => romdata <= X"AC38FF17";
    when 16#0070A# => romdata <= X"7081FF06";
    when 16#0070B# => romdata <= X"585580C4";
    when 16#0070C# => romdata <= X"CD3FB008";
    when 16#0070D# => romdata <= X"802EFEB6";
    when 16#0070E# => romdata <= X"38FEC239";
    when 16#0070F# => romdata <= X"FF177081";
    when 16#00710# => romdata <= X"FF065855";
    when 16#00711# => romdata <= X"D039FF17";
    when 16#00712# => romdata <= X"7081FF06";
    when 16#00713# => romdata <= X"5854FFA5";
    when 16#00714# => romdata <= X"3981960B";
    when 16#00715# => romdata <= X"81CEF408";
    when 16#00716# => romdata <= X"84110884";
    when 16#00717# => romdata <= X"0A078412";
    when 16#00718# => romdata <= X"0C5657A8";
    when 16#00719# => romdata <= X"C83F8052";
    when 16#0071A# => romdata <= X"81C39451";
    when 16#0071B# => romdata <= X"AB923F80";
    when 16#0071C# => romdata <= X"C48C3FB0";
    when 16#0071D# => romdata <= X"08802EFD";
    when 16#0071E# => romdata <= X"F538FE81";
    when 16#0071F# => romdata <= X"39819676";
    when 16#00720# => romdata <= X"822A8306";
    when 16#00721# => romdata <= X"53768306";
    when 16#00722# => romdata <= X"5257F4D3";
    when 16#00723# => romdata <= X"3FFEB239";
    when 16#00724# => romdata <= X"FE3D0D81";
    when 16#00725# => romdata <= X"5195CB3F";
    when 16#00726# => romdata <= X"B00881FF";
    when 16#00727# => romdata <= X"06538251";
    when 16#00728# => romdata <= X"95C03FB0";
    when 16#00729# => romdata <= X"0881FF06";
    when 16#0072A# => romdata <= X"527251F4";
    when 16#0072B# => romdata <= X"B23F800B";
    when 16#0072C# => romdata <= X"B00C843D";
    when 16#0072D# => romdata <= X"0D04F93D";
    when 16#0072E# => romdata <= X"0D815195";
    when 16#0072F# => romdata <= X"A53FB008";
    when 16#00730# => romdata <= X"81FF0681";
    when 16#00731# => romdata <= X"BCC45257";
    when 16#00732# => romdata <= X"BFC23F81";
    when 16#00733# => romdata <= X"BCD851BF";
    when 16#00734# => romdata <= X"BB3FF880";
    when 16#00735# => romdata <= X"809A8054";
    when 16#00736# => romdata <= X"80557370";
    when 16#00737# => romdata <= X"84055508";
    when 16#00738# => romdata <= X"74708405";
    when 16#00739# => romdata <= X"56085456";
    when 16#0073A# => romdata <= X"72A03881";
    when 16#0073B# => romdata <= X"157081FF";
    when 16#0073C# => romdata <= X"06565687";
    when 16#0073D# => romdata <= X"7527E338";
    when 16#0073E# => romdata <= X"76812E80";
    when 16#0073F# => romdata <= X"D9388A51";
    when 16#00740# => romdata <= X"BEF03F76";
    when 16#00741# => romdata <= X"B00C893D";
    when 16#00742# => romdata <= X"0D048A51";
    when 16#00743# => romdata <= X"BEE43F72";
    when 16#00744# => romdata <= X"5180C0C2";
    when 16#00745# => romdata <= X"3FB00881";
    when 16#00746# => romdata <= X"FF065372";
    when 16#00747# => romdata <= X"8C279338";
    when 16#00748# => romdata <= X"A051BECE";
    when 16#00749# => romdata <= X"3F811370";
    when 16#0074A# => romdata <= X"81FF0651";
    when 16#0074B# => romdata <= X"538C7326";
    when 16#0074C# => romdata <= X"EF3881BC";
    when 16#0074D# => romdata <= X"F051BED4";
    when 16#0074E# => romdata <= X"3F7552A0";
    when 16#0074F# => romdata <= X"51BEF03F";
    when 16#00750# => romdata <= X"7551D9C1";
    when 16#00751# => romdata <= X"3F811570";
    when 16#00752# => romdata <= X"81FF0656";
    when 16#00753# => romdata <= X"56877527";
    when 16#00754# => romdata <= X"FF8838FF";
    when 16#00755# => romdata <= X"A339F880";
    when 16#00756# => romdata <= X"809A8054";
    when 16#00757# => romdata <= X"80538074";
    when 16#00758# => romdata <= X"70840556";
    when 16#00759# => romdata <= X"0C807470";
    when 16#0075A# => romdata <= X"8405560C";
    when 16#0075B# => romdata <= X"81137081";
    when 16#0075C# => romdata <= X"FF065455";
    when 16#0075D# => romdata <= X"728726FF";
    when 16#0075E# => romdata <= X"85388074";
    when 16#0075F# => romdata <= X"70840556";
    when 16#00760# => romdata <= X"0C807470";
    when 16#00761# => romdata <= X"8405560C";
    when 16#00762# => romdata <= X"81137081";
    when 16#00763# => romdata <= X"FF065455";
    when 16#00764# => romdata <= X"877327CA";
    when 16#00765# => romdata <= X"38FEE739";
    when 16#00766# => romdata <= X"FE3D0D81";
    when 16#00767# => romdata <= X"5193C33F";
    when 16#00768# => romdata <= X"B00881FF";
    when 16#00769# => romdata <= X"0681CEB4";
    when 16#0076A# => romdata <= X"08718812";
    when 16#0076B# => romdata <= X"0C53B00C";
    when 16#0076C# => romdata <= X"843D0D04";
    when 16#0076D# => romdata <= X"803D0D81";
    when 16#0076E# => romdata <= X"5194D93F";
    when 16#0076F# => romdata <= X"B00883FF";
    when 16#00770# => romdata <= X"FF0651D2";
    when 16#00771# => romdata <= X"EE3FB008";
    when 16#00772# => romdata <= X"83FFFF06";
    when 16#00773# => romdata <= X"B00C823D";
    when 16#00774# => romdata <= X"0D04803D";
    when 16#00775# => romdata <= X"0D815193";
    when 16#00776# => romdata <= X"893FB008";
    when 16#00777# => romdata <= X"81FF0651";
    when 16#00778# => romdata <= X"9E863F80";
    when 16#00779# => romdata <= X"0BB00C82";
    when 16#0077A# => romdata <= X"3D0D0480";
    when 16#0077B# => romdata <= X"3D0D81CF";
    when 16#0077C# => romdata <= X"800851F8";
    when 16#0077D# => romdata <= X"BB9586A1";
    when 16#0077E# => romdata <= X"710C810B";
    when 16#0077F# => romdata <= X"B00C823D";
    when 16#00780# => romdata <= X"0D04FC3D";
    when 16#00781# => romdata <= X"0D815192";
    when 16#00782# => romdata <= X"D93FB008";
    when 16#00783# => romdata <= X"81FF0654";
    when 16#00784# => romdata <= X"825192CE";
    when 16#00785# => romdata <= X"3FB00881";
    when 16#00786# => romdata <= X"FF0681CE";
    when 16#00787# => romdata <= X"F4088411";
    when 16#00788# => romdata <= X"0870FE8F";
    when 16#00789# => romdata <= X"0A067798";
    when 16#0078A# => romdata <= X"2B075154";
    when 16#0078B# => romdata <= X"56537280";
    when 16#0078C# => romdata <= X"2E863871";
    when 16#0078D# => romdata <= X"810A0752";
    when 16#0078E# => romdata <= X"7184160C";
    when 16#0078F# => romdata <= X"71B00C86";
    when 16#00790# => romdata <= X"3D0D04FD";
    when 16#00791# => romdata <= X"3D0D81CE";
    when 16#00792# => romdata <= X"F4088411";
    when 16#00793# => romdata <= X"08555381";
    when 16#00794# => romdata <= X"51928F3F";
    when 16#00795# => romdata <= X"B00881FF";
    when 16#00796# => romdata <= X"0674DFFF";
    when 16#00797# => romdata <= X"FF065452";
    when 16#00798# => romdata <= X"71802E87";
    when 16#00799# => romdata <= X"3873A080";
    when 16#0079A# => romdata <= X"80075382";
    when 16#0079B# => romdata <= X"5191F33F";
    when 16#0079C# => romdata <= X"B00881FF";
    when 16#0079D# => romdata <= X"0673EFFF";
    when 16#0079E# => romdata <= X"0A065552";
    when 16#0079F# => romdata <= X"71802E87";
    when 16#007A0# => romdata <= X"38729080";
    when 16#007A1# => romdata <= X"0A075483";
    when 16#007A2# => romdata <= X"5191D73F";
    when 16#007A3# => romdata <= X"B00881FF";
    when 16#007A4# => romdata <= X"0674F7FF";
    when 16#007A5# => romdata <= X"0A065452";
    when 16#007A6# => romdata <= X"71802E87";
    when 16#007A7# => romdata <= X"38738880";
    when 16#007A8# => romdata <= X"0A075384";
    when 16#007A9# => romdata <= X"5191BB3F";
    when 16#007AA# => romdata <= X"B00881FF";
    when 16#007AB# => romdata <= X"0673FBFF";
    when 16#007AC# => romdata <= X"0A065552";
    when 16#007AD# => romdata <= X"71802E87";
    when 16#007AE# => romdata <= X"38728480";
    when 16#007AF# => romdata <= X"0A075485";
    when 16#007B0# => romdata <= X"51919F3F";
    when 16#007B1# => romdata <= X"B00881FF";
    when 16#007B2# => romdata <= X"0674FDFF";
    when 16#007B3# => romdata <= X"0A065452";
    when 16#007B4# => romdata <= X"71802E87";
    when 16#007B5# => romdata <= X"38738280";
    when 16#007B6# => romdata <= X"0A075381";
    when 16#007B7# => romdata <= X"CEF40873";
    when 16#007B8# => romdata <= X"84120C54";
    when 16#007B9# => romdata <= X"72B00C85";
    when 16#007BA# => romdata <= X"3D0D04FA";
    when 16#007BB# => romdata <= X"3D0D880A";
    when 16#007BC# => romdata <= X"0B81CEB8";
    when 16#007BD# => romdata <= X"088C1108";
    when 16#007BE# => romdata <= X"59555681";
    when 16#007BF# => romdata <= X"5190E33F";
    when 16#007C0# => romdata <= X"B008902B";
    when 16#007C1# => romdata <= X"70902C56";
    when 16#007C2# => romdata <= X"53807727";
    when 16#007C3# => romdata <= X"99388077";
    when 16#007C4# => romdata <= X"54547383";
    when 16#007C5# => romdata <= X"FFFF0676";
    when 16#007C6# => romdata <= X"70840558";
    when 16#007C7# => romdata <= X"0CFF1375";
    when 16#007C8# => romdata <= X"15555372";
    when 16#007C9# => romdata <= X"ED38800B";
    when 16#007CA# => romdata <= X"B00C883D";
    when 16#007CB# => romdata <= X"0D04FC3D";
    when 16#007CC# => romdata <= X"0D81BCF8";
    when 16#007CD# => romdata <= X"51BAD53F";
    when 16#007CE# => romdata <= X"81CEF408";
    when 16#007CF# => romdata <= X"7008709E";
    when 16#007D0# => romdata <= X"2A708106";
    when 16#007D1# => romdata <= X"51545454";
    when 16#007D2# => romdata <= X"81537183";
    when 16#007D3# => romdata <= X"38715372";
    when 16#007D4# => romdata <= X"802E80D2";
    when 16#007D5# => romdata <= X"3881BD88";
    when 16#007D6# => romdata <= X"51BAB13F";
    when 16#007D7# => romdata <= X"81519082";
    when 16#007D8# => romdata <= X"3FB00881";
    when 16#007D9# => romdata <= X"FF0681BC";
    when 16#007DA# => romdata <= X"F85255BA";
    when 16#007DB# => romdata <= X"9F3F7480";
    when 16#007DC# => romdata <= X"2EAB3881";
    when 16#007DD# => romdata <= X"BD9051BA";
    when 16#007DE# => romdata <= X"933F81CE";
    when 16#007DF# => romdata <= X"F4088411";
    when 16#007E0# => romdata <= X"0870FD0A";
    when 16#007E1# => romdata <= X"06545454";
    when 16#007E2# => romdata <= X"74802E86";
    when 16#007E3# => romdata <= X"3872820A";
    when 16#007E4# => romdata <= X"07527184";
    when 16#007E5# => romdata <= X"150C71B0";
    when 16#007E6# => romdata <= X"0C863D0D";
    when 16#007E7# => romdata <= X"0481B2B8";
    when 16#007E8# => romdata <= X"51B9E93F";
    when 16#007E9# => romdata <= X"CE3981B2";
    when 16#007EA# => romdata <= X"B851B9E0";
    when 16#007EB# => romdata <= X"3F81BD88";
    when 16#007EC# => romdata <= X"51B9D93F";
    when 16#007ED# => romdata <= X"81518FAA";
    when 16#007EE# => romdata <= X"3FB00881";
    when 16#007EF# => romdata <= X"FF0681BC";
    when 16#007F0# => romdata <= X"F85255B9";
    when 16#007F1# => romdata <= X"C73F74FF";
    when 16#007F2# => romdata <= X"AA38D239";
    when 16#007F3# => romdata <= X"FD3D0D81";
    when 16#007F4# => romdata <= X"518F8F3F";
    when 16#007F5# => romdata <= X"B00881FF";
    when 16#007F6# => romdata <= X"0681BD9C";
    when 16#007F7# => romdata <= X"5254B9AC";
    when 16#007F8# => romdata <= X"3F73A438";
    when 16#007F9# => romdata <= X"81B2B051";
    when 16#007FA# => romdata <= X"B9A23F81";
    when 16#007FB# => romdata <= X"CEF40884";
    when 16#007FC# => romdata <= X"110870FB";
    when 16#007FD# => romdata <= X"0A068413";
    when 16#007FE# => romdata <= X"0C53538A";
    when 16#007FF# => romdata <= X"51B8F33F";
    when 16#00800# => romdata <= X"73B00C85";
    when 16#00801# => romdata <= X"3D0D0481";
    when 16#00802# => romdata <= X"AED851B8";
    when 16#00803# => romdata <= X"FF3F81CE";
    when 16#00804# => romdata <= X"F4088411";
    when 16#00805# => romdata <= X"0870840A";
    when 16#00806# => romdata <= X"0784130C";
    when 16#00807# => romdata <= X"53538A51";
    when 16#00808# => romdata <= X"B8D03F73";
    when 16#00809# => romdata <= X"B00C853D";
    when 16#0080A# => romdata <= X"0D04FD3D";
    when 16#0080B# => romdata <= X"0D81DECC";
    when 16#0080C# => romdata <= X"0852F881";
    when 16#0080D# => romdata <= X"C08E800B";
    when 16#0080E# => romdata <= X"81CEF408";
    when 16#0080F# => romdata <= X"55537180";
    when 16#00810# => romdata <= X"2E80F738";
    when 16#00811# => romdata <= X"7281FF06";
    when 16#00812# => romdata <= X"84150C81";
    when 16#00813# => romdata <= X"CEB03370";
    when 16#00814# => romdata <= X"81FF0651";
    when 16#00815# => romdata <= X"5271802E";
    when 16#00816# => romdata <= X"80C23872";
    when 16#00817# => romdata <= X"9F2A7310";
    when 16#00818# => romdata <= X"075381DE";
    when 16#00819# => romdata <= X"D0337081";
    when 16#0081A# => romdata <= X"FF065152";
    when 16#0081B# => romdata <= X"71802ED4";
    when 16#0081C# => romdata <= X"38800B81";
    when 16#0081D# => romdata <= X"DED03491";
    when 16#0081E# => romdata <= X"ED3F81CE";
    when 16#0081F# => romdata <= X"C0335473";
    when 16#00820# => romdata <= X"80E23881";
    when 16#00821# => romdata <= X"CEF40873";
    when 16#00822# => romdata <= X"81FF0684";
    when 16#00823# => romdata <= X"120C81CE";
    when 16#00824# => romdata <= X"B0337081";
    when 16#00825# => romdata <= X"FF065153";
    when 16#00826# => romdata <= X"5471C038";
    when 16#00827# => romdata <= X"72812A73";
    when 16#00828# => romdata <= X"9F2B0753";
    when 16#00829# => romdata <= X"FFBC3972";
    when 16#0082A# => romdata <= X"812A739F";
    when 16#0082B# => romdata <= X"2B075380";
    when 16#0082C# => romdata <= X"FD51BAEB";
    when 16#0082D# => romdata <= X"3F81CEF4";
    when 16#0082E# => romdata <= X"08547281";
    when 16#0082F# => romdata <= X"FF068415";
    when 16#00830# => romdata <= X"0C81CEB0";
    when 16#00831# => romdata <= X"337081FF";
    when 16#00832# => romdata <= X"06535471";
    when 16#00833# => romdata <= X"802ED838";
    when 16#00834# => romdata <= X"729F2A73";
    when 16#00835# => romdata <= X"10075380";
    when 16#00836# => romdata <= X"FD51BAC3";
    when 16#00837# => romdata <= X"3F81CEF4";
    when 16#00838# => romdata <= X"0854D739";
    when 16#00839# => romdata <= X"800BB00C";
    when 16#0083A# => romdata <= X"853D0D04";
    when 16#0083B# => romdata <= X"F73D0D85";
    when 16#0083C# => romdata <= X"3D549653";
    when 16#0083D# => romdata <= X"81BDB052";
    when 16#0083E# => romdata <= X"7351BE85";
    when 16#0083F# => romdata <= X"3FA09F3F";
    when 16#00840# => romdata <= X"81518CDE";
    when 16#00841# => romdata <= X"3F805280";
    when 16#00842# => romdata <= X"519DFF3F";
    when 16#00843# => romdata <= X"73538052";
    when 16#00844# => romdata <= X"81C39451";
    when 16#00845# => romdata <= X"B2BE3F80";
    when 16#00846# => romdata <= X"5281519D";
    when 16#00847# => romdata <= X"ED3F7353";
    when 16#00848# => romdata <= X"825281C3";
    when 16#00849# => romdata <= X"9451B2AC";
    when 16#0084A# => romdata <= X"3F805282";
    when 16#0084B# => romdata <= X"519DDB3F";
    when 16#0084C# => romdata <= X"73538152";
    when 16#0084D# => romdata <= X"81C39451";
    when 16#0084E# => romdata <= X"B29A3F80";
    when 16#0084F# => romdata <= X"5284519D";
    when 16#00850# => romdata <= X"C93F7353";
    when 16#00851# => romdata <= X"845281C3";
    when 16#00852# => romdata <= X"9451B288";
    when 16#00853# => romdata <= X"3F805285";
    when 16#00854# => romdata <= X"519DB73F";
    when 16#00855# => romdata <= X"73539052";
    when 16#00856# => romdata <= X"81C39451";
    when 16#00857# => romdata <= X"B1F63F80";
    when 16#00858# => romdata <= X"5286519D";
    when 16#00859# => romdata <= X"A53F7353";
    when 16#0085A# => romdata <= X"835281C3";
    when 16#0085B# => romdata <= X"9451B1E4";
    when 16#0085C# => romdata <= X"3F8B3D0D";
    when 16#0085D# => romdata <= X"04FEF53F";
    when 16#0085E# => romdata <= X"800BB00C";
    when 16#0085F# => romdata <= X"04FC3D0D";
    when 16#00860# => romdata <= X"81A1D854";
    when 16#00861# => romdata <= X"80558452";
    when 16#00862# => romdata <= X"74519CFE";
    when 16#00863# => romdata <= X"3F805373";
    when 16#00864# => romdata <= X"70810555";
    when 16#00865# => romdata <= X"33519DF8";
    when 16#00866# => romdata <= X"3F811370";
    when 16#00867# => romdata <= X"81FF0651";
    when 16#00868# => romdata <= X"5380DC73";
    when 16#00869# => romdata <= X"27E93881";
    when 16#0086A# => romdata <= X"157081FF";
    when 16#0086B# => romdata <= X"06565387";
    when 16#0086C# => romdata <= X"7527D338";
    when 16#0086D# => romdata <= X"800BB00C";
    when 16#0086E# => romdata <= X"863D0D04";
    when 16#0086F# => romdata <= X"FD3D0D81";
    when 16#00870# => romdata <= X"CEB03370";
    when 16#00871# => romdata <= X"81FF0654";
    when 16#00872# => romdata <= X"5472BF26";
    when 16#00873# => romdata <= X"AC3881CE";
    when 16#00874# => romdata <= X"B0337081";
    when 16#00875# => romdata <= X"FF0681CE";
    when 16#00876# => romdata <= X"B4085288";
    when 16#00877# => romdata <= X"120C5480";
    when 16#00878# => romdata <= X"E45280C3";
    when 16#00879# => romdata <= X"BC518FDE";
    when 16#0087A# => romdata <= X"3F81CEB0";
    when 16#0087B# => romdata <= X"33810553";
    when 16#0087C# => romdata <= X"7281CEB0";
    when 16#0087D# => romdata <= X"34853D0D";
    when 16#0087E# => romdata <= X"0480E452";
    when 16#0087F# => romdata <= X"80C49351";
    when 16#00880# => romdata <= X"8FC43F81";
    when 16#00881# => romdata <= X"CEB03381";
    when 16#00882# => romdata <= X"05537281";
    when 16#00883# => romdata <= X"CEB03485";
    when 16#00884# => romdata <= X"3D0D04FD";
    when 16#00885# => romdata <= X"3D0D81CE";
    when 16#00886# => romdata <= X"B0337081";
    when 16#00887# => romdata <= X"FF065454";
    when 16#00888# => romdata <= X"72BF2680";
    when 16#00889# => romdata <= X"C93881CE";
    when 16#0088A# => romdata <= X"B0337081";
    when 16#0088B# => romdata <= X"FF0681CE";
    when 16#0088C# => romdata <= X"B4085688";
    when 16#0088D# => romdata <= X"160C5381";
    when 16#0088E# => romdata <= X"CEB03370";
    when 16#0088F# => romdata <= X"81FF0655";
    when 16#00890# => romdata <= X"5373BF2E";
    when 16#00891# => romdata <= X"80D13880";
    when 16#00892# => romdata <= X"E45280C4";
    when 16#00893# => romdata <= X"93518EF6";
    when 16#00894# => romdata <= X"3F81CEB0";
    when 16#00895# => romdata <= X"33810553";
    when 16#00896# => romdata <= X"7281CEB0";
    when 16#00897# => romdata <= X"3481CEB0";
    when 16#00898# => romdata <= X"3380FF06";
    when 16#00899# => romdata <= X"537281CE";
    when 16#0089A# => romdata <= X"B034853D";
    when 16#0089B# => romdata <= X"0D0481CE";
    when 16#0089C# => romdata <= X"B0337081";
    when 16#0089D# => romdata <= X"FF0680FF";
    when 16#0089E# => romdata <= X"713181CE";
    when 16#0089F# => romdata <= X"B4085288";
    when 16#008A0# => romdata <= X"120C5553";
    when 16#008A1# => romdata <= X"81CEB033";
    when 16#008A2# => romdata <= X"7081FF06";
    when 16#008A3# => romdata <= X"555373BF";
    when 16#008A4# => romdata <= X"2E098106";
    when 16#008A5# => romdata <= X"FFB13880";
    when 16#008A6# => romdata <= X"CE905280";
    when 16#008A7# => romdata <= X"C493518E";
    when 16#008A8# => romdata <= X"A53F81CE";
    when 16#008A9# => romdata <= X"B0338105";
    when 16#008AA# => romdata <= X"537281CE";
    when 16#008AB# => romdata <= X"B03481CE";
    when 16#008AC# => romdata <= X"B03380FF";
    when 16#008AD# => romdata <= X"06537281";
    when 16#008AE# => romdata <= X"CEB03485";
    when 16#008AF# => romdata <= X"3D0D0481";
    when 16#008B0# => romdata <= X"0B81CEC0";
    when 16#008B1# => romdata <= X"3404FE3D";
    when 16#008B2# => romdata <= X"0D81CEF8";
    when 16#008B3# => romdata <= X"08981108";
    when 16#008B4# => romdata <= X"70842A70";
    when 16#008B5# => romdata <= X"81065153";
    when 16#008B6# => romdata <= X"53537080";
    when 16#008B7# => romdata <= X"2E8D3871";
    when 16#008B8# => romdata <= X"EF069814";
    when 16#008B9# => romdata <= X"0C810B81";
    when 16#008BA# => romdata <= X"DED03484";
    when 16#008BB# => romdata <= X"3D0D04FB";
    when 16#008BC# => romdata <= X"3D0D81CE";
    when 16#008BD# => romdata <= X"F4087008";
    when 16#008BE# => romdata <= X"810A0681";
    when 16#008BF# => romdata <= X"DECC0C54";
    when 16#008C0# => romdata <= X"B6C03FB6";
    when 16#008C1# => romdata <= X"E33F8EFB";
    when 16#008C2# => romdata <= X"3F81CEF8";
    when 16#008C3# => romdata <= X"08981108";
    when 16#008C4# => romdata <= X"88079812";
    when 16#008C5# => romdata <= X"0C5481DE";
    when 16#008C6# => romdata <= X"CC0880F8";
    when 16#008C7# => romdata <= X"DC555372";
    when 16#008C8# => romdata <= X"84388880";
    when 16#008C9# => romdata <= X"547381F2";
    when 16#008CA# => romdata <= X"D40C7280";
    when 16#008CB# => romdata <= X"2E849A38";
    when 16#008CC# => romdata <= X"81A8A451";
    when 16#008CD# => romdata <= X"B2D63F8C";
    when 16#008CE# => romdata <= X"51B2B73F";
    when 16#008CF# => romdata <= X"81BDB051";
    when 16#008D0# => romdata <= X"B2CA3F81";
    when 16#008D1# => romdata <= X"DECC0880";
    when 16#008D2# => romdata <= X"2E81D238";
    when 16#008D3# => romdata <= X"81BDC851";
    when 16#008D4# => romdata <= X"B2BA3F81";
    when 16#008D5# => romdata <= X"DECC0854";
    when 16#008D6# => romdata <= X"73802E82";
    when 16#008D7# => romdata <= X"BD3881CE";
    when 16#008D8# => romdata <= X"B8085481";
    when 16#008D9# => romdata <= X"740C81CE";
    when 16#008DA# => romdata <= X"F4088411";
    when 16#008DB# => romdata <= X"08705657";
    when 16#008DC# => romdata <= X"55805373";
    when 16#008DD# => romdata <= X"FE8F0A06";
    when 16#008DE# => romdata <= X"73982B07";
    when 16#008DF# => romdata <= X"7084170C";
    when 16#008E0# => romdata <= X"81147081";
    when 16#008E1# => romdata <= X"FF065154";
    when 16#008E2# => romdata <= X"548F7327";
    when 16#008E3# => romdata <= X"E6387584";
    when 16#008E4# => romdata <= X"160C81CE";
    when 16#008E5# => romdata <= X"BC085480";
    when 16#008E6# => romdata <= X"0BB8150C";
    when 16#008E7# => romdata <= X"825280C5";
    when 16#008E8# => romdata <= X"BF518CA2";
    when 16#008E9# => romdata <= X"3FF881C0";
    when 16#008EA# => romdata <= X"8E800B81";
    when 16#008EB# => romdata <= X"CEF40856";
    when 16#008EC# => romdata <= X"5481DECC";
    when 16#008ED# => romdata <= X"08802E81";
    when 16#008EE# => romdata <= X"B7387381";
    when 16#008EF# => romdata <= X"FF068416";
    when 16#008F0# => romdata <= X"0C81CEB0";
    when 16#008F1# => romdata <= X"337081FF";
    when 16#008F2# => romdata <= X"06545672";
    when 16#008F3# => romdata <= X"802E80C2";
    when 16#008F4# => romdata <= X"38739F2A";
    when 16#008F5# => romdata <= X"74100754";
    when 16#008F6# => romdata <= X"81DED033";
    when 16#008F7# => romdata <= X"7081FF06";
    when 16#008F8# => romdata <= X"57537580";
    when 16#008F9# => romdata <= X"2ED43880";
    when 16#008FA# => romdata <= X"0B81DED0";
    when 16#008FB# => romdata <= X"348AF73F";
    when 16#008FC# => romdata <= X"81CEC033";
    when 16#008FD# => romdata <= X"557482E2";
    when 16#008FE# => romdata <= X"3881CEF4";
    when 16#008FF# => romdata <= X"087481FF";
    when 16#00900# => romdata <= X"0684120C";
    when 16#00901# => romdata <= X"81CEB033";
    when 16#00902# => romdata <= X"7081FF06";
    when 16#00903# => romdata <= X"55575572";
    when 16#00904# => romdata <= X"C0387381";
    when 16#00905# => romdata <= X"2A749F2B";
    when 16#00906# => romdata <= X"0754FFBC";
    when 16#00907# => romdata <= X"3981BDD4";
    when 16#00908# => romdata <= X"51B0E93F";
    when 16#00909# => romdata <= X"810A51B0";
    when 16#0090A# => romdata <= X"E33F81BD";
    when 16#0090B# => romdata <= X"E851B0DC";
    when 16#0090C# => romdata <= X"3F81BE90";
    when 16#0090D# => romdata <= X"51B0D53F";
    when 16#0090E# => romdata <= X"B451B29A";
    when 16#0090F# => romdata <= X"3F81BEA4";
    when 16#00910# => romdata <= X"51B0C93F";
    when 16#00911# => romdata <= X"81BEAC51";
    when 16#00912# => romdata <= X"B0C23F81";
    when 16#00913# => romdata <= X"BEB851B0";
    when 16#00914# => romdata <= X"BB3F81DE";
    when 16#00915# => romdata <= X"CC085473";
    when 16#00916# => romdata <= X"FE8438BE";
    when 16#00917# => romdata <= X"3973812A";
    when 16#00918# => romdata <= X"749F2B07";
    when 16#00919# => romdata <= X"5480FD51";
    when 16#0091A# => romdata <= X"B3B53F81";
    when 16#0091B# => romdata <= X"CEF40855";
    when 16#0091C# => romdata <= X"7381FF06";
    when 16#0091D# => romdata <= X"84160C81";
    when 16#0091E# => romdata <= X"CEB03370";
    when 16#0091F# => romdata <= X"81FF0656";
    when 16#00920# => romdata <= X"5674802E";
    when 16#00921# => romdata <= X"D838739F";
    when 16#00922# => romdata <= X"2A741007";
    when 16#00923# => romdata <= X"5480FD51";
    when 16#00924# => romdata <= X"B38D3F81";
    when 16#00925# => romdata <= X"CEF40855";
    when 16#00926# => romdata <= X"D73981CE";
    when 16#00927# => romdata <= X"BC0874B4";
    when 16#00928# => romdata <= X"120C5681";
    when 16#00929# => romdata <= X"8051C58B";
    when 16#0092A# => romdata <= X"3F828051";
    when 16#0092B# => romdata <= X"C5853F84";
    when 16#0092C# => romdata <= X"8351C4FF";
    when 16#0092D# => romdata <= X"3F86F151";
    when 16#0092E# => romdata <= X"C4F93F88";
    when 16#0092F# => romdata <= X"8351C4F3";
    when 16#00930# => romdata <= X"3F81CEF4";
    when 16#00931# => romdata <= X"08700870";
    when 16#00932# => romdata <= X"9E2A7081";
    when 16#00933# => romdata <= X"06515556";
    when 16#00934# => romdata <= X"54815572";
    when 16#00935# => romdata <= X"802E80FD";
    when 16#00936# => romdata <= X"387481FF";
    when 16#00937# => romdata <= X"06841508";
    when 16#00938# => romdata <= X"70FD0A06";
    when 16#00939# => romdata <= X"58565372";
    when 16#0093A# => romdata <= X"802E8638";
    when 16#0093B# => romdata <= X"74820A07";
    when 16#0093C# => romdata <= X"56758415";
    when 16#0093D# => romdata <= X"0C841408";
    when 16#0093E# => romdata <= X"BE800A07";
    when 16#0093F# => romdata <= X"84150C84";
    when 16#00940# => romdata <= X"1408840A";
    when 16#00941# => romdata <= X"0784150C";
    when 16#00942# => romdata <= X"81CEBC08";
    when 16#00943# => romdata <= X"55800BB8";
    when 16#00944# => romdata <= X"160C81CE";
    when 16#00945# => romdata <= X"B8085481";
    when 16#00946# => romdata <= X"740C93C4";
    when 16#00947# => romdata <= X"5280C2FD";
    when 16#00948# => romdata <= X"5189A33F";
    when 16#00949# => romdata <= X"87E85280";
    when 16#0094A# => romdata <= X"C3BC5189";
    when 16#0094B# => romdata <= X"993FE8E9";
    when 16#0094C# => romdata <= X"3F81CEB8";
    when 16#0094D# => romdata <= X"08548174";
    when 16#0094E# => romdata <= X"0C81CEF4";
    when 16#0094F# => romdata <= X"08841108";
    when 16#00950# => romdata <= X"70565755";
    when 16#00951# => romdata <= X"8053FCAB";
    when 16#00952# => romdata <= X"39B3B83F";
    when 16#00953# => romdata <= X"93C43F97";
    when 16#00954# => romdata <= X"CD3FFBDC";
    when 16#00955# => romdata <= X"397255FF";
    when 16#00956# => romdata <= X"8039B598";
    when 16#00957# => romdata <= X"3F800B81";
    when 16#00958# => romdata <= X"F1E83480";
    when 16#00959# => romdata <= X"0B81F1E4";
    when 16#0095A# => romdata <= X"34800B81";
    when 16#0095B# => romdata <= X"F1EC0C04";
    when 16#0095C# => romdata <= X"FC3D0D76";
    when 16#0095D# => romdata <= X"5281F1E4";
    when 16#0095E# => romdata <= X"33701010";
    when 16#0095F# => romdata <= X"10711005";
    when 16#00960# => romdata <= X"81DED405";
    when 16#00961# => romdata <= X"5254BA87";
    when 16#00962# => romdata <= X"3F775281";
    when 16#00963# => romdata <= X"F1E43370";
    when 16#00964# => romdata <= X"90297131";
    when 16#00965# => romdata <= X"70101081";
    when 16#00966# => romdata <= X"E1940553";
    when 16#00967# => romdata <= X"5555B9EF";
    when 16#00968# => romdata <= X"3F81F1E4";
    when 16#00969# => romdata <= X"33701010";
    when 16#0096A# => romdata <= X"81F09405";
    when 16#0096B# => romdata <= X"7A710C54";
    when 16#0096C# => romdata <= X"81055372";
    when 16#0096D# => romdata <= X"81F1E434";
    when 16#0096E# => romdata <= X"863D0D04";
    when 16#0096F# => romdata <= X"803D0D81";
    when 16#00970# => romdata <= X"BEFC51AD";
    when 16#00971# => romdata <= X"C73F823D";
    when 16#00972# => romdata <= X"0D04FE3D";
    when 16#00973# => romdata <= X"0D81F1EC";
    when 16#00974# => romdata <= X"08537285";
    when 16#00975# => romdata <= X"38843D0D";
    when 16#00976# => romdata <= X"04722DB0";
    when 16#00977# => romdata <= X"0853800B";
    when 16#00978# => romdata <= X"81F1EC0C";
    when 16#00979# => romdata <= X"B0088C38";
    when 16#0097A# => romdata <= X"81BEFC51";
    when 16#0097B# => romdata <= X"AD9E3F84";
    when 16#0097C# => romdata <= X"3D0D0481";
    when 16#0097D# => romdata <= X"C2C051AD";
    when 16#0097E# => romdata <= X"933F7283";
    when 16#0097F# => romdata <= X"FFFF26AA";
    when 16#00980# => romdata <= X"3881FF73";
    when 16#00981# => romdata <= X"27963872";
    when 16#00982# => romdata <= X"529051AD";
    when 16#00983# => romdata <= X"A23F8A51";
    when 16#00984# => romdata <= X"ACE03F81";
    when 16#00985# => romdata <= X"BEFC51AC";
    when 16#00986# => romdata <= X"F33FD439";
    when 16#00987# => romdata <= X"72528851";
    when 16#00988# => romdata <= X"AD8D3F8A";
    when 16#00989# => romdata <= X"51ACCB3F";
    when 16#0098A# => romdata <= X"EA397252";
    when 16#0098B# => romdata <= X"A051ACFF";
    when 16#0098C# => romdata <= X"3F8A51AC";
    when 16#0098D# => romdata <= X"BD3FDC39";
    when 16#0098E# => romdata <= X"FA3D0D02";
    when 16#0098F# => romdata <= X"A3053356";
    when 16#00990# => romdata <= X"758D2E80";
    when 16#00991# => romdata <= X"F4387588";
    when 16#00992# => romdata <= X"32703077";
    when 16#00993# => romdata <= X"80FF3270";
    when 16#00994# => romdata <= X"30728025";
    when 16#00995# => romdata <= X"71802507";
    when 16#00996# => romdata <= X"54515658";
    when 16#00997# => romdata <= X"55749538";
    when 16#00998# => romdata <= X"9F76278C";
    when 16#00999# => romdata <= X"3881F1E8";
    when 16#0099A# => romdata <= X"335580CE";
    when 16#0099B# => romdata <= X"7527AE38";
    when 16#0099C# => romdata <= X"883D0D04";
    when 16#0099D# => romdata <= X"81F1E833";
    when 16#0099E# => romdata <= X"5675802E";
    when 16#0099F# => romdata <= X"F3388851";
    when 16#009A0# => romdata <= X"ABF03FA0";
    when 16#009A1# => romdata <= X"51ABEB3F";
    when 16#009A2# => romdata <= X"8851ABE6";
    when 16#009A3# => romdata <= X"3F81F1E8";
    when 16#009A4# => romdata <= X"33FF0557";
    when 16#009A5# => romdata <= X"7681F1E8";
    when 16#009A6# => romdata <= X"34883D0D";
    when 16#009A7# => romdata <= X"047551AB";
    when 16#009A8# => romdata <= X"D13F81F1";
    when 16#009A9# => romdata <= X"E8338111";
    when 16#009AA# => romdata <= X"55577381";
    when 16#009AB# => romdata <= X"F1E83475";
    when 16#009AC# => romdata <= X"81F19418";
    when 16#009AD# => romdata <= X"34883D0D";
    when 16#009AE# => romdata <= X"048A51AB";
    when 16#009AF# => romdata <= X"B53F81F1";
    when 16#009B0# => romdata <= X"E8338111";
    when 16#009B1# => romdata <= X"56547481";
    when 16#009B2# => romdata <= X"F1E83480";
    when 16#009B3# => romdata <= X"0B81F194";
    when 16#009B4# => romdata <= X"15348056";
    when 16#009B5# => romdata <= X"800B81F1";
    when 16#009B6# => romdata <= X"94173356";
    when 16#009B7# => romdata <= X"5474A02E";
    when 16#009B8# => romdata <= X"83388154";
    when 16#009B9# => romdata <= X"74802E90";
    when 16#009BA# => romdata <= X"3873802E";
    when 16#009BB# => romdata <= X"8B388116";
    when 16#009BC# => romdata <= X"7081FF06";
    when 16#009BD# => romdata <= X"5757DD39";
    when 16#009BE# => romdata <= X"75802EBF";
    when 16#009BF# => romdata <= X"38800B81";
    when 16#009C0# => romdata <= X"F1E43355";
    when 16#009C1# => romdata <= X"55747427";
    when 16#009C2# => romdata <= X"AB387357";
    when 16#009C3# => romdata <= X"74101010";
    when 16#009C4# => romdata <= X"75100576";
    when 16#009C5# => romdata <= X"5481F194";
    when 16#009C6# => romdata <= X"5381DED4";
    when 16#009C7# => romdata <= X"0551B8BB";
    when 16#009C8# => romdata <= X"3FB00880";
    when 16#009C9# => romdata <= X"2EA63881";
    when 16#009CA# => romdata <= X"157081FF";
    when 16#009CB# => romdata <= X"06565476";
    when 16#009CC# => romdata <= X"7526D938";
    when 16#009CD# => romdata <= X"81BF8051";
    when 16#009CE# => romdata <= X"AAD23F81";
    when 16#009CF# => romdata <= X"BEFC51AA";
    when 16#009D0# => romdata <= X"CB3F800B";
    when 16#009D1# => romdata <= X"81F1E834";
    when 16#009D2# => romdata <= X"883D0D04";
    when 16#009D3# => romdata <= X"74101081";
    when 16#009D4# => romdata <= X"F0940570";
    when 16#009D5# => romdata <= X"0881F1EC";
    when 16#009D6# => romdata <= X"0C56800B";
    when 16#009D7# => romdata <= X"81F1E834";
    when 16#009D8# => romdata <= X"E739F73D";
    when 16#009D9# => romdata <= X"0D02AF05";
    when 16#009DA# => romdata <= X"3359800B";
    when 16#009DB# => romdata <= X"81F19433";
    when 16#009DC# => romdata <= X"81F19459";
    when 16#009DD# => romdata <= X"555673A0";
    when 16#009DE# => romdata <= X"2E098106";
    when 16#009DF# => romdata <= X"96388116";
    when 16#009E0# => romdata <= X"7081FF06";
    when 16#009E1# => romdata <= X"81F19411";
    when 16#009E2# => romdata <= X"70335359";
    when 16#009E3# => romdata <= X"575473A0";
    when 16#009E4# => romdata <= X"2EEC3880";
    when 16#009E5# => romdata <= X"58777927";
    when 16#009E6# => romdata <= X"80EA3880";
    when 16#009E7# => romdata <= X"77335654";
    when 16#009E8# => romdata <= X"74742E83";
    when 16#009E9# => romdata <= X"38815474";
    when 16#009EA# => romdata <= X"A02E9A38";
    when 16#009EB# => romdata <= X"7380C538";
    when 16#009EC# => romdata <= X"74A02E91";
    when 16#009ED# => romdata <= X"38811870";
    when 16#009EE# => romdata <= X"81FF0659";
    when 16#009EF# => romdata <= X"55787826";
    when 16#009F0# => romdata <= X"DA3880C0";
    when 16#009F1# => romdata <= X"39811670";
    when 16#009F2# => romdata <= X"81FF0681";
    when 16#009F3# => romdata <= X"F1941170";
    when 16#009F4# => romdata <= X"33575257";
    when 16#009F5# => romdata <= X"5773A02E";
    when 16#009F6# => romdata <= X"098106D9";
    when 16#009F7# => romdata <= X"38811670";
    when 16#009F8# => romdata <= X"81FF0681";
    when 16#009F9# => romdata <= X"F1941170";
    when 16#009FA# => romdata <= X"33575257";
    when 16#009FB# => romdata <= X"5773A02E";
    when 16#009FC# => romdata <= X"D438C239";
    when 16#009FD# => romdata <= X"81167081";
    when 16#009FE# => romdata <= X"FF0681F1";
    when 16#009FF# => romdata <= X"94115957";
    when 16#00A00# => romdata <= X"55FF9839";
    when 16#00A01# => romdata <= X"8A538B3D";
    when 16#00A02# => romdata <= X"FC055276";
    when 16#00A03# => romdata <= X"51BB913F";
    when 16#00A04# => romdata <= X"8B3D0D04";
    when 16#00A05# => romdata <= X"F73D0D02";
    when 16#00A06# => romdata <= X"AF053359";
    when 16#00A07# => romdata <= X"800B81F1";
    when 16#00A08# => romdata <= X"943381F1";
    when 16#00A09# => romdata <= X"94595556";
    when 16#00A0A# => romdata <= X"73A02E09";
    when 16#00A0B# => romdata <= X"81069638";
    when 16#00A0C# => romdata <= X"81167081";
    when 16#00A0D# => romdata <= X"FF0681F1";
    when 16#00A0E# => romdata <= X"94117033";
    when 16#00A0F# => romdata <= X"53595754";
    when 16#00A10# => romdata <= X"73A02EEC";
    when 16#00A11# => romdata <= X"38805877";
    when 16#00A12# => romdata <= X"792780EA";
    when 16#00A13# => romdata <= X"38807733";
    when 16#00A14# => romdata <= X"56547474";
    when 16#00A15# => romdata <= X"2E833881";
    when 16#00A16# => romdata <= X"5474A02E";
    when 16#00A17# => romdata <= X"9A387380";
    when 16#00A18# => romdata <= X"C53874A0";
    when 16#00A19# => romdata <= X"2E913881";
    when 16#00A1A# => romdata <= X"187081FF";
    when 16#00A1B# => romdata <= X"06595578";
    when 16#00A1C# => romdata <= X"7826DA38";
    when 16#00A1D# => romdata <= X"80C03981";
    when 16#00A1E# => romdata <= X"167081FF";
    when 16#00A1F# => romdata <= X"0681F194";
    when 16#00A20# => romdata <= X"11703357";
    when 16#00A21# => romdata <= X"52575773";
    when 16#00A22# => romdata <= X"A02E0981";
    when 16#00A23# => romdata <= X"06D93881";
    when 16#00A24# => romdata <= X"167081FF";
    when 16#00A25# => romdata <= X"0681F194";
    when 16#00A26# => romdata <= X"11703357";
    when 16#00A27# => romdata <= X"52575773";
    when 16#00A28# => romdata <= X"A02ED438";
    when 16#00A29# => romdata <= X"C2398116";
    when 16#00A2A# => romdata <= X"7081FF06";
    when 16#00A2B# => romdata <= X"81F19411";
    when 16#00A2C# => romdata <= X"595755FF";
    when 16#00A2D# => romdata <= X"98399053";
    when 16#00A2E# => romdata <= X"8B3DFC05";
    when 16#00A2F# => romdata <= X"527651BC";
    when 16#00A30# => romdata <= X"FC3F8B3D";
    when 16#00A31# => romdata <= X"0D04FC3D";
    when 16#00A32# => romdata <= X"0D8A51A7";
    when 16#00A33# => romdata <= X"A53F81BF";
    when 16#00A34# => romdata <= X"9451A7B8";
    when 16#00A35# => romdata <= X"3F800B81";
    when 16#00A36# => romdata <= X"F1E43353";
    when 16#00A37# => romdata <= X"53727227";
    when 16#00A38# => romdata <= X"80F53872";
    when 16#00A39# => romdata <= X"10101073";
    when 16#00A3A# => romdata <= X"100581DE";
    when 16#00A3B# => romdata <= X"D4057052";
    when 16#00A3C# => romdata <= X"54A7993F";
    when 16#00A3D# => romdata <= X"72842B70";
    when 16#00A3E# => romdata <= X"7431822B";
    when 16#00A3F# => romdata <= X"81E19411";
    when 16#00A40# => romdata <= X"33515355";
    when 16#00A41# => romdata <= X"71802EB7";
    when 16#00A42# => romdata <= X"387351B3";
    when 16#00A43# => romdata <= X"EF3FB008";
    when 16#00A44# => romdata <= X"81FF0652";
    when 16#00A45# => romdata <= X"71892693";
    when 16#00A46# => romdata <= X"38A051A6";
    when 16#00A47# => romdata <= X"D53F8112";
    when 16#00A48# => romdata <= X"7081FF06";
    when 16#00A49# => romdata <= X"53548972";
    when 16#00A4A# => romdata <= X"27EF3881";
    when 16#00A4B# => romdata <= X"BFAC51A6";
    when 16#00A4C# => romdata <= X"DB3F7473";
    when 16#00A4D# => romdata <= X"31822B81";
    when 16#00A4E# => romdata <= X"E1940551";
    when 16#00A4F# => romdata <= X"A6CE3F8A";
    when 16#00A50# => romdata <= X"51A6AF3F";
    when 16#00A51# => romdata <= X"81137081";
    when 16#00A52# => romdata <= X"FF0681F1";
    when 16#00A53# => romdata <= X"E4335454";
    when 16#00A54# => romdata <= X"55717326";
    when 16#00A55# => romdata <= X"FF8D388A";
    when 16#00A56# => romdata <= X"51A6973F";
    when 16#00A57# => romdata <= X"81F1E433";
    when 16#00A58# => romdata <= X"B00C863D";
    when 16#00A59# => romdata <= X"0D04FE3D";
    when 16#00A5A# => romdata <= X"0D81F2C4";
    when 16#00A5B# => romdata <= X"22FF0551";
    when 16#00A5C# => romdata <= X"7081F2C4";
    when 16#00A5D# => romdata <= X"237083FF";
    when 16#00A5E# => romdata <= X"FF065170";
    when 16#00A5F# => romdata <= X"80C43881";
    when 16#00A60# => romdata <= X"F2C83351";
    when 16#00A61# => romdata <= X"7081FF2E";
    when 16#00A62# => romdata <= X"B9387010";
    when 16#00A63# => romdata <= X"101081F1";
    when 16#00A64# => romdata <= X"F4055271";
    when 16#00A65# => romdata <= X"3381F2C8";
    when 16#00A66# => romdata <= X"34FE7234";
    when 16#00A67# => romdata <= X"81F2C833";
    when 16#00A68# => romdata <= X"70101010";
    when 16#00A69# => romdata <= X"81F1F405";
    when 16#00A6A# => romdata <= X"52538211";
    when 16#00A6B# => romdata <= X"2281F2C4";
    when 16#00A6C# => romdata <= X"23841208";
    when 16#00A6D# => romdata <= X"53722D81";
    when 16#00A6E# => romdata <= X"F2C42251";
    when 16#00A6F# => romdata <= X"70802EFF";
    when 16#00A70# => romdata <= X"BE38843D";
    when 16#00A71# => romdata <= X"0D04F93D";
    when 16#00A72# => romdata <= X"0D02AA05";
    when 16#00A73# => romdata <= X"22568055";
    when 16#00A74# => romdata <= X"74101010";
    when 16#00A75# => romdata <= X"81F1F405";
    when 16#00A76# => romdata <= X"70335252";
    when 16#00A77# => romdata <= X"7081FE2E";
    when 16#00A78# => romdata <= X"99388115";
    when 16#00A79# => romdata <= X"7081FF06";
    when 16#00A7A# => romdata <= X"5652748A";
    when 16#00A7B# => romdata <= X"2E098106";
    when 16#00A7C# => romdata <= X"DF38810B";
    when 16#00A7D# => romdata <= X"B00C893D";
    when 16#00A7E# => romdata <= X"0D0481F2";
    when 16#00A7F# => romdata <= X"C8337081";
    when 16#00A80# => romdata <= X"FF0681F2";
    when 16#00A81# => romdata <= X"C4225354";
    when 16#00A82# => romdata <= X"587281FF";
    when 16#00A83# => romdata <= X"2EB03872";
    when 16#00A84# => romdata <= X"832B5470";
    when 16#00A85# => romdata <= X"762780DE";
    when 16#00A86# => romdata <= X"38757131";
    when 16#00A87# => romdata <= X"7083FFFF";
    when 16#00A88# => romdata <= X"067481F1";
    when 16#00A89# => romdata <= X"F4173370";
    when 16#00A8A# => romdata <= X"832B81F1";
    when 16#00A8B# => romdata <= X"F6112256";
    when 16#00A8C# => romdata <= X"58565257";
    when 16#00A8D# => romdata <= X"577281FF";
    when 16#00A8E# => romdata <= X"2E098106";
    when 16#00A8F# => romdata <= X"D6387272";
    when 16#00A90# => romdata <= X"34758213";
    when 16#00A91# => romdata <= X"23798413";
    when 16#00A92# => romdata <= X"0C7781FF";
    when 16#00A93# => romdata <= X"06547373";
    when 16#00A94# => romdata <= X"2E963876";
    when 16#00A95# => romdata <= X"10101081";
    when 16#00A96# => romdata <= X"F1F40553";
    when 16#00A97# => romdata <= X"74733480";
    when 16#00A98# => romdata <= X"5170B00C";
    when 16#00A99# => romdata <= X"893D0D04";
    when 16#00A9A# => romdata <= X"7481F2C8";
    when 16#00A9B# => romdata <= X"347581F2";
    when 16#00A9C# => romdata <= X"C4238051";
    when 16#00A9D# => romdata <= X"EC397076";
    when 16#00A9E# => romdata <= X"31517081";
    when 16#00A9F# => romdata <= X"F1F61523";
    when 16#00AA0# => romdata <= X"FFBC39FF";
    when 16#00AA1# => romdata <= X"3D0D8A52";
    when 16#00AA2# => romdata <= X"71101010";
    when 16#00AA3# => romdata <= X"81F1EC05";
    when 16#00AA4# => romdata <= X"51FE7134";
    when 16#00AA5# => romdata <= X"FF127081";
    when 16#00AA6# => romdata <= X"FF065351";
    when 16#00AA7# => romdata <= X"71EA38FF";
    when 16#00AA8# => romdata <= X"0B81F2C8";
    when 16#00AA9# => romdata <= X"34833D0D";
    when 16#00AAA# => romdata <= X"04FE3D0D";
    when 16#00AAB# => romdata <= X"02930533";
    when 16#00AAC# => romdata <= X"02840597";
    when 16#00AAD# => romdata <= X"05335452";
    when 16#00AAE# => romdata <= X"71812E92";
    when 16#00AAF# => romdata <= X"387180D5";
    when 16#00AB0# => romdata <= X"2EBB3881";
    when 16#00AB1# => romdata <= X"BFB051A3";
    when 16#00AB2# => romdata <= X"C33F843D";
    when 16#00AB3# => romdata <= X"0D0481BF";
    when 16#00AB4# => romdata <= X"BC51A3B8";
    when 16#00AB5# => romdata <= X"3F72912E";
    when 16#00AB6# => romdata <= X"81EF3872";
    when 16#00AB7# => romdata <= X"9124B538";
    when 16#00AB8# => romdata <= X"728C2E81";
    when 16#00AB9# => romdata <= X"FA38728C";
    when 16#00ABA# => romdata <= X"2480DC38";
    when 16#00ABB# => romdata <= X"72862E81";
    when 16#00ABC# => romdata <= X"CD3881BF";
    when 16#00ABD# => romdata <= X"C851A394";
    when 16#00ABE# => romdata <= X"3F843D0D";
    when 16#00ABF# => romdata <= X"0481BFD8";
    when 16#00AC0# => romdata <= X"51A3893F";
    when 16#00AC1# => romdata <= X"728926EA";
    when 16#00AC2# => romdata <= X"38721010";
    when 16#00AC3# => romdata <= X"81C2EC05";
    when 16#00AC4# => romdata <= X"52710804";
    when 16#00AC5# => romdata <= X"72A82E81";
    when 16#00AC6# => romdata <= X"BB3872A8";
    when 16#00AC7# => romdata <= X"24943872";
    when 16#00AC8# => romdata <= X"9A2E0981";
    when 16#00AC9# => romdata <= X"06CC3881";
    when 16#00ACA# => romdata <= X"BFE451A2";
    when 16#00ACB# => romdata <= X"DF3F843D";
    when 16#00ACC# => romdata <= X"0D047280";
    when 16#00ACD# => romdata <= X"E12E0981";
    when 16#00ACE# => romdata <= X"06FFB738";
    when 16#00ACF# => romdata <= X"81C08051";
    when 16#00AD0# => romdata <= X"A2CA3F84";
    when 16#00AD1# => romdata <= X"3D0D0472";
    when 16#00AD2# => romdata <= X"8F2E0981";
    when 16#00AD3# => romdata <= X"06FFA338";
    when 16#00AD4# => romdata <= X"81C09051";
    when 16#00AD5# => romdata <= X"A2B63F84";
    when 16#00AD6# => romdata <= X"3D0D0481";
    when 16#00AD7# => romdata <= X"C0AC51A2";
    when 16#00AD8# => romdata <= X"AB3F843D";
    when 16#00AD9# => romdata <= X"0D0481BD";
    when 16#00ADA# => romdata <= X"B051A2A0";
    when 16#00ADB# => romdata <= X"3F843D0D";
    when 16#00ADC# => romdata <= X"0481C0C4";
    when 16#00ADD# => romdata <= X"51A2953F";
    when 16#00ADE# => romdata <= X"843D0D04";
    when 16#00ADF# => romdata <= X"81C0D851";
    when 16#00AE0# => romdata <= X"A28A3F84";
    when 16#00AE1# => romdata <= X"3D0D0481";
    when 16#00AE2# => romdata <= X"C0E851A1";
    when 16#00AE3# => romdata <= X"FF3F843D";
    when 16#00AE4# => romdata <= X"0D0481C0";
    when 16#00AE5# => romdata <= X"FC51A1F4";
    when 16#00AE6# => romdata <= X"3F843D0D";
    when 16#00AE7# => romdata <= X"0481C198";
    when 16#00AE8# => romdata <= X"51A1E93F";
    when 16#00AE9# => romdata <= X"843D0D04";
    when 16#00AEA# => romdata <= X"81C1B051";
    when 16#00AEB# => romdata <= X"A1DE3F84";
    when 16#00AEC# => romdata <= X"3D0D0481";
    when 16#00AED# => romdata <= X"C1C451A1";
    when 16#00AEE# => romdata <= X"D33F843D";
    when 16#00AEF# => romdata <= X"0D0481C1";
    when 16#00AF0# => romdata <= X"D451A1C8";
    when 16#00AF1# => romdata <= X"3F843D0D";
    when 16#00AF2# => romdata <= X"0481C1E4";
    when 16#00AF3# => romdata <= X"51A1BD3F";
    when 16#00AF4# => romdata <= X"843D0D04";
    when 16#00AF5# => romdata <= X"81C1F851";
    when 16#00AF6# => romdata <= X"A1B23F84";
    when 16#00AF7# => romdata <= X"3D0D0481";
    when 16#00AF8# => romdata <= X"C29851A1";
    when 16#00AF9# => romdata <= X"A73F843D";
    when 16#00AFA# => romdata <= X"0D04F73D";
    when 16#00AFB# => romdata <= X"0D02B305";
    when 16#00AFC# => romdata <= X"337C7008";
    when 16#00AFD# => romdata <= X"C0808006";
    when 16#00AFE# => romdata <= X"59545A80";
    when 16#00AFF# => romdata <= X"5675832B";
    when 16#00B00# => romdata <= X"7707BFE0";
    when 16#00B01# => romdata <= X"80077070";
    when 16#00B02# => romdata <= X"84055208";
    when 16#00B03# => romdata <= X"71088C2A";
    when 16#00B04# => romdata <= X"BFFE8006";
    when 16#00B05# => romdata <= X"79077198";
    when 16#00B06# => romdata <= X"2A728C2A";
    when 16#00B07# => romdata <= X"9FFF0673";
    when 16#00B08# => romdata <= X"852A708F";
    when 16#00B09# => romdata <= X"06759F06";
    when 16#00B0A# => romdata <= X"5651585D";
    when 16#00B0B# => romdata <= X"58525558";
    when 16#00B0C# => romdata <= X"748D3881";
    when 16#00B0D# => romdata <= X"16568F76";
    when 16#00B0E# => romdata <= X"27C3388B";
    when 16#00B0F# => romdata <= X"3D0D0481";
    when 16#00B10# => romdata <= X"C2A851A0";
    when 16#00B11# => romdata <= X"C73F7551";
    when 16#00B12# => romdata <= X"A28C3F84";
    when 16#00B13# => romdata <= X"52B00851";
    when 16#00B14# => romdata <= X"FFBB873F";
    when 16#00B15# => romdata <= X"81C2B451";
    when 16#00B16# => romdata <= X"A0B23F74";
    when 16#00B17# => romdata <= X"528851A0";
    when 16#00B18# => romdata <= X"CE3F8452";
    when 16#00B19# => romdata <= X"B00851FF";
    when 16#00B1A# => romdata <= X"BAF03F81";
    when 16#00B1B# => romdata <= X"C2BC51A0";
    when 16#00B1C# => romdata <= X"9B3F7852";
    when 16#00B1D# => romdata <= X"9051A0B7";
    when 16#00B1E# => romdata <= X"3F8652B0";
    when 16#00B1F# => romdata <= X"0851FFBA";
    when 16#00B20# => romdata <= X"D93F81C2";
    when 16#00B21# => romdata <= X"C451A084";
    when 16#00B22# => romdata <= X"3F7251A1";
    when 16#00B23# => romdata <= X"C93F8452";
    when 16#00B24# => romdata <= X"B00851FF";
    when 16#00B25# => romdata <= X"BAC43F81";
    when 16#00B26# => romdata <= X"C2CC519F";
    when 16#00B27# => romdata <= X"EF3F7351";
    when 16#00B28# => romdata <= X"A1B43F84";
    when 16#00B29# => romdata <= X"52B00851";
    when 16#00B2A# => romdata <= X"FFBAAF3F";
    when 16#00B2B# => romdata <= X"81C2D451";
    when 16#00B2C# => romdata <= X"9FDA3F77";
    when 16#00B2D# => romdata <= X"52A0519F";
    when 16#00B2E# => romdata <= X"F63F8A52";
    when 16#00B2F# => romdata <= X"B00851FF";
    when 16#00B30# => romdata <= X"BA983F79";
    when 16#00B31# => romdata <= X"92388A51";
    when 16#00B32# => romdata <= X"9FA83F81";
    when 16#00B33# => romdata <= X"16568F76";
    when 16#00B34# => romdata <= X"27FEAA38";
    when 16#00B35# => romdata <= X"FEE53978";
    when 16#00B36# => romdata <= X"81FF0652";
    when 16#00B37# => romdata <= X"7451FBC9";
    when 16#00B38# => romdata <= X"3F8A519F";
    when 16#00B39# => romdata <= X"8D3FE439";
    when 16#00B3A# => romdata <= X"F83D0D02";
    when 16#00B3B# => romdata <= X"AB053359";
    when 16#00B3C# => romdata <= X"80567585";
    when 16#00B3D# => romdata <= X"2BE09011";
    when 16#00B3E# => romdata <= X"E0801208";
    when 16#00B3F# => romdata <= X"70982A71";
    when 16#00B40# => romdata <= X"8C2A9FFF";
    when 16#00B41# => romdata <= X"0672852A";
    when 16#00B42# => romdata <= X"708F0674";
    when 16#00B43# => romdata <= X"9F065551";
    when 16#00B44# => romdata <= X"585B5356";
    when 16#00B45# => romdata <= X"59557480";
    when 16#00B46# => romdata <= X"2E81A738";
    when 16#00B47# => romdata <= X"75BF2681";
    when 16#00B48# => romdata <= X"AF3881C2";
    when 16#00B49# => romdata <= X"DC519EE4";
    when 16#00B4A# => romdata <= X"3F7551A0";
    when 16#00B4B# => romdata <= X"A93F8652";
    when 16#00B4C# => romdata <= X"B00851FF";
    when 16#00B4D# => romdata <= X"B9A43F81";
    when 16#00B4E# => romdata <= X"C2B4519E";
    when 16#00B4F# => romdata <= X"CF3F7452";
    when 16#00B50# => romdata <= X"88519EEB";
    when 16#00B51# => romdata <= X"3F8452B0";
    when 16#00B52# => romdata <= X"0851FFB9";
    when 16#00B53# => romdata <= X"8D3F81C2";
    when 16#00B54# => romdata <= X"BC519EB8";
    when 16#00B55# => romdata <= X"3F765290";
    when 16#00B56# => romdata <= X"519ED43F";
    when 16#00B57# => romdata <= X"8652B008";
    when 16#00B58# => romdata <= X"51FFB8F6";
    when 16#00B59# => romdata <= X"3F81C2C4";
    when 16#00B5A# => romdata <= X"519EA13F";
    when 16#00B5B# => romdata <= X"72519FE6";
    when 16#00B5C# => romdata <= X"3F8452B0";
    when 16#00B5D# => romdata <= X"0851FFB8";
    when 16#00B5E# => romdata <= X"E13F81C2";
    when 16#00B5F# => romdata <= X"CC519E8C";
    when 16#00B60# => romdata <= X"3F73519F";
    when 16#00B61# => romdata <= X"D13F8452";
    when 16#00B62# => romdata <= X"B00851FF";
    when 16#00B63# => romdata <= X"B8CC3F81";
    when 16#00B64# => romdata <= X"C2D4519D";
    when 16#00B65# => romdata <= X"F73F7708";
    when 16#00B66# => romdata <= X"C0808006";
    when 16#00B67# => romdata <= X"52A0519E";
    when 16#00B68# => romdata <= X"8E3F8A52";
    when 16#00B69# => romdata <= X"B00851FF";
    when 16#00B6A# => romdata <= X"B8B03F78";
    when 16#00B6B# => romdata <= X"81B2388A";
    when 16#00B6C# => romdata <= X"519DBF3F";
    when 16#00B6D# => romdata <= X"80537481";
    when 16#00B6E# => romdata <= X"2E81DF38";
    when 16#00B6F# => romdata <= X"76862E81";
    when 16#00B70# => romdata <= X"BB388116";
    when 16#00B71# => romdata <= X"5680FF76";
    when 16#00B72# => romdata <= X"27FEA738";
    when 16#00B73# => romdata <= X"8A3D0D04";
    when 16#00B74# => romdata <= X"81C2E451";
    when 16#00B75# => romdata <= X"9DB63FC0";
    when 16#00B76# => romdata <= X"16519EFA";
    when 16#00B77# => romdata <= X"3F8652B0";
    when 16#00B78# => romdata <= X"0851FFB7";
    when 16#00B79# => romdata <= X"F53F81C2";
    when 16#00B7A# => romdata <= X"B4519DA0";
    when 16#00B7B# => romdata <= X"3F745288";
    when 16#00B7C# => romdata <= X"519DBC3F";
    when 16#00B7D# => romdata <= X"8452B008";
    when 16#00B7E# => romdata <= X"51FFB7DE";
    when 16#00B7F# => romdata <= X"3F81C2BC";
    when 16#00B80# => romdata <= X"519D893F";
    when 16#00B81# => romdata <= X"76529051";
    when 16#00B82# => romdata <= X"9DA53F86";
    when 16#00B83# => romdata <= X"52B00851";
    when 16#00B84# => romdata <= X"FFB7C73F";
    when 16#00B85# => romdata <= X"81C2C451";
    when 16#00B86# => romdata <= X"9CF23F72";
    when 16#00B87# => romdata <= X"519EB73F";
    when 16#00B88# => romdata <= X"8452B008";
    when 16#00B89# => romdata <= X"51FFB7B2";
    when 16#00B8A# => romdata <= X"3F81C2CC";
    when 16#00B8B# => romdata <= X"519CDD3F";
    when 16#00B8C# => romdata <= X"73519EA2";
    when 16#00B8D# => romdata <= X"3F8452B0";
    when 16#00B8E# => romdata <= X"0851FFB7";
    when 16#00B8F# => romdata <= X"9D3F81C2";
    when 16#00B90# => romdata <= X"D4519CC8";
    when 16#00B91# => romdata <= X"3F7708C0";
    when 16#00B92# => romdata <= X"80800652";
    when 16#00B93# => romdata <= X"A0519CDF";
    when 16#00B94# => romdata <= X"3F8A52B0";
    when 16#00B95# => romdata <= X"0851FFB7";
    when 16#00B96# => romdata <= X"813F7880";
    when 16#00B97# => romdata <= X"2EFED038";
    when 16#00B98# => romdata <= X"7681FF06";
    when 16#00B99# => romdata <= X"527451F8";
    when 16#00B9A# => romdata <= X"C03F8A51";
    when 16#00B9B# => romdata <= X"9C843F80";
    when 16#00B9C# => romdata <= X"5374812E";
    when 16#00B9D# => romdata <= X"098106FE";
    when 16#00B9E# => romdata <= X"C3389F39";
    when 16#00B9F# => romdata <= X"72810657";
    when 16#00BA0# => romdata <= X"76802EFE";
    when 16#00BA1# => romdata <= X"BD387852";
    when 16#00BA2# => romdata <= X"7751FADE";
    when 16#00BA3# => romdata <= X"3F811656";
    when 16#00BA4# => romdata <= X"80FF7627";
    when 16#00BA5# => romdata <= X"FCDC38FE";
    when 16#00BA6# => romdata <= X"B3397453";
    when 16#00BA7# => romdata <= X"76862E09";
    when 16#00BA8# => romdata <= X"8106FE9E";
    when 16#00BA9# => romdata <= X"38D63980";
    when 16#00BAA# => romdata <= X"3D0D81CE";
    when 16#00BAB# => romdata <= X"EC085199";
    when 16#00BAC# => romdata <= X"710C8180";
    when 16#00BAD# => romdata <= X"0B84120C";
    when 16#00BAE# => romdata <= X"81CEE808";
    when 16#00BAF# => romdata <= X"5199710C";
    when 16#00BB0# => romdata <= X"81800B84";
    when 16#00BB1# => romdata <= X"120C823D";
    when 16#00BB2# => romdata <= X"0D04FE3D";
    when 16#00BB3# => romdata <= X"0D740284";
    when 16#00BB4# => romdata <= X"05970533";
    when 16#00BB5# => romdata <= X"0288059B";
    when 16#00BB6# => romdata <= X"05338813";
    when 16#00BB7# => romdata <= X"0C8C120C";
    when 16#00BB8# => romdata <= X"538C1308";
    when 16#00BB9# => romdata <= X"70812A81";
    when 16#00BBA# => romdata <= X"06515271";
    when 16#00BBB# => romdata <= X"F4388C13";
    when 16#00BBC# => romdata <= X"087081FF";
    when 16#00BBD# => romdata <= X"06B00C51";
    when 16#00BBE# => romdata <= X"843D0D04";
    when 16#00BBF# => romdata <= X"803D0D72";
    when 16#00BC0# => romdata <= X"8C110870";
    when 16#00BC1# => romdata <= X"872A8132";
    when 16#00BC2# => romdata <= X"8106B00C";
    when 16#00BC3# => romdata <= X"5151823D";
    when 16#00BC4# => romdata <= X"0D04FE3D";
    when 16#00BC5# => romdata <= X"0DFF903F";
    when 16#00BC6# => romdata <= X"81EC5381";
    when 16#00BC7# => romdata <= X"905281CE";
    when 16#00BC8# => romdata <= X"EC0851FF";
    when 16#00BC9# => romdata <= X"A53F9D53";
    when 16#00BCA# => romdata <= X"905281CE";
    when 16#00BCB# => romdata <= X"EC0851FF";
    when 16#00BCC# => romdata <= X"993F80C5";
    when 16#00BCD# => romdata <= X"5380D052";
    when 16#00BCE# => romdata <= X"81CEEC08";
    when 16#00BCF# => romdata <= X"51FF8B3F";
    when 16#00BD0# => romdata <= X"81EC5381";
    when 16#00BD1# => romdata <= X"905281CE";
    when 16#00BD2# => romdata <= X"EC0851FE";
    when 16#00BD3# => romdata <= X"FD3FA153";
    when 16#00BD4# => romdata <= X"905281CE";
    when 16#00BD5# => romdata <= X"EC0851FE";
    when 16#00BD6# => romdata <= X"F13F8953";
    when 16#00BD7# => romdata <= X"80D05281";
    when 16#00BD8# => romdata <= X"CEEC0851";
    when 16#00BD9# => romdata <= X"FEE43F81";
    when 16#00BDA# => romdata <= X"EC538190";
    when 16#00BDB# => romdata <= X"5281CEEC";
    when 16#00BDC# => romdata <= X"0851FED6";
    when 16#00BDD# => romdata <= X"3FB35390";
    when 16#00BDE# => romdata <= X"5281CEEC";
    when 16#00BDF# => romdata <= X"0851FECA";
    when 16#00BE0# => romdata <= X"3F885380";
    when 16#00BE1# => romdata <= X"D05281CE";
    when 16#00BE2# => romdata <= X"EC0851FE";
    when 16#00BE3# => romdata <= X"BD3F81EC";
    when 16#00BE4# => romdata <= X"53819052";
    when 16#00BE5# => romdata <= X"81CEEC08";
    when 16#00BE6# => romdata <= X"51FEAF3F";
    when 16#00BE7# => romdata <= X"B4539052";
    when 16#00BE8# => romdata <= X"81CEEC08";
    when 16#00BE9# => romdata <= X"51FEA33F";
    when 16#00BEA# => romdata <= X"965380D0";
    when 16#00BEB# => romdata <= X"5281CEEC";
    when 16#00BEC# => romdata <= X"0851FE96";
    when 16#00BED# => romdata <= X"3F81EC53";
    when 16#00BEE# => romdata <= X"81905281";
    when 16#00BEF# => romdata <= X"CEEC0851";
    when 16#00BF0# => romdata <= X"FE883FB6";
    when 16#00BF1# => romdata <= X"53905281";
    when 16#00BF2# => romdata <= X"CEEC0851";
    when 16#00BF3# => romdata <= X"FDFC3F80";
    when 16#00BF4# => romdata <= X"E05380D0";
    when 16#00BF5# => romdata <= X"5281CEEC";
    when 16#00BF6# => romdata <= X"0851FDEE";
    when 16#00BF7# => romdata <= X"3F81EC53";
    when 16#00BF8# => romdata <= X"81905281";
    when 16#00BF9# => romdata <= X"CEEC0851";
    when 16#00BFA# => romdata <= X"FDE03F80";
    when 16#00BFB# => romdata <= X"C9539052";
    when 16#00BFC# => romdata <= X"81CEEC08";
    when 16#00BFD# => romdata <= X"51FDD33F";
    when 16#00BFE# => romdata <= X"81C05380";
    when 16#00BFF# => romdata <= X"D05281CE";
    when 16#00C00# => romdata <= X"EC0851FD";
    when 16#00C01# => romdata <= X"C53F843D";
    when 16#00C02# => romdata <= X"0D04FD3D";
    when 16#00C03# => romdata <= X"0D029705";
    when 16#00C04# => romdata <= X"33028405";
    when 16#00C05# => romdata <= X"9B053371";
    when 16#00C06# => romdata <= X"81B00781";
    when 16#00C07# => romdata <= X"BF065354";
    when 16#00C08# => romdata <= X"54F88080";
    when 16#00C09# => romdata <= X"98807171";
    when 16#00C0A# => romdata <= X"0C73842A";
    when 16#00C0B# => romdata <= X"9007710C";
    when 16#00C0C# => romdata <= X"738F0671";
    when 16#00C0D# => romdata <= X"0C527281";
    when 16#00C0E# => romdata <= X"CEC83473";
    when 16#00C0F# => romdata <= X"81CECC34";
    when 16#00C10# => romdata <= X"853D0D04";
    when 16#00C11# => romdata <= X"FD3D0D02";
    when 16#00C12# => romdata <= X"97053381";
    when 16#00C13# => romdata <= X"CECC3354";
    when 16#00C14# => romdata <= X"73058706";
    when 16#00C15# => romdata <= X"0284059A";
    when 16#00C16# => romdata <= X"052281CE";
    when 16#00C17# => romdata <= X"C8335473";
    when 16#00C18# => romdata <= X"057081FF";
    when 16#00C19# => romdata <= X"067281B0";
    when 16#00C1A# => romdata <= X"07545154";
    when 16#00C1B# => romdata <= X"54F88080";
    when 16#00C1C# => romdata <= X"98807171";
    when 16#00C1D# => romdata <= X"0C73842A";
    when 16#00C1E# => romdata <= X"9007710C";
    when 16#00C1F# => romdata <= X"738F0671";
    when 16#00C20# => romdata <= X"0C527281";
    when 16#00C21# => romdata <= X"CEC83473";
    when 16#00C22# => romdata <= X"81CECC34";
    when 16#00C23# => romdata <= X"853D0D04";
    when 16#00C24# => romdata <= X"FF3D0D02";
    when 16#00C25# => romdata <= X"8F0533F8";
    when 16#00C26# => romdata <= X"80809884";
    when 16#00C27# => romdata <= X"0C81CEC8";
    when 16#00C28# => romdata <= X"33810551";
    when 16#00C29# => romdata <= X"7081CEC8";
    when 16#00C2A# => romdata <= X"34833D0D";
    when 16#00C2B# => romdata <= X"04FF3D0D";
    when 16#00C2C# => romdata <= X"80527181";
    when 16#00C2D# => romdata <= X"B00781BF";
    when 16#00C2E# => romdata <= X"06F88080";
    when 16#00C2F# => romdata <= X"98800C90";
    when 16#00C30# => romdata <= X"0BF88080";
    when 16#00C31# => romdata <= X"98800C80";
    when 16#00C32# => romdata <= X"0BF88080";
    when 16#00C33# => romdata <= X"98800C80";
    when 16#00C34# => romdata <= X"51800BF8";
    when 16#00C35# => romdata <= X"80809884";
    when 16#00C36# => romdata <= X"0C811170";
    when 16#00C37# => romdata <= X"81FF0651";
    when 16#00C38# => romdata <= X"5180E571";
    when 16#00C39# => romdata <= X"27EB3881";
    when 16#00C3A# => romdata <= X"127081FF";
    when 16#00C3B# => romdata <= X"06535187";
    when 16#00C3C# => romdata <= X"7227FFBE";
    when 16#00C3D# => romdata <= X"3881B00B";
    when 16#00C3E# => romdata <= X"F8808098";
    when 16#00C3F# => romdata <= X"800C900B";
    when 16#00C40# => romdata <= X"F8808098";
    when 16#00C41# => romdata <= X"800C800B";
    when 16#00C42# => romdata <= X"F8808098";
    when 16#00C43# => romdata <= X"800C800B";
    when 16#00C44# => romdata <= X"81CEC834";
    when 16#00C45# => romdata <= X"800B81CE";
    when 16#00C46# => romdata <= X"CC34833D";
    when 16#00C47# => romdata <= X"0D04FF3D";
    when 16#00C48# => romdata <= X"0D80C00B";
    when 16#00C49# => romdata <= X"F8808098";
    when 16#00C4A# => romdata <= X"800C81A1";
    when 16#00C4B# => romdata <= X"0BF88080";
    when 16#00C4C# => romdata <= X"98800C81";
    when 16#00C4D# => romdata <= X"C00BF880";
    when 16#00C4E# => romdata <= X"8098800C";
    when 16#00C4F# => romdata <= X"81A40BF8";
    when 16#00C50# => romdata <= X"80809880";
    when 16#00C51# => romdata <= X"0C81A60B";
    when 16#00C52# => romdata <= X"F8808098";
    when 16#00C53# => romdata <= X"800C81A2";
    when 16#00C54# => romdata <= X"0BF88080";
    when 16#00C55# => romdata <= X"98800CAF";
    when 16#00C56# => romdata <= X"0BF88080";
    when 16#00C57# => romdata <= X"98800CA5";
    when 16#00C58# => romdata <= X"0BF88080";
    when 16#00C59# => romdata <= X"98800C81";
    when 16#00C5A# => romdata <= X"810BF880";
    when 16#00C5B# => romdata <= X"8098800C";
    when 16#00C5C# => romdata <= X"9D0BF880";
    when 16#00C5D# => romdata <= X"8098800C";
    when 16#00C5E# => romdata <= X"81FA0BF8";
    when 16#00C5F# => romdata <= X"80809880";
    when 16#00C60# => romdata <= X"0C800BF8";
    when 16#00C61# => romdata <= X"80809880";
    when 16#00C62# => romdata <= X"0C805271";
    when 16#00C63# => romdata <= X"81B00781";
    when 16#00C64# => romdata <= X"BF06F880";
    when 16#00C65# => romdata <= X"8098800C";
    when 16#00C66# => romdata <= X"900BF880";
    when 16#00C67# => romdata <= X"8098800C";
    when 16#00C68# => romdata <= X"800BF880";
    when 16#00C69# => romdata <= X"8098800C";
    when 16#00C6A# => romdata <= X"8051800B";
    when 16#00C6B# => romdata <= X"F8808098";
    when 16#00C6C# => romdata <= X"840C8111";
    when 16#00C6D# => romdata <= X"7081FF06";
    when 16#00C6E# => romdata <= X"515180E5";
    when 16#00C6F# => romdata <= X"7127EB38";
    when 16#00C70# => romdata <= X"81127081";
    when 16#00C71# => romdata <= X"FF065351";
    when 16#00C72# => romdata <= X"877227FF";
    when 16#00C73# => romdata <= X"BE3881B0";
    when 16#00C74# => romdata <= X"0BF88080";
    when 16#00C75# => romdata <= X"98800C90";
    when 16#00C76# => romdata <= X"0BF88080";
    when 16#00C77# => romdata <= X"98800C80";
    when 16#00C78# => romdata <= X"0BF88080";
    when 16#00C79# => romdata <= X"98800C80";
    when 16#00C7A# => romdata <= X"0B81CEC8";
    when 16#00C7B# => romdata <= X"34800B81";
    when 16#00C7C# => romdata <= X"CECC3481";
    when 16#00C7D# => romdata <= X"AF0BF880";
    when 16#00C7E# => romdata <= X"8098800C";
    when 16#00C7F# => romdata <= X"833D0D04";
    when 16#00C80# => romdata <= X"803D0D02";
    when 16#00C81# => romdata <= X"8F053373";
    when 16#00C82# => romdata <= X"81F2CC0C";
    when 16#00C83# => romdata <= X"517081F2";
    when 16#00C84# => romdata <= X"D034823D";
    when 16#00C85# => romdata <= X"0D04EE3D";
    when 16#00C86# => romdata <= X"0D640284";
    when 16#00C87# => romdata <= X"0580D705";
    when 16#00C88# => romdata <= X"33028805";
    when 16#00C89# => romdata <= X"80DB0533";
    when 16#00C8A# => romdata <= X"59575980";
    when 16#00C8B# => romdata <= X"76810677";
    when 16#00C8C# => romdata <= X"812A8106";
    when 16#00C8D# => romdata <= X"78832B81";
    when 16#00C8E# => romdata <= X"80067982";
    when 16#00C8F# => romdata <= X"2A810657";
    when 16#00C90# => romdata <= X"5E415F5D";
    when 16#00C91# => romdata <= X"81FF4272";
    when 16#00C92# => romdata <= X"7D2E0981";
    when 16#00C93# => romdata <= X"0683387C";
    when 16#00C94# => romdata <= X"42768A2E";
    when 16#00C95# => romdata <= X"83B93888";
    when 16#00C96# => romdata <= X"19085574";
    when 16#00C97# => romdata <= X"802E83A4";
    when 16#00C98# => romdata <= X"38851933";
    when 16#00C99# => romdata <= X"5AFF5376";
    when 16#00C9A# => romdata <= X"7A268E38";
    when 16#00C9B# => romdata <= X"84193354";
    when 16#00C9C# => romdata <= X"73772685";
    when 16#00C9D# => romdata <= X"38767431";
    when 16#00C9E# => romdata <= X"53741370";
    when 16#00C9F# => romdata <= X"33545872";
    when 16#00CA0# => romdata <= X"81FF0683";
    when 16#00CA1# => romdata <= X"1A337098";
    when 16#00CA2# => romdata <= X"2B81FF0A";
    when 16#00CA3# => romdata <= X"119B2A81";
    when 16#00CA4# => romdata <= X"055B4542";
    when 16#00CA5# => romdata <= X"40815374";
    when 16#00CA6# => romdata <= X"83387453";
    when 16#00CA7# => romdata <= X"7281FF06";
    when 16#00CA8# => romdata <= X"43807A81";
    when 16#00CA9# => romdata <= X"FF06545C";
    when 16#00CAA# => romdata <= X"FF547673";
    when 16#00CAB# => romdata <= X"268B3884";
    when 16#00CAC# => romdata <= X"19335376";
    when 16#00CAD# => romdata <= X"732783F4";
    when 16#00CAE# => romdata <= X"38737481";
    when 16#00CAF# => romdata <= X"FF065553";
    when 16#00CB0# => romdata <= X"805A7973";
    when 16#00CB1# => romdata <= X"24AB3874";
    when 16#00CB2# => romdata <= X"7A2E0981";
    when 16#00CB3# => romdata <= X"0682E138";
    when 16#00CB4# => romdata <= X"60982B81";
    when 16#00CB5# => romdata <= X"FF0A119B";
    when 16#00CB6# => romdata <= X"2A821B33";
    when 16#00CB7# => romdata <= X"71712911";
    when 16#00CB8# => romdata <= X"7081FF06";
    when 16#00CB9# => romdata <= X"7871298C";
    when 16#00CBA# => romdata <= X"1F080552";
    when 16#00CBB# => romdata <= X"455D575D";
    when 16#00CBC# => romdata <= X"537F6305";
    when 16#00CBD# => romdata <= X"7081FF06";
    when 16#00CBE# => romdata <= X"70612B70";
    when 16#00CBF# => romdata <= X"81FF067B";
    when 16#00CC0# => romdata <= X"622B7081";
    when 16#00CC1# => romdata <= X"FF067B83";
    when 16#00CC2# => romdata <= X"2A81065F";
    when 16#00CC3# => romdata <= X"5358525E";
    when 16#00CC4# => romdata <= X"42557880";
    when 16#00CC5# => romdata <= X"2E8F3881";
    when 16#00CC6# => romdata <= X"CEC83361";
    when 16#00CC7# => romdata <= X"05567580";
    when 16#00CC8# => romdata <= X"E62483C5";
    when 16#00CC9# => romdata <= X"387F7829";
    when 16#00CCA# => romdata <= X"61304157";
    when 16#00CCB# => romdata <= X"7C7E2C98";
    when 16#00CCC# => romdata <= X"2B70982C";
    when 16#00CCD# => romdata <= X"55557377";
    when 16#00CCE# => romdata <= X"25818238";
    when 16#00CCF# => romdata <= X"FF1C7D81";
    when 16#00CD0# => romdata <= X"065A537C";
    when 16#00CD1# => romdata <= X"732E83C4";
    when 16#00CD2# => romdata <= X"387E86A6";
    when 16#00CD3# => romdata <= X"386184EB";
    when 16#00CD4# => romdata <= X"387D802E";
    when 16#00CD5# => romdata <= X"82A43879";
    when 16#00CD6# => romdata <= X"14703370";
    when 16#00CD7# => romdata <= X"58545580";
    when 16#00CD8# => romdata <= X"5578752E";
    when 16#00CD9# => romdata <= X"85387284";
    when 16#00CDA# => romdata <= X"2A567583";
    when 16#00CDB# => romdata <= X"2A708106";
    when 16#00CDC# => romdata <= X"51537280";
    when 16#00CDD# => romdata <= X"2E843881";
    when 16#00CDE# => romdata <= X"C0557582";
    when 16#00CDF# => romdata <= X"2A708106";
    when 16#00CE0# => romdata <= X"51537280";
    when 16#00CE1# => romdata <= X"2E853874";
    when 16#00CE2# => romdata <= X"B0075575";
    when 16#00CE3# => romdata <= X"812A7081";
    when 16#00CE4# => romdata <= X"06515372";
    when 16#00CE5# => romdata <= X"802E8538";
    when 16#00CE6# => romdata <= X"748C0755";
    when 16#00CE7# => romdata <= X"75810653";
    when 16#00CE8# => romdata <= X"72802E85";
    when 16#00CE9# => romdata <= X"38748307";
    when 16#00CEA# => romdata <= X"557451F9";
    when 16#00CEB# => romdata <= X"E33F7714";
    when 16#00CEC# => romdata <= X"982B7098";
    when 16#00CED# => romdata <= X"2C555676";
    when 16#00CEE# => romdata <= X"7424FF9B";
    when 16#00CEF# => romdata <= X"3862802E";
    when 16#00CF0# => romdata <= X"953861FF";
    when 16#00CF1# => romdata <= X"1D54547C";
    when 16#00CF2# => romdata <= X"732E81FB";
    when 16#00CF3# => romdata <= X"387351F9";
    when 16#00CF4# => romdata <= X"BF3F7E81";
    when 16#00CF5# => romdata <= X"EA387F52";
    when 16#00CF6# => romdata <= X"8151F8E8";
    when 16#00CF7# => romdata <= X"3F811D70";
    when 16#00CF8# => romdata <= X"81FF065E";
    when 16#00CF9# => romdata <= X"547B7D26";
    when 16#00CFA# => romdata <= X"FEC23860";
    when 16#00CFB# => romdata <= X"527B3070";
    when 16#00CFC# => romdata <= X"982B7098";
    when 16#00CFD# => romdata <= X"2C53585B";
    when 16#00CFE# => romdata <= X"F8CA3F60";
    when 16#00CFF# => romdata <= X"5372B00C";
    when 16#00D00# => romdata <= X"943D0D04";
    when 16#00D01# => romdata <= X"82193385";
    when 16#00D02# => romdata <= X"1A335B53";
    when 16#00D03# => romdata <= X"FCF13981";
    when 16#00D04# => romdata <= X"CECC3353";
    when 16#00D05# => romdata <= X"72872681";
    when 16#00D06# => romdata <= X"9A388113";
    when 16#00D07# => romdata <= X"56805275";
    when 16#00D08# => romdata <= X"81FF0651";
    when 16#00D09# => romdata <= X"F7E43F80";
    when 16#00D0A# => romdata <= X"5372B00C";
    when 16#00D0B# => romdata <= X"943D0D04";
    when 16#00D0C# => romdata <= X"73802EAF";
    when 16#00D0D# => romdata <= X"38FF1470";
    when 16#00D0E# => romdata <= X"81FF0655";
    when 16#00D0F# => romdata <= X"5A7381FF";
    when 16#00D10# => romdata <= X"2EA13874";
    when 16#00D11# => romdata <= X"70810556";
    when 16#00D12# => romdata <= X"337C0570";
    when 16#00D13# => romdata <= X"83FFFF06";
    when 16#00D14# => romdata <= X"FF167081";
    when 16#00D15# => romdata <= X"FF06575C";
    when 16#00D16# => romdata <= X"5D537381";
    when 16#00D17# => romdata <= X"FF2E0981";
    when 16#00D18# => romdata <= X"06E13860";
    when 16#00D19# => romdata <= X"982B81FF";
    when 16#00D1A# => romdata <= X"0A119B2A";
    when 16#00D1B# => romdata <= X"707E291E";
    when 16#00D1C# => romdata <= X"8C1C0805";
    when 16#00D1D# => romdata <= X"5C4255FC";
    when 16#00D1E# => romdata <= X"F8397914";
    when 16#00D1F# => romdata <= X"70335259";
    when 16#00D20# => romdata <= X"F88E3F77";
    when 16#00D21# => romdata <= X"14982B70";
    when 16#00D22# => romdata <= X"982C5556";
    when 16#00D23# => romdata <= X"737725FE";
    when 16#00D24# => romdata <= X"AC387914";
    when 16#00D25# => romdata <= X"70335259";
    when 16#00D26# => romdata <= X"F7F63F77";
    when 16#00D27# => romdata <= X"14982B70";
    when 16#00D28# => romdata <= X"982C5556";
    when 16#00D29# => romdata <= X"767424D2";
    when 16#00D2A# => romdata <= X"38FE9239";
    when 16#00D2B# => romdata <= X"76733154";
    when 16#00D2C# => romdata <= X"FC873980";
    when 16#00D2D# => romdata <= X"528051F6";
    when 16#00D2E# => romdata <= X"D13F8053";
    when 16#00D2F# => romdata <= X"FEEB3973";
    when 16#00D30# => romdata <= X"51F7CD3F";
    when 16#00D31# => romdata <= X"FE903961";
    when 16#00D32# => romdata <= X"7B327081";
    when 16#00D33# => romdata <= X"FF065555";
    when 16#00D34# => romdata <= X"7D802EFD";
    when 16#00D35# => romdata <= X"F8387A81";
    when 16#00D36# => romdata <= X"2A743270";
    when 16#00D37# => romdata <= X"5254F7B0";
    when 16#00D38# => romdata <= X"3F7E802E";
    when 16#00D39# => romdata <= X"FDF038D7";
    when 16#00D3A# => romdata <= X"3981CECC";
    when 16#00D3B# => romdata <= X"337C0553";
    when 16#00D3C# => romdata <= X"80527281";
    when 16#00D3D# => romdata <= X"FF0651F6";
    when 16#00D3E# => romdata <= X"913F8053";
    when 16#00D3F# => romdata <= X"76A02EFD";
    when 16#00D40# => romdata <= X"FC387F78";
    when 16#00D41# => romdata <= X"29613041";
    when 16#00D42# => romdata <= X"57FCA139";
    when 16#00D43# => romdata <= X"7E87AD38";
    when 16#00D44# => romdata <= X"6185EB38";
    when 16#00D45# => romdata <= X"7D802E80";
    when 16#00D46# => romdata <= X"EC387914";
    when 16#00D47# => romdata <= X"70337C07";
    when 16#00D48# => romdata <= X"70525456";
    when 16#00D49# => romdata <= X"80557875";
    when 16#00D4A# => romdata <= X"2E853872";
    when 16#00D4B# => romdata <= X"842A5675";
    when 16#00D4C# => romdata <= X"832A7081";
    when 16#00D4D# => romdata <= X"06515372";
    when 16#00D4E# => romdata <= X"802E8438";
    when 16#00D4F# => romdata <= X"81C05575";
    when 16#00D50# => romdata <= X"822A7081";
    when 16#00D51# => romdata <= X"06515372";
    when 16#00D52# => romdata <= X"802E8538";
    when 16#00D53# => romdata <= X"74B00755";
    when 16#00D54# => romdata <= X"75812A70";
    when 16#00D55# => romdata <= X"81065153";
    when 16#00D56# => romdata <= X"72802E85";
    when 16#00D57# => romdata <= X"38748C07";
    when 16#00D58# => romdata <= X"55758106";
    when 16#00D59# => romdata <= X"5372802E";
    when 16#00D5A# => romdata <= X"85387483";
    when 16#00D5B# => romdata <= X"07557451";
    when 16#00D5C# => romdata <= X"F69E3F77";
    when 16#00D5D# => romdata <= X"14982B70";
    when 16#00D5E# => romdata <= X"982C5553";
    when 16#00D5F# => romdata <= X"767424FF";
    when 16#00D60# => romdata <= X"9938FCB9";
    when 16#00D61# => romdata <= X"39791470";
    when 16#00D62# => romdata <= X"337C0752";
    when 16#00D63# => romdata <= X"56F6813F";
    when 16#00D64# => romdata <= X"7714982B";
    when 16#00D65# => romdata <= X"70982C55";
    when 16#00D66# => romdata <= X"59737725";
    when 16#00D67# => romdata <= X"FC9F3879";
    when 16#00D68# => romdata <= X"1470337C";
    when 16#00D69# => romdata <= X"075256F5";
    when 16#00D6A# => romdata <= X"E73F7714";
    when 16#00D6B# => romdata <= X"982B7098";
    when 16#00D6C# => romdata <= X"2C555976";
    when 16#00D6D# => romdata <= X"7424CE38";
    when 16#00D6E# => romdata <= X"FC83397D";
    when 16#00D6F# => romdata <= X"802E80F0";
    when 16#00D70# => romdata <= X"38791470";
    when 16#00D71# => romdata <= X"33705854";
    when 16#00D72# => romdata <= X"55805578";
    when 16#00D73# => romdata <= X"752E8538";
    when 16#00D74# => romdata <= X"72842A56";
    when 16#00D75# => romdata <= X"75832A70";
    when 16#00D76# => romdata <= X"81065153";
    when 16#00D77# => romdata <= X"72802E84";
    when 16#00D78# => romdata <= X"3881C055";
    when 16#00D79# => romdata <= X"75822A70";
    when 16#00D7A# => romdata <= X"81065153";
    when 16#00D7B# => romdata <= X"72802E85";
    when 16#00D7C# => romdata <= X"3874B007";
    when 16#00D7D# => romdata <= X"5575812A";
    when 16#00D7E# => romdata <= X"70810651";
    when 16#00D7F# => romdata <= X"5372802E";
    when 16#00D80# => romdata <= X"8538748C";
    when 16#00D81# => romdata <= X"07557581";
    when 16#00D82# => romdata <= X"06537280";
    when 16#00D83# => romdata <= X"2E853874";
    when 16#00D84# => romdata <= X"83075574";
    when 16#00D85# => romdata <= X"097081FF";
    when 16#00D86# => romdata <= X"065253F4";
    when 16#00D87# => romdata <= X"F33F7714";
    when 16#00D88# => romdata <= X"982B7098";
    when 16#00D89# => romdata <= X"2C555676";
    when 16#00D8A# => romdata <= X"7424FF95";
    when 16#00D8B# => romdata <= X"38FB8E39";
    when 16#00D8C# => romdata <= X"79147033";
    when 16#00D8D# => romdata <= X"70097081";
    when 16#00D8E# => romdata <= X"FF065458";
    when 16#00D8F# => romdata <= X"5455F4D0";
    when 16#00D90# => romdata <= X"3F771498";
    when 16#00D91# => romdata <= X"2B70982C";
    when 16#00D92# => romdata <= X"55597377";
    when 16#00D93# => romdata <= X"25FAEE38";
    when 16#00D94# => romdata <= X"79147033";
    when 16#00D95# => romdata <= X"70097081";
    when 16#00D96# => romdata <= X"FF065458";
    when 16#00D97# => romdata <= X"5455F4B0";
    when 16#00D98# => romdata <= X"3F771498";
    when 16#00D99# => romdata <= X"2B70982C";
    when 16#00D9A# => romdata <= X"55597674";
    when 16#00D9B# => romdata <= X"24C238FA";
    when 16#00D9C# => romdata <= X"CC396180";
    when 16#00D9D# => romdata <= X"2E81CE38";
    when 16#00D9E# => romdata <= X"7D802E80";
    when 16#00D9F# => romdata <= X"F7387914";
    when 16#00DA0# => romdata <= X"70337058";
    when 16#00DA1# => romdata <= X"54558055";
    when 16#00DA2# => romdata <= X"78752E85";
    when 16#00DA3# => romdata <= X"3872842A";
    when 16#00DA4# => romdata <= X"5675832A";
    when 16#00DA5# => romdata <= X"70810651";
    when 16#00DA6# => romdata <= X"5372802E";
    when 16#00DA7# => romdata <= X"843881C0";
    when 16#00DA8# => romdata <= X"5575822A";
    when 16#00DA9# => romdata <= X"70810651";
    when 16#00DAA# => romdata <= X"5372802E";
    when 16#00DAB# => romdata <= X"853874B0";
    when 16#00DAC# => romdata <= X"07557581";
    when 16#00DAD# => romdata <= X"2A708106";
    when 16#00DAE# => romdata <= X"51537280";
    when 16#00DAF# => romdata <= X"2E853874";
    when 16#00DB0# => romdata <= X"8C075575";
    when 16#00DB1# => romdata <= X"81065372";
    when 16#00DB2# => romdata <= X"802E8538";
    when 16#00DB3# => romdata <= X"74830755";
    when 16#00DB4# => romdata <= X"74097081";
    when 16#00DB5# => romdata <= X"FF067053";
    when 16#00DB6# => romdata <= X"5753F3B4";
    when 16#00DB7# => romdata <= X"3F7551F3";
    when 16#00DB8# => romdata <= X"AF3F7714";
    when 16#00DB9# => romdata <= X"982B7098";
    when 16#00DBA# => romdata <= X"2C555576";
    when 16#00DBB# => romdata <= X"7424FF8E";
    when 16#00DBC# => romdata <= X"38F9CA39";
    when 16#00DBD# => romdata <= X"79147033";
    when 16#00DBE# => romdata <= X"70097081";
    when 16#00DBF# => romdata <= X"FF067055";
    when 16#00DC0# => romdata <= X"59555659";
    when 16#00DC1# => romdata <= X"F38A3F75";
    when 16#00DC2# => romdata <= X"51F3853F";
    when 16#00DC3# => romdata <= X"7714982B";
    when 16#00DC4# => romdata <= X"70982C55";
    when 16#00DC5# => romdata <= X"59737725";
    when 16#00DC6# => romdata <= X"F9A33879";
    when 16#00DC7# => romdata <= X"14703370";
    when 16#00DC8# => romdata <= X"097081FF";
    when 16#00DC9# => romdata <= X"06705559";
    when 16#00DCA# => romdata <= X"555659F2";
    when 16#00DCB# => romdata <= X"E33F7551";
    when 16#00DCC# => romdata <= X"F2DE3F77";
    when 16#00DCD# => romdata <= X"14982B70";
    when 16#00DCE# => romdata <= X"982C5559";
    when 16#00DCF# => romdata <= X"767424FF";
    when 16#00DD0# => romdata <= X"B338F8F9";
    when 16#00DD1# => romdata <= X"397D802E";
    when 16#00DD2# => romdata <= X"80F43879";
    when 16#00DD3# => romdata <= X"14703370";
    when 16#00DD4# => romdata <= X"58545580";
    when 16#00DD5# => romdata <= X"5578752E";
    when 16#00DD6# => romdata <= X"85387284";
    when 16#00DD7# => romdata <= X"2A567583";
    when 16#00DD8# => romdata <= X"2A708106";
    when 16#00DD9# => romdata <= X"51537280";
    when 16#00DDA# => romdata <= X"2E843881";
    when 16#00DDB# => romdata <= X"C0557582";
    when 16#00DDC# => romdata <= X"2A708106";
    when 16#00DDD# => romdata <= X"51537280";
    when 16#00DDE# => romdata <= X"2E853874";
    when 16#00DDF# => romdata <= X"B0075575";
    when 16#00DE0# => romdata <= X"812A7081";
    when 16#00DE1# => romdata <= X"06515372";
    when 16#00DE2# => romdata <= X"802E8538";
    when 16#00DE3# => romdata <= X"748C0755";
    when 16#00DE4# => romdata <= X"75810653";
    when 16#00DE5# => romdata <= X"72802E85";
    when 16#00DE6# => romdata <= X"38748307";
    when 16#00DE7# => romdata <= X"557481FF";
    when 16#00DE8# => romdata <= X"06705256";
    when 16#00DE9# => romdata <= X"F1EA3F75";
    when 16#00DEA# => romdata <= X"51F1E53F";
    when 16#00DEB# => romdata <= X"7714982B";
    when 16#00DEC# => romdata <= X"70982C55";
    when 16#00DED# => romdata <= X"55767424";
    when 16#00DEE# => romdata <= X"FF9138F8";
    when 16#00DEF# => romdata <= X"80397914";
    when 16#00DF0# => romdata <= X"70337053";
    when 16#00DF1# => romdata <= X"5753F1C8";
    when 16#00DF2# => romdata <= X"3F7551F1";
    when 16#00DF3# => romdata <= X"C33F7714";
    when 16#00DF4# => romdata <= X"982B7098";
    when 16#00DF5# => romdata <= X"2C555973";
    when 16#00DF6# => romdata <= X"7725F7E1";
    when 16#00DF7# => romdata <= X"38791470";
    when 16#00DF8# => romdata <= X"33705357";
    when 16#00DF9# => romdata <= X"53F1A93F";
    when 16#00DFA# => romdata <= X"7551F1A4";
    when 16#00DFB# => romdata <= X"3F771498";
    when 16#00DFC# => romdata <= X"2B70982C";
    when 16#00DFD# => romdata <= X"55597674";
    when 16#00DFE# => romdata <= X"24C438F7";
    when 16#00DFF# => romdata <= X"C0397D80";
    when 16#00E00# => romdata <= X"2E80F238";
    when 16#00E01# => romdata <= X"79147033";
    when 16#00E02# => romdata <= X"7C077052";
    when 16#00E03# => romdata <= X"54568055";
    when 16#00E04# => romdata <= X"78752E85";
    when 16#00E05# => romdata <= X"3872842A";
    when 16#00E06# => romdata <= X"5675832A";
    when 16#00E07# => romdata <= X"70810651";
    when 16#00E08# => romdata <= X"5372802E";
    when 16#00E09# => romdata <= X"843881C0";
    when 16#00E0A# => romdata <= X"5575822A";
    when 16#00E0B# => romdata <= X"70810651";
    when 16#00E0C# => romdata <= X"5372802E";
    when 16#00E0D# => romdata <= X"853874B0";
    when 16#00E0E# => romdata <= X"07557581";
    when 16#00E0F# => romdata <= X"2A708106";
    when 16#00E10# => romdata <= X"51537280";
    when 16#00E11# => romdata <= X"2E853874";
    when 16#00E12# => romdata <= X"8C075575";
    when 16#00E13# => romdata <= X"81065372";
    when 16#00E14# => romdata <= X"802E8538";
    when 16#00E15# => romdata <= X"74830755";
    when 16#00E16# => romdata <= X"74097081";
    when 16#00E17# => romdata <= X"FF065256";
    when 16#00E18# => romdata <= X"F0AE3F77";
    when 16#00E19# => romdata <= X"14982B70";
    when 16#00E1A# => romdata <= X"982C5553";
    when 16#00E1B# => romdata <= X"767424FF";
    when 16#00E1C# => romdata <= X"9338F6C9";
    when 16#00E1D# => romdata <= X"39791470";
    when 16#00E1E# => romdata <= X"337C0770";
    when 16#00E1F# => romdata <= X"097081FF";
    when 16#00E20# => romdata <= X"06545556";
    when 16#00E21# => romdata <= X"59F0893F";
    when 16#00E22# => romdata <= X"7714982B";
    when 16#00E23# => romdata <= X"70982C55";
    when 16#00E24# => romdata <= X"59737725";
    when 16#00E25# => romdata <= X"F6A73879";
    when 16#00E26# => romdata <= X"1470337C";
    when 16#00E27# => romdata <= X"07700970";
    when 16#00E28# => romdata <= X"81FF0654";
    when 16#00E29# => romdata <= X"555659EF";
    when 16#00E2A# => romdata <= X"E73F7714";
    when 16#00E2B# => romdata <= X"982B7098";
    when 16#00E2C# => romdata <= X"2C555976";
    when 16#00E2D# => romdata <= X"7424FFBD";
    when 16#00E2E# => romdata <= X"38F68239";
    when 16#00E2F# => romdata <= X"61802E81";
    when 16#00E30# => romdata <= X"D4387D80";
    when 16#00E31# => romdata <= X"2E80F938";
    when 16#00E32# => romdata <= X"79147033";
    when 16#00E33# => romdata <= X"7C077052";
    when 16#00E34# => romdata <= X"54568055";
    when 16#00E35# => romdata <= X"78752E85";
    when 16#00E36# => romdata <= X"3872842A";
    when 16#00E37# => romdata <= X"5675832A";
    when 16#00E38# => romdata <= X"70810651";
    when 16#00E39# => romdata <= X"5372802E";
    when 16#00E3A# => romdata <= X"843881C0";
    when 16#00E3B# => romdata <= X"5575822A";
    when 16#00E3C# => romdata <= X"70810651";
    when 16#00E3D# => romdata <= X"5372802E";
    when 16#00E3E# => romdata <= X"853874B0";
    when 16#00E3F# => romdata <= X"07557581";
    when 16#00E40# => romdata <= X"2A708106";
    when 16#00E41# => romdata <= X"51537280";
    when 16#00E42# => romdata <= X"2E853874";
    when 16#00E43# => romdata <= X"8C075575";
    when 16#00E44# => romdata <= X"81065372";
    when 16#00E45# => romdata <= X"802E8538";
    when 16#00E46# => romdata <= X"74830755";
    when 16#00E47# => romdata <= X"74097081";
    when 16#00E48# => romdata <= X"FF067053";
    when 16#00E49# => romdata <= X"5456EEE8";
    when 16#00E4A# => romdata <= X"3F7251EE";
    when 16#00E4B# => romdata <= X"E33F7714";
    when 16#00E4C# => romdata <= X"982B7098";
    when 16#00E4D# => romdata <= X"2C555676";
    when 16#00E4E# => romdata <= X"7424FF8C";
    when 16#00E4F# => romdata <= X"38F4FE39";
    when 16#00E50# => romdata <= X"79147033";
    when 16#00E51# => romdata <= X"7C077009";
    when 16#00E52# => romdata <= X"7081FF06";
    when 16#00E53# => romdata <= X"70555357";
    when 16#00E54# => romdata <= X"5753EEBC";
    when 16#00E55# => romdata <= X"3F7251EE";
    when 16#00E56# => romdata <= X"B73F7714";
    when 16#00E57# => romdata <= X"982B7098";
    when 16#00E58# => romdata <= X"2C555973";
    when 16#00E59# => romdata <= X"7725F4D5";
    when 16#00E5A# => romdata <= X"38791470";
    when 16#00E5B# => romdata <= X"337C0770";
    when 16#00E5C# => romdata <= X"097081FF";
    when 16#00E5D# => romdata <= X"06705553";
    when 16#00E5E# => romdata <= X"575753EE";
    when 16#00E5F# => romdata <= X"933F7251";
    when 16#00E60# => romdata <= X"EE8E3F77";
    when 16#00E61# => romdata <= X"14982B70";
    when 16#00E62# => romdata <= X"982C5559";
    when 16#00E63# => romdata <= X"767424FF";
    when 16#00E64# => romdata <= X"AF38F4A9";
    when 16#00E65# => romdata <= X"397D802E";
    when 16#00E66# => romdata <= X"80F63879";
    when 16#00E67# => romdata <= X"1470337C";
    when 16#00E68# => romdata <= X"07705254";
    when 16#00E69# => romdata <= X"56805578";
    when 16#00E6A# => romdata <= X"752E8538";
    when 16#00E6B# => romdata <= X"72842A56";
    when 16#00E6C# => romdata <= X"75832A70";
    when 16#00E6D# => romdata <= X"81065153";
    when 16#00E6E# => romdata <= X"72802E84";
    when 16#00E6F# => romdata <= X"3881C055";
    when 16#00E70# => romdata <= X"75822A70";
    when 16#00E71# => romdata <= X"81065153";
    when 16#00E72# => romdata <= X"72802E85";
    when 16#00E73# => romdata <= X"3874B007";
    when 16#00E74# => romdata <= X"5575812A";
    when 16#00E75# => romdata <= X"70810651";
    when 16#00E76# => romdata <= X"5372802E";
    when 16#00E77# => romdata <= X"8538748C";
    when 16#00E78# => romdata <= X"07557581";
    when 16#00E79# => romdata <= X"06537280";
    when 16#00E7A# => romdata <= X"2E853874";
    when 16#00E7B# => romdata <= X"83075574";
    when 16#00E7C# => romdata <= X"81FF0670";
    when 16#00E7D# => romdata <= X"5256ED98";
    when 16#00E7E# => romdata <= X"3F7551ED";
    when 16#00E7F# => romdata <= X"933F7714";
    when 16#00E80# => romdata <= X"982B7098";
    when 16#00E81# => romdata <= X"2C555376";
    when 16#00E82# => romdata <= X"7424FF8F";
    when 16#00E83# => romdata <= X"38F3AE39";
    when 16#00E84# => romdata <= X"79147033";
    when 16#00E85# => romdata <= X"7C077053";
    when 16#00E86# => romdata <= X"5456ECF4";
    when 16#00E87# => romdata <= X"3F7251EC";
    when 16#00E88# => romdata <= X"EF3F7714";
    when 16#00E89# => romdata <= X"982B7098";
    when 16#00E8A# => romdata <= X"2C555973";
    when 16#00E8B# => romdata <= X"7725F38D";
    when 16#00E8C# => romdata <= X"38791470";
    when 16#00E8D# => romdata <= X"337C0770";
    when 16#00E8E# => romdata <= X"535456EC";
    when 16#00E8F# => romdata <= X"D33F7251";
    when 16#00E90# => romdata <= X"ECCE3F77";
    when 16#00E91# => romdata <= X"14982B70";
    when 16#00E92# => romdata <= X"982C5559";
    when 16#00E93# => romdata <= X"767424C0";
    when 16#00E94# => romdata <= X"38F2EA39";
    when 16#00E95# => romdata <= X"F83D0D7A";
    when 16#00E96# => romdata <= X"7D028805";
    when 16#00E97# => romdata <= X"AF05335A";
    when 16#00E98# => romdata <= X"55598074";
    when 16#00E99# => romdata <= X"70810556";
    when 16#00E9A# => romdata <= X"33755856";
    when 16#00E9B# => romdata <= X"5774772E";
    when 16#00E9C# => romdata <= X"09810688";
    when 16#00E9D# => romdata <= X"3876B00C";
    when 16#00E9E# => romdata <= X"8A3D0D04";
    when 16#00E9F# => romdata <= X"74537752";
    when 16#00EA0# => romdata <= X"7851EF92";
    when 16#00EA1# => romdata <= X"3FB00881";
    when 16#00EA2# => romdata <= X"FF067705";
    when 16#00EA3# => romdata <= X"7083FFFF";
    when 16#00EA4# => romdata <= X"06777081";
    when 16#00EA5# => romdata <= X"05593352";
    when 16#00EA6# => romdata <= X"58557480";
    when 16#00EA7# => romdata <= X"2ED73874";
    when 16#00EA8# => romdata <= X"53775278";
    when 16#00EA9# => romdata <= X"51EEEF3F";
    when 16#00EAA# => romdata <= X"B00881FF";
    when 16#00EAB# => romdata <= X"06770570";
    when 16#00EAC# => romdata <= X"83FFFF06";
    when 16#00EAD# => romdata <= X"77708105";
    when 16#00EAE# => romdata <= X"59335258";
    when 16#00EAF# => romdata <= X"5574FFBC";
    when 16#00EB0# => romdata <= X"38FFB239";
    when 16#00EB1# => romdata <= X"FE3D0D02";
    when 16#00EB2# => romdata <= X"93053353";
    when 16#00EB3# => romdata <= X"81F2D033";
    when 16#00EB4# => romdata <= X"5281F2CC";
    when 16#00EB5# => romdata <= X"0851EEBE";
    when 16#00EB6# => romdata <= X"3FB00881";
    when 16#00EB7# => romdata <= X"FF06B00C";
    when 16#00EB8# => romdata <= X"843D0D04";
    when 16#00EB9# => romdata <= X"D0893F04";
    when 16#00EBA# => romdata <= X"FB3D0D77";
    when 16#00EBB# => romdata <= X"79555580";
    when 16#00EBC# => romdata <= X"56757524";
    when 16#00EBD# => romdata <= X"AB388074";
    when 16#00EBE# => romdata <= X"249D3880";
    when 16#00EBF# => romdata <= X"53735274";
    when 16#00EC0# => romdata <= X"5180E13F";
    when 16#00EC1# => romdata <= X"B0085475";
    when 16#00EC2# => romdata <= X"802E8538";
    when 16#00EC3# => romdata <= X"B0083054";
    when 16#00EC4# => romdata <= X"73B00C87";
    when 16#00EC5# => romdata <= X"3D0D0473";
    when 16#00EC6# => romdata <= X"30768132";
    when 16#00EC7# => romdata <= X"5754DC39";
    when 16#00EC8# => romdata <= X"74305581";
    when 16#00EC9# => romdata <= X"56738025";
    when 16#00ECA# => romdata <= X"D238EC39";
    when 16#00ECB# => romdata <= X"FA3D0D78";
    when 16#00ECC# => romdata <= X"7A575580";
    when 16#00ECD# => romdata <= X"57767524";
    when 16#00ECE# => romdata <= X"A438759F";
    when 16#00ECF# => romdata <= X"2C548153";
    when 16#00ED0# => romdata <= X"75743274";
    when 16#00ED1# => romdata <= X"31527451";
    when 16#00ED2# => romdata <= X"9B3FB008";
    when 16#00ED3# => romdata <= X"5476802E";
    when 16#00ED4# => romdata <= X"8538B008";
    when 16#00ED5# => romdata <= X"305473B0";
    when 16#00ED6# => romdata <= X"0C883D0D";
    when 16#00ED7# => romdata <= X"04743055";
    when 16#00ED8# => romdata <= X"8157D739";
    when 16#00ED9# => romdata <= X"FC3D0D76";
    when 16#00EDA# => romdata <= X"78535481";
    when 16#00EDB# => romdata <= X"53807473";
    when 16#00EDC# => romdata <= X"26525572";
    when 16#00EDD# => romdata <= X"802E9838";
    when 16#00EDE# => romdata <= X"70802EA9";
    when 16#00EDF# => romdata <= X"38807224";
    when 16#00EE0# => romdata <= X"A4387110";
    when 16#00EE1# => romdata <= X"73107572";
    when 16#00EE2# => romdata <= X"26535452";
    when 16#00EE3# => romdata <= X"72EA3873";
    when 16#00EE4# => romdata <= X"51788338";
    when 16#00EE5# => romdata <= X"745170B0";
    when 16#00EE6# => romdata <= X"0C863D0D";
    when 16#00EE7# => romdata <= X"0472812A";
    when 16#00EE8# => romdata <= X"72812A53";
    when 16#00EE9# => romdata <= X"5372802E";
    when 16#00EEA# => romdata <= X"E6387174";
    when 16#00EEB# => romdata <= X"26EF3873";
    when 16#00EEC# => romdata <= X"72317574";
    when 16#00EED# => romdata <= X"0774812A";
    when 16#00EEE# => romdata <= X"74812A55";
    when 16#00EEF# => romdata <= X"555654E5";
    when 16#00EF0# => romdata <= X"39101010";
    when 16#00EF1# => romdata <= X"10101010";
    when 16#00EF2# => romdata <= X"10101010";
    when 16#00EF3# => romdata <= X"10101010";
    when 16#00EF4# => romdata <= X"10101010";
    when 16#00EF5# => romdata <= X"10101010";
    when 16#00EF6# => romdata <= X"10101010";
    when 16#00EF7# => romdata <= X"10101010";
    when 16#00EF8# => romdata <= X"53510473";
    when 16#00EF9# => romdata <= X"81FF0673";
    when 16#00EFA# => romdata <= X"83060981";
    when 16#00EFB# => romdata <= X"05830510";
    when 16#00EFC# => romdata <= X"10102B07";
    when 16#00EFD# => romdata <= X"72FC060C";
    when 16#00EFE# => romdata <= X"5151043C";
    when 16#00EFF# => romdata <= X"04727280";
    when 16#00F00# => romdata <= X"728106FF";
    when 16#00F01# => romdata <= X"05097206";
    when 16#00F02# => romdata <= X"05711052";
    when 16#00F03# => romdata <= X"720A100A";
    when 16#00F04# => romdata <= X"5372ED38";
    when 16#00F05# => romdata <= X"51515351";
    when 16#00F06# => romdata <= X"04B008B4";
    when 16#00F07# => romdata <= X"08B80875";
    when 16#00F08# => romdata <= X"7580F6AC";
    when 16#00F09# => romdata <= X"2D5050B0";
    when 16#00F0A# => romdata <= X"0856B80C";
    when 16#00F0B# => romdata <= X"B40CB00C";
    when 16#00F0C# => romdata <= X"5104B008";
    when 16#00F0D# => romdata <= X"B408B808";
    when 16#00F0E# => romdata <= X"757580F5";
    when 16#00F0F# => romdata <= X"E82D5050";
    when 16#00F10# => romdata <= X"B00856B8";
    when 16#00F11# => romdata <= X"0CB40CB0";
    when 16#00F12# => romdata <= X"0C5104B0";
    when 16#00F13# => romdata <= X"08B408B8";
    when 16#00F14# => romdata <= X"0880C5C6";
    when 16#00F15# => romdata <= X"2DB80CB4";
    when 16#00F16# => romdata <= X"0CB00C04";
    when 16#00F17# => romdata <= X"FF3D0D02";
    when 16#00F18# => romdata <= X"8F053381";
    when 16#00F19# => romdata <= X"CF840852";
    when 16#00F1A# => romdata <= X"710C800B";
    when 16#00F1B# => romdata <= X"B00C833D";
    when 16#00F1C# => romdata <= X"0D04FF3D";
    when 16#00F1D# => romdata <= X"0D028F05";
    when 16#00F1E# => romdata <= X"335181F2";
    when 16#00F1F# => romdata <= X"D4085271";
    when 16#00F20# => romdata <= X"2DB00881";
    when 16#00F21# => romdata <= X"FF06B00C";
    when 16#00F22# => romdata <= X"833D0D04";
    when 16#00F23# => romdata <= X"FE3D0D74";
    when 16#00F24# => romdata <= X"70335353";
    when 16#00F25# => romdata <= X"71802E93";
    when 16#00F26# => romdata <= X"38811372";
    when 16#00F27# => romdata <= X"5281F2D4";
    when 16#00F28# => romdata <= X"08535371";
    when 16#00F29# => romdata <= X"2D723352";
    when 16#00F2A# => romdata <= X"71EF3884";
    when 16#00F2B# => romdata <= X"3D0D04F4";
    when 16#00F2C# => romdata <= X"3D0D7F02";
    when 16#00F2D# => romdata <= X"8405BB05";
    when 16#00F2E# => romdata <= X"33555788";
    when 16#00F2F# => romdata <= X"0B8C3D5B";
    when 16#00F30# => romdata <= X"59895381";
    when 16#00F31# => romdata <= X"CC9C5279";
    when 16#00F32# => romdata <= X"5186B63F";
    when 16#00F33# => romdata <= X"73792E80";
    when 16#00F34# => romdata <= X"FF387856";
    when 16#00F35# => romdata <= X"73902E80";
    when 16#00F36# => romdata <= X"EC3802A7";
    when 16#00F37# => romdata <= X"0558768F";
    when 16#00F38# => romdata <= X"06547389";
    when 16#00F39# => romdata <= X"2680C238";
    when 16#00F3A# => romdata <= X"7518B015";
    when 16#00F3B# => romdata <= X"55557375";
    when 16#00F3C# => romdata <= X"3476842A";
    when 16#00F3D# => romdata <= X"FF177081";
    when 16#00F3E# => romdata <= X"FF065855";
    when 16#00F3F# => romdata <= X"5775DF38";
    when 16#00F40# => romdata <= X"781A5575";
    when 16#00F41# => romdata <= X"75347970";
    when 16#00F42# => romdata <= X"33555573";
    when 16#00F43# => romdata <= X"802E9338";
    when 16#00F44# => romdata <= X"81157452";
    when 16#00F45# => romdata <= X"81F2D408";
    when 16#00F46# => romdata <= X"5755752D";
    when 16#00F47# => romdata <= X"74335473";
    when 16#00F48# => romdata <= X"EF3878B0";
    when 16#00F49# => romdata <= X"0C8E3D0D";
    when 16#00F4A# => romdata <= X"047518B7";
    when 16#00F4B# => romdata <= X"15555573";
    when 16#00F4C# => romdata <= X"75347684";
    when 16#00F4D# => romdata <= X"2AFF1770";
    when 16#00F4E# => romdata <= X"81FF0658";
    when 16#00F4F# => romdata <= X"555775FF";
    when 16#00F50# => romdata <= X"9D38FFBC";
    when 16#00F51# => romdata <= X"39847057";
    when 16#00F52# => romdata <= X"5902A705";
    when 16#00F53# => romdata <= X"58FF8F39";
    when 16#00F54# => romdata <= X"82705759";
    when 16#00F55# => romdata <= X"F439F13D";
    when 16#00F56# => romdata <= X"0D618D3D";
    when 16#00F57# => romdata <= X"705B5C5A";
    when 16#00F58# => romdata <= X"807A5657";
    when 16#00F59# => romdata <= X"767A2481";
    when 16#00F5A# => romdata <= X"85387817";
    when 16#00F5B# => romdata <= X"548A5274";
    when 16#00F5C# => romdata <= X"5184DC3F";
    when 16#00F5D# => romdata <= X"B008B005";
    when 16#00F5E# => romdata <= X"53727434";
    when 16#00F5F# => romdata <= X"8117578A";
    when 16#00F60# => romdata <= X"52745184";
    when 16#00F61# => romdata <= X"A53FB008";
    when 16#00F62# => romdata <= X"55B008DE";
    when 16#00F63# => romdata <= X"38B00877";
    when 16#00F64# => romdata <= X"9F2A1870";
    when 16#00F65# => romdata <= X"812C5A56";
    when 16#00F66# => romdata <= X"56807825";
    when 16#00F67# => romdata <= X"9E387817";
    when 16#00F68# => romdata <= X"FF055575";
    when 16#00F69# => romdata <= X"19703355";
    when 16#00F6A# => romdata <= X"53743373";
    when 16#00F6B# => romdata <= X"34737534";
    when 16#00F6C# => romdata <= X"8116FF16";
    when 16#00F6D# => romdata <= X"56567776";
    when 16#00F6E# => romdata <= X"24E93876";
    when 16#00F6F# => romdata <= X"19588078";
    when 16#00F70# => romdata <= X"34807A24";
    when 16#00F71# => romdata <= X"177081FF";
    when 16#00F72# => romdata <= X"067C7033";
    when 16#00F73# => romdata <= X"56575556";
    when 16#00F74# => romdata <= X"72802E93";
    when 16#00F75# => romdata <= X"38811573";
    when 16#00F76# => romdata <= X"5281F2D4";
    when 16#00F77# => romdata <= X"08585576";
    when 16#00F78# => romdata <= X"2D743353";
    when 16#00F79# => romdata <= X"72EF3873";
    when 16#00F7A# => romdata <= X"B00C913D";
    when 16#00F7B# => romdata <= X"0D04AD7B";
    when 16#00F7C# => romdata <= X"3402AD05";
    when 16#00F7D# => romdata <= X"7A307119";
    when 16#00F7E# => romdata <= X"5656598A";
    when 16#00F7F# => romdata <= X"52745183";
    when 16#00F80# => romdata <= X"CE3FB008";
    when 16#00F81# => romdata <= X"B0055372";
    when 16#00F82# => romdata <= X"74348117";
    when 16#00F83# => romdata <= X"578A5274";
    when 16#00F84# => romdata <= X"5183973F";
    when 16#00F85# => romdata <= X"B00855B0";
    when 16#00F86# => romdata <= X"08FECF38";
    when 16#00F87# => romdata <= X"FEEF39FD";
    when 16#00F88# => romdata <= X"3D0D81CE";
    when 16#00F89# => romdata <= X"F80876B2";
    when 16#00F8A# => romdata <= X"E4299412";
    when 16#00F8B# => romdata <= X"0C54850B";
    when 16#00F8C# => romdata <= X"98150C98";
    when 16#00F8D# => romdata <= X"14087081";
    when 16#00F8E# => romdata <= X"06515372";
    when 16#00F8F# => romdata <= X"F638853D";
    when 16#00F90# => romdata <= X"0D04803D";
    when 16#00F91# => romdata <= X"0D81CEF8";
    when 16#00F92# => romdata <= X"0851870B";
    when 16#00F93# => romdata <= X"84120CFF";
    when 16#00F94# => romdata <= X"0BA4120C";
    when 16#00F95# => romdata <= X"A70BA812";
    when 16#00F96# => romdata <= X"0CB2E40B";
    when 16#00F97# => romdata <= X"94120C87";
    when 16#00F98# => romdata <= X"0B98120C";
    when 16#00F99# => romdata <= X"823D0D04";
    when 16#00F9A# => romdata <= X"803D0D81";
    when 16#00F9B# => romdata <= X"CEFC0851";
    when 16#00F9C# => romdata <= X"B80B8C12";
    when 16#00F9D# => romdata <= X"0C830B88";
    when 16#00F9E# => romdata <= X"120C823D";
    when 16#00F9F# => romdata <= X"0D04803D";
    when 16#00FA0# => romdata <= X"0D81CEFC";
    when 16#00FA1# => romdata <= X"08841108";
    when 16#00FA2# => romdata <= X"8106B00C";
    when 16#00FA3# => romdata <= X"51823D0D";
    when 16#00FA4# => romdata <= X"04FF3D0D";
    when 16#00FA5# => romdata <= X"81CEFC08";
    when 16#00FA6# => romdata <= X"52841208";
    when 16#00FA7# => romdata <= X"70810651";
    when 16#00FA8# => romdata <= X"5170802E";
    when 16#00FA9# => romdata <= X"F4387108";
    when 16#00FAA# => romdata <= X"7081FF06";
    when 16#00FAB# => romdata <= X"B00C5183";
    when 16#00FAC# => romdata <= X"3D0D04FE";
    when 16#00FAD# => romdata <= X"3D0D0293";
    when 16#00FAE# => romdata <= X"05335372";
    when 16#00FAF# => romdata <= X"8A2E9C38";
    when 16#00FB0# => romdata <= X"81CEFC08";
    when 16#00FB1# => romdata <= X"52841208";
    when 16#00FB2# => romdata <= X"70892A70";
    when 16#00FB3# => romdata <= X"81065151";
    when 16#00FB4# => romdata <= X"5170F238";
    when 16#00FB5# => romdata <= X"72720C84";
    when 16#00FB6# => romdata <= X"3D0D0481";
    when 16#00FB7# => romdata <= X"CEFC0852";
    when 16#00FB8# => romdata <= X"84120870";
    when 16#00FB9# => romdata <= X"892A7081";
    when 16#00FBA# => romdata <= X"06515151";
    when 16#00FBB# => romdata <= X"70F2388D";
    when 16#00FBC# => romdata <= X"720C8412";
    when 16#00FBD# => romdata <= X"0870892A";
    when 16#00FBE# => romdata <= X"70810651";
    when 16#00FBF# => romdata <= X"515170C5";
    when 16#00FC0# => romdata <= X"38D23980";
    when 16#00FC1# => romdata <= X"3D0D81CE";
    when 16#00FC2# => romdata <= X"F0085180";
    when 16#00FC3# => romdata <= X"0B84120C";
    when 16#00FC4# => romdata <= X"83FE800B";
    when 16#00FC5# => romdata <= X"88120C80";
    when 16#00FC6# => romdata <= X"0B81F2D8";
    when 16#00FC7# => romdata <= X"34800B81";
    when 16#00FC8# => romdata <= X"F2DC3482";
    when 16#00FC9# => romdata <= X"3D0D04FA";
    when 16#00FCA# => romdata <= X"3D0D02A3";
    when 16#00FCB# => romdata <= X"053381CE";
    when 16#00FCC# => romdata <= X"F00881F2";
    when 16#00FCD# => romdata <= X"D8337081";
    when 16#00FCE# => romdata <= X"FF067010";
    when 16#00FCF# => romdata <= X"101181F2";
    when 16#00FD0# => romdata <= X"DC337081";
    when 16#00FD1# => romdata <= X"FF067290";
    when 16#00FD2# => romdata <= X"29117088";
    when 16#00FD3# => romdata <= X"2B780777";
    when 16#00FD4# => romdata <= X"0C535B5B";
    when 16#00FD5# => romdata <= X"55555954";
    when 16#00FD6# => romdata <= X"54738A2E";
    when 16#00FD7# => romdata <= X"98387480";
    when 16#00FD8# => romdata <= X"CF2E9238";
    when 16#00FD9# => romdata <= X"738C2EA4";
    when 16#00FDA# => romdata <= X"38811653";
    when 16#00FDB# => romdata <= X"7281F2DC";
    when 16#00FDC# => romdata <= X"34883D0D";
    when 16#00FDD# => romdata <= X"0471A326";
    when 16#00FDE# => romdata <= X"A3388117";
    when 16#00FDF# => romdata <= X"527181F2";
    when 16#00FE0# => romdata <= X"D834800B";
    when 16#00FE1# => romdata <= X"81F2DC34";
    when 16#00FE2# => romdata <= X"883D0D04";
    when 16#00FE3# => romdata <= X"80527188";
    when 16#00FE4# => romdata <= X"2B730C81";
    when 16#00FE5# => romdata <= X"12529790";
    when 16#00FE6# => romdata <= X"7226F338";
    when 16#00FE7# => romdata <= X"800B81F2";
    when 16#00FE8# => romdata <= X"D834800B";
    when 16#00FE9# => romdata <= X"81F2DC34";
    when 16#00FEA# => romdata <= X"DF39BC08";
    when 16#00FEB# => romdata <= X"02BC0CFD";
    when 16#00FEC# => romdata <= X"3D0D8053";
    when 16#00FED# => romdata <= X"BC088C05";
    when 16#00FEE# => romdata <= X"0852BC08";
    when 16#00FEF# => romdata <= X"88050851";
    when 16#00FF0# => romdata <= X"F7A23FB0";
    when 16#00FF1# => romdata <= X"0870B00C";
    when 16#00FF2# => romdata <= X"54853D0D";
    when 16#00FF3# => romdata <= X"BC0C04BC";
    when 16#00FF4# => romdata <= X"0802BC0C";
    when 16#00FF5# => romdata <= X"FD3D0D81";
    when 16#00FF6# => romdata <= X"53BC088C";
    when 16#00FF7# => romdata <= X"050852BC";
    when 16#00FF8# => romdata <= X"08880508";
    when 16#00FF9# => romdata <= X"51F6FD3F";
    when 16#00FFA# => romdata <= X"B00870B0";
    when 16#00FFB# => romdata <= X"0C54853D";
    when 16#00FFC# => romdata <= X"0DBC0C04";
    when 16#00FFD# => romdata <= X"803D0D86";
    when 16#00FFE# => romdata <= X"5184963F";
    when 16#00FFF# => romdata <= X"8151A1D3";
    when 16#01000# => romdata <= X"3FFC3D0D";
    when 16#01001# => romdata <= X"7670797B";
    when 16#01002# => romdata <= X"55555555";
    when 16#01003# => romdata <= X"8F72278C";
    when 16#01004# => romdata <= X"38727507";
    when 16#01005# => romdata <= X"83065170";
    when 16#01006# => romdata <= X"802EA738";
    when 16#01007# => romdata <= X"FF125271";
    when 16#01008# => romdata <= X"FF2E9838";
    when 16#01009# => romdata <= X"72708105";
    when 16#0100A# => romdata <= X"54337470";
    when 16#0100B# => romdata <= X"81055634";
    when 16#0100C# => romdata <= X"FF125271";
    when 16#0100D# => romdata <= X"FF2E0981";
    when 16#0100E# => romdata <= X"06EA3874";
    when 16#0100F# => romdata <= X"B00C863D";
    when 16#01010# => romdata <= X"0D047451";
    when 16#01011# => romdata <= X"72708405";
    when 16#01012# => romdata <= X"54087170";
    when 16#01013# => romdata <= X"8405530C";
    when 16#01014# => romdata <= X"72708405";
    when 16#01015# => romdata <= X"54087170";
    when 16#01016# => romdata <= X"8405530C";
    when 16#01017# => romdata <= X"72708405";
    when 16#01018# => romdata <= X"54087170";
    when 16#01019# => romdata <= X"8405530C";
    when 16#0101A# => romdata <= X"72708405";
    when 16#0101B# => romdata <= X"54087170";
    when 16#0101C# => romdata <= X"8405530C";
    when 16#0101D# => romdata <= X"F0125271";
    when 16#0101E# => romdata <= X"8F26C938";
    when 16#0101F# => romdata <= X"83722795";
    when 16#01020# => romdata <= X"38727084";
    when 16#01021# => romdata <= X"05540871";
    when 16#01022# => romdata <= X"70840553";
    when 16#01023# => romdata <= X"0CFC1252";
    when 16#01024# => romdata <= X"718326ED";
    when 16#01025# => romdata <= X"387054FF";
    when 16#01026# => romdata <= X"8339FD3D";
    when 16#01027# => romdata <= X"0D755384";
    when 16#01028# => romdata <= X"D8130880";
    when 16#01029# => romdata <= X"2E8A3880";
    when 16#0102A# => romdata <= X"5372B00C";
    when 16#0102B# => romdata <= X"853D0D04";
    when 16#0102C# => romdata <= X"81805272";
    when 16#0102D# => romdata <= X"518D9B3F";
    when 16#0102E# => romdata <= X"B00884D8";
    when 16#0102F# => romdata <= X"140CFF53";
    when 16#01030# => romdata <= X"B008802E";
    when 16#01031# => romdata <= X"E438B008";
    when 16#01032# => romdata <= X"549F5380";
    when 16#01033# => romdata <= X"74708405";
    when 16#01034# => romdata <= X"560CFF13";
    when 16#01035# => romdata <= X"53807324";
    when 16#01036# => romdata <= X"CE388074";
    when 16#01037# => romdata <= X"70840556";
    when 16#01038# => romdata <= X"0CFF1353";
    when 16#01039# => romdata <= X"728025E3";
    when 16#0103A# => romdata <= X"38FFBC39";
    when 16#0103B# => romdata <= X"FD3D0D75";
    when 16#0103C# => romdata <= X"7755539F";
    when 16#0103D# => romdata <= X"74278D38";
    when 16#0103E# => romdata <= X"96730CFF";
    when 16#0103F# => romdata <= X"5271B00C";
    when 16#01040# => romdata <= X"853D0D04";
    when 16#01041# => romdata <= X"84D81308";
    when 16#01042# => romdata <= X"5271802E";
    when 16#01043# => romdata <= X"93387310";
    when 16#01044# => romdata <= X"10127008";
    when 16#01045# => romdata <= X"79720C51";
    when 16#01046# => romdata <= X"5271B00C";
    when 16#01047# => romdata <= X"853D0D04";
    when 16#01048# => romdata <= X"7251FEF6";
    when 16#01049# => romdata <= X"3FFF52B0";
    when 16#0104A# => romdata <= X"08D33884";
    when 16#0104B# => romdata <= X"D8130874";
    when 16#0104C# => romdata <= X"10101170";
    when 16#0104D# => romdata <= X"087A720C";
    when 16#0104E# => romdata <= X"515152DD";
    when 16#0104F# => romdata <= X"39F93D0D";
    when 16#01050# => romdata <= X"797B5856";
    when 16#01051# => romdata <= X"769F2680";
    when 16#01052# => romdata <= X"E83884D8";
    when 16#01053# => romdata <= X"16085473";
    when 16#01054# => romdata <= X"802EAA38";
    when 16#01055# => romdata <= X"76101014";
    when 16#01056# => romdata <= X"70085555";
    when 16#01057# => romdata <= X"73802EBA";
    when 16#01058# => romdata <= X"38805873";
    when 16#01059# => romdata <= X"812E8F38";
    when 16#0105A# => romdata <= X"73FF2EA3";
    when 16#0105B# => romdata <= X"3880750C";
    when 16#0105C# => romdata <= X"7651732D";
    when 16#0105D# => romdata <= X"805877B0";
    when 16#0105E# => romdata <= X"0C893D0D";
    when 16#0105F# => romdata <= X"047551FE";
    when 16#01060# => romdata <= X"993FFF58";
    when 16#01061# => romdata <= X"B008EF38";
    when 16#01062# => romdata <= X"84D81608";
    when 16#01063# => romdata <= X"54C63996";
    when 16#01064# => romdata <= X"760C810B";
    when 16#01065# => romdata <= X"B00C893D";
    when 16#01066# => romdata <= X"0D047551";
    when 16#01067# => romdata <= X"81ED3F76";
    when 16#01068# => romdata <= X"53B00852";
    when 16#01069# => romdata <= X"755181AD";
    when 16#0106A# => romdata <= X"3FB008B0";
    when 16#0106B# => romdata <= X"0C893D0D";
    when 16#0106C# => romdata <= X"0496760C";
    when 16#0106D# => romdata <= X"FF0BB00C";
    when 16#0106E# => romdata <= X"893D0D04";
    when 16#0106F# => romdata <= X"FC3D0D76";
    when 16#01070# => romdata <= X"785653FF";
    when 16#01071# => romdata <= X"54749F26";
    when 16#01072# => romdata <= X"B13884D8";
    when 16#01073# => romdata <= X"13085271";
    when 16#01074# => romdata <= X"802EAE38";
    when 16#01075# => romdata <= X"74101012";
    when 16#01076# => romdata <= X"70085353";
    when 16#01077# => romdata <= X"81547180";
    when 16#01078# => romdata <= X"2E983882";
    when 16#01079# => romdata <= X"5471FF2E";
    when 16#0107A# => romdata <= X"91388354";
    when 16#0107B# => romdata <= X"71812E8A";
    when 16#0107C# => romdata <= X"3880730C";
    when 16#0107D# => romdata <= X"7451712D";
    when 16#0107E# => romdata <= X"805473B0";
    when 16#0107F# => romdata <= X"0C863D0D";
    when 16#01080# => romdata <= X"047251FD";
    when 16#01081# => romdata <= X"953FB008";
    when 16#01082# => romdata <= X"F13884D8";
    when 16#01083# => romdata <= X"130852C4";
    when 16#01084# => romdata <= X"39FF3D0D";
    when 16#01085# => romdata <= X"735281CF";
    when 16#01086# => romdata <= X"880851FE";
    when 16#01087# => romdata <= X"A03F833D";
    when 16#01088# => romdata <= X"0D04FE3D";
    when 16#01089# => romdata <= X"0D755374";
    when 16#0108A# => romdata <= X"5281CF88";
    when 16#0108B# => romdata <= X"0851FDBC";
    when 16#0108C# => romdata <= X"3F843D0D";
    when 16#0108D# => romdata <= X"04803D0D";
    when 16#0108E# => romdata <= X"81CF8808";
    when 16#0108F# => romdata <= X"51FCDB3F";
    when 16#01090# => romdata <= X"823D0D04";
    when 16#01091# => romdata <= X"FF3D0D73";
    when 16#01092# => romdata <= X"5281CF88";
    when 16#01093# => romdata <= X"0851FEEC";
    when 16#01094# => romdata <= X"3F833D0D";
    when 16#01095# => romdata <= X"04FC3D0D";
    when 16#01096# => romdata <= X"800B81F2";
    when 16#01097# => romdata <= X"E40C7852";
    when 16#01098# => romdata <= X"77519CAA";
    when 16#01099# => romdata <= X"3FB00854";
    when 16#0109A# => romdata <= X"B008FF2E";
    when 16#0109B# => romdata <= X"883873B0";
    when 16#0109C# => romdata <= X"0C863D0D";
    when 16#0109D# => romdata <= X"0481F2E4";
    when 16#0109E# => romdata <= X"08557480";
    when 16#0109F# => romdata <= X"2EF03876";
    when 16#010A0# => romdata <= X"75710C53";
    when 16#010A1# => romdata <= X"73B00C86";
    when 16#010A2# => romdata <= X"3D0D049B";
    when 16#010A3# => romdata <= X"FC3F04FC";
    when 16#010A4# => romdata <= X"3D0D7670";
    when 16#010A5# => romdata <= X"79707307";
    when 16#010A6# => romdata <= X"83065454";
    when 16#010A7# => romdata <= X"54557080";
    when 16#010A8# => romdata <= X"C3387170";
    when 16#010A9# => romdata <= X"08700970";
    when 16#010AA# => romdata <= X"F7FBFDFF";
    when 16#010AB# => romdata <= X"130670F8";
    when 16#010AC# => romdata <= X"84828180";
    when 16#010AD# => romdata <= X"06515153";
    when 16#010AE# => romdata <= X"535470A6";
    when 16#010AF# => romdata <= X"38841472";
    when 16#010B0# => romdata <= X"74708405";
    when 16#010B1# => romdata <= X"560C7008";
    when 16#010B2# => romdata <= X"700970F7";
    when 16#010B3# => romdata <= X"FBFDFF13";
    when 16#010B4# => romdata <= X"0670F884";
    when 16#010B5# => romdata <= X"82818006";
    when 16#010B6# => romdata <= X"51515353";
    when 16#010B7# => romdata <= X"5470802E";
    when 16#010B8# => romdata <= X"DC387352";
    when 16#010B9# => romdata <= X"71708105";
    when 16#010BA# => romdata <= X"53335170";
    when 16#010BB# => romdata <= X"73708105";
    when 16#010BC# => romdata <= X"553470F0";
    when 16#010BD# => romdata <= X"3874B00C";
    when 16#010BE# => romdata <= X"863D0D04";
    when 16#010BF# => romdata <= X"FD3D0D75";
    when 16#010C0# => romdata <= X"70718306";
    when 16#010C1# => romdata <= X"53555270";
    when 16#010C2# => romdata <= X"B8387170";
    when 16#010C3# => romdata <= X"087009F7";
    when 16#010C4# => romdata <= X"FBFDFF12";
    when 16#010C5# => romdata <= X"0670F884";
    when 16#010C6# => romdata <= X"82818006";
    when 16#010C7# => romdata <= X"51515253";
    when 16#010C8# => romdata <= X"709D3884";
    when 16#010C9# => romdata <= X"13700870";
    when 16#010CA# => romdata <= X"09F7FBFD";
    when 16#010CB# => romdata <= X"FF120670";
    when 16#010CC# => romdata <= X"F8848281";
    when 16#010CD# => romdata <= X"80065151";
    when 16#010CE# => romdata <= X"52537080";
    when 16#010CF# => romdata <= X"2EE53872";
    when 16#010D0# => romdata <= X"52713351";
    when 16#010D1# => romdata <= X"70802E8A";
    when 16#010D2# => romdata <= X"38811270";
    when 16#010D3# => romdata <= X"33525270";
    when 16#010D4# => romdata <= X"F8387174";
    when 16#010D5# => romdata <= X"31B00C85";
    when 16#010D6# => romdata <= X"3D0D04FA";
    when 16#010D7# => romdata <= X"3D0D787A";
    when 16#010D8# => romdata <= X"7C705455";
    when 16#010D9# => romdata <= X"55527280";
    when 16#010DA# => romdata <= X"2E80D938";
    when 16#010DB# => romdata <= X"71740783";
    when 16#010DC# => romdata <= X"06517080";
    when 16#010DD# => romdata <= X"2E80D438";
    when 16#010DE# => romdata <= X"FF135372";
    when 16#010DF# => romdata <= X"FF2EB138";
    when 16#010E0# => romdata <= X"71337433";
    when 16#010E1# => romdata <= X"56517471";
    when 16#010E2# => romdata <= X"2E098106";
    when 16#010E3# => romdata <= X"A9387280";
    when 16#010E4# => romdata <= X"2E818738";
    when 16#010E5# => romdata <= X"7081FF06";
    when 16#010E6# => romdata <= X"5170802E";
    when 16#010E7# => romdata <= X"80FC3881";
    when 16#010E8# => romdata <= X"128115FF";
    when 16#010E9# => romdata <= X"15555552";
    when 16#010EA# => romdata <= X"72FF2E09";
    when 16#010EB# => romdata <= X"8106D138";
    when 16#010EC# => romdata <= X"71337433";
    when 16#010ED# => romdata <= X"56517081";
    when 16#010EE# => romdata <= X"FF067581";
    when 16#010EF# => romdata <= X"FF067171";
    when 16#010F0# => romdata <= X"31515252";
    when 16#010F1# => romdata <= X"70B00C88";
    when 16#010F2# => romdata <= X"3D0D0471";
    when 16#010F3# => romdata <= X"74575583";
    when 16#010F4# => romdata <= X"73278838";
    when 16#010F5# => romdata <= X"71087408";
    when 16#010F6# => romdata <= X"2E883874";
    when 16#010F7# => romdata <= X"765552FF";
    when 16#010F8# => romdata <= X"9739FC13";
    when 16#010F9# => romdata <= X"5372802E";
    when 16#010FA# => romdata <= X"B1387408";
    when 16#010FB# => romdata <= X"7009F7FB";
    when 16#010FC# => romdata <= X"FDFF1206";
    when 16#010FD# => romdata <= X"70F88482";
    when 16#010FE# => romdata <= X"81800651";
    when 16#010FF# => romdata <= X"5151709A";
    when 16#01100# => romdata <= X"38841584";
    when 16#01101# => romdata <= X"17575583";
    when 16#01102# => romdata <= X"7327D038";
    when 16#01103# => romdata <= X"74087608";
    when 16#01104# => romdata <= X"2ED03874";
    when 16#01105# => romdata <= X"765552FE";
    when 16#01106# => romdata <= X"DF39800B";
    when 16#01107# => romdata <= X"B00C883D";
    when 16#01108# => romdata <= X"0D04F33D";
    when 16#01109# => romdata <= X"0D606264";
    when 16#0110A# => romdata <= X"725A5A5E";
    when 16#0110B# => romdata <= X"5E805C76";
    when 16#0110C# => romdata <= X"70810558";
    when 16#0110D# => romdata <= X"3381CCA9";
    when 16#0110E# => romdata <= X"11337083";
    when 16#0110F# => romdata <= X"2A708106";
    when 16#01110# => romdata <= X"51555556";
    when 16#01111# => romdata <= X"72E93875";
    when 16#01112# => romdata <= X"AD2E8288";
    when 16#01113# => romdata <= X"3875AB2E";
    when 16#01114# => romdata <= X"82843877";
    when 16#01115# => romdata <= X"30707907";
    when 16#01116# => romdata <= X"80257990";
    when 16#01117# => romdata <= X"32703070";
    when 16#01118# => romdata <= X"72078025";
    when 16#01119# => romdata <= X"73075357";
    when 16#0111A# => romdata <= X"57515372";
    when 16#0111B# => romdata <= X"802E8738";
    when 16#0111C# => romdata <= X"75B02E81";
    when 16#0111D# => romdata <= X"EB38778A";
    when 16#0111E# => romdata <= X"38885875";
    when 16#0111F# => romdata <= X"B02E8338";
    when 16#01120# => romdata <= X"8A58810A";
    when 16#01121# => romdata <= X"5A7B8438";
    when 16#01122# => romdata <= X"FE0A5A77";
    when 16#01123# => romdata <= X"527951F6";
    when 16#01124# => romdata <= X"BE3FB008";
    when 16#01125# => romdata <= X"78537A52";
    when 16#01126# => romdata <= X"5BF68F3F";
    when 16#01127# => romdata <= X"B0085A80";
    when 16#01128# => romdata <= X"7081CCA9";
    when 16#01129# => romdata <= X"18337082";
    when 16#0112A# => romdata <= X"2A708106";
    when 16#0112B# => romdata <= X"5156565A";
    when 16#0112C# => romdata <= X"5572802E";
    when 16#0112D# => romdata <= X"80C138D0";
    when 16#0112E# => romdata <= X"16567578";
    when 16#0112F# => romdata <= X"2580D738";
    when 16#01130# => romdata <= X"80792475";
    when 16#01131# => romdata <= X"7B260753";
    when 16#01132# => romdata <= X"72933874";
    when 16#01133# => romdata <= X"7A2E80EB";
    when 16#01134# => romdata <= X"387A7625";
    when 16#01135# => romdata <= X"80ED3872";
    when 16#01136# => romdata <= X"802E80E7";
    when 16#01137# => romdata <= X"38FF7770";
    when 16#01138# => romdata <= X"81055933";
    when 16#01139# => romdata <= X"575981CC";
    when 16#0113A# => romdata <= X"A9163370";
    when 16#0113B# => romdata <= X"822A7081";
    when 16#0113C# => romdata <= X"06515454";
    when 16#0113D# => romdata <= X"72C13873";
    when 16#0113E# => romdata <= X"83065372";
    when 16#0113F# => romdata <= X"802E9738";
    when 16#01140# => romdata <= X"738106C9";
    when 16#01141# => romdata <= X"17555372";
    when 16#01142# => romdata <= X"8538FFA9";
    when 16#01143# => romdata <= X"16547356";
    when 16#01144# => romdata <= X"777624FF";
    when 16#01145# => romdata <= X"AB388079";
    when 16#01146# => romdata <= X"2480F038";
    when 16#01147# => romdata <= X"7B802E84";
    when 16#01148# => romdata <= X"38743055";
    when 16#01149# => romdata <= X"7C802E8C";
    when 16#0114A# => romdata <= X"38FF1753";
    when 16#0114B# => romdata <= X"7883387D";
    when 16#0114C# => romdata <= X"53727D0C";
    when 16#0114D# => romdata <= X"74B00C8F";
    when 16#0114E# => romdata <= X"3D0D0481";
    when 16#0114F# => romdata <= X"53757B24";
    when 16#01150# => romdata <= X"FF953881";
    when 16#01151# => romdata <= X"75792917";
    when 16#01152# => romdata <= X"78708105";
    when 16#01153# => romdata <= X"5A335856";
    when 16#01154# => romdata <= X"59FF9339";
    when 16#01155# => romdata <= X"815C7670";
    when 16#01156# => romdata <= X"81055833";
    when 16#01157# => romdata <= X"56FDF439";
    when 16#01158# => romdata <= X"80773354";
    when 16#01159# => romdata <= X"547280F8";
    when 16#0115A# => romdata <= X"2EB23872";
    when 16#0115B# => romdata <= X"80D83270";
    when 16#0115C# => romdata <= X"30708025";
    when 16#0115D# => romdata <= X"76075151";
    when 16#0115E# => romdata <= X"5372802E";
    when 16#0115F# => romdata <= X"FDF83881";
    when 16#01160# => romdata <= X"17338218";
    when 16#01161# => romdata <= X"58569058";
    when 16#01162# => romdata <= X"FDF83981";
    when 16#01163# => romdata <= X"0A557B84";
    when 16#01164# => romdata <= X"38FE0A55";
    when 16#01165# => romdata <= X"7F53A273";
    when 16#01166# => romdata <= X"0CFF8939";
    when 16#01167# => romdata <= X"8154CC39";
    when 16#01168# => romdata <= X"FD3D0D77";
    when 16#01169# => romdata <= X"54765375";
    when 16#0116A# => romdata <= X"5281CF88";
    when 16#0116B# => romdata <= X"0851FCF2";
    when 16#0116C# => romdata <= X"3F853D0D";
    when 16#0116D# => romdata <= X"04F33D0D";
    when 16#0116E# => romdata <= X"60626472";
    when 16#0116F# => romdata <= X"5A5A5D5D";
    when 16#01170# => romdata <= X"805E7670";
    when 16#01171# => romdata <= X"81055833";
    when 16#01172# => romdata <= X"81CCA911";
    when 16#01173# => romdata <= X"3370832A";
    when 16#01174# => romdata <= X"70810651";
    when 16#01175# => romdata <= X"55555672";
    when 16#01176# => romdata <= X"E93875AD";
    when 16#01177# => romdata <= X"2E81FF38";
    when 16#01178# => romdata <= X"75AB2E81";
    when 16#01179# => romdata <= X"FB387730";
    when 16#0117A# => romdata <= X"70790780";
    when 16#0117B# => romdata <= X"25799032";
    when 16#0117C# => romdata <= X"70307072";
    when 16#0117D# => romdata <= X"07802573";
    when 16#0117E# => romdata <= X"07535757";
    when 16#0117F# => romdata <= X"51537280";
    when 16#01180# => romdata <= X"2E873875";
    when 16#01181# => romdata <= X"B02E81E2";
    when 16#01182# => romdata <= X"38778A38";
    when 16#01183# => romdata <= X"885875B0";
    when 16#01184# => romdata <= X"2E83388A";
    when 16#01185# => romdata <= X"587752FF";
    when 16#01186# => romdata <= X"51F38F3F";
    when 16#01187# => romdata <= X"B0087853";
    when 16#01188# => romdata <= X"5AFF51F3";
    when 16#01189# => romdata <= X"AA3FB008";
    when 16#0118A# => romdata <= X"5B80705A";
    when 16#0118B# => romdata <= X"5581CCA9";
    when 16#0118C# => romdata <= X"16337082";
    when 16#0118D# => romdata <= X"2A708106";
    when 16#0118E# => romdata <= X"51545472";
    when 16#0118F# => romdata <= X"802E80C1";
    when 16#01190# => romdata <= X"38D01656";
    when 16#01191# => romdata <= X"75782580";
    when 16#01192# => romdata <= X"D7388079";
    when 16#01193# => romdata <= X"24757B26";
    when 16#01194# => romdata <= X"07537293";
    when 16#01195# => romdata <= X"38747A2E";
    when 16#01196# => romdata <= X"80EB387A";
    when 16#01197# => romdata <= X"762580ED";
    when 16#01198# => romdata <= X"3872802E";
    when 16#01199# => romdata <= X"80E738FF";
    when 16#0119A# => romdata <= X"77708105";
    when 16#0119B# => romdata <= X"59335759";
    when 16#0119C# => romdata <= X"81CCA916";
    when 16#0119D# => romdata <= X"3370822A";
    when 16#0119E# => romdata <= X"70810651";
    when 16#0119F# => romdata <= X"545472C1";
    when 16#011A0# => romdata <= X"38738306";
    when 16#011A1# => romdata <= X"5372802E";
    when 16#011A2# => romdata <= X"97387381";
    when 16#011A3# => romdata <= X"06C91755";
    when 16#011A4# => romdata <= X"53728538";
    when 16#011A5# => romdata <= X"FFA91654";
    when 16#011A6# => romdata <= X"73567776";
    when 16#011A7# => romdata <= X"24FFAB38";
    when 16#011A8# => romdata <= X"80792481";
    when 16#011A9# => romdata <= X"89387D80";
    when 16#011AA# => romdata <= X"2E843874";
    when 16#011AB# => romdata <= X"30557B80";
    when 16#011AC# => romdata <= X"2E8C38FF";
    when 16#011AD# => romdata <= X"17537883";
    when 16#011AE# => romdata <= X"387C5372";
    when 16#011AF# => romdata <= X"7C0C74B0";
    when 16#011B0# => romdata <= X"0C8F3D0D";
    when 16#011B1# => romdata <= X"04815375";
    when 16#011B2# => romdata <= X"7B24FF95";
    when 16#011B3# => romdata <= X"38817579";
    when 16#011B4# => romdata <= X"29177870";
    when 16#011B5# => romdata <= X"81055A33";
    when 16#011B6# => romdata <= X"585659FF";
    when 16#011B7# => romdata <= X"9339815E";
    when 16#011B8# => romdata <= X"76708105";
    when 16#011B9# => romdata <= X"583356FD";
    when 16#011BA# => romdata <= X"FD398077";
    when 16#011BB# => romdata <= X"33545472";
    when 16#011BC# => romdata <= X"80F82E80";
    when 16#011BD# => romdata <= X"C3387280";
    when 16#011BE# => romdata <= X"D8327030";
    when 16#011BF# => romdata <= X"70802576";
    when 16#011C0# => romdata <= X"07515153";
    when 16#011C1# => romdata <= X"72802EFE";
    when 16#011C2# => romdata <= X"80388117";
    when 16#011C3# => romdata <= X"33821858";
    when 16#011C4# => romdata <= X"56907053";
    when 16#011C5# => romdata <= X"58FF51F1";
    when 16#011C6# => romdata <= X"913FB008";
    when 16#011C7# => romdata <= X"78535AFF";
    when 16#011C8# => romdata <= X"51F1AC3F";
    when 16#011C9# => romdata <= X"B0085B80";
    when 16#011CA# => romdata <= X"705A55FE";
    when 16#011CB# => romdata <= X"8039FF60";
    when 16#011CC# => romdata <= X"5455A273";
    when 16#011CD# => romdata <= X"0CFEF739";
    when 16#011CE# => romdata <= X"8154FFBA";
    when 16#011CF# => romdata <= X"39FD3D0D";
    when 16#011D0# => romdata <= X"77547653";
    when 16#011D1# => romdata <= X"755281CF";
    when 16#011D2# => romdata <= X"880851FC";
    when 16#011D3# => romdata <= X"E83F853D";
    when 16#011D4# => romdata <= X"0D04F33D";
    when 16#011D5# => romdata <= X"0D7F618B";
    when 16#011D6# => romdata <= X"1170F806";
    when 16#011D7# => romdata <= X"5C55555E";
    when 16#011D8# => romdata <= X"72962683";
    when 16#011D9# => romdata <= X"38905980";
    when 16#011DA# => romdata <= X"7924747A";
    when 16#011DB# => romdata <= X"26075380";
    when 16#011DC# => romdata <= X"5472742E";
    when 16#011DD# => romdata <= X"09810680";
    when 16#011DE# => romdata <= X"CB387D51";
    when 16#011DF# => romdata <= X"8BCA3F78";
    when 16#011E0# => romdata <= X"83F72680";
    when 16#011E1# => romdata <= X"C6387883";
    when 16#011E2# => romdata <= X"2A701010";
    when 16#011E3# => romdata <= X"1081D6C4";
    when 16#011E4# => romdata <= X"058C1108";
    when 16#011E5# => romdata <= X"59595A76";
    when 16#011E6# => romdata <= X"782E83B0";
    when 16#011E7# => romdata <= X"38841708";
    when 16#011E8# => romdata <= X"FC06568C";
    when 16#011E9# => romdata <= X"17088818";
    when 16#011EA# => romdata <= X"08718C12";
    when 16#011EB# => romdata <= X"0C88120C";
    when 16#011EC# => romdata <= X"58751784";
    when 16#011ED# => romdata <= X"11088107";
    when 16#011EE# => romdata <= X"84120C53";
    when 16#011EF# => romdata <= X"7D518B89";
    when 16#011F0# => romdata <= X"3F881754";
    when 16#011F1# => romdata <= X"73B00C8F";
    when 16#011F2# => romdata <= X"3D0D0478";
    when 16#011F3# => romdata <= X"892A7983";
    when 16#011F4# => romdata <= X"2A5B5372";
    when 16#011F5# => romdata <= X"802EBF38";
    when 16#011F6# => romdata <= X"78862AB8";
    when 16#011F7# => romdata <= X"055A8473";
    when 16#011F8# => romdata <= X"27B43880";
    when 16#011F9# => romdata <= X"DB135A94";
    when 16#011FA# => romdata <= X"7327AB38";
    when 16#011FB# => romdata <= X"788C2A80";
    when 16#011FC# => romdata <= X"EE055A80";
    when 16#011FD# => romdata <= X"D473279E";
    when 16#011FE# => romdata <= X"38788F2A";
    when 16#011FF# => romdata <= X"80F7055A";
    when 16#01200# => romdata <= X"82D47327";
    when 16#01201# => romdata <= X"91387892";
    when 16#01202# => romdata <= X"2A80FC05";
    when 16#01203# => romdata <= X"5A8AD473";
    when 16#01204# => romdata <= X"27843880";
    when 16#01205# => romdata <= X"FE5A7910";
    when 16#01206# => romdata <= X"101081D6";
    when 16#01207# => romdata <= X"C4058C11";
    when 16#01208# => romdata <= X"08585576";
    when 16#01209# => romdata <= X"752EA338";
    when 16#0120A# => romdata <= X"841708FC";
    when 16#0120B# => romdata <= X"06707A31";
    when 16#0120C# => romdata <= X"5556738F";
    when 16#0120D# => romdata <= X"2488D538";
    when 16#0120E# => romdata <= X"738025FE";
    when 16#0120F# => romdata <= X"E6388C17";
    when 16#01210# => romdata <= X"08577675";
    when 16#01211# => romdata <= X"2E098106";
    when 16#01212# => romdata <= X"DF38811A";
    when 16#01213# => romdata <= X"5A81D6D4";
    when 16#01214# => romdata <= X"08577681";
    when 16#01215# => romdata <= X"D6CC2E82";
    when 16#01216# => romdata <= X"C0388417";
    when 16#01217# => romdata <= X"08FC0670";
    when 16#01218# => romdata <= X"7A315556";
    when 16#01219# => romdata <= X"738F2481";
    when 16#0121A# => romdata <= X"F93881D6";
    when 16#0121B# => romdata <= X"CC0B81D6";
    when 16#0121C# => romdata <= X"D80C81D6";
    when 16#0121D# => romdata <= X"CC0B81D6";
    when 16#0121E# => romdata <= X"D40C7380";
    when 16#0121F# => romdata <= X"25FEB238";
    when 16#01220# => romdata <= X"83FF7627";
    when 16#01221# => romdata <= X"83DF3875";
    when 16#01222# => romdata <= X"892A7683";
    when 16#01223# => romdata <= X"2A555372";
    when 16#01224# => romdata <= X"802EBF38";
    when 16#01225# => romdata <= X"75862AB8";
    when 16#01226# => romdata <= X"05548473";
    when 16#01227# => romdata <= X"27B43880";
    when 16#01228# => romdata <= X"DB135494";
    when 16#01229# => romdata <= X"7327AB38";
    when 16#0122A# => romdata <= X"758C2A80";
    when 16#0122B# => romdata <= X"EE055480";
    when 16#0122C# => romdata <= X"D473279E";
    when 16#0122D# => romdata <= X"38758F2A";
    when 16#0122E# => romdata <= X"80F70554";
    when 16#0122F# => romdata <= X"82D47327";
    when 16#01230# => romdata <= X"91387592";
    when 16#01231# => romdata <= X"2A80FC05";
    when 16#01232# => romdata <= X"548AD473";
    when 16#01233# => romdata <= X"27843880";
    when 16#01234# => romdata <= X"FE547310";
    when 16#01235# => romdata <= X"101081D6";
    when 16#01236# => romdata <= X"C4058811";
    when 16#01237# => romdata <= X"08565874";
    when 16#01238# => romdata <= X"782E86CF";
    when 16#01239# => romdata <= X"38841508";
    when 16#0123A# => romdata <= X"FC065375";
    when 16#0123B# => romdata <= X"73278D38";
    when 16#0123C# => romdata <= X"88150855";
    when 16#0123D# => romdata <= X"74782E09";
    when 16#0123E# => romdata <= X"8106EA38";
    when 16#0123F# => romdata <= X"8C150881";
    when 16#01240# => romdata <= X"D6C40B84";
    when 16#01241# => romdata <= X"0508718C";
    when 16#01242# => romdata <= X"1A0C7688";
    when 16#01243# => romdata <= X"1A0C7888";
    when 16#01244# => romdata <= X"130C788C";
    when 16#01245# => romdata <= X"180C5D58";
    when 16#01246# => romdata <= X"7953807A";
    when 16#01247# => romdata <= X"2483E638";
    when 16#01248# => romdata <= X"72822C81";
    when 16#01249# => romdata <= X"712B5C53";
    when 16#0124A# => romdata <= X"7A7C2681";
    when 16#0124B# => romdata <= X"98387B7B";
    when 16#0124C# => romdata <= X"06537282";
    when 16#0124D# => romdata <= X"F13879FC";
    when 16#0124E# => romdata <= X"0684055A";
    when 16#0124F# => romdata <= X"7A10707D";
    when 16#01250# => romdata <= X"06545B72";
    when 16#01251# => romdata <= X"82E03884";
    when 16#01252# => romdata <= X"1A5AF139";
    when 16#01253# => romdata <= X"88178C11";
    when 16#01254# => romdata <= X"08585876";
    when 16#01255# => romdata <= X"782E0981";
    when 16#01256# => romdata <= X"06FCC238";
    when 16#01257# => romdata <= X"821A5AFD";
    when 16#01258# => romdata <= X"EC397817";
    when 16#01259# => romdata <= X"79810784";
    when 16#0125A# => romdata <= X"190C7081";
    when 16#0125B# => romdata <= X"D6D80C70";
    when 16#0125C# => romdata <= X"81D6D40C";
    when 16#0125D# => romdata <= X"81D6CC0B";
    when 16#0125E# => romdata <= X"8C120C8C";
    when 16#0125F# => romdata <= X"11088812";
    when 16#01260# => romdata <= X"0C748107";
    when 16#01261# => romdata <= X"84120C74";
    when 16#01262# => romdata <= X"1175710C";
    when 16#01263# => romdata <= X"51537D51";
    when 16#01264# => romdata <= X"87B73F88";
    when 16#01265# => romdata <= X"1754FCAC";
    when 16#01266# => romdata <= X"3981D6C4";
    when 16#01267# => romdata <= X"0B840508";
    when 16#01268# => romdata <= X"7A545C79";
    when 16#01269# => romdata <= X"8025FEF8";
    when 16#0126A# => romdata <= X"3882DA39";
    when 16#0126B# => romdata <= X"7A097C06";
    when 16#0126C# => romdata <= X"7081D6C4";
    when 16#0126D# => romdata <= X"0B84050C";
    when 16#0126E# => romdata <= X"5C7A105B";
    when 16#0126F# => romdata <= X"7A7C2685";
    when 16#01270# => romdata <= X"387A85B8";
    when 16#01271# => romdata <= X"3881D6C4";
    when 16#01272# => romdata <= X"0B880508";
    when 16#01273# => romdata <= X"70841208";
    when 16#01274# => romdata <= X"FC06707C";
    when 16#01275# => romdata <= X"317C7226";
    when 16#01276# => romdata <= X"8F722507";
    when 16#01277# => romdata <= X"57575C5D";
    when 16#01278# => romdata <= X"5572802E";
    when 16#01279# => romdata <= X"80DB3879";
    when 16#0127A# => romdata <= X"7A1681D6";
    when 16#0127B# => romdata <= X"BC081B90";
    when 16#0127C# => romdata <= X"115A5557";
    when 16#0127D# => romdata <= X"5B81D6B8";
    when 16#0127E# => romdata <= X"08FF2E88";
    when 16#0127F# => romdata <= X"38A08F13";
    when 16#01280# => romdata <= X"E0800657";
    when 16#01281# => romdata <= X"76527D51";
    when 16#01282# => romdata <= X"86C03FB0";
    when 16#01283# => romdata <= X"0854B008";
    when 16#01284# => romdata <= X"FF2E9038";
    when 16#01285# => romdata <= X"B0087627";
    when 16#01286# => romdata <= X"82993874";
    when 16#01287# => romdata <= X"81D6C42E";
    when 16#01288# => romdata <= X"82913881";
    when 16#01289# => romdata <= X"D6C40B88";
    when 16#0128A# => romdata <= X"05085584";
    when 16#0128B# => romdata <= X"1508FC06";
    when 16#0128C# => romdata <= X"707A317A";
    when 16#0128D# => romdata <= X"72268F72";
    when 16#0128E# => romdata <= X"25075255";
    when 16#0128F# => romdata <= X"537283E6";
    when 16#01290# => romdata <= X"38747981";
    when 16#01291# => romdata <= X"0784170C";
    when 16#01292# => romdata <= X"79167081";
    when 16#01293# => romdata <= X"D6C40B88";
    when 16#01294# => romdata <= X"050C7581";
    when 16#01295# => romdata <= X"0784120C";
    when 16#01296# => romdata <= X"547E5257";
    when 16#01297# => romdata <= X"85EB3F88";
    when 16#01298# => romdata <= X"1754FAE0";
    when 16#01299# => romdata <= X"3975832A";
    when 16#0129A# => romdata <= X"70545480";
    when 16#0129B# => romdata <= X"7424819B";
    when 16#0129C# => romdata <= X"3872822C";
    when 16#0129D# => romdata <= X"81712B81";
    when 16#0129E# => romdata <= X"D6C80807";
    when 16#0129F# => romdata <= X"7081D6C4";
    when 16#012A0# => romdata <= X"0B84050C";
    when 16#012A1# => romdata <= X"75101010";
    when 16#012A2# => romdata <= X"81D6C405";
    when 16#012A3# => romdata <= X"88110858";
    when 16#012A4# => romdata <= X"5A5D5377";
    when 16#012A5# => romdata <= X"8C180C74";
    when 16#012A6# => romdata <= X"88180C76";
    when 16#012A7# => romdata <= X"88190C76";
    when 16#012A8# => romdata <= X"8C160CFC";
    when 16#012A9# => romdata <= X"F339797A";
    when 16#012AA# => romdata <= X"10101081";
    when 16#012AB# => romdata <= X"D6C40570";
    when 16#012AC# => romdata <= X"57595D8C";
    when 16#012AD# => romdata <= X"15085776";
    when 16#012AE# => romdata <= X"752EA338";
    when 16#012AF# => romdata <= X"841708FC";
    when 16#012B0# => romdata <= X"06707A31";
    when 16#012B1# => romdata <= X"5556738F";
    when 16#012B2# => romdata <= X"2483CA38";
    when 16#012B3# => romdata <= X"73802584";
    when 16#012B4# => romdata <= X"81388C17";
    when 16#012B5# => romdata <= X"08577675";
    when 16#012B6# => romdata <= X"2E098106";
    when 16#012B7# => romdata <= X"DF388815";
    when 16#012B8# => romdata <= X"811B7083";
    when 16#012B9# => romdata <= X"06555B55";
    when 16#012BA# => romdata <= X"72C9387C";
    when 16#012BB# => romdata <= X"83065372";
    when 16#012BC# => romdata <= X"802EFDB8";
    when 16#012BD# => romdata <= X"38FF1DF8";
    when 16#012BE# => romdata <= X"19595D88";
    when 16#012BF# => romdata <= X"1808782E";
    when 16#012C0# => romdata <= X"EA38FDB5";
    when 16#012C1# => romdata <= X"39831A53";
    when 16#012C2# => romdata <= X"FC963983";
    when 16#012C3# => romdata <= X"1470822C";
    when 16#012C4# => romdata <= X"81712B81";
    when 16#012C5# => romdata <= X"D6C80807";
    when 16#012C6# => romdata <= X"7081D6C4";
    when 16#012C7# => romdata <= X"0B84050C";
    when 16#012C8# => romdata <= X"76101010";
    when 16#012C9# => romdata <= X"81D6C405";
    when 16#012CA# => romdata <= X"88110859";
    when 16#012CB# => romdata <= X"5B5E5153";
    when 16#012CC# => romdata <= X"FEE13981";
    when 16#012CD# => romdata <= X"D6880817";
    when 16#012CE# => romdata <= X"58B00876";
    when 16#012CF# => romdata <= X"2E818D38";
    when 16#012D0# => romdata <= X"81D6B808";
    when 16#012D1# => romdata <= X"FF2E83EC";
    when 16#012D2# => romdata <= X"38737631";
    when 16#012D3# => romdata <= X"1881D688";
    when 16#012D4# => romdata <= X"0C738706";
    when 16#012D5# => romdata <= X"70575372";
    when 16#012D6# => romdata <= X"802E8838";
    when 16#012D7# => romdata <= X"88733170";
    when 16#012D8# => romdata <= X"15555676";
    when 16#012D9# => romdata <= X"149FFF06";
    when 16#012DA# => romdata <= X"A0807131";
    when 16#012DB# => romdata <= X"1770547F";
    when 16#012DC# => romdata <= X"53575383";
    when 16#012DD# => romdata <= X"D53FB008";
    when 16#012DE# => romdata <= X"53B008FF";
    when 16#012DF# => romdata <= X"2E81A038";
    when 16#012E0# => romdata <= X"81D68808";
    when 16#012E1# => romdata <= X"167081D6";
    when 16#012E2# => romdata <= X"880C7475";
    when 16#012E3# => romdata <= X"81D6C40B";
    when 16#012E4# => romdata <= X"88050C74";
    when 16#012E5# => romdata <= X"76311870";
    when 16#012E6# => romdata <= X"81075155";
    when 16#012E7# => romdata <= X"56587B81";
    when 16#012E8# => romdata <= X"D6C42E83";
    when 16#012E9# => romdata <= X"9C38798F";
    when 16#012EA# => romdata <= X"2682CB38";
    when 16#012EB# => romdata <= X"810B8415";
    when 16#012EC# => romdata <= X"0C841508";
    when 16#012ED# => romdata <= X"FC06707A";
    when 16#012EE# => romdata <= X"317A7226";
    when 16#012EF# => romdata <= X"8F722507";
    when 16#012F0# => romdata <= X"52555372";
    when 16#012F1# => romdata <= X"802EFCF9";
    when 16#012F2# => romdata <= X"3880DB39";
    when 16#012F3# => romdata <= X"B0089FFF";
    when 16#012F4# => romdata <= X"065372FE";
    when 16#012F5# => romdata <= X"EB387781";
    when 16#012F6# => romdata <= X"D6880C81";
    when 16#012F7# => romdata <= X"D6C40B88";
    when 16#012F8# => romdata <= X"05087B18";
    when 16#012F9# => romdata <= X"81078412";
    when 16#012FA# => romdata <= X"0C5581D6";
    when 16#012FB# => romdata <= X"B4087827";
    when 16#012FC# => romdata <= X"86387781";
    when 16#012FD# => romdata <= X"D6B40C81";
    when 16#012FE# => romdata <= X"D6B00878";
    when 16#012FF# => romdata <= X"27FCAC38";
    when 16#01300# => romdata <= X"7781D6B0";
    when 16#01301# => romdata <= X"0C841508";
    when 16#01302# => romdata <= X"FC06707A";
    when 16#01303# => romdata <= X"317A7226";
    when 16#01304# => romdata <= X"8F722507";
    when 16#01305# => romdata <= X"52555372";
    when 16#01306# => romdata <= X"802EFCA5";
    when 16#01307# => romdata <= X"38883980";
    when 16#01308# => romdata <= X"745456FE";
    when 16#01309# => romdata <= X"DB397D51";
    when 16#0130A# => romdata <= X"829F3F80";
    when 16#0130B# => romdata <= X"0BB00C8F";
    when 16#0130C# => romdata <= X"3D0D0473";
    when 16#0130D# => romdata <= X"53807424";
    when 16#0130E# => romdata <= X"A9387282";
    when 16#0130F# => romdata <= X"2C81712B";
    when 16#01310# => romdata <= X"81D6C808";
    when 16#01311# => romdata <= X"077081D6";
    when 16#01312# => romdata <= X"C40B8405";
    when 16#01313# => romdata <= X"0C5D5377";
    when 16#01314# => romdata <= X"8C180C74";
    when 16#01315# => romdata <= X"88180C76";
    when 16#01316# => romdata <= X"88190C76";
    when 16#01317# => romdata <= X"8C160CF9";
    when 16#01318# => romdata <= X"B7398314";
    when 16#01319# => romdata <= X"70822C81";
    when 16#0131A# => romdata <= X"712B81D6";
    when 16#0131B# => romdata <= X"C8080770";
    when 16#0131C# => romdata <= X"81D6C40B";
    when 16#0131D# => romdata <= X"84050C5E";
    when 16#0131E# => romdata <= X"5153D439";
    when 16#0131F# => romdata <= X"7B7B0653";
    when 16#01320# => romdata <= X"72FCA338";
    when 16#01321# => romdata <= X"841A7B10";
    when 16#01322# => romdata <= X"5C5AF139";
    when 16#01323# => romdata <= X"FF1A8111";
    when 16#01324# => romdata <= X"515AF7B9";
    when 16#01325# => romdata <= X"39781779";
    when 16#01326# => romdata <= X"81078419";
    when 16#01327# => romdata <= X"0C8C1808";
    when 16#01328# => romdata <= X"88190871";
    when 16#01329# => romdata <= X"8C120C88";
    when 16#0132A# => romdata <= X"120C5970";
    when 16#0132B# => romdata <= X"81D6D80C";
    when 16#0132C# => romdata <= X"7081D6D4";
    when 16#0132D# => romdata <= X"0C81D6CC";
    when 16#0132E# => romdata <= X"0B8C120C";
    when 16#0132F# => romdata <= X"8C110888";
    when 16#01330# => romdata <= X"120C7481";
    when 16#01331# => romdata <= X"0784120C";
    when 16#01332# => romdata <= X"74117571";
    when 16#01333# => romdata <= X"0C5153F9";
    when 16#01334# => romdata <= X"BD397517";
    when 16#01335# => romdata <= X"84110881";
    when 16#01336# => romdata <= X"0784120C";
    when 16#01337# => romdata <= X"538C1708";
    when 16#01338# => romdata <= X"88180871";
    when 16#01339# => romdata <= X"8C120C88";
    when 16#0133A# => romdata <= X"120C587D";
    when 16#0133B# => romdata <= X"5180DA3F";
    when 16#0133C# => romdata <= X"881754F5";
    when 16#0133D# => romdata <= X"CF397284";
    when 16#0133E# => romdata <= X"150CF41A";
    when 16#0133F# => romdata <= X"F8067084";
    when 16#01340# => romdata <= X"1E088106";
    when 16#01341# => romdata <= X"07841E0C";
    when 16#01342# => romdata <= X"701D545B";
    when 16#01343# => romdata <= X"850B8414";
    when 16#01344# => romdata <= X"0C850B88";
    when 16#01345# => romdata <= X"140C8F7B";
    when 16#01346# => romdata <= X"27FDCF38";
    when 16#01347# => romdata <= X"881C527D";
    when 16#01348# => romdata <= X"5182903F";
    when 16#01349# => romdata <= X"81D6C40B";
    when 16#0134A# => romdata <= X"88050881";
    when 16#0134B# => romdata <= X"D6880859";
    when 16#0134C# => romdata <= X"55FDB739";
    when 16#0134D# => romdata <= X"7781D688";
    when 16#0134E# => romdata <= X"0C7381D6";
    when 16#0134F# => romdata <= X"B80CFC91";
    when 16#01350# => romdata <= X"39728415";
    when 16#01351# => romdata <= X"0CFDA339";
    when 16#01352# => romdata <= X"0404FD3D";
    when 16#01353# => romdata <= X"0D800B81";
    when 16#01354# => romdata <= X"F2E40C76";
    when 16#01355# => romdata <= X"5186CB3F";
    when 16#01356# => romdata <= X"B00853B0";
    when 16#01357# => romdata <= X"08FF2E88";
    when 16#01358# => romdata <= X"3872B00C";
    when 16#01359# => romdata <= X"853D0D04";
    when 16#0135A# => romdata <= X"81F2E408";
    when 16#0135B# => romdata <= X"5473802E";
    when 16#0135C# => romdata <= X"F0387574";
    when 16#0135D# => romdata <= X"710C5272";
    when 16#0135E# => romdata <= X"B00C853D";
    when 16#0135F# => romdata <= X"0D04FB3D";
    when 16#01360# => romdata <= X"0D777052";
    when 16#01361# => romdata <= X"56C23F81";
    when 16#01362# => romdata <= X"D6C40B88";
    when 16#01363# => romdata <= X"05088411";
    when 16#01364# => romdata <= X"08FC0670";
    when 16#01365# => romdata <= X"7B319FEF";
    when 16#01366# => romdata <= X"05E08006";
    when 16#01367# => romdata <= X"E0800556";
    when 16#01368# => romdata <= X"5653A080";
    when 16#01369# => romdata <= X"74249438";
    when 16#0136A# => romdata <= X"80527551";
    when 16#0136B# => romdata <= X"FF9C3F81";
    when 16#0136C# => romdata <= X"D6CC0815";
    when 16#0136D# => romdata <= X"5372B008";
    when 16#0136E# => romdata <= X"2E8F3875";
    when 16#0136F# => romdata <= X"51FF8A3F";
    when 16#01370# => romdata <= X"805372B0";
    when 16#01371# => romdata <= X"0C873D0D";
    when 16#01372# => romdata <= X"04733052";
    when 16#01373# => romdata <= X"7551FEFA";
    when 16#01374# => romdata <= X"3FB008FF";
    when 16#01375# => romdata <= X"2EA83881";
    when 16#01376# => romdata <= X"D6C40B88";
    when 16#01377# => romdata <= X"05087575";
    when 16#01378# => romdata <= X"31810784";
    when 16#01379# => romdata <= X"120C5381";
    when 16#0137A# => romdata <= X"D6880874";
    when 16#0137B# => romdata <= X"3181D688";
    when 16#0137C# => romdata <= X"0C7551FE";
    when 16#0137D# => romdata <= X"D43F810B";
    when 16#0137E# => romdata <= X"B00C873D";
    when 16#0137F# => romdata <= X"0D048052";
    when 16#01380# => romdata <= X"7551FEC6";
    when 16#01381# => romdata <= X"3F81D6C4";
    when 16#01382# => romdata <= X"0B880508";
    when 16#01383# => romdata <= X"B0087131";
    when 16#01384# => romdata <= X"56538F75";
    when 16#01385# => romdata <= X"25FFA438";
    when 16#01386# => romdata <= X"B00881D6";
    when 16#01387# => romdata <= X"B8083181";
    when 16#01388# => romdata <= X"D6880C74";
    when 16#01389# => romdata <= X"81078414";
    when 16#0138A# => romdata <= X"0C7551FE";
    when 16#0138B# => romdata <= X"9C3F8053";
    when 16#0138C# => romdata <= X"FF9039F6";
    when 16#0138D# => romdata <= X"3D0D7C7E";
    when 16#0138E# => romdata <= X"545B7280";
    when 16#0138F# => romdata <= X"2E828338";
    when 16#01390# => romdata <= X"7A51FE84";
    when 16#01391# => romdata <= X"3FF81384";
    when 16#01392# => romdata <= X"110870FE";
    when 16#01393# => romdata <= X"06701384";
    when 16#01394# => romdata <= X"1108FC06";
    when 16#01395# => romdata <= X"5D585954";
    when 16#01396# => romdata <= X"5881D6CC";
    when 16#01397# => romdata <= X"08752E82";
    when 16#01398# => romdata <= X"DE387884";
    when 16#01399# => romdata <= X"160C8073";
    when 16#0139A# => romdata <= X"8106545A";
    when 16#0139B# => romdata <= X"727A2E81";
    when 16#0139C# => romdata <= X"D5387815";
    when 16#0139D# => romdata <= X"84110881";
    when 16#0139E# => romdata <= X"06515372";
    when 16#0139F# => romdata <= X"A0387817";
    when 16#013A0# => romdata <= X"577981E6";
    when 16#013A1# => romdata <= X"38881508";
    when 16#013A2# => romdata <= X"537281D6";
    when 16#013A3# => romdata <= X"CC2E82F9";
    when 16#013A4# => romdata <= X"388C1508";
    when 16#013A5# => romdata <= X"708C150C";
    when 16#013A6# => romdata <= X"7388120C";
    when 16#013A7# => romdata <= X"56768107";
    when 16#013A8# => romdata <= X"84190C76";
    when 16#013A9# => romdata <= X"1877710C";
    when 16#013AA# => romdata <= X"53798191";
    when 16#013AB# => romdata <= X"3883FF77";
    when 16#013AC# => romdata <= X"2781C838";
    when 16#013AD# => romdata <= X"76892A77";
    when 16#013AE# => romdata <= X"832A5653";
    when 16#013AF# => romdata <= X"72802EBF";
    when 16#013B0# => romdata <= X"3876862A";
    when 16#013B1# => romdata <= X"B8055584";
    when 16#013B2# => romdata <= X"7327B438";
    when 16#013B3# => romdata <= X"80DB1355";
    when 16#013B4# => romdata <= X"947327AB";
    when 16#013B5# => romdata <= X"38768C2A";
    when 16#013B6# => romdata <= X"80EE0555";
    when 16#013B7# => romdata <= X"80D47327";
    when 16#013B8# => romdata <= X"9E38768F";
    when 16#013B9# => romdata <= X"2A80F705";
    when 16#013BA# => romdata <= X"5582D473";
    when 16#013BB# => romdata <= X"27913876";
    when 16#013BC# => romdata <= X"922A80FC";
    when 16#013BD# => romdata <= X"05558AD4";
    when 16#013BE# => romdata <= X"73278438";
    when 16#013BF# => romdata <= X"80FE5574";
    when 16#013C0# => romdata <= X"10101081";
    when 16#013C1# => romdata <= X"D6C40588";
    when 16#013C2# => romdata <= X"11085556";
    when 16#013C3# => romdata <= X"73762E82";
    when 16#013C4# => romdata <= X"B3388414";
    when 16#013C5# => romdata <= X"08FC0653";
    when 16#013C6# => romdata <= X"7673278D";
    when 16#013C7# => romdata <= X"38881408";
    when 16#013C8# => romdata <= X"5473762E";
    when 16#013C9# => romdata <= X"098106EA";
    when 16#013CA# => romdata <= X"388C1408";
    when 16#013CB# => romdata <= X"708C1A0C";
    when 16#013CC# => romdata <= X"74881A0C";
    when 16#013CD# => romdata <= X"7888120C";
    when 16#013CE# => romdata <= X"56778C15";
    when 16#013CF# => romdata <= X"0C7A51FC";
    when 16#013D0# => romdata <= X"883F8C3D";
    when 16#013D1# => romdata <= X"0D047708";
    when 16#013D2# => romdata <= X"78713159";
    when 16#013D3# => romdata <= X"77058819";
    when 16#013D4# => romdata <= X"08545772";
    when 16#013D5# => romdata <= X"81D6CC2E";
    when 16#013D6# => romdata <= X"80E0388C";
    when 16#013D7# => romdata <= X"1808708C";
    when 16#013D8# => romdata <= X"150C7388";
    when 16#013D9# => romdata <= X"120C56FE";
    when 16#013DA# => romdata <= X"89398815";
    when 16#013DB# => romdata <= X"088C1608";
    when 16#013DC# => romdata <= X"708C130C";
    when 16#013DD# => romdata <= X"5788170C";
    when 16#013DE# => romdata <= X"FEA33976";
    when 16#013DF# => romdata <= X"832A7054";
    when 16#013E0# => romdata <= X"55807524";
    when 16#013E1# => romdata <= X"81983872";
    when 16#013E2# => romdata <= X"822C8171";
    when 16#013E3# => romdata <= X"2B81D6C8";
    when 16#013E4# => romdata <= X"080781D6";
    when 16#013E5# => romdata <= X"C40B8405";
    when 16#013E6# => romdata <= X"0C537410";
    when 16#013E7# => romdata <= X"101081D6";
    when 16#013E8# => romdata <= X"C4058811";
    when 16#013E9# => romdata <= X"08555675";
    when 16#013EA# => romdata <= X"8C190C73";
    when 16#013EB# => romdata <= X"88190C77";
    when 16#013EC# => romdata <= X"88170C77";
    when 16#013ED# => romdata <= X"8C150CFF";
    when 16#013EE# => romdata <= X"8439815A";
    when 16#013EF# => romdata <= X"FDB43978";
    when 16#013F0# => romdata <= X"17738106";
    when 16#013F1# => romdata <= X"54577298";
    when 16#013F2# => romdata <= X"38770878";
    when 16#013F3# => romdata <= X"71315977";
    when 16#013F4# => romdata <= X"058C1908";
    when 16#013F5# => romdata <= X"881A0871";
    when 16#013F6# => romdata <= X"8C120C88";
    when 16#013F7# => romdata <= X"120C5757";
    when 16#013F8# => romdata <= X"76810784";
    when 16#013F9# => romdata <= X"190C7781";
    when 16#013FA# => romdata <= X"D6C40B88";
    when 16#013FB# => romdata <= X"050C81D6";
    when 16#013FC# => romdata <= X"C0087726";
    when 16#013FD# => romdata <= X"FEC73881";
    when 16#013FE# => romdata <= X"D6BC0852";
    when 16#013FF# => romdata <= X"7A51FAFE";
    when 16#01400# => romdata <= X"3F7A51FA";
    when 16#01401# => romdata <= X"C43FFEBA";
    when 16#01402# => romdata <= X"3981788C";
    when 16#01403# => romdata <= X"150C7888";
    when 16#01404# => romdata <= X"150C738C";
    when 16#01405# => romdata <= X"1A0C7388";
    when 16#01406# => romdata <= X"1A0C5AFD";
    when 16#01407# => romdata <= X"80398315";
    when 16#01408# => romdata <= X"70822C81";
    when 16#01409# => romdata <= X"712B81D6";
    when 16#0140A# => romdata <= X"C8080781";
    when 16#0140B# => romdata <= X"D6C40B84";
    when 16#0140C# => romdata <= X"050C5153";
    when 16#0140D# => romdata <= X"74101010";
    when 16#0140E# => romdata <= X"81D6C405";
    when 16#0140F# => romdata <= X"88110855";
    when 16#01410# => romdata <= X"56FEE439";
    when 16#01411# => romdata <= X"74538075";
    when 16#01412# => romdata <= X"24A73872";
    when 16#01413# => romdata <= X"822C8171";
    when 16#01414# => romdata <= X"2B81D6C8";
    when 16#01415# => romdata <= X"080781D6";
    when 16#01416# => romdata <= X"C40B8405";
    when 16#01417# => romdata <= X"0C53758C";
    when 16#01418# => romdata <= X"190C7388";
    when 16#01419# => romdata <= X"190C7788";
    when 16#0141A# => romdata <= X"170C778C";
    when 16#0141B# => romdata <= X"150CFDCD";
    when 16#0141C# => romdata <= X"39831570";
    when 16#0141D# => romdata <= X"822C8171";
    when 16#0141E# => romdata <= X"2B81D6C8";
    when 16#0141F# => romdata <= X"080781D6";
    when 16#01420# => romdata <= X"C40B8405";
    when 16#01421# => romdata <= X"0C5153D6";
    when 16#01422# => romdata <= X"39810BB0";
    when 16#01423# => romdata <= X"0C04803D";
    when 16#01424# => romdata <= X"0D72812E";
    when 16#01425# => romdata <= X"8938800B";
    when 16#01426# => romdata <= X"B00C823D";
    when 16#01427# => romdata <= X"0D047351";
    when 16#01428# => romdata <= X"B23FFE3D";
    when 16#01429# => romdata <= X"0D81F2E0";
    when 16#0142A# => romdata <= X"0851708A";
    when 16#0142B# => romdata <= X"3881F2E8";
    when 16#0142C# => romdata <= X"7081F2E0";
    when 16#0142D# => romdata <= X"0C517075";
    when 16#0142E# => romdata <= X"125252FF";
    when 16#0142F# => romdata <= X"537087FB";
    when 16#01430# => romdata <= X"80802688";
    when 16#01431# => romdata <= X"387081F2";
    when 16#01432# => romdata <= X"E00C7153";
    when 16#01433# => romdata <= X"72B00C84";
    when 16#01434# => romdata <= X"3D0D0400";
    when 16#01435# => romdata <= X"FF390000";
    when 16#01436# => romdata <= X"00000000";
    when 16#01437# => romdata <= X"00000000";
    when 16#01438# => romdata <= X"00000000";
    when 16#01439# => romdata <= X"00000000";
    when 16#0143A# => romdata <= X"00CAC5CA";
    when 16#0143B# => romdata <= X"C5C0C0C0";
    when 16#0143C# => romdata <= X"C0C0C0C0";
    when 16#0143D# => romdata <= X"C0C0C0CF";
    when 16#0143E# => romdata <= X"CFCFCF00";
    when 16#0143F# => romdata <= X"00000F0F";
    when 16#01440# => romdata <= X"0F0F8F8F";
    when 16#01441# => romdata <= X"CFCFCFCF";
    when 16#01442# => romdata <= X"CFCF4F0F";
    when 16#01443# => romdata <= X"0F0F0000";
    when 16#01444# => romdata <= X"CFCFCFCF";
    when 16#01445# => romdata <= X"0F0F0F0F";
    when 16#01446# => romdata <= X"0F0F0F0F";
    when 16#01447# => romdata <= X"0F0FFEFE";
    when 16#01448# => romdata <= X"FEFC0000";
    when 16#01449# => romdata <= X"CFCFCFCF";
    when 16#0144A# => romdata <= X"CFCFCFCF";
    when 16#0144B# => romdata <= X"CFCFCFCF";
    when 16#0144C# => romdata <= X"CFFFFF7E";
    when 16#0144D# => romdata <= X"7E000000";
    when 16#0144E# => romdata <= X"00000000";
    when 16#0144F# => romdata <= X"00000000";
    when 16#01450# => romdata <= X"00000000";
    when 16#01451# => romdata <= X"00003F3F";
    when 16#01452# => romdata <= X"3F3F0101";
    when 16#01453# => romdata <= X"01010101";
    when 16#01454# => romdata <= X"01010101";
    when 16#01455# => romdata <= X"3F3F3F3F";
    when 16#01456# => romdata <= X"0000383C";
    when 16#01457# => romdata <= X"3E3E3F3F";
    when 16#01458# => romdata <= X"3F3B3B39";
    when 16#01459# => romdata <= X"39383838";
    when 16#0145A# => romdata <= X"38383800";
    when 16#0145B# => romdata <= X"003F3F3F";
    when 16#0145C# => romdata <= X"3F383838";
    when 16#0145D# => romdata <= X"38383838";
    when 16#0145E# => romdata <= X"38383C3F";
    when 16#0145F# => romdata <= X"3F1F0F00";
    when 16#01460# => romdata <= X"003F3F3F";
    when 16#01461# => romdata <= X"3F030303";
    when 16#01462# => romdata <= X"03030303";
    when 16#01463# => romdata <= X"03033F3F";
    when 16#01464# => romdata <= X"3F3E0000";
    when 16#01465# => romdata <= X"00000000";
    when 16#01466# => romdata <= X"00000000";
    when 16#01467# => romdata <= X"00000000";
    when 16#01468# => romdata <= X"00000000";
    when 16#01469# => romdata <= X"00000000";
    when 16#0146A# => romdata <= X"00000000";
    when 16#0146B# => romdata <= X"00000000";
    when 16#0146C# => romdata <= X"00000000";
    when 16#0146D# => romdata <= X"00000000";
    when 16#0146E# => romdata <= X"00000000";
    when 16#0146F# => romdata <= X"00000000";
    when 16#01470# => romdata <= X"00000000";
    when 16#01471# => romdata <= X"00000000";
    when 16#01472# => romdata <= X"00000000";
    when 16#01473# => romdata <= X"00000000";
    when 16#01474# => romdata <= X"00000000";
    when 16#01475# => romdata <= X"00000000";
    when 16#01476# => romdata <= X"00000000";
    when 16#01477# => romdata <= X"00000000";
    when 16#01478# => romdata <= X"00000000";
    when 16#01479# => romdata <= X"00000000";
    when 16#0147A# => romdata <= X"00000000";
    when 16#0147B# => romdata <= X"00000000";
    when 16#0147C# => romdata <= X"00000000";
    when 16#0147D# => romdata <= X"8080C0C0";
    when 16#0147E# => romdata <= X"E0E06000";
    when 16#0147F# => romdata <= X"00000000";
    when 16#01480# => romdata <= X"00000000";
    when 16#01481# => romdata <= X"00000000";
    when 16#01482# => romdata <= X"00000000";
    when 16#01483# => romdata <= X"00000000";
    when 16#01484# => romdata <= X"00000000";
    when 16#01485# => romdata <= X"00000000";
    when 16#01486# => romdata <= X"00000000";
    when 16#01487# => romdata <= X"00000000";
    when 16#01488# => romdata <= X"00000000";
    when 16#01489# => romdata <= X"00000000";
    when 16#0148A# => romdata <= X"00000000";
    when 16#0148B# => romdata <= X"00000000";
    when 16#0148C# => romdata <= X"00000000";
    when 16#0148D# => romdata <= X"00000000";
    when 16#0148E# => romdata <= X"00000000";
    when 16#0148F# => romdata <= X"00000000";
    when 16#01490# => romdata <= X"00000000";
    when 16#01491# => romdata <= X"00000000";
    when 16#01492# => romdata <= X"00000000";
    when 16#01493# => romdata <= X"806098EE";
    when 16#01494# => romdata <= X"77BBDDEC";
    when 16#01495# => romdata <= X"EE6E0200";
    when 16#01496# => romdata <= X"00000000";
    when 16#01497# => romdata <= X"00E08080";
    when 16#01498# => romdata <= X"E00000E0";
    when 16#01499# => romdata <= X"A0A00000";
    when 16#0149A# => romdata <= X"E0000000";
    when 16#0149B# => romdata <= X"00E0C000";
    when 16#0149C# => romdata <= X"C0E00000";
    when 16#0149D# => romdata <= X"E08080E0";
    when 16#0149E# => romdata <= X"0000C020";
    when 16#0149F# => romdata <= X"20C00000";
    when 16#014A0# => romdata <= X"E0000000";
    when 16#014A1# => romdata <= X"20E02000";
    when 16#014A2# => romdata <= X"0020A060";
    when 16#014A3# => romdata <= X"20000000";
    when 16#014A4# => romdata <= X"00000000";
    when 16#014A5# => romdata <= X"00000000";
    when 16#014A6# => romdata <= X"00000000";
    when 16#014A7# => romdata <= X"00000000";
    when 16#014A8# => romdata <= X"00000000";
    when 16#014A9# => romdata <= X"00000000";
    when 16#014AA# => romdata <= X"00030007";
    when 16#014AB# => romdata <= X"00070701";
    when 16#014AC# => romdata <= X"00000000";
    when 16#014AD# => romdata <= X"00000000";
    when 16#014AE# => romdata <= X"00000300";
    when 16#014AF# => romdata <= X"C0030000";
    when 16#014B0# => romdata <= X"034242C0";
    when 16#014B1# => romdata <= X"00C34242";
    when 16#014B2# => romdata <= X"0000C380";
    when 16#014B3# => romdata <= X"01C00340";
    when 16#014B4# => romdata <= X"C04300C0";
    when 16#014B5# => romdata <= X"43408001";
    when 16#014B6# => romdata <= X"C20201C0";
    when 16#014B7# => romdata <= X"00C38202";
    when 16#014B8# => romdata <= X"80C00300";
    when 16#014B9# => romdata <= X"00C04342";
    when 16#014BA# => romdata <= X"8202C040";
    when 16#014BB# => romdata <= X"40800000";
    when 16#014BC# => romdata <= X"C0404000";
    when 16#014BD# => romdata <= X"80404000";
    when 16#014BE# => romdata <= X"00C04040";
    when 16#014BF# => romdata <= X"8000C040";
    when 16#014C0# => romdata <= X"4000C080";
    when 16#014C1# => romdata <= X"00C00000";
    when 16#014C2# => romdata <= X"00000000";
    when 16#014C3# => romdata <= X"00000000";
    when 16#014C4# => romdata <= X"00000000";
    when 16#014C5# => romdata <= X"00000000";
    when 16#014C6# => romdata <= X"00FF0000";
    when 16#014C7# => romdata <= X"0000C645";
    when 16#014C8# => romdata <= X"44800785";
    when 16#014C9# => romdata <= X"45408007";
    when 16#014CA# => romdata <= X"80424700";
    when 16#014CB# => romdata <= X"80474000";
    when 16#014CC# => romdata <= X"07C14344";
    when 16#014CD# => romdata <= X"00C38404";
    when 16#014CE# => romdata <= X"C30007C1";
    when 16#014CF# => romdata <= X"42418700";
    when 16#014D0# => romdata <= X"80404784";
    when 16#014D1# => romdata <= X"04C34047";
    when 16#014D2# => romdata <= X"8101C640";
    when 16#014D3# => romdata <= X"40070505";
    when 16#014D4# => romdata <= X"00040502";
    when 16#014D5# => romdata <= X"00000704";
    when 16#014D6# => romdata <= X"04030007";
    when 16#014D7# => romdata <= X"05050007";
    when 16#014D8# => romdata <= X"00020700";
    when 16#014D9# => romdata <= X"00000000";
    when 16#014DA# => romdata <= X"00000000";
    when 16#014DB# => romdata <= X"00000000";
    when 16#014DC# => romdata <= X"00000000";
    when 16#014DD# => romdata <= X"0000FF00";
    when 16#014DE# => romdata <= X"00000007";
    when 16#014DF# => romdata <= X"01030500";
    when 16#014E0# => romdata <= X"03040403";
    when 16#014E1# => romdata <= X"00040502";
    when 16#014E2# => romdata <= X"00040502";
    when 16#014E3# => romdata <= X"00000705";
    when 16#014E4# => romdata <= X"05000700";
    when 16#014E5# => romdata <= X"02070000";
    when 16#014E6# => romdata <= X"07040403";
    when 16#014E7# => romdata <= X"00030404";
    when 16#014E8# => romdata <= X"03000701";
    when 16#014E9# => romdata <= X"03050007";
    when 16#014EA# => romdata <= X"01010000";
    when 16#014EB# => romdata <= X"00000000";
    when 16#014EC# => romdata <= X"00000000";
    when 16#014ED# => romdata <= X"00000000";
    when 16#014EE# => romdata <= X"00000000";
    when 16#014EF# => romdata <= X"00000000";
    when 16#014F0# => romdata <= X"71756974";
    when 16#014F1# => romdata <= X"00000000";
    when 16#014F2# => romdata <= X"68656C70";
    when 16#014F3# => romdata <= X"00000000";
    when 16#014F4# => romdata <= X"0A307800";
    when 16#014F5# => romdata <= X"69326320";
    when 16#014F6# => romdata <= X"464D430A";
    when 16#014F7# => romdata <= X"00000000";
    when 16#014F8# => romdata <= X"61646472";
    when 16#014F9# => romdata <= X"6573733A";
    when 16#014FA# => romdata <= X"20307800";
    when 16#014FB# => romdata <= X"2020202D";
    when 16#014FC# => romdata <= X"2D3E2020";
    when 16#014FD# => romdata <= X"2041434B";
    when 16#014FE# => romdata <= X"0A000000";
    when 16#014FF# => romdata <= X"72656164";
    when 16#01500# => romdata <= X"20646174";
    when 16#01501# => romdata <= X"61202800";
    when 16#01502# => romdata <= X"20627974";
    when 16#01503# => romdata <= X"65732920";
    when 16#01504# => romdata <= X"66726F6D";
    when 16#01505# => romdata <= X"20493243";
    when 16#01506# => romdata <= X"2D616464";
    when 16#01507# => romdata <= X"72657373";
    when 16#01508# => romdata <= X"20307800";
    when 16#01509# => romdata <= X"0A0A0000";
    when 16#0150A# => romdata <= X"6E6F6163";
    when 16#0150B# => romdata <= X"6B200000";
    when 16#0150C# => romdata <= X"6368726F";
    when 16#0150D# => romdata <= X"6E74656C";
    when 16#0150E# => romdata <= X"20726567";
    when 16#0150F# => romdata <= X"20307800";
    when 16#01510# => romdata <= X"3A203078";
    when 16#01511# => romdata <= X"00000000";
    when 16#01512# => romdata <= X"206E6163";
    when 16#01513# => romdata <= X"6B000000";
    when 16#01514# => romdata <= X"6572726F";
    when 16#01515# => romdata <= X"7220286E";
    when 16#01516# => romdata <= X"61636B29";
    when 16#01517# => romdata <= X"0A000000";
    when 16#01518# => romdata <= X"0A202063";
    when 16#01519# => romdata <= X"68616E6E";
    when 16#0151A# => romdata <= X"656C2033";
    when 16#0151B# => romdata <= X"20696E70";
    when 16#0151C# => romdata <= X"7574206F";
    when 16#0151D# => romdata <= X"76657266";
    when 16#0151E# => romdata <= X"6C6F7700";
    when 16#0151F# => romdata <= X"0A202063";
    when 16#01520# => romdata <= X"68616E6E";
    when 16#01521# => romdata <= X"656C2032";
    when 16#01522# => romdata <= X"20696E70";
    when 16#01523# => romdata <= X"7574206F";
    when 16#01524# => romdata <= X"76657266";
    when 16#01525# => romdata <= X"6C6F7700";
    when 16#01526# => romdata <= X"0A202063";
    when 16#01527# => romdata <= X"68616E6E";
    when 16#01528# => romdata <= X"656C2031";
    when 16#01529# => romdata <= X"20696E70";
    when 16#0152A# => romdata <= X"7574206F";
    when 16#0152B# => romdata <= X"76657266";
    when 16#0152C# => romdata <= X"6C6F7700";
    when 16#0152D# => romdata <= X"0A202063";
    when 16#0152E# => romdata <= X"68616E6E";
    when 16#0152F# => romdata <= X"656C2030";
    when 16#01530# => romdata <= X"20696E70";
    when 16#01531# => romdata <= X"7574206F";
    when 16#01532# => romdata <= X"76657266";
    when 16#01533# => romdata <= X"6C6F7700";
    when 16#01534# => romdata <= X"0A202063";
    when 16#01535# => romdata <= X"68616E6E";
    when 16#01536# => romdata <= X"656C2033";
    when 16#01537# => romdata <= X"20717561";
    when 16#01538# => romdata <= X"6473756D";
    when 16#01539# => romdata <= X"206F7665";
    when 16#0153A# => romdata <= X"72666C6F";
    when 16#0153B# => romdata <= X"77000000";
    when 16#0153C# => romdata <= X"0A202063";
    when 16#0153D# => romdata <= X"68616E6E";
    when 16#0153E# => romdata <= X"656C2032";
    when 16#0153F# => romdata <= X"20717561";
    when 16#01540# => romdata <= X"6473756D";
    when 16#01541# => romdata <= X"206F7665";
    when 16#01542# => romdata <= X"72666C6F";
    when 16#01543# => romdata <= X"77000000";
    when 16#01544# => romdata <= X"0A202063";
    when 16#01545# => romdata <= X"68616E6E";
    when 16#01546# => romdata <= X"656C2031";
    when 16#01547# => romdata <= X"20717561";
    when 16#01548# => romdata <= X"6473756D";
    when 16#01549# => romdata <= X"206F7665";
    when 16#0154A# => romdata <= X"72666C6F";
    when 16#0154B# => romdata <= X"77000000";
    when 16#0154C# => romdata <= X"0A202063";
    when 16#0154D# => romdata <= X"68616E6E";
    when 16#0154E# => romdata <= X"656C2030";
    when 16#0154F# => romdata <= X"20717561";
    when 16#01550# => romdata <= X"6473756D";
    when 16#01551# => romdata <= X"206F7665";
    when 16#01552# => romdata <= X"72666C6F";
    when 16#01553# => romdata <= X"77000000";
    when 16#01554# => romdata <= X"0A202073";
    when 16#01555# => romdata <= X"756D2076";
    when 16#01556# => romdata <= X"616C7565";
    when 16#01557# => romdata <= X"20637574";
    when 16#01558# => romdata <= X"74656400";
    when 16#01559# => romdata <= X"0A202063";
    when 16#0155A# => romdata <= X"68616E6E";
    when 16#0155B# => romdata <= X"656C2033";
    when 16#0155C# => romdata <= X"20646976";
    when 16#0155D# => romdata <= X"6964656E";
    when 16#0155E# => romdata <= X"64206375";
    when 16#0155F# => romdata <= X"74746564";
    when 16#01560# => romdata <= X"00000000";
    when 16#01561# => romdata <= X"0A202063";
    when 16#01562# => romdata <= X"68616E6E";
    when 16#01563# => romdata <= X"656C2033";
    when 16#01564# => romdata <= X"206E6F69";
    when 16#01565# => romdata <= X"73652063";
    when 16#01566# => romdata <= X"6F6D7065";
    when 16#01567# => romdata <= X"6E736174";
    when 16#01568# => romdata <= X"696F6E20";
    when 16#01569# => romdata <= X"746F2062";
    when 16#0156A# => romdata <= X"69670000";
    when 16#0156B# => romdata <= X"0A202063";
    when 16#0156C# => romdata <= X"68616E6E";
    when 16#0156D# => romdata <= X"656C2033";
    when 16#0156E# => romdata <= X"206E6F69";
    when 16#0156F# => romdata <= X"73652076";
    when 16#01570# => romdata <= X"616C7565";
    when 16#01571# => romdata <= X"20637574";
    when 16#01572# => romdata <= X"74656400";
    when 16#01573# => romdata <= X"0A202063";
    when 16#01574# => romdata <= X"68616E6E";
    when 16#01575# => romdata <= X"656C2032";
    when 16#01576# => romdata <= X"20646976";
    when 16#01577# => romdata <= X"6964656E";
    when 16#01578# => romdata <= X"64206375";
    when 16#01579# => romdata <= X"74746564";
    when 16#0157A# => romdata <= X"00000000";
    when 16#0157B# => romdata <= X"0A202063";
    when 16#0157C# => romdata <= X"68616E6E";
    when 16#0157D# => romdata <= X"656C2032";
    when 16#0157E# => romdata <= X"206E6F69";
    when 16#0157F# => romdata <= X"73652063";
    when 16#01580# => romdata <= X"6F6D7065";
    when 16#01581# => romdata <= X"6E736174";
    when 16#01582# => romdata <= X"696F6E20";
    when 16#01583# => romdata <= X"746F2062";
    when 16#01584# => romdata <= X"69670000";
    when 16#01585# => romdata <= X"0A202063";
    when 16#01586# => romdata <= X"68616E6E";
    when 16#01587# => romdata <= X"656C2032";
    when 16#01588# => romdata <= X"206E6F69";
    when 16#01589# => romdata <= X"73652076";
    when 16#0158A# => romdata <= X"616C7565";
    when 16#0158B# => romdata <= X"20637574";
    when 16#0158C# => romdata <= X"74656400";
    when 16#0158D# => romdata <= X"0A202063";
    when 16#0158E# => romdata <= X"68616E6E";
    when 16#0158F# => romdata <= X"656C2031";
    when 16#01590# => romdata <= X"20646976";
    when 16#01591# => romdata <= X"6964656E";
    when 16#01592# => romdata <= X"64206375";
    when 16#01593# => romdata <= X"74746564";
    when 16#01594# => romdata <= X"00000000";
    when 16#01595# => romdata <= X"0A202063";
    when 16#01596# => romdata <= X"68616E6E";
    when 16#01597# => romdata <= X"656C2031";
    when 16#01598# => romdata <= X"206E6F69";
    when 16#01599# => romdata <= X"73652063";
    when 16#0159A# => romdata <= X"6F6D7065";
    when 16#0159B# => romdata <= X"6E736174";
    when 16#0159C# => romdata <= X"696F6E20";
    when 16#0159D# => romdata <= X"746F2062";
    when 16#0159E# => romdata <= X"69670000";
    when 16#0159F# => romdata <= X"0A202063";
    when 16#015A0# => romdata <= X"68616E6E";
    when 16#015A1# => romdata <= X"656C2031";
    when 16#015A2# => romdata <= X"206E6F69";
    when 16#015A3# => romdata <= X"73652076";
    when 16#015A4# => romdata <= X"616C7565";
    when 16#015A5# => romdata <= X"20637574";
    when 16#015A6# => romdata <= X"74656400";
    when 16#015A7# => romdata <= X"0A202063";
    when 16#015A8# => romdata <= X"68616E6E";
    when 16#015A9# => romdata <= X"656C2030";
    when 16#015AA# => romdata <= X"20646976";
    when 16#015AB# => romdata <= X"6964656E";
    when 16#015AC# => romdata <= X"64206375";
    when 16#015AD# => romdata <= X"74746564";
    when 16#015AE# => romdata <= X"00000000";
    when 16#015AF# => romdata <= X"0A202063";
    when 16#015B0# => romdata <= X"68616E6E";
    when 16#015B1# => romdata <= X"656C2030";
    when 16#015B2# => romdata <= X"206E6F69";
    when 16#015B3# => romdata <= X"73652063";
    when 16#015B4# => romdata <= X"6F6D7065";
    when 16#015B5# => romdata <= X"6E736174";
    when 16#015B6# => romdata <= X"696F6E20";
    when 16#015B7# => romdata <= X"746F2062";
    when 16#015B8# => romdata <= X"69670000";
    when 16#015B9# => romdata <= X"0A202063";
    when 16#015BA# => romdata <= X"68616E6E";
    when 16#015BB# => romdata <= X"656C2030";
    when 16#015BC# => romdata <= X"206E6F69";
    when 16#015BD# => romdata <= X"73652076";
    when 16#015BE# => romdata <= X"616C7565";
    when 16#015BF# => romdata <= X"20637574";
    when 16#015C0# => romdata <= X"74656400";
    when 16#015C1# => romdata <= X"0A202073";
    when 16#015C2# => romdata <= X"6F667477";
    when 16#015C3# => romdata <= X"61726520";
    when 16#015C4# => romdata <= X"6572726F";
    when 16#015C5# => romdata <= X"72000000";
    when 16#015C6# => romdata <= X"0A657874";
    when 16#015C7# => romdata <= X"65726E61";
    when 16#015C8# => romdata <= X"6C20636C";
    when 16#015C9# => romdata <= X"6F636B20";
    when 16#015CA# => romdata <= X"20202020";
    when 16#015CB# => romdata <= X"2020203A";
    when 16#015CC# => romdata <= X"20000000";
    when 16#015CD# => romdata <= X"61637469";
    when 16#015CE# => romdata <= X"76650000";
    when 16#015CF# => romdata <= X"0A6D6963";
    when 16#015D0# => romdata <= X"726F7075";
    when 16#015D1# => romdata <= X"6C736520";
    when 16#015D2# => romdata <= X"736F7572";
    when 16#015D3# => romdata <= X"63652020";
    when 16#015D4# => romdata <= X"2020203A";
    when 16#015D5# => romdata <= X"20000000";
    when 16#015D6# => romdata <= X"65787465";
    when 16#015D7# => romdata <= X"726E616C";
    when 16#015D8# => romdata <= X"00000000";
    when 16#015D9# => romdata <= X"0A6D6963";
    when 16#015DA# => romdata <= X"726F7075";
    when 16#015DB# => romdata <= X"6C736520";
    when 16#015DC# => romdata <= X"6576656E";
    when 16#015DD# => romdata <= X"74206C69";
    when 16#015DE# => romdata <= X"6D69743A";
    when 16#015DF# => romdata <= X"20000000";
    when 16#015E0# => romdata <= X"0A6D6561";
    when 16#015E1# => romdata <= X"73757265";
    when 16#015E2# => romdata <= X"6D656E74";
    when 16#015E3# => romdata <= X"206C656E";
    when 16#015E4# => romdata <= X"67746820";
    when 16#015E5# => romdata <= X"2020203A";
    when 16#015E6# => romdata <= X"20000000";
    when 16#015E7# => romdata <= X"0A626561";
    when 16#015E8# => romdata <= X"6D20706F";
    when 16#015E9# => romdata <= X"73697469";
    when 16#015EA# => romdata <= X"6F6E206D";
    when 16#015EB# => romdata <= X"6F6E6974";
    when 16#015EC# => romdata <= X"6F722072";
    when 16#015ED# => romdata <= X"65676973";
    when 16#015EE# => romdata <= X"74657273";
    when 16#015EF# => romdata <= X"00000000";
    when 16#015F0# => romdata <= X"0A202020";
    when 16#015F1# => romdata <= X"20202020";
    when 16#015F2# => romdata <= X"20202020";
    when 16#015F3# => romdata <= X"20202020";
    when 16#015F4# => romdata <= X"20202020";
    when 16#015F5# => romdata <= X"20202020";
    when 16#015F6# => romdata <= X"20636861";
    when 16#015F7# => romdata <= X"6E6E656C";
    when 16#015F8# => romdata <= X"20302020";
    when 16#015F9# => romdata <= X"20636861";
    when 16#015FA# => romdata <= X"6E6E656C";
    when 16#015FB# => romdata <= X"20312020";
    when 16#015FC# => romdata <= X"20636861";
    when 16#015FD# => romdata <= X"6E6E656C";
    when 16#015FE# => romdata <= X"20322020";
    when 16#015FF# => romdata <= X"20636861";
    when 16#01600# => romdata <= X"6E6E656C";
    when 16#01601# => romdata <= X"20330000";
    when 16#01602# => romdata <= X"0A202020";
    when 16#01603# => romdata <= X"20202020";
    when 16#01604# => romdata <= X"20202020";
    when 16#01605# => romdata <= X"20202020";
    when 16#01606# => romdata <= X"20202020";
    when 16#01607# => romdata <= X"20202020";
    when 16#01608# => romdata <= X"202D2D2D";
    when 16#01609# => romdata <= X"2D20686F";
    when 16#0160A# => romdata <= X"72697A6F";
    when 16#0160B# => romdata <= X"6E74616C";
    when 16#0160C# => romdata <= X"202D2D2D";
    when 16#0160D# => romdata <= X"2D2D2020";
    when 16#0160E# => romdata <= X"202D2D2D";
    when 16#0160F# => romdata <= X"2D2D2D20";
    when 16#01610# => romdata <= X"76657274";
    when 16#01611# => romdata <= X"6963616C";
    when 16#01612# => romdata <= X"202D2D2D";
    when 16#01613# => romdata <= X"2D2D0000";
    when 16#01614# => romdata <= X"0A736361";
    when 16#01615# => romdata <= X"6C657220";
    when 16#01616# => romdata <= X"76616C75";
    when 16#01617# => romdata <= X"65732020";
    when 16#01618# => romdata <= X"20202020";
    when 16#01619# => romdata <= X"20202020";
    when 16#0161A# => romdata <= X"20000000";
    when 16#0161B# => romdata <= X"0A6E6F69";
    when 16#0161C# => romdata <= X"73652063";
    when 16#0161D# => romdata <= X"6F6D7065";
    when 16#0161E# => romdata <= X"6E736174";
    when 16#0161F# => romdata <= X"696F6E20";
    when 16#01620# => romdata <= X"20202020";
    when 16#01621# => romdata <= X"20000000";
    when 16#01622# => romdata <= X"0A6D6561";
    when 16#01623# => romdata <= X"73757265";
    when 16#01624# => romdata <= X"6D656E74";
    when 16#01625# => romdata <= X"20202020";
    when 16#01626# => romdata <= X"20202020";
    when 16#01627# => romdata <= X"20202020";
    when 16#01628# => romdata <= X"20000000";
    when 16#01629# => romdata <= X"0A73616D";
    when 16#0162A# => romdata <= X"706C6573";
    when 16#0162B# => romdata <= X"20286469";
    when 16#0162C# => romdata <= X"7629203A";
    when 16#0162D# => romdata <= X"20000000";
    when 16#0162E# => romdata <= X"0A73756D";
    when 16#0162F# => romdata <= X"20636861";
    when 16#01630# => romdata <= X"6E6E656C";
    when 16#01631# => romdata <= X"2020203A";
    when 16#01632# => romdata <= X"20000000";
    when 16#01633# => romdata <= X"0A0A706F";
    when 16#01634# => romdata <= X"73697469";
    when 16#01635# => romdata <= X"6F6E2063";
    when 16#01636# => romdata <= X"6F6D7075";
    when 16#01637# => romdata <= X"74617469";
    when 16#01638# => romdata <= X"6F6E0000";
    when 16#01639# => romdata <= X"0A202073";
    when 16#0163A# => romdata <= X"63616C65";
    when 16#0163B# => romdata <= X"72207661";
    when 16#0163C# => romdata <= X"6C756573";
    when 16#0163D# => romdata <= X"20202020";
    when 16#0163E# => romdata <= X"20202020";
    when 16#0163F# => romdata <= X"20000000";
    when 16#01640# => romdata <= X"0A20206F";
    when 16#01641# => romdata <= X"66667365";
    when 16#01642# => romdata <= X"74202020";
    when 16#01643# => romdata <= X"20202020";
    when 16#01644# => romdata <= X"20202020";
    when 16#01645# => romdata <= X"20202020";
    when 16#01646# => romdata <= X"20000000";
    when 16#01647# => romdata <= X"0A6F7574";
    when 16#01648# => romdata <= X"70757420";
    when 16#01649# => romdata <= X"73656C65";
    when 16#0164A# => romdata <= X"6374203A";
    when 16#0164B# => romdata <= X"20000000";
    when 16#0164C# => romdata <= X"74657374";
    when 16#0164D# => romdata <= X"67656E00";
    when 16#0164E# => romdata <= X"4E4F5420";
    when 16#0164F# => romdata <= X"00000000";
    when 16#01650# => romdata <= X"6368616E";
    when 16#01651# => romdata <= X"6E656C20";
    when 16#01652# => romdata <= X"30000000";
    when 16#01653# => romdata <= X"0A63616C";
    when 16#01654# => romdata <= X"63207374";
    when 16#01655# => romdata <= X"61746520";
    when 16#01656# => romdata <= X"2020203A";
    when 16#01657# => romdata <= X"20307800";
    when 16#01658# => romdata <= X"76657274";
    when 16#01659# => romdata <= X"6963616C";
    when 16#0165A# => romdata <= X"00000000";
    when 16#0165B# => romdata <= X"686F7269";
    when 16#0165C# => romdata <= X"7A6F6E74";
    when 16#0165D# => romdata <= X"616C0000";
    when 16#0165E# => romdata <= X"73756D00";
    when 16#0165F# => romdata <= X"6368616E";
    when 16#01660# => romdata <= X"6E656C20";
    when 16#01661# => romdata <= X"33000000";
    when 16#01662# => romdata <= X"6368616E";
    when 16#01663# => romdata <= X"6E656C20";
    when 16#01664# => romdata <= X"32000000";
    when 16#01665# => romdata <= X"6368616E";
    when 16#01666# => romdata <= X"6E656C20";
    when 16#01667# => romdata <= X"31000000";
    when 16#01668# => romdata <= X"786D6F64";
    when 16#01669# => romdata <= X"656D2074";
    when 16#0166A# => romdata <= X"72616E73";
    when 16#0166B# => romdata <= X"6D69742E";
    when 16#0166C# => romdata <= X"2E2E0A00";
    when 16#0166D# => romdata <= X"20627974";
    when 16#0166E# => romdata <= X"65732074";
    when 16#0166F# => romdata <= X"72616E73";
    when 16#01670# => romdata <= X"6D697474";
    when 16#01671# => romdata <= X"65640A00";
    when 16#01672# => romdata <= X"63616E63";
    when 16#01673# => romdata <= X"656C0A00";
    when 16#01674# => romdata <= X"72657472";
    when 16#01675# => romdata <= X"79206F75";
    when 16#01676# => romdata <= X"740A0000";
    when 16#01677# => romdata <= X"786D6F64";
    when 16#01678# => romdata <= X"656D2072";
    when 16#01679# => romdata <= X"65636569";
    when 16#0167A# => romdata <= X"76652E2E";
    when 16#0167B# => romdata <= X"2E0A0000";
    when 16#0167C# => romdata <= X"20627974";
    when 16#0167D# => romdata <= X"65732072";
    when 16#0167E# => romdata <= X"65636569";
    when 16#0167F# => romdata <= X"7665640A";
    when 16#01680# => romdata <= X"00000000";
    when 16#01681# => romdata <= X"72782062";
    when 16#01682# => romdata <= X"75666665";
    when 16#01683# => romdata <= X"72206675";
    when 16#01684# => romdata <= X"6C6C0A00";
    when 16#01685# => romdata <= X"74696D65";
    when 16#01686# => romdata <= X"206F7574";
    when 16#01687# => romdata <= X"0A000000";
    when 16#01688# => romdata <= X"64656275";
    when 16#01689# => romdata <= X"67207265";
    when 16#0168A# => romdata <= X"67697374";
    when 16#0168B# => romdata <= X"65727300";
    when 16#0168C# => romdata <= X"0A6D6F64";
    when 16#0168D# => romdata <= X"65202020";
    when 16#0168E# => romdata <= X"20202020";
    when 16#0168F# => romdata <= X"203A2000";
    when 16#01690# => romdata <= X"0A616464";
    when 16#01691# => romdata <= X"72657373";
    when 16#01692# => romdata <= X"20302020";
    when 16#01693# => romdata <= X"203A2030";
    when 16#01694# => romdata <= X"78000000";
    when 16#01695# => romdata <= X"0A616464";
    when 16#01696# => romdata <= X"72657373";
    when 16#01697# => romdata <= X"20312020";
    when 16#01698# => romdata <= X"203A2030";
    when 16#01699# => romdata <= X"78000000";
    when 16#0169A# => romdata <= X"0A627566";
    when 16#0169B# => romdata <= X"66657220";
    when 16#0169C# => romdata <= X"73697A65";
    when 16#0169D# => romdata <= X"203A2000";
    when 16#0169E# => romdata <= X"6D61783A";
    when 16#0169F# => romdata <= X"20000000";
    when 16#016A0# => romdata <= X"6D696E3A";
    when 16#016A1# => romdata <= X"20000000";
    when 16#016A2# => romdata <= X"63683A20";
    when 16#016A3# => romdata <= X"00000000";
    when 16#016A4# => romdata <= X"73706C3A";
    when 16#016A5# => romdata <= X"20000000";
    when 16#016A6# => romdata <= X"73686F77";
    when 16#016A7# => romdata <= X"2042504D";
    when 16#016A8# => romdata <= X"20726567";
    when 16#016A9# => romdata <= X"69737465";
    when 16#016AA# => romdata <= X"72730000";
    when 16#016AB# => romdata <= X"62706D00";
    when 16#016AC# => romdata <= X"73656C65";
    when 16#016AD# => romdata <= X"6374206F";
    when 16#016AE# => romdata <= X"75747075";
    when 16#016AF# => romdata <= X"74206368";
    when 16#016B0# => romdata <= X"616E6E65";
    when 16#016B1# => romdata <= X"6C202830";
    when 16#016B2# => romdata <= X"2E2E3320";
    when 16#016B3# => romdata <= X"73756D20";
    when 16#016B4# => romdata <= X"68207629";
    when 16#016B5# => romdata <= X"00000000";
    when 16#016B6# => romdata <= X"73656C65";
    when 16#016B7# => romdata <= X"63740000";
    when 16#016B8# => romdata <= X"73797374";
    when 16#016B9# => romdata <= X"656D2072";
    when 16#016BA# => romdata <= X"65736574";
    when 16#016BB# => romdata <= X"00000000";
    when 16#016BC# => romdata <= X"72657365";
    when 16#016BD# => romdata <= X"74000000";
    when 16#016BE# => romdata <= X"73686F77";
    when 16#016BF# => romdata <= X"20737973";
    when 16#016C0# => romdata <= X"74656D20";
    when 16#016C1# => romdata <= X"696E666F";
    when 16#016C2# => romdata <= X"203C7665";
    when 16#016C3# => romdata <= X"72626F73";
    when 16#016C4# => romdata <= X"653E0000";
    when 16#016C5# => romdata <= X"73797369";
    when 16#016C6# => romdata <= X"6E666F00";
    when 16#016C7# => romdata <= X"73686F77";
    when 16#016C8# => romdata <= X"2F736574";
    when 16#016C9# => romdata <= X"20646562";
    when 16#016CA# => romdata <= X"75672072";
    when 16#016CB# => romdata <= X"65676973";
    when 16#016CC# => romdata <= X"74657273";
    when 16#016CD# => romdata <= X"203C7365";
    when 16#016CE# => romdata <= X"74206D6F";
    when 16#016CF# => romdata <= X"64653E00";
    when 16#016D0# => romdata <= X"64656275";
    when 16#016D1# => romdata <= X"67000000";
    when 16#016D2# => romdata <= X"636C6B20";
    when 16#016D3# => romdata <= X"736F7572";
    when 16#016D4# => romdata <= X"63653A20";
    when 16#016D5# => romdata <= X"2030203D";
    when 16#016D6# => romdata <= X"20696E74";
    when 16#016D7# => romdata <= X"2C203120";
    when 16#016D8# => romdata <= X"3D206578";
    when 16#016D9# => romdata <= X"74000000";
    when 16#016DA# => romdata <= X"636C6B00";
    when 16#016DB# => romdata <= X"6D696372";
    when 16#016DC# => romdata <= X"6F70756C";
    when 16#016DD# => romdata <= X"73652073";
    when 16#016DE# => romdata <= X"6F757263";
    when 16#016DF# => romdata <= X"653A2030";
    when 16#016E0# => romdata <= X"203D2069";
    when 16#016E1# => romdata <= X"6E742C20";
    when 16#016E2# => romdata <= X"31203D20";
    when 16#016E3# => romdata <= X"65787400";
    when 16#016E4# => romdata <= X"6D696372";
    when 16#016E5# => romdata <= X"6F000000";
    when 16#016E6# => romdata <= X"74657374";
    when 16#016E7# => romdata <= X"67656E65";
    when 16#016E8# => romdata <= X"7261746F";
    when 16#016E9# => romdata <= X"72203C73";
    when 16#016EA# => romdata <= X"63616C65";
    when 16#016EB# => romdata <= X"723E203C";
    when 16#016EC# => romdata <= X"72657374";
    when 16#016ED# => romdata <= X"6172743E";
    when 16#016EE# => romdata <= X"00000000";
    when 16#016EF# => romdata <= X"3C6D7574";
    when 16#016F0# => romdata <= X"655F6E3E";
    when 16#016F1# => romdata <= X"203C7273";
    when 16#016F2# => romdata <= X"745F6E3E";
    when 16#016F3# => romdata <= X"203C6270";
    when 16#016F4# => romdata <= X"625F6E3E";
    when 16#016F5# => romdata <= X"203C6F73";
    when 16#016F6# => romdata <= X"72313E20";
    when 16#016F7# => romdata <= X"3C6F7372";
    when 16#016F8# => romdata <= X"323E0000";
    when 16#016F9# => romdata <= X"64616363";
    when 16#016FA# => romdata <= X"6F6E6600";
    when 16#016FB# => romdata <= X"3C6D756C";
    when 16#016FC# => romdata <= X"7469706C";
    when 16#016FD# => romdata <= X"6965723E";
    when 16#016FE# => romdata <= X"20696E69";
    when 16#016FF# => romdata <= X"7469616C";
    when 16#01700# => romdata <= X"697A6520";
    when 16#01701# => romdata <= X"62756666";
    when 16#01702# => romdata <= X"65720000";
    when 16#01703# => romdata <= X"64616374";
    when 16#01704# => romdata <= X"65737400";
    when 16#01705# => romdata <= X"72657365";
    when 16#01706# => romdata <= X"74206361";
    when 16#01707# => romdata <= X"6C63756C";
    when 16#01708# => romdata <= X"6174696F";
    when 16#01709# => romdata <= X"6E206572";
    when 16#0170A# => romdata <= X"726F7273";
    when 16#0170B# => romdata <= X"00000000";
    when 16#0170C# => romdata <= X"63616C63";
    when 16#0170D# => romdata <= X"72657300";
    when 16#0170E# => romdata <= X"73686F77";
    when 16#0170F# => romdata <= X"20646562";
    when 16#01710# => romdata <= X"75672062";
    when 16#01711# => romdata <= X"75666665";
    when 16#01712# => romdata <= X"72203C6C";
    when 16#01713# => romdata <= X"656E6774";
    when 16#01714# => romdata <= X"683E0000";
    when 16#01715# => romdata <= X"636C6561";
    when 16#01716# => romdata <= X"72206465";
    when 16#01717# => romdata <= X"62756720";
    when 16#01718# => romdata <= X"62756666";
    when 16#01719# => romdata <= X"65720000";
    when 16#0171A# => romdata <= X"62636C65";
    when 16#0171B# => romdata <= X"61720000";
    when 16#0171C# => romdata <= X"62756666";
    when 16#0171D# => romdata <= X"6572206F";
    when 16#0171E# => romdata <= X"6E204C43";
    when 16#0171F# => romdata <= X"44203C63";
    when 16#01720# => romdata <= X"683E203C";
    when 16#01721# => romdata <= X"636F6D62";
    when 16#01722# => romdata <= X"3E000000";
    when 16#01723# => romdata <= X"73636F70";
    when 16#01724# => romdata <= X"65000000";
    when 16#01725# => romdata <= X"64656275";
    when 16#01726# => romdata <= X"67207472";
    when 16#01727# => romdata <= X"61636520";
    when 16#01728# => romdata <= X"3C636C65";
    when 16#01729# => romdata <= X"61723E00";
    when 16#0172A# => romdata <= X"74726163";
    when 16#0172B# => romdata <= X"65000000";
    when 16#0172C# => romdata <= X"73657475";
    when 16#0172D# => romdata <= X"70206368";
    when 16#0172E# => romdata <= X"616E6E65";
    when 16#0172F# => romdata <= X"6C207465";
    when 16#01730# => romdata <= X"7374203C";
    when 16#01731# => romdata <= X"63683E20";
    when 16#01732# => romdata <= X"3C76616C";
    when 16#01733# => romdata <= X"302E2E37";
    when 16#01734# => romdata <= X"3E000000";
    when 16#01735# => romdata <= X"63687465";
    when 16#01736# => romdata <= X"73740000";
    when 16#01737# => romdata <= X"72756E6E";
    when 16#01738# => romdata <= X"696E6720";
    when 16#01739# => romdata <= X"6C696768";
    when 16#0173A# => romdata <= X"74000000";
    when 16#0173B# => romdata <= X"72756E00";
    when 16#0173C# => romdata <= X"72756E20";
    when 16#0173D# => romdata <= X"64697370";
    when 16#0173E# => romdata <= X"6C617920";
    when 16#0173F# => romdata <= X"74657374";
    when 16#01740# => romdata <= X"2066756E";
    when 16#01741# => romdata <= X"6374696F";
    when 16#01742# => romdata <= X"6E000000";
    when 16#01743# => romdata <= X"64697370";
    when 16#01744# => romdata <= X"6C617900";
    when 16#01745# => romdata <= X"73657420";
    when 16#01746# => romdata <= X"6261636B";
    when 16#01747# => romdata <= X"6C696768";
    when 16#01748# => romdata <= X"74203C30";
    when 16#01749# => romdata <= X"2E2E3331";
    when 16#0174A# => romdata <= X"3E000000";
    when 16#0174B# => romdata <= X"6261636B";
    when 16#0174C# => romdata <= X"00000000";
    when 16#0174D# => romdata <= X"73686F77";
    when 16#0174E# => romdata <= X"206C6F67";
    when 16#0174F# => romdata <= X"6F206F6E";
    when 16#01750# => romdata <= X"20676C63";
    when 16#01751# => romdata <= X"64000000";
    when 16#01752# => romdata <= X"6C6F676F";
    when 16#01753# => romdata <= X"00000000";
    when 16#01754# => romdata <= X"63686563";
    when 16#01755# => romdata <= X"6B204932";
    when 16#01756# => romdata <= X"43206164";
    when 16#01757# => romdata <= X"64726573";
    when 16#01758# => romdata <= X"73000000";
    when 16#01759# => romdata <= X"69326300";
    when 16#0175A# => romdata <= X"72656164";
    when 16#0175B# => romdata <= X"20454550";
    when 16#0175C# => romdata <= X"524F4D20";
    when 16#0175D# => romdata <= X"3C627573";
    when 16#0175E# => romdata <= X"3E203C69";
    when 16#0175F# => romdata <= X"32635F61";
    when 16#01760# => romdata <= X"6464723E";
    when 16#01761# => romdata <= X"203C6C65";
    when 16#01762# => romdata <= X"6E677468";
    when 16#01763# => romdata <= X"3E000000";
    when 16#01764# => romdata <= X"65657072";
    when 16#01765# => romdata <= X"6F6D0000";
    when 16#01766# => romdata <= X"41444320";
    when 16#01767# => romdata <= X"72656769";
    when 16#01768# => romdata <= X"73746572";
    when 16#01769# => romdata <= X"20747261";
    when 16#0176A# => romdata <= X"6E736665";
    when 16#0176B# => romdata <= X"72203C76";
    when 16#0176C# => romdata <= X"616C7565";
    when 16#0176D# => romdata <= X"3E000000";
    when 16#0176E# => romdata <= X"61747261";
    when 16#0176F# => romdata <= X"6E730000";
    when 16#01770# => romdata <= X"696E6974";
    when 16#01771# => romdata <= X"20414443";
    when 16#01772# => romdata <= X"20726567";
    when 16#01773# => romdata <= X"69737465";
    when 16#01774# => romdata <= X"72730000";
    when 16#01775# => romdata <= X"61696E69";
    when 16#01776# => romdata <= X"74000000";
    when 16#01777# => romdata <= X"616C6961";
    when 16#01778# => romdata <= X"7320666F";
    when 16#01779# => romdata <= X"72207800";
    when 16#0177A# => romdata <= X"6D656D00";
    when 16#0177B# => romdata <= X"77726974";
    when 16#0177C# => romdata <= X"6520776F";
    when 16#0177D# => romdata <= X"7264203C";
    when 16#0177E# => romdata <= X"61646472";
    when 16#0177F# => romdata <= X"3E203C6C";
    when 16#01780# => romdata <= X"656E6774";
    when 16#01781# => romdata <= X"683E203C";
    when 16#01782# => romdata <= X"76616C75";
    when 16#01783# => romdata <= X"65287329";
    when 16#01784# => romdata <= X"3E000000";
    when 16#01785# => romdata <= X"776D656D";
    when 16#01786# => romdata <= X"00000000";
    when 16#01787# => romdata <= X"6558616D";
    when 16#01788# => romdata <= X"696E6520";
    when 16#01789# => romdata <= X"6D656D6F";
    when 16#0178A# => romdata <= X"72790000";
    when 16#0178B# => romdata <= X"636C6561";
    when 16#0178C# => romdata <= X"72207363";
    when 16#0178D# => romdata <= X"7265656E";
    when 16#0178E# => romdata <= X"00000000";
    when 16#0178F# => romdata <= X"636C6561";
    when 16#01790# => romdata <= X"72000000";
    when 16#01791# => romdata <= X"0A646562";
    when 16#01792# => romdata <= X"75672074";
    when 16#01793# => romdata <= X"72616365";
    when 16#01794# => romdata <= X"206D656D";
    when 16#01795# => romdata <= X"6F727900";
    when 16#01796# => romdata <= X"0A74696D";
    when 16#01797# => romdata <= X"65207374";
    when 16#01798# => romdata <= X"616D7020";
    when 16#01799# => romdata <= X"20202073";
    when 16#0179A# => romdata <= X"74617465";
    when 16#0179B# => romdata <= X"00000000";
    when 16#0179C# => romdata <= X"20203078";
    when 16#0179D# => romdata <= X"00000000";
    when 16#0179E# => romdata <= X"65787465";
    when 16#0179F# => romdata <= X"726E616C";
    when 16#017A0# => romdata <= X"20636C6F";
    when 16#017A1# => romdata <= X"636B2000";
    when 16#017A2# => romdata <= X"61637469";
    when 16#017A3# => romdata <= X"76650A00";
    when 16#017A4# => romdata <= X"73656C65";
    when 16#017A5# => romdata <= X"63746564";
    when 16#017A6# => romdata <= X"0A000000";
    when 16#017A7# => romdata <= X"6D696372";
    when 16#017A8# => romdata <= X"6F70756C";
    when 16#017A9# => romdata <= X"73652073";
    when 16#017AA# => romdata <= X"6F757263";
    when 16#017AB# => romdata <= X"653A2000";
    when 16#017AC# => romdata <= X"6265616D";
    when 16#017AD# => romdata <= X"20706F73";
    when 16#017AE# => romdata <= X"6974696F";
    when 16#017AF# => romdata <= X"6E206D6F";
    when 16#017B0# => romdata <= X"6E69746F";
    when 16#017B1# => romdata <= X"72000000";
    when 16#017B2# => romdata <= X"20286F6E";
    when 16#017B3# => romdata <= X"2073696D";
    when 16#017B4# => romdata <= X"290A0000";
    when 16#017B5# => romdata <= X"0A485720";
    when 16#017B6# => romdata <= X"73796E74";
    when 16#017B7# => romdata <= X"68657369";
    when 16#017B8# => romdata <= X"7A65643A";
    when 16#017B9# => romdata <= X"20000000";
    when 16#017BA# => romdata <= X"0A535720";
    when 16#017BB# => romdata <= X"636F6D70";
    when 16#017BC# => romdata <= X"696C6564";
    when 16#017BD# => romdata <= X"2020203A";
    when 16#017BE# => romdata <= X"20417567";
    when 16#017BF# => romdata <= X"20313120";
    when 16#017C0# => romdata <= X"32303131";
    when 16#017C1# => romdata <= X"20203131";
    when 16#017C2# => romdata <= X"3A30353A";
    when 16#017C3# => romdata <= X"32370000";
    when 16#017C4# => romdata <= X"0A737973";
    when 16#017C5# => romdata <= X"74656D20";
    when 16#017C6# => romdata <= X"636C6F63";
    when 16#017C7# => romdata <= X"6B20203A";
    when 16#017C8# => romdata <= X"20000000";
    when 16#017C9# => romdata <= X"204D487A";
    when 16#017CA# => romdata <= X"0A000000";
    when 16#017CB# => romdata <= X"44454255";
    when 16#017CC# => romdata <= X"47204D4F";
    when 16#017CD# => romdata <= X"44450000";
    when 16#017CE# => romdata <= X"204F4E0A";
    when 16#017CF# => romdata <= X"00000000";
    when 16#017D0# => romdata <= X"0000117B";
    when 16#017D1# => romdata <= X"000011E4";
    when 16#017D2# => romdata <= X"000011D9";
    when 16#017D3# => romdata <= X"000011CE";
    when 16#017D4# => romdata <= X"000011C3";
    when 16#017D5# => romdata <= X"000011B9";
    when 16#017D6# => romdata <= X"000011AF";
    when 16#017D7# => romdata <= X"000002C2";
    when 16#017D8# => romdata <= X"FC1902C4";
    when 16#017D9# => romdata <= X"FFFEFD3F";
    when 16#017DA# => romdata <= X"03E7FD3B";
    when 16#017DB# => romdata <= X"0000485D";
    when 16#017DC# => romdata <= X"999B4888";
    when 16#017DD# => romdata <= X"FFC4B7CE";
    when 16#017DE# => romdata <= X"6665B74E";
    when 16#017DF# => romdata <= X"3E200000";
    when 16#017E0# => romdata <= X"636F6D6D";
    when 16#017E1# => romdata <= X"616E6420";
    when 16#017E2# => romdata <= X"6E6F7420";
    when 16#017E3# => romdata <= X"666F756E";
    when 16#017E4# => romdata <= X"642E0A00";
    when 16#017E5# => romdata <= X"73757070";
    when 16#017E6# => romdata <= X"6F727465";
    when 16#017E7# => romdata <= X"6420636F";
    when 16#017E8# => romdata <= X"6D6D616E";
    when 16#017E9# => romdata <= X"64733A0A";
    when 16#017EA# => romdata <= X"0A000000";
    when 16#017EB# => romdata <= X"202D2000";
    when 16#017EC# => romdata <= X"76656E64";
    when 16#017ED# => romdata <= X"6F723F20";
    when 16#017EE# => romdata <= X"20000000";
    when 16#017EF# => romdata <= X"67616973";
    when 16#017F0# => romdata <= X"6C657220";
    when 16#017F1# => romdata <= X"20000000";
    when 16#017F2# => romdata <= X"756E6B6E";
    when 16#017F3# => romdata <= X"6F776E20";
    when 16#017F4# => romdata <= X"64657669";
    when 16#017F5# => romdata <= X"63650000";
    when 16#017F6# => romdata <= X"485A4452";
    when 16#017F7# => romdata <= X"20202020";
    when 16#017F8# => romdata <= X"20000000";
    when 16#017F9# => romdata <= X"47656E65";
    when 16#017FA# => romdata <= X"72616C20";
    when 16#017FB# => romdata <= X"50757270";
    when 16#017FC# => romdata <= X"6F736520";
    when 16#017FD# => romdata <= X"492F4F20";
    when 16#017FE# => romdata <= X"706F7274";
    when 16#017FF# => romdata <= X"00000000";
    when 16#01800# => romdata <= X"56474120";
    when 16#01801# => romdata <= X"636F6E74";
    when 16#01802# => romdata <= X"726F6C6C";
    when 16#01803# => romdata <= X"65720000";
    when 16#01804# => romdata <= X"4475616C";
    when 16#01805# => romdata <= X"2D706F72";
    when 16#01806# => romdata <= X"74204148";
    when 16#01807# => romdata <= X"42205352";
    when 16#01808# => romdata <= X"414D206D";
    when 16#01809# => romdata <= X"6F64756C";
    when 16#0180A# => romdata <= X"65000000";
    when 16#0180B# => romdata <= X"64656275";
    when 16#0180C# => romdata <= X"67206275";
    when 16#0180D# => romdata <= X"66666572";
    when 16#0180E# => romdata <= X"20636F6E";
    when 16#0180F# => romdata <= X"74726F6C";
    when 16#01810# => romdata <= X"00000000";
    when 16#01811# => romdata <= X"74726967";
    when 16#01812# => romdata <= X"67657220";
    when 16#01813# => romdata <= X"67656E65";
    when 16#01814# => romdata <= X"7261746F";
    when 16#01815# => romdata <= X"72000000";
    when 16#01816# => romdata <= X"64656275";
    when 16#01817# => romdata <= X"6720636F";
    when 16#01818# => romdata <= X"6E736F6C";
    when 16#01819# => romdata <= X"65000000";
    when 16#0181A# => romdata <= X"64656275";
    when 16#0181B# => romdata <= X"67207472";
    when 16#0181C# => romdata <= X"61636572";
    when 16#0181D# => romdata <= X"206D656D";
    when 16#0181E# => romdata <= X"6F727900";
    when 16#0181F# => romdata <= X"4541444F";
    when 16#01820# => romdata <= X"47533130";
    when 16#01821# => romdata <= X"32206469";
    when 16#01822# => romdata <= X"73706C61";
    when 16#01823# => romdata <= X"79206472";
    when 16#01824# => romdata <= X"69766572";
    when 16#01825# => romdata <= X"00000000";
    when 16#01826# => romdata <= X"44434D20";
    when 16#01827# => romdata <= X"70686173";
    when 16#01828# => romdata <= X"65207368";
    when 16#01829# => romdata <= X"69667420";
    when 16#0182A# => romdata <= X"636F6E74";
    when 16#0182B# => romdata <= X"726F6C00";
    when 16#0182C# => romdata <= X"5A505520";
    when 16#0182D# => romdata <= X"4D656D6F";
    when 16#0182E# => romdata <= X"72792077";
    when 16#0182F# => romdata <= X"72617070";
    when 16#01830# => romdata <= X"65720000";
    when 16#01831# => romdata <= X"5A505520";
    when 16#01832# => romdata <= X"41484220";
    when 16#01833# => romdata <= X"57726170";
    when 16#01834# => romdata <= X"70657200";
    when 16#01835# => romdata <= X"4148422F";
    when 16#01836# => romdata <= X"41504220";
    when 16#01837# => romdata <= X"42726964";
    when 16#01838# => romdata <= X"67650000";
    when 16#01839# => romdata <= X"4D6F6475";
    when 16#0183A# => romdata <= X"6C617220";
    when 16#0183B# => romdata <= X"54696D65";
    when 16#0183C# => romdata <= X"7220556E";
    when 16#0183D# => romdata <= X"69740000";
    when 16#0183E# => romdata <= X"414D4241";
    when 16#0183F# => romdata <= X"20577261";
    when 16#01840# => romdata <= X"70706572";
    when 16#01841# => romdata <= X"20666F72";
    when 16#01842# => romdata <= X"204F4320";
    when 16#01843# => romdata <= X"4932432D";
    when 16#01844# => romdata <= X"6D617374";
    when 16#01845# => romdata <= X"65720000";
    when 16#01846# => romdata <= X"47656E65";
    when 16#01847# => romdata <= X"72696320";
    when 16#01848# => romdata <= X"55415254";
    when 16#01849# => romdata <= X"00000000";
    when 16#0184A# => romdata <= X"20206170";
    when 16#0184B# => romdata <= X"62736C76";
    when 16#0184C# => romdata <= X"00000000";
    when 16#0184D# => romdata <= X"76656E64";
    when 16#0184E# => romdata <= X"20307800";
    when 16#0184F# => romdata <= X"64657620";
    when 16#01850# => romdata <= X"30780000";
    when 16#01851# => romdata <= X"76657220";
    when 16#01852# => romdata <= X"00000000";
    when 16#01853# => romdata <= X"69727120";
    when 16#01854# => romdata <= X"00000000";
    when 16#01855# => romdata <= X"61646472";
    when 16#01856# => romdata <= X"20307800";
    when 16#01857# => romdata <= X"6168626D";
    when 16#01858# => romdata <= X"73740000";
    when 16#01859# => romdata <= X"61686273";
    when 16#0185A# => romdata <= X"6C760000";
    when 16#0185B# => romdata <= X"00002AF2";
    when 16#0185C# => romdata <= X"00002BB3";
    when 16#0185D# => romdata <= X"00002BA8";
    when 16#0185E# => romdata <= X"00002B9D";
    when 16#0185F# => romdata <= X"00002B7C";
    when 16#01860# => romdata <= X"00002B71";
    when 16#01861# => romdata <= X"00002B66";
    when 16#01862# => romdata <= X"00002B5B";
    when 16#01863# => romdata <= X"00002B92";
    when 16#01864# => romdata <= X"00002B87";
    when 16#01865# => romdata <= X"04580808";
    when 16#01866# => romdata <= X"20FF0000";
    when 16#01867# => romdata <= X"000061A4";
    when 16#01868# => romdata <= X"00006284";
    when 16#01869# => romdata <= X"02010305";
    when 16#0186A# => romdata <= X"05070501";
    when 16#0186B# => romdata <= X"03030505";
    when 16#0186C# => romdata <= X"02030104";
    when 16#0186D# => romdata <= X"05050505";
    when 16#0186E# => romdata <= X"05050505";
    when 16#0186F# => romdata <= X"05050101";
    when 16#01870# => romdata <= X"04050404";
    when 16#01871# => romdata <= X"07050505";
    when 16#01872# => romdata <= X"05050505";
    when 16#01873# => romdata <= X"05030405";
    when 16#01874# => romdata <= X"05050505";
    when 16#01875# => romdata <= X"05050505";
    when 16#01876# => romdata <= X"05050505";
    when 16#01877# => romdata <= X"05050503";
    when 16#01878# => romdata <= X"04030505";
    when 16#01879# => romdata <= X"02050504";
    when 16#0187A# => romdata <= X"05050405";
    when 16#0187B# => romdata <= X"04010204";
    when 16#0187C# => romdata <= X"02050404";
    when 16#0187D# => romdata <= X"05050404";
    when 16#0187E# => romdata <= X"04040507";
    when 16#0187F# => romdata <= X"05040404";
    when 16#01880# => romdata <= X"02040500";
    when 16#01881# => romdata <= X"04050200";
    when 16#01882# => romdata <= X"04080303";
    when 16#01883# => romdata <= X"04090003";
    when 16#01884# => romdata <= X"06000000";
    when 16#01885# => romdata <= X"00020204";
    when 16#01886# => romdata <= X"04040400";
    when 16#01887# => romdata <= X"04060003";
    when 16#01888# => romdata <= X"05000000";
    when 16#01889# => romdata <= X"00000404";
    when 16#0188A# => romdata <= X"05050204";
    when 16#0188B# => romdata <= X"05060305";
    when 16#0188C# => romdata <= X"04030705";
    when 16#0188D# => romdata <= X"04050303";
    when 16#0188E# => romdata <= X"02040502";
    when 16#0188F# => romdata <= X"03020405";
    when 16#01890# => romdata <= X"06060604";
    when 16#01891# => romdata <= X"05050505";
    when 16#01892# => romdata <= X"05050504";
    when 16#01893# => romdata <= X"04040404";
    when 16#01894# => romdata <= X"03030303";
    when 16#01895# => romdata <= X"05050505";
    when 16#01896# => romdata <= X"05050505";
    when 16#01897# => romdata <= X"05040404";
    when 16#01898# => romdata <= X"04050404";
    when 16#01899# => romdata <= X"04040404";
    when 16#0189A# => romdata <= X"04040503";
    when 16#0189B# => romdata <= X"04040404";
    when 16#0189C# => romdata <= X"02020303";
    when 16#0189D# => romdata <= X"04040404";
    when 16#0189E# => romdata <= X"04040405";
    when 16#0189F# => romdata <= X"04040404";
    when 16#018A0# => romdata <= X"04030303";
    when 16#018A1# => romdata <= X"00005F07";
    when 16#018A2# => romdata <= X"0007741C";
    when 16#018A3# => romdata <= X"771C172E";
    when 16#018A4# => romdata <= X"6A3E2B3A";
    when 16#018A5# => romdata <= X"06493608";
    when 16#018A6# => romdata <= X"36493036";
    when 16#018A7# => romdata <= X"49597648";
    when 16#018A8# => romdata <= X"073C4281";
    when 16#018A9# => romdata <= X"81423C0A";
    when 16#018AA# => romdata <= X"041F040A";
    when 16#018AB# => romdata <= X"08083E08";
    when 16#018AC# => romdata <= X"08806008";
    when 16#018AD# => romdata <= X"080840C0";
    when 16#018AE# => romdata <= X"300C033E";
    when 16#018AF# => romdata <= X"4141413E";
    when 16#018B0# => romdata <= X"44427F40";
    when 16#018B1# => romdata <= X"40466151";
    when 16#018B2# => romdata <= X"49462241";
    when 16#018B3# => romdata <= X"49493618";
    when 16#018B4# => romdata <= X"14127F10";
    when 16#018B5# => romdata <= X"27454545";
    when 16#018B6# => romdata <= X"393E4949";
    when 16#018B7# => romdata <= X"49300101";
    when 16#018B8# => romdata <= X"710D0336";
    when 16#018B9# => romdata <= X"49494936";
    when 16#018BA# => romdata <= X"06494929";
    when 16#018BB# => romdata <= X"1E36D008";
    when 16#018BC# => romdata <= X"14224114";
    when 16#018BD# => romdata <= X"14141414";
    when 16#018BE# => romdata <= X"41221408";
    when 16#018BF# => romdata <= X"02510906";
    when 16#018C0# => romdata <= X"3C4299A5";
    when 16#018C1# => romdata <= X"BD421C7C";
    when 16#018C2# => romdata <= X"1211127C";
    when 16#018C3# => romdata <= X"7F494949";
    when 16#018C4# => romdata <= X"363E4141";
    when 16#018C5# => romdata <= X"41227F41";
    when 16#018C6# => romdata <= X"41413E7F";
    when 16#018C7# => romdata <= X"49494941";
    when 16#018C8# => romdata <= X"7F090909";
    when 16#018C9# => romdata <= X"013E4149";
    when 16#018CA# => romdata <= X"497A7F08";
    when 16#018CB# => romdata <= X"08087F41";
    when 16#018CC# => romdata <= X"7F414041";
    when 16#018CD# => romdata <= X"413F7F08";
    when 16#018CE# => romdata <= X"1422417F";
    when 16#018CF# => romdata <= X"40404040";
    when 16#018D0# => romdata <= X"7F060C06";
    when 16#018D1# => romdata <= X"7F7F0608";
    when 16#018D2# => romdata <= X"307F3E41";
    when 16#018D3# => romdata <= X"41413E7F";
    when 16#018D4# => romdata <= X"09090906";
    when 16#018D5# => romdata <= X"3E4161C1";
    when 16#018D6# => romdata <= X"BE7F0919";
    when 16#018D7# => romdata <= X"29462649";
    when 16#018D8# => romdata <= X"49493201";
    when 16#018D9# => romdata <= X"017F0101";
    when 16#018DA# => romdata <= X"3F404040";
    when 16#018DB# => romdata <= X"3F073840";
    when 16#018DC# => romdata <= X"38071F60";
    when 16#018DD# => romdata <= X"1F601F63";
    when 16#018DE# => romdata <= X"14081463";
    when 16#018DF# => romdata <= X"01067806";
    when 16#018E0# => romdata <= X"01615149";
    when 16#018E1# => romdata <= X"45437F41";
    when 16#018E2# => romdata <= X"41030C30";
    when 16#018E3# => romdata <= X"C041417F";
    when 16#018E4# => romdata <= X"04020102";
    when 16#018E5# => romdata <= X"04808080";
    when 16#018E6# => romdata <= X"80800102";
    when 16#018E7# => romdata <= X"20545454";
    when 16#018E8# => romdata <= X"787F4444";
    when 16#018E9# => romdata <= X"44383844";
    when 16#018EA# => romdata <= X"44443844";
    when 16#018EB# => romdata <= X"44447F38";
    when 16#018EC# => romdata <= X"54545458";
    when 16#018ED# => romdata <= X"087E0901";
    when 16#018EE# => romdata <= X"18A4A4A4";
    when 16#018EF# => romdata <= X"787F0404";
    when 16#018F0# => romdata <= X"787D807D";
    when 16#018F1# => romdata <= X"7F102844";
    when 16#018F2# => romdata <= X"3F407C04";
    when 16#018F3# => romdata <= X"7804787C";
    when 16#018F4# => romdata <= X"04047838";
    when 16#018F5# => romdata <= X"444438FC";
    when 16#018F6# => romdata <= X"24242418";
    when 16#018F7# => romdata <= X"18242424";
    when 16#018F8# => romdata <= X"FC7C0804";
    when 16#018F9# => romdata <= X"04485454";
    when 16#018FA# => romdata <= X"24043F44";
    when 16#018FB# => romdata <= X"403C4040";
    when 16#018FC# => romdata <= X"7C1C2040";
    when 16#018FD# => romdata <= X"201C1C60";
    when 16#018FE# => romdata <= X"601C6060";
    when 16#018FF# => romdata <= X"1C442810";
    when 16#01900# => romdata <= X"28449CA0";
    when 16#01901# => romdata <= X"601C6454";
    when 16#01902# => romdata <= X"544C187E";
    when 16#01903# => romdata <= X"8181FFFF";
    when 16#01904# => romdata <= X"81817E18";
    when 16#01905# => romdata <= X"18040810";
    when 16#01906# => romdata <= X"0C143E55";
    when 16#01907# => romdata <= X"55FF8181";
    when 16#01908# => romdata <= X"81FF8060";
    when 16#01909# => romdata <= X"80608060";
    when 16#0190A# => romdata <= X"60600060";
    when 16#0190B# => romdata <= X"60006060";
    when 16#0190C# => romdata <= X"047F0414";
    when 16#0190D# => romdata <= X"7F140201";
    when 16#0190E# => romdata <= X"01024629";
    when 16#0190F# => romdata <= X"1608344A";
    when 16#01910# => romdata <= X"31483000";
    when 16#01911# => romdata <= X"18243E41";
    when 16#01912# => romdata <= X"227F4941";
    when 16#01913# => romdata <= X"03040403";
    when 16#01914# => romdata <= X"03040304";
    when 16#01915# => romdata <= X"04030403";
    when 16#01916# => romdata <= X"183C3C18";
    when 16#01917# => romdata <= X"08080808";
    when 16#01918# => romdata <= X"03010203";
    when 16#01919# => romdata <= X"020E020E";
    when 16#0191A# => romdata <= X"060E0048";
    when 16#0191B# => romdata <= X"30384438";
    when 16#0191C# => romdata <= X"54483844";
    when 16#0191D# => romdata <= X"FE44487E";
    when 16#0191E# => romdata <= X"49014438";
    when 16#0191F# => romdata <= X"28384403";
    when 16#01920# => romdata <= X"147C1403";
    when 16#01921# => romdata <= X"E7E74E55";
    when 16#01922# => romdata <= X"55390101";
    when 16#01923# => romdata <= X"0001011C";
    when 16#01924# => romdata <= X"2A555522";
    when 16#01925# => romdata <= X"1C1D151E";
    when 16#01926# => romdata <= X"18240018";
    when 16#01927# => romdata <= X"24080808";
    when 16#01928# => romdata <= X"18080808";
    when 16#01929# => romdata <= X"3C42BD95";
    when 16#0192A# => romdata <= X"A9423C01";
    when 16#0192B# => romdata <= X"01010101";
    when 16#0192C# => romdata <= X"06090906";
    when 16#0192D# => romdata <= X"44445F44";
    when 16#0192E# => romdata <= X"44191512";
    when 16#0192F# => romdata <= X"15150A02";
    when 16#01930# => romdata <= X"01FC2020";
    when 16#01931# => romdata <= X"1C0E7F01";
    when 16#01932# => romdata <= X"7F011818";
    when 16#01933# => romdata <= X"00804002";
    when 16#01934# => romdata <= X"1F060909";
    when 16#01935# => romdata <= X"06241800";
    when 16#01936# => romdata <= X"2418824F";
    when 16#01937# => romdata <= X"304C62F1";
    when 16#01938# => romdata <= X"824F300C";
    when 16#01939# => romdata <= X"D2B1955F";
    when 16#0193A# => romdata <= X"304C62F1";
    when 16#0193B# => romdata <= X"30484520";
    when 16#0193C# => romdata <= X"60392E38";
    when 16#0193D# => romdata <= X"6060382E";
    when 16#0193E# => romdata <= X"3960701D";
    when 16#0193F# => romdata <= X"131D7072";
    when 16#01940# => romdata <= X"1D121E71";
    when 16#01941# => romdata <= X"701D121D";
    when 16#01942# => romdata <= X"70603B25";
    when 16#01943# => romdata <= X"3B607E11";
    when 16#01944# => romdata <= X"7F49411E";
    when 16#01945# => romdata <= X"2161927C";
    when 16#01946# => romdata <= X"5556447C";
    when 16#01947# => romdata <= X"5655447C";
    when 16#01948# => romdata <= X"5655467D";
    when 16#01949# => romdata <= X"54544545";
    when 16#0194A# => romdata <= X"7E44447E";
    when 16#0194B# => romdata <= X"45467D46";
    when 16#0194C# => romdata <= X"457C4508";
    when 16#0194D# => romdata <= X"7F49413E";
    when 16#0194E# => romdata <= X"7E091222";
    when 16#0194F# => romdata <= X"7D384546";
    when 16#01950# => romdata <= X"44383844";
    when 16#01951# => romdata <= X"46453838";
    when 16#01952# => romdata <= X"46454638";
    when 16#01953# => romdata <= X"3A454546";
    when 16#01954# => romdata <= X"39384544";
    when 16#01955# => romdata <= X"45382214";
    when 16#01956# => romdata <= X"081422BC";
    when 16#01957# => romdata <= X"625A463D";
    when 16#01958# => romdata <= X"3C41423C";
    when 16#01959# => romdata <= X"3C42413C";
    when 16#0195A# => romdata <= X"3C42413E";
    when 16#0195B# => romdata <= X"3D40403D";
    when 16#0195C# => romdata <= X"0608F209";
    when 16#0195D# => romdata <= X"067F2222";
    when 16#0195E# => romdata <= X"1CFE0989";
    when 16#0195F# => romdata <= X"76205556";
    when 16#01960# => romdata <= X"78205655";
    when 16#01961# => romdata <= X"78225555";
    when 16#01962# => romdata <= X"7A235556";
    when 16#01963# => romdata <= X"7B205554";
    when 16#01964# => romdata <= X"79275557";
    when 16#01965# => romdata <= X"78205438";
    when 16#01966# => romdata <= X"54483844";
    when 16#01967# => romdata <= X"C4385556";
    when 16#01968# => romdata <= X"58385655";
    when 16#01969# => romdata <= X"583A5555";
    when 16#0196A# => romdata <= X"5A395454";
    when 16#0196B# => romdata <= X"59017A7A";
    when 16#0196C# => romdata <= X"01027902";
    when 16#0196D# => romdata <= X"02780260";
    when 16#0196E# => romdata <= X"91927C7B";
    when 16#0196F# => romdata <= X"090A7338";
    when 16#01970# => romdata <= X"45463838";
    when 16#01971# => romdata <= X"4645383A";
    when 16#01972# => romdata <= X"45453A3B";
    when 16#01973# => romdata <= X"45463B39";
    when 16#01974# => romdata <= X"44443908";
    when 16#01975# => romdata <= X"082A0808";
    when 16#01976# => romdata <= X"B8644C3A";
    when 16#01977# => romdata <= X"3C41427C";
    when 16#01978# => romdata <= X"3C42417C";
    when 16#01979# => romdata <= X"3A41417A";
    when 16#0197A# => romdata <= X"3D40407D";
    when 16#0197B# => romdata <= X"986219FF";
    when 16#0197C# => romdata <= X"423C9A60";
    when 16#0197D# => romdata <= X"1A000000";
    when 16#0197E# => romdata <= X"30622020";
    when 16#0197F# => romdata <= X"20202020";
    when 16#01980# => romdata <= X"20202020";
    when 16#01981# => romdata <= X"20202020";
    when 16#01982# => romdata <= X"20202020";
    when 16#01983# => romdata <= X"20202020";
    when 16#01984# => romdata <= X"20202020";
    when 16#01985# => romdata <= X"20202020";
    when 16#01986# => romdata <= X"20200000";
    when 16#01987# => romdata <= X"20202020";
    when 16#01988# => romdata <= X"20202020";
    when 16#01989# => romdata <= X"00000000";
    when 16#0198A# => romdata <= X"00202020";
    when 16#0198B# => romdata <= X"20202020";
    when 16#0198C# => romdata <= X"20202828";
    when 16#0198D# => romdata <= X"28282820";
    when 16#0198E# => romdata <= X"20202020";
    when 16#0198F# => romdata <= X"20202020";
    when 16#01990# => romdata <= X"20202020";
    when 16#01991# => romdata <= X"20202020";
    when 16#01992# => romdata <= X"20881010";
    when 16#01993# => romdata <= X"10101010";
    when 16#01994# => romdata <= X"10101010";
    when 16#01995# => romdata <= X"10101010";
    when 16#01996# => romdata <= X"10040404";
    when 16#01997# => romdata <= X"04040404";
    when 16#01998# => romdata <= X"04040410";
    when 16#01999# => romdata <= X"10101010";
    when 16#0199A# => romdata <= X"10104141";
    when 16#0199B# => romdata <= X"41414141";
    when 16#0199C# => romdata <= X"01010101";
    when 16#0199D# => romdata <= X"01010101";
    when 16#0199E# => romdata <= X"01010101";
    when 16#0199F# => romdata <= X"01010101";
    when 16#019A0# => romdata <= X"01010101";
    when 16#019A1# => romdata <= X"10101010";
    when 16#019A2# => romdata <= X"10104242";
    when 16#019A3# => romdata <= X"42424242";
    when 16#019A4# => romdata <= X"02020202";
    when 16#019A5# => romdata <= X"02020202";
    when 16#019A6# => romdata <= X"02020202";
    when 16#019A7# => romdata <= X"02020202";
    when 16#019A8# => romdata <= X"02020202";
    when 16#019A9# => romdata <= X"10101010";
    when 16#019AA# => romdata <= X"20000000";
    when 16#019AB# => romdata <= X"00000000";
    when 16#019AC# => romdata <= X"00000000";
    when 16#019AD# => romdata <= X"00000000";
    when 16#019AE# => romdata <= X"00000000";
    when 16#019AF# => romdata <= X"00000000";
    when 16#019B0# => romdata <= X"00000000";
    when 16#019B1# => romdata <= X"00000000";
    when 16#019B2# => romdata <= X"00000000";
    when 16#019B3# => romdata <= X"00000000";
    when 16#019B4# => romdata <= X"00000000";
    when 16#019B5# => romdata <= X"00000000";
    when 16#019B6# => romdata <= X"00000000";
    when 16#019B7# => romdata <= X"00000000";
    when 16#019B8# => romdata <= X"00000000";
    when 16#019B9# => romdata <= X"00000000";
    when 16#019BA# => romdata <= X"00000000";
    when 16#019BB# => romdata <= X"00000000";
    when 16#019BC# => romdata <= X"00000000";
    when 16#019BD# => romdata <= X"00000000";
    when 16#019BE# => romdata <= X"00000000";
    when 16#019BF# => romdata <= X"00000000";
    when 16#019C0# => romdata <= X"00000000";
    when 16#019C1# => romdata <= X"00000000";
    when 16#019C2# => romdata <= X"00000000";
    when 16#019C3# => romdata <= X"00000000";
    when 16#019C4# => romdata <= X"00000000";
    when 16#019C5# => romdata <= X"00000000";
    when 16#019C6# => romdata <= X"00000000";
    when 16#019C7# => romdata <= X"00000000";
    when 16#019C8# => romdata <= X"00000000";
    when 16#019C9# => romdata <= X"00000000";
    when 16#019CA# => romdata <= X"00000000";
    when 16#019CB# => romdata <= X"43000000";
    when 16#019CC# => romdata <= X"00000000";
    when 16#019CD# => romdata <= X"80000C00";
    when 16#019CE# => romdata <= X"80000B00";
    when 16#019CF# => romdata <= X"80000800";
    when 16#019D0# => romdata <= X"00000000";
    when 16#019D1# => romdata <= X"FF000000";
    when 16#019D2# => romdata <= X"00000000";
    when 16#019D3# => romdata <= X"00000000";
    when 16#019D4# => romdata <= X"00FFFFFF";
    when 16#019D5# => romdata <= X"FF00FFFF";
    when 16#019D6# => romdata <= X"FFFF00FF";
    when 16#019D7# => romdata <= X"FFFFFF00";
    when 16#019D8# => romdata <= X"00000000";
    when 16#019D9# => romdata <= X"00000000";
    when 16#019DA# => romdata <= X"80000A00";
    when 16#019DB# => romdata <= X"80000700";
    when 16#019DC# => romdata <= X"80000600";
    when 16#019DD# => romdata <= X"80000400";
    when 16#019DE# => romdata <= X"80000200";
    when 16#019DF# => romdata <= X"80000100";
    when 16#019E0# => romdata <= X"80000004";
    when 16#019E1# => romdata <= X"80000000";
    when 16#019E2# => romdata <= X"0000678C";
    when 16#019E3# => romdata <= X"00000000";
    when 16#019E4# => romdata <= X"000069F4";
    when 16#019E5# => romdata <= X"00006A50";
    when 16#019E6# => romdata <= X"00006AAC";
    when 16#019E7# => romdata <= X"00000000";
    when 16#019E8# => romdata <= X"00000000";
    when 16#019E9# => romdata <= X"00000000";
    when 16#019EA# => romdata <= X"00000000";
    when 16#019EB# => romdata <= X"00000000";
    when 16#019EC# => romdata <= X"00000000";
    when 16#019ED# => romdata <= X"00000000";
    when 16#019EE# => romdata <= X"00000000";
    when 16#019EF# => romdata <= X"00000000";
    when 16#019F0# => romdata <= X"0000672C";
    when 16#019F1# => romdata <= X"00000000";
    when 16#019F2# => romdata <= X"00000000";
    when 16#019F3# => romdata <= X"00000000";
    when 16#019F4# => romdata <= X"00000000";
    when 16#019F5# => romdata <= X"00000000";
    when 16#019F6# => romdata <= X"00000000";
    when 16#019F7# => romdata <= X"00000000";
    when 16#019F8# => romdata <= X"00000000";
    when 16#019F9# => romdata <= X"00000000";
    when 16#019FA# => romdata <= X"00000000";
    when 16#019FB# => romdata <= X"00000000";
    when 16#019FC# => romdata <= X"00000000";
    when 16#019FD# => romdata <= X"00000000";
    when 16#019FE# => romdata <= X"00000000";
    when 16#019FF# => romdata <= X"00000000";
    when 16#01A00# => romdata <= X"00000000";
    when 16#01A01# => romdata <= X"00000000";
    when 16#01A02# => romdata <= X"00000000";
    when 16#01A03# => romdata <= X"00000000";
    when 16#01A04# => romdata <= X"00000000";
    when 16#01A05# => romdata <= X"00000000";
    when 16#01A06# => romdata <= X"00000000";
    when 16#01A07# => romdata <= X"00000000";
    when 16#01A08# => romdata <= X"00000000";
    when 16#01A09# => romdata <= X"00000000";
    when 16#01A0A# => romdata <= X"00000000";
    when 16#01A0B# => romdata <= X"00000000";
    when 16#01A0C# => romdata <= X"00000000";
    when 16#01A0D# => romdata <= X"00000001";
    when 16#01A0E# => romdata <= X"330EABCD";
    when 16#01A0F# => romdata <= X"1234E66D";
    when 16#01A10# => romdata <= X"DEEC0005";
    when 16#01A11# => romdata <= X"000B0000";
    when 16#01A12# => romdata <= X"00000000";
    when 16#01A13# => romdata <= X"00000000";
    when 16#01A14# => romdata <= X"00000000";
    when 16#01A15# => romdata <= X"00000000";
    when 16#01A16# => romdata <= X"00000000";
    when 16#01A17# => romdata <= X"00000000";
    when 16#01A18# => romdata <= X"00000000";
    when 16#01A19# => romdata <= X"00000000";
    when 16#01A1A# => romdata <= X"00000000";
    when 16#01A1B# => romdata <= X"00000000";
    when 16#01A1C# => romdata <= X"00000000";
    when 16#01A1D# => romdata <= X"00000000";
    when 16#01A1E# => romdata <= X"00000000";
    when 16#01A1F# => romdata <= X"00000000";
    when 16#01A20# => romdata <= X"00000000";
    when 16#01A21# => romdata <= X"00000000";
    when 16#01A22# => romdata <= X"00000000";
    when 16#01A23# => romdata <= X"00000000";
    when 16#01A24# => romdata <= X"00000000";
    when 16#01A25# => romdata <= X"00000000";
    when 16#01A26# => romdata <= X"00000000";
    when 16#01A27# => romdata <= X"00000000";
    when 16#01A28# => romdata <= X"00000000";
    when 16#01A29# => romdata <= X"00000000";
    when 16#01A2A# => romdata <= X"00000000";
    when 16#01A2B# => romdata <= X"00000000";
    when 16#01A2C# => romdata <= X"00000000";
    when 16#01A2D# => romdata <= X"00000000";
    when 16#01A2E# => romdata <= X"00000000";
    when 16#01A2F# => romdata <= X"00000000";
    when 16#01A30# => romdata <= X"00000000";
    when 16#01A31# => romdata <= X"00000000";
    when 16#01A32# => romdata <= X"00000000";
    when 16#01A33# => romdata <= X"00000000";
    when 16#01A34# => romdata <= X"00000000";
    when 16#01A35# => romdata <= X"00000000";
    when 16#01A36# => romdata <= X"00000000";
    when 16#01A37# => romdata <= X"00000000";
    when 16#01A38# => romdata <= X"00000000";
    when 16#01A39# => romdata <= X"00000000";
    when 16#01A3A# => romdata <= X"00000000";
    when 16#01A3B# => romdata <= X"00000000";
    when 16#01A3C# => romdata <= X"00000000";
    when 16#01A3D# => romdata <= X"00000000";
    when 16#01A3E# => romdata <= X"00000000";
    when 16#01A3F# => romdata <= X"00000000";
    when 16#01A40# => romdata <= X"00000000";
    when 16#01A41# => romdata <= X"00000000";
    when 16#01A42# => romdata <= X"00000000";
    when 16#01A43# => romdata <= X"00000000";
    when 16#01A44# => romdata <= X"00000000";
    when 16#01A45# => romdata <= X"00000000";
    when 16#01A46# => romdata <= X"00000000";
    when 16#01A47# => romdata <= X"00000000";
    when 16#01A48# => romdata <= X"00000000";
    when 16#01A49# => romdata <= X"00000000";
    when 16#01A4A# => romdata <= X"00000000";
    when 16#01A4B# => romdata <= X"00000000";
    when 16#01A4C# => romdata <= X"00000000";
    when 16#01A4D# => romdata <= X"00000000";
    when 16#01A4E# => romdata <= X"00000000";
    when 16#01A4F# => romdata <= X"00000000";
    when 16#01A50# => romdata <= X"00000000";
    when 16#01A51# => romdata <= X"00000000";
    when 16#01A52# => romdata <= X"00000000";
    when 16#01A53# => romdata <= X"00000000";
    when 16#01A54# => romdata <= X"00000000";
    when 16#01A55# => romdata <= X"00000000";
    when 16#01A56# => romdata <= X"00000000";
    when 16#01A57# => romdata <= X"00000000";
    when 16#01A58# => romdata <= X"00000000";
    when 16#01A59# => romdata <= X"00000000";
    when 16#01A5A# => romdata <= X"00000000";
    when 16#01A5B# => romdata <= X"00000000";
    when 16#01A5C# => romdata <= X"00000000";
    when 16#01A5D# => romdata <= X"00000000";
    when 16#01A5E# => romdata <= X"00000000";
    when 16#01A5F# => romdata <= X"00000000";
    when 16#01A60# => romdata <= X"00000000";
    when 16#01A61# => romdata <= X"00000000";
    when 16#01A62# => romdata <= X"00000000";
    when 16#01A63# => romdata <= X"00000000";
    when 16#01A64# => romdata <= X"00000000";
    when 16#01A65# => romdata <= X"00000000";
    when 16#01A66# => romdata <= X"00000000";
    when 16#01A67# => romdata <= X"00000000";
    when 16#01A68# => romdata <= X"00000000";
    when 16#01A69# => romdata <= X"00000000";
    when 16#01A6A# => romdata <= X"00000000";
    when 16#01A6B# => romdata <= X"00000000";
    when 16#01A6C# => romdata <= X"00000000";
    when 16#01A6D# => romdata <= X"00000000";
    when 16#01A6E# => romdata <= X"00000000";
    when 16#01A6F# => romdata <= X"00000000";
    when 16#01A70# => romdata <= X"00000000";
    when 16#01A71# => romdata <= X"00000000";
    when 16#01A72# => romdata <= X"00000000";
    when 16#01A73# => romdata <= X"00000000";
    when 16#01A74# => romdata <= X"00000000";
    when 16#01A75# => romdata <= X"00000000";
    when 16#01A76# => romdata <= X"00000000";
    when 16#01A77# => romdata <= X"00000000";
    when 16#01A78# => romdata <= X"00000000";
    when 16#01A79# => romdata <= X"00000000";
    when 16#01A7A# => romdata <= X"00000000";
    when 16#01A7B# => romdata <= X"00000000";
    when 16#01A7C# => romdata <= X"00000000";
    when 16#01A7D# => romdata <= X"00000000";
    when 16#01A7E# => romdata <= X"00000000";
    when 16#01A7F# => romdata <= X"00000000";
    when 16#01A80# => romdata <= X"00000000";
    when 16#01A81# => romdata <= X"00000000";
    when 16#01A82# => romdata <= X"00000000";
    when 16#01A83# => romdata <= X"00000000";
    when 16#01A84# => romdata <= X"00000000";
    when 16#01A85# => romdata <= X"00000000";
    when 16#01A86# => romdata <= X"00000000";
    when 16#01A87# => romdata <= X"00000000";
    when 16#01A88# => romdata <= X"00000000";
    when 16#01A89# => romdata <= X"00000000";
    when 16#01A8A# => romdata <= X"00000000";
    when 16#01A8B# => romdata <= X"00000000";
    when 16#01A8C# => romdata <= X"00000000";
    when 16#01A8D# => romdata <= X"00000000";
    when 16#01A8E# => romdata <= X"00000000";
    when 16#01A8F# => romdata <= X"00000000";
    when 16#01A90# => romdata <= X"00000000";
    when 16#01A91# => romdata <= X"00000000";
    when 16#01A92# => romdata <= X"00000000";
    when 16#01A93# => romdata <= X"00000000";
    when 16#01A94# => romdata <= X"00000000";
    when 16#01A95# => romdata <= X"00000000";
    when 16#01A96# => romdata <= X"00000000";
    when 16#01A97# => romdata <= X"00000000";
    when 16#01A98# => romdata <= X"00000000";
    when 16#01A99# => romdata <= X"00000000";
    when 16#01A9A# => romdata <= X"00000000";
    when 16#01A9B# => romdata <= X"00000000";
    when 16#01A9C# => romdata <= X"00000000";
    when 16#01A9D# => romdata <= X"00000000";
    when 16#01A9E# => romdata <= X"00000000";
    when 16#01A9F# => romdata <= X"00000000";
    when 16#01AA0# => romdata <= X"00000000";
    when 16#01AA1# => romdata <= X"00000000";
    when 16#01AA2# => romdata <= X"00000000";
    when 16#01AA3# => romdata <= X"00000000";
    when 16#01AA4# => romdata <= X"00000000";
    when 16#01AA5# => romdata <= X"00000000";
    when 16#01AA6# => romdata <= X"00000000";
    when 16#01AA7# => romdata <= X"00000000";
    when 16#01AA8# => romdata <= X"00000000";
    when 16#01AA9# => romdata <= X"00000000";
    when 16#01AAA# => romdata <= X"00000000";
    when 16#01AAB# => romdata <= X"00000000";
    when 16#01AAC# => romdata <= X"00000000";
    when 16#01AAD# => romdata <= X"00000000";
    when 16#01AAE# => romdata <= X"00000000";
    when 16#01AAF# => romdata <= X"00000000";
    when 16#01AB0# => romdata <= X"00000000";
    when 16#01AB1# => romdata <= X"00000000";
    when 16#01AB2# => romdata <= X"00000000";
    when 16#01AB3# => romdata <= X"00000000";
    when 16#01AB4# => romdata <= X"00000000";
    when 16#01AB5# => romdata <= X"00000000";
    when 16#01AB6# => romdata <= X"00000000";
    when 16#01AB7# => romdata <= X"00000000";
    when 16#01AB8# => romdata <= X"00000000";
    when 16#01AB9# => romdata <= X"00000000";
    when 16#01ABA# => romdata <= X"00000000";
    when 16#01ABB# => romdata <= X"00000000";
    when 16#01ABC# => romdata <= X"00000000";
    when 16#01ABD# => romdata <= X"00000000";
    when 16#01ABE# => romdata <= X"00000000";
    when 16#01ABF# => romdata <= X"00000000";
    when 16#01AC0# => romdata <= X"00000000";
    when 16#01AC1# => romdata <= X"00000000";
    when 16#01AC2# => romdata <= X"00000000";
    when 16#01AC3# => romdata <= X"00000000";
    when 16#01AC4# => romdata <= X"00000000";
    when 16#01AC5# => romdata <= X"00000000";
    when 16#01AC6# => romdata <= X"00000000";
    when 16#01AC7# => romdata <= X"00000000";
    when 16#01AC8# => romdata <= X"00000000";
    when 16#01AC9# => romdata <= X"00000000";
    when 16#01ACA# => romdata <= X"00000000";
    when 16#01ACB# => romdata <= X"00000000";
    when 16#01ACC# => romdata <= X"00000000";
    when 16#01ACD# => romdata <= X"00000000";
    when 16#01ACE# => romdata <= X"FFFFFFFF";
    when 16#01ACF# => romdata <= X"00000000";
    when 16#01AD0# => romdata <= X"00020000";
    when 16#01AD1# => romdata <= X"00000000";
    when 16#01AD2# => romdata <= X"00000000";
    when 16#01AD3# => romdata <= X"00006B44";
    when 16#01AD4# => romdata <= X"00006B44";
    when 16#01AD5# => romdata <= X"00006B4C";
    when 16#01AD6# => romdata <= X"00006B4C";
    when 16#01AD7# => romdata <= X"00006B54";
    when 16#01AD8# => romdata <= X"00006B54";
    when 16#01AD9# => romdata <= X"00006B5C";
    when 16#01ADA# => romdata <= X"00006B5C";
    when 16#01ADB# => romdata <= X"00006B64";
    when 16#01ADC# => romdata <= X"00006B64";
    when 16#01ADD# => romdata <= X"00006B6C";
    when 16#01ADE# => romdata <= X"00006B6C";
    when 16#01ADF# => romdata <= X"00006B74";
    when 16#01AE0# => romdata <= X"00006B74";
    when 16#01AE1# => romdata <= X"00006B7C";
    when 16#01AE2# => romdata <= X"00006B7C";
    when 16#01AE3# => romdata <= X"00006B84";
    when 16#01AE4# => romdata <= X"00006B84";
    when 16#01AE5# => romdata <= X"00006B8C";
    when 16#01AE6# => romdata <= X"00006B8C";
    when 16#01AE7# => romdata <= X"00006B94";
    when 16#01AE8# => romdata <= X"00006B94";
    when 16#01AE9# => romdata <= X"00006B9C";
    when 16#01AEA# => romdata <= X"00006B9C";
    when 16#01AEB# => romdata <= X"00006BA4";
    when 16#01AEC# => romdata <= X"00006BA4";
    when 16#01AED# => romdata <= X"00006BAC";
    when 16#01AEE# => romdata <= X"00006BAC";
    when 16#01AEF# => romdata <= X"00006BB4";
    when 16#01AF0# => romdata <= X"00006BB4";
    when 16#01AF1# => romdata <= X"00006BBC";
    when 16#01AF2# => romdata <= X"00006BBC";
    when 16#01AF3# => romdata <= X"00006BC4";
    when 16#01AF4# => romdata <= X"00006BC4";
    when 16#01AF5# => romdata <= X"00006BCC";
    when 16#01AF6# => romdata <= X"00006BCC";
    when 16#01AF7# => romdata <= X"00006BD4";
    when 16#01AF8# => romdata <= X"00006BD4";
    when 16#01AF9# => romdata <= X"00006BDC";
    when 16#01AFA# => romdata <= X"00006BDC";
    when 16#01AFB# => romdata <= X"00006BE4";
    when 16#01AFC# => romdata <= X"00006BE4";
    when 16#01AFD# => romdata <= X"00006BEC";
    when 16#01AFE# => romdata <= X"00006BEC";
    when 16#01AFF# => romdata <= X"00006BF4";
    when 16#01B00# => romdata <= X"00006BF4";
    when 16#01B01# => romdata <= X"00006BFC";
    when 16#01B02# => romdata <= X"00006BFC";
    when 16#01B03# => romdata <= X"00006C04";
    when 16#01B04# => romdata <= X"00006C04";
    when 16#01B05# => romdata <= X"00006C0C";
    when 16#01B06# => romdata <= X"00006C0C";
    when 16#01B07# => romdata <= X"00006C14";
    when 16#01B08# => romdata <= X"00006C14";
    when 16#01B09# => romdata <= X"00006C1C";
    when 16#01B0A# => romdata <= X"00006C1C";
    when 16#01B0B# => romdata <= X"00006C24";
    when 16#01B0C# => romdata <= X"00006C24";
    when 16#01B0D# => romdata <= X"00006C2C";
    when 16#01B0E# => romdata <= X"00006C2C";
    when 16#01B0F# => romdata <= X"00006C34";
    when 16#01B10# => romdata <= X"00006C34";
    when 16#01B11# => romdata <= X"00006C3C";
    when 16#01B12# => romdata <= X"00006C3C";
    when 16#01B13# => romdata <= X"00006C44";
    when 16#01B14# => romdata <= X"00006C44";
    when 16#01B15# => romdata <= X"00006C4C";
    when 16#01B16# => romdata <= X"00006C4C";
    when 16#01B17# => romdata <= X"00006C54";
    when 16#01B18# => romdata <= X"00006C54";
    when 16#01B19# => romdata <= X"00006C5C";
    when 16#01B1A# => romdata <= X"00006C5C";
    when 16#01B1B# => romdata <= X"00006C64";
    when 16#01B1C# => romdata <= X"00006C64";
    when 16#01B1D# => romdata <= X"00006C6C";
    when 16#01B1E# => romdata <= X"00006C6C";
    when 16#01B1F# => romdata <= X"00006C74";
    when 16#01B20# => romdata <= X"00006C74";
    when 16#01B21# => romdata <= X"00006C7C";
    when 16#01B22# => romdata <= X"00006C7C";
    when 16#01B23# => romdata <= X"00006C84";
    when 16#01B24# => romdata <= X"00006C84";
    when 16#01B25# => romdata <= X"00006C8C";
    when 16#01B26# => romdata <= X"00006C8C";
    when 16#01B27# => romdata <= X"00006C94";
    when 16#01B28# => romdata <= X"00006C94";
    when 16#01B29# => romdata <= X"00006C9C";
    when 16#01B2A# => romdata <= X"00006C9C";
    when 16#01B2B# => romdata <= X"00006CA4";
    when 16#01B2C# => romdata <= X"00006CA4";
    when 16#01B2D# => romdata <= X"00006CAC";
    when 16#01B2E# => romdata <= X"00006CAC";
    when 16#01B2F# => romdata <= X"00006CB4";
    when 16#01B30# => romdata <= X"00006CB4";
    when 16#01B31# => romdata <= X"00006CBC";
    when 16#01B32# => romdata <= X"00006CBC";
    when 16#01B33# => romdata <= X"00006CC4";
    when 16#01B34# => romdata <= X"00006CC4";
    when 16#01B35# => romdata <= X"00006CCC";
    when 16#01B36# => romdata <= X"00006CCC";
    when 16#01B37# => romdata <= X"00006CD4";
    when 16#01B38# => romdata <= X"00006CD4";
    when 16#01B39# => romdata <= X"00006CDC";
    when 16#01B3A# => romdata <= X"00006CDC";
    when 16#01B3B# => romdata <= X"00006CE4";
    when 16#01B3C# => romdata <= X"00006CE4";
    when 16#01B3D# => romdata <= X"00006CEC";
    when 16#01B3E# => romdata <= X"00006CEC";
    when 16#01B3F# => romdata <= X"00006CF4";
    when 16#01B40# => romdata <= X"00006CF4";
    when 16#01B41# => romdata <= X"00006CFC";
    when 16#01B42# => romdata <= X"00006CFC";
    when 16#01B43# => romdata <= X"00006D04";
    when 16#01B44# => romdata <= X"00006D04";
    when 16#01B45# => romdata <= X"00006D0C";
    when 16#01B46# => romdata <= X"00006D0C";
    when 16#01B47# => romdata <= X"00006D14";
    when 16#01B48# => romdata <= X"00006D14";
    when 16#01B49# => romdata <= X"00006D1C";
    when 16#01B4A# => romdata <= X"00006D1C";
    when 16#01B4B# => romdata <= X"00006D24";
    when 16#01B4C# => romdata <= X"00006D24";
    when 16#01B4D# => romdata <= X"00006D2C";
    when 16#01B4E# => romdata <= X"00006D2C";
    when 16#01B4F# => romdata <= X"00006D34";
    when 16#01B50# => romdata <= X"00006D34";
    when 16#01B51# => romdata <= X"00006D3C";
    when 16#01B52# => romdata <= X"00006D3C";
    when 16#01B53# => romdata <= X"00006D44";
    when 16#01B54# => romdata <= X"00006D44";
    when 16#01B55# => romdata <= X"00006D4C";
    when 16#01B56# => romdata <= X"00006D4C";
    when 16#01B57# => romdata <= X"00006D54";
    when 16#01B58# => romdata <= X"00006D54";
    when 16#01B59# => romdata <= X"00006D5C";
    when 16#01B5A# => romdata <= X"00006D5C";
    when 16#01B5B# => romdata <= X"00006D64";
    when 16#01B5C# => romdata <= X"00006D64";
    when 16#01B5D# => romdata <= X"00006D6C";
    when 16#01B5E# => romdata <= X"00006D6C";
    when 16#01B5F# => romdata <= X"00006D74";
    when 16#01B60# => romdata <= X"00006D74";
    when 16#01B61# => romdata <= X"00006D7C";
    when 16#01B62# => romdata <= X"00006D7C";
    when 16#01B63# => romdata <= X"00006D84";
    when 16#01B64# => romdata <= X"00006D84";
    when 16#01B65# => romdata <= X"00006D8C";
    when 16#01B66# => romdata <= X"00006D8C";
    when 16#01B67# => romdata <= X"00006D94";
    when 16#01B68# => romdata <= X"00006D94";
    when 16#01B69# => romdata <= X"00006D9C";
    when 16#01B6A# => romdata <= X"00006D9C";
    when 16#01B6B# => romdata <= X"00006DA4";
    when 16#01B6C# => romdata <= X"00006DA4";
    when 16#01B6D# => romdata <= X"00006DAC";
    when 16#01B6E# => romdata <= X"00006DAC";
    when 16#01B6F# => romdata <= X"00006DB4";
    when 16#01B70# => romdata <= X"00006DB4";
    when 16#01B71# => romdata <= X"00006DBC";
    when 16#01B72# => romdata <= X"00006DBC";
    when 16#01B73# => romdata <= X"00006DC4";
    when 16#01B74# => romdata <= X"00006DC4";
    when 16#01B75# => romdata <= X"00006DCC";
    when 16#01B76# => romdata <= X"00006DCC";
    when 16#01B77# => romdata <= X"00006DD4";
    when 16#01B78# => romdata <= X"00006DD4";
    when 16#01B79# => romdata <= X"00006DDC";
    when 16#01B7A# => romdata <= X"00006DDC";
    when 16#01B7B# => romdata <= X"00006DE4";
    when 16#01B7C# => romdata <= X"00006DE4";
    when 16#01B7D# => romdata <= X"00006DEC";
    when 16#01B7E# => romdata <= X"00006DEC";
    when 16#01B7F# => romdata <= X"00006DF4";
    when 16#01B80# => romdata <= X"00006DF4";
    when 16#01B81# => romdata <= X"00006DFC";
    when 16#01B82# => romdata <= X"00006DFC";
    when 16#01B83# => romdata <= X"00006E04";
    when 16#01B84# => romdata <= X"00006E04";
    when 16#01B85# => romdata <= X"00006E0C";
    when 16#01B86# => romdata <= X"00006E0C";
    when 16#01B87# => romdata <= X"00006E14";
    when 16#01B88# => romdata <= X"00006E14";
    when 16#01B89# => romdata <= X"00006E1C";
    when 16#01B8A# => romdata <= X"00006E1C";
    when 16#01B8B# => romdata <= X"00006E24";
    when 16#01B8C# => romdata <= X"00006E24";
    when 16#01B8D# => romdata <= X"00006E2C";
    when 16#01B8E# => romdata <= X"00006E2C";
    when 16#01B8F# => romdata <= X"00006E34";
    when 16#01B90# => romdata <= X"00006E34";
    when 16#01B91# => romdata <= X"00006E3C";
    when 16#01B92# => romdata <= X"00006E3C";
    when 16#01B93# => romdata <= X"00006E44";
    when 16#01B94# => romdata <= X"00006E44";
    when 16#01B95# => romdata <= X"00006E4C";
    when 16#01B96# => romdata <= X"00006E4C";
    when 16#01B97# => romdata <= X"00006E54";
    when 16#01B98# => romdata <= X"00006E54";
    when 16#01B99# => romdata <= X"00006E5C";
    when 16#01B9A# => romdata <= X"00006E5C";
    when 16#01B9B# => romdata <= X"00006E64";
    when 16#01B9C# => romdata <= X"00006E64";
    when 16#01B9D# => romdata <= X"00006E6C";
    when 16#01B9E# => romdata <= X"00006E6C";
    when 16#01B9F# => romdata <= X"00006E74";
    when 16#01BA0# => romdata <= X"00006E74";
    when 16#01BA1# => romdata <= X"00006E7C";
    when 16#01BA2# => romdata <= X"00006E7C";
    when 16#01BA3# => romdata <= X"00006E84";
    when 16#01BA4# => romdata <= X"00006E84";
    when 16#01BA5# => romdata <= X"00006E8C";
    when 16#01BA6# => romdata <= X"00006E8C";
    when 16#01BA7# => romdata <= X"00006E94";
    when 16#01BA8# => romdata <= X"00006E94";
    when 16#01BA9# => romdata <= X"00006E9C";
    when 16#01BAA# => romdata <= X"00006E9C";
    when 16#01BAB# => romdata <= X"00006EA4";
    when 16#01BAC# => romdata <= X"00006EA4";
    when 16#01BAD# => romdata <= X"00006EAC";
    when 16#01BAE# => romdata <= X"00006EAC";
    when 16#01BAF# => romdata <= X"00006EB4";
    when 16#01BB0# => romdata <= X"00006EB4";
    when 16#01BB1# => romdata <= X"00006EBC";
    when 16#01BB2# => romdata <= X"00006EBC";
    when 16#01BB3# => romdata <= X"00006EC4";
    when 16#01BB4# => romdata <= X"00006EC4";
    when 16#01BB5# => romdata <= X"00006ECC";
    when 16#01BB6# => romdata <= X"00006ECC";
    when 16#01BB7# => romdata <= X"00006ED4";
    when 16#01BB8# => romdata <= X"00006ED4";
    when 16#01BB9# => romdata <= X"00006EDC";
    when 16#01BBA# => romdata <= X"00006EDC";
    when 16#01BBB# => romdata <= X"00006EE4";
    when 16#01BBC# => romdata <= X"00006EE4";
    when 16#01BBD# => romdata <= X"00006EEC";
    when 16#01BBE# => romdata <= X"00006EEC";
    when 16#01BBF# => romdata <= X"00006EF4";
    when 16#01BC0# => romdata <= X"00006EF4";
    when 16#01BC1# => romdata <= X"00006EFC";
    when 16#01BC2# => romdata <= X"00006EFC";
    when 16#01BC3# => romdata <= X"00006F04";
    when 16#01BC4# => romdata <= X"00006F04";
    when 16#01BC5# => romdata <= X"00006F0C";
    when 16#01BC6# => romdata <= X"00006F0C";
    when 16#01BC7# => romdata <= X"00006F14";
    when 16#01BC8# => romdata <= X"00006F14";
    when 16#01BC9# => romdata <= X"00006F1C";
    when 16#01BCA# => romdata <= X"00006F1C";
    when 16#01BCB# => romdata <= X"00006F24";
    when 16#01BCC# => romdata <= X"00006F24";
    when 16#01BCD# => romdata <= X"00006F2C";
    when 16#01BCE# => romdata <= X"00006F2C";
    when 16#01BCF# => romdata <= X"00006F34";
    when 16#01BD0# => romdata <= X"00006F34";
    when 16#01BD1# => romdata <= X"00006F3C";
    when 16#01BD2# => romdata <= X"00006F3C";
    when 16#01BD3# => romdata <= X"00006F3C";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
