-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
	--others => x"00dead00" -- mask for mem check
	others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
