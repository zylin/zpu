-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80d9800c",
     3 => x"3a0b0b80",
     4 => x"d0c70400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0b89",
     9 => x"90040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80d8",
   162 => x"ec738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0b88",
   169 => x"f8040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0b88",
   177 => x"e0040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80d8fc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82c23f80",
   257 => x"cab13f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80088408",
   281 => x"88087575",
   282 => x"b0d32d50",
   283 => x"50800856",
   284 => x"880c840c",
   285 => x"800c5104",
   286 => x"80088408",
   287 => x"88087575",
   288 => x"afa12d50",
   289 => x"50800856",
   290 => x"880c840c",
   291 => x"800c5104",
   292 => x"80088408",
   293 => x"880880d1",
   294 => x"902d880c",
   295 => x"840c800c",
   296 => x"0480d8fc",
   297 => x"08802ea4",
   298 => x"3880d980",
   299 => x"08822ebd",
   300 => x"38838080",
   301 => x"0b0b0b80",
   302 => x"e9800c82",
   303 => x"a0800b80",
   304 => x"e9840c82",
   305 => x"90800b80",
   306 => x"e9880c04",
   307 => x"f8808080",
   308 => x"a40b0b0b",
   309 => x"80e9800c",
   310 => x"f8808082",
   311 => x"800b80e9",
   312 => x"840cf880",
   313 => x"8084800b",
   314 => x"80e9880c",
   315 => x"0480c0a8",
   316 => x"808c0b0b",
   317 => x"0b80e980",
   318 => x"0c80c0a8",
   319 => x"80940b80",
   320 => x"e9840c0b",
   321 => x"0b80d2e4",
   322 => x"0b80e988",
   323 => x"0c04ff3d",
   324 => x"0d80e98c",
   325 => x"335170a7",
   326 => x"3880d988",
   327 => x"08700852",
   328 => x"5270802e",
   329 => x"94388412",
   330 => x"80d9880c",
   331 => x"702d80d9",
   332 => x"88087008",
   333 => x"525270ee",
   334 => x"38810b80",
   335 => x"e98c3483",
   336 => x"3d0d0404",
   337 => x"803d0d0b",
   338 => x"0b80e8fc",
   339 => x"08802e8e",
   340 => x"380b0b0b",
   341 => x"0b800b80",
   342 => x"2e098106",
   343 => x"8538823d",
   344 => x"0d040b0b",
   345 => x"80e8fc51",
   346 => x"0b0b0bf5",
   347 => x"933f823d",
   348 => x"0d0404fd",
   349 => x"3d0d80d9",
   350 => x"94088811",
   351 => x"0883de80",
   352 => x"0788120c",
   353 => x"841108fc",
   354 => x"a1ff0684",
   355 => x"120c538f",
   356 => x"51a0df3f",
   357 => x"80d99408",
   358 => x"841108e1",
   359 => x"ff068412",
   360 => x"0c841108",
   361 => x"86800784",
   362 => x"120c8411",
   363 => x"0880c080",
   364 => x"0784120c",
   365 => x"538151a0",
   366 => x"943f80d9",
   367 => x"94088411",
   368 => x"08ffbfff",
   369 => x"0684120c",
   370 => x"538551a0",
   371 => x"a53f80d9",
   372 => x"94088411",
   373 => x"0880c080",
   374 => x"0784120c",
   375 => x"5381519f",
   376 => x"ec3f80d9",
   377 => x"94088411",
   378 => x"08ffbfff",
   379 => x"0684120c",
   380 => x"5381519f",
   381 => x"fd3f80d9",
   382 => x"94088411",
   383 => x"0880c080",
   384 => x"0784120c",
   385 => x"5381519f",
   386 => x"c43f80d9",
   387 => x"94088411",
   388 => x"08ffbfff",
   389 => x"0684120c",
   390 => x"5381519f",
   391 => x"d53f80d9",
   392 => x"94088411",
   393 => x"08e1ff06",
   394 => x"84120c53",
   395 => x"84800b84",
   396 => x"14087072",
   397 => x"0784160c",
   398 => x"53841408",
   399 => x"7080c080",
   400 => x"0784160c",
   401 => x"53548151",
   402 => x"9f833f80",
   403 => x"d9940884",
   404 => x"110870ff",
   405 => x"bfff0684",
   406 => x"130c5353",
   407 => x"85519f92",
   408 => x"3f80d994",
   409 => x"08841108",
   410 => x"70feffff",
   411 => x"0684130c",
   412 => x"53841108",
   413 => x"70e1ff06",
   414 => x"84130c53",
   415 => x"84110870",
   416 => x"76078413",
   417 => x"0c538411",
   418 => x"0880c080",
   419 => x"0784120c",
   420 => x"5381519e",
   421 => x"b83f80d9",
   422 => x"94088411",
   423 => x"08ffbfff",
   424 => x"0684120c",
   425 => x"841108e1",
   426 => x"ff068412",
   427 => x"0c841108",
   428 => x"90800784",
   429 => x"120c8411",
   430 => x"0880c080",
   431 => x"0784120c",
   432 => x"5481519e",
   433 => x"883f80d9",
   434 => x"94088411",
   435 => x"08ffbfff",
   436 => x"0684120c",
   437 => x"54aa519d",
   438 => x"f43f80d9",
   439 => x"94088411",
   440 => x"08feffff",
   441 => x"0684120c",
   442 => x"841108e1",
   443 => x"ff068412",
   444 => x"0c841108",
   445 => x"84120c84",
   446 => x"110880c0",
   447 => x"80078412",
   448 => x"0c548151",
   449 => x"9dc73f80",
   450 => x"d9940884",
   451 => x"1108ffbf",
   452 => x"ff068412",
   453 => x"0c841108",
   454 => x"e1ff0684",
   455 => x"120c8411",
   456 => x"08988007",
   457 => x"84120c84",
   458 => x"110880c0",
   459 => x"80078412",
   460 => x"0c548151",
   461 => x"9d973f80",
   462 => x"d9940884",
   463 => x"1108ffbf",
   464 => x"ff068412",
   465 => x"0c54aa51",
   466 => x"9d833f80",
   467 => x"d9940884",
   468 => x"1108feff",
   469 => x"ff068412",
   470 => x"0c841108",
   471 => x"e1ff0684",
   472 => x"120c8411",
   473 => x"0884120c",
   474 => x"84110880",
   475 => x"c0800784",
   476 => x"120c5481",
   477 => x"519cd63f",
   478 => x"80d99408",
   479 => x"841108ff",
   480 => x"bfff0684",
   481 => x"120c8411",
   482 => x"08e1ff06",
   483 => x"84120c84",
   484 => x"11088c80",
   485 => x"0784120c",
   486 => x"84110880",
   487 => x"c0800784",
   488 => x"120c5481",
   489 => x"519ca63f",
   490 => x"80d99408",
   491 => x"841108ff",
   492 => x"bfff0684",
   493 => x"120c54aa",
   494 => x"519c923f",
   495 => x"810b80d9",
   496 => x"94088411",
   497 => x"0870feff",
   498 => x"ff068413",
   499 => x"0c548411",
   500 => x"0870e1ff",
   501 => x"0684130c",
   502 => x"54841108",
   503 => x"84120c84",
   504 => x"11087080",
   505 => x"c0800784",
   506 => x"130c5454",
   507 => x"7052549b",
   508 => x"dc3f80d9",
   509 => x"94088411",
   510 => x"0870ffbf",
   511 => x"ff068413",
   512 => x"0c538411",
   513 => x"0870e1ff",
   514 => x"0684130c",
   515 => x"53841108",
   516 => x"70828007",
   517 => x"84130c53",
   518 => x"84110870",
   519 => x"80c08007",
   520 => x"84130c53",
   521 => x"5373519b",
   522 => x"a43f80d9",
   523 => x"94088411",
   524 => x"08ffbfff",
   525 => x"0684120c",
   526 => x"53aa519b",
   527 => x"903f8251",
   528 => x"9bb03f85",
   529 => x"3d0d04fc",
   530 => x"3d0d029b",
   531 => x"05330284",
   532 => x"059f0533",
   533 => x"54527282",
   534 => x"2e81ad38",
   535 => x"82732591",
   536 => x"3872832e",
   537 => x"83bc3872",
   538 => x"842e82a9",
   539 => x"38863d0d",
   540 => x"0472812e",
   541 => x"098106f5",
   542 => x"38ff8012",
   543 => x"7081ff06",
   544 => x"80d99408",
   545 => x"841108fe",
   546 => x"ffff0684",
   547 => x"120c8411",
   548 => x"08e1ff06",
   549 => x"84120c71",
   550 => x"842b9e80",
   551 => x"06841208",
   552 => x"70720784",
   553 => x"140c5484",
   554 => x"120880c0",
   555 => x"80078413",
   556 => x"0c575556",
   557 => x"5281519a",
   558 => x"943f80d9",
   559 => x"94088411",
   560 => x"08ffbfff",
   561 => x"0684120c",
   562 => x"841108e1",
   563 => x"ff068412",
   564 => x"0c75882b",
   565 => x"9e800684",
   566 => x"12087107",
   567 => x"84130c84",
   568 => x"120880c0",
   569 => x"80078413",
   570 => x"0c555381",
   571 => x"5199de3f",
   572 => x"80d99408",
   573 => x"841108ff",
   574 => x"bfff0684",
   575 => x"120c53aa",
   576 => x"5199ca3f",
   577 => x"863d0d04",
   578 => x"c0127081",
   579 => x"ff0680d9",
   580 => x"94088411",
   581 => x"08feffff",
   582 => x"0684120c",
   583 => x"841108e1",
   584 => x"ff068412",
   585 => x"0c71842b",
   586 => x"9e800684",
   587 => x"12087072",
   588 => x"0784140c",
   589 => x"54841208",
   590 => x"80c08007",
   591 => x"84130c57",
   592 => x"55565281",
   593 => x"5199863f",
   594 => x"80d99408",
   595 => x"841108ff",
   596 => x"bfff0684",
   597 => x"120c8411",
   598 => x"08e1ff06",
   599 => x"84120c75",
   600 => x"882b9e80",
   601 => x"06841208",
   602 => x"71078413",
   603 => x"0c841208",
   604 => x"80c08007",
   605 => x"84130c55",
   606 => x"53815198",
   607 => x"d03f80d9",
   608 => x"94088411",
   609 => x"08ffbfff",
   610 => x"0684120c",
   611 => x"53aa5198",
   612 => x"bc3ffef0",
   613 => x"39d01270",
   614 => x"81ff0680",
   615 => x"d9940884",
   616 => x"1108feff",
   617 => x"ff068412",
   618 => x"0c841108",
   619 => x"e1ff0684",
   620 => x"120c7184",
   621 => x"2b9e8006",
   622 => x"84120870",
   623 => x"72078414",
   624 => x"0c548412",
   625 => x"0880c080",
   626 => x"0784130c",
   627 => x"57555652",
   628 => x"815197f9",
   629 => x"3f80d994",
   630 => x"08841108",
   631 => x"ffbfff06",
   632 => x"84120c84",
   633 => x"1108e1ff",
   634 => x"0684120c",
   635 => x"75882b9e",
   636 => x"80068412",
   637 => x"08710784",
   638 => x"130c8412",
   639 => x"0880c080",
   640 => x"0784130c",
   641 => x"55538151",
   642 => x"97c33f80",
   643 => x"d9940884",
   644 => x"1108ffbf",
   645 => x"ff068412",
   646 => x"0c53aa51",
   647 => x"97af3ffd",
   648 => x"e339ff90",
   649 => x"127081ff",
   650 => x"0680d994",
   651 => x"08841108",
   652 => x"feffff06",
   653 => x"84120c84",
   654 => x"1108e1ff",
   655 => x"0684120c",
   656 => x"71842b9e",
   657 => x"80068412",
   658 => x"08707207",
   659 => x"84140c54",
   660 => x"84120880",
   661 => x"c0800784",
   662 => x"130c5755",
   663 => x"56528151",
   664 => x"96eb3f80",
   665 => x"d9940884",
   666 => x"1108ffbf",
   667 => x"ff068412",
   668 => x"0c841108",
   669 => x"e1ff0684",
   670 => x"120c7588",
   671 => x"2b9e8006",
   672 => x"84120871",
   673 => x"0784130c",
   674 => x"84120880",
   675 => x"c0800784",
   676 => x"130c5553",
   677 => x"815196b5",
   678 => x"3f80d994",
   679 => x"08841108",
   680 => x"ffbfff06",
   681 => x"84120c53",
   682 => x"aa5196a1",
   683 => x"3ffcd539",
   684 => x"fb3d0d77",
   685 => x"70335356",
   686 => x"71802e81",
   687 => x"8f387155",
   688 => x"811680d9",
   689 => x"94088411",
   690 => x"08818080",
   691 => x"0784120c",
   692 => x"841108e1",
   693 => x"ff068412",
   694 => x"0c76842b",
   695 => x"9e800684",
   696 => x"12087072",
   697 => x"0784140c",
   698 => x"55841208",
   699 => x"80c08007",
   700 => x"84130c56",
   701 => x"54568151",
   702 => x"95d33f80",
   703 => x"d9940884",
   704 => x"1108ffbf",
   705 => x"ff068412",
   706 => x"0c841108",
   707 => x"e1ff0684",
   708 => x"120c7588",
   709 => x"2b9e8006",
   710 => x"84120871",
   711 => x"0784130c",
   712 => x"84120880",
   713 => x"c0800784",
   714 => x"130c5553",
   715 => x"8151959d",
   716 => x"3f80d994",
   717 => x"08841108",
   718 => x"ffbfff06",
   719 => x"84120c53",
   720 => x"ae519589",
   721 => x"3f753355",
   722 => x"74fef538",
   723 => x"873d0d04",
   724 => x"ff3d0d02",
   725 => x"8f053370",
   726 => x"52529684",
   727 => x"3f715196",
   728 => x"f33f7180",
   729 => x"0c833d0d",
   730 => x"04fa3d0d",
   731 => x"02a30533",
   732 => x"56758d2e",
   733 => x"80f43875",
   734 => x"88327030",
   735 => x"7780ff32",
   736 => x"70307280",
   737 => x"25718025",
   738 => x"07545156",
   739 => x"58557495",
   740 => x"389f7627",
   741 => x"8c3880f0",
   742 => x"c8335580",
   743 => x"ce7527ae",
   744 => x"38883d0d",
   745 => x"0480f0c8",
   746 => x"33567580",
   747 => x"2ef33888",
   748 => x"5192a13f",
   749 => x"a051929c",
   750 => x"3f885192",
   751 => x"973f80f0",
   752 => x"c833ff05",
   753 => x"577680f0",
   754 => x"c834883d",
   755 => x"0d047551",
   756 => x"92823f80",
   757 => x"f0c83381",
   758 => x"11555773",
   759 => x"80f0c834",
   760 => x"7580eff4",
   761 => x"1834883d",
   762 => x"0d048a51",
   763 => x"91e63f80",
   764 => x"f0c83381",
   765 => x"11565474",
   766 => x"80f0c834",
   767 => x"800b80ef",
   768 => x"f4153480",
   769 => x"56800b80",
   770 => x"eff41733",
   771 => x"565474a0",
   772 => x"2e833881",
   773 => x"5474802e",
   774 => x"90387380",
   775 => x"2e8b3881",
   776 => x"167081ff",
   777 => x"065757dd",
   778 => x"3975802e",
   779 => x"bf38800b",
   780 => x"80f0c433",
   781 => x"55557474",
   782 => x"27ab3873",
   783 => x"57741010",
   784 => x"10751005",
   785 => x"765480ef",
   786 => x"f45380e9",
   787 => x"940551a0",
   788 => x"9a3f8008",
   789 => x"802ea638",
   790 => x"81157081",
   791 => x"ff065654",
   792 => x"767526d9",
   793 => x"3880d2ec",
   794 => x"5191833f",
   795 => x"80d2e851",
   796 => x"90fc3f80",
   797 => x"0b80f0c8",
   798 => x"34883d0d",
   799 => x"04741010",
   800 => x"80efb405",
   801 => x"700880f0",
   802 => x"cc0c5680",
   803 => x"0b80f0c8",
   804 => x"34e739fc",
   805 => x"3d0d8a51",
   806 => x"90ba3f80",
   807 => x"0b80f0c8",
   808 => x"34800b80",
   809 => x"f0c43480",
   810 => x"0b80f0cc",
   811 => x"0c80d380",
   812 => x"5280e994",
   813 => x"519de83f",
   814 => x"80d38452",
   815 => x"80f0c433",
   816 => x"70101011",
   817 => x"70101010",
   818 => x"80eab405",
   819 => x"5356549d",
   820 => x"ce3f80f0",
   821 => x"c4337010",
   822 => x"1080efb4",
   823 => x"059fe071",
   824 => x"0c548111",
   825 => x"51557480",
   826 => x"f0c43480",
   827 => x"d3ac5274",
   828 => x"81ff0670",
   829 => x"8a2980e9",
   830 => x"94055253",
   831 => x"9da13f80",
   832 => x"d3b45280",
   833 => x"f0c43370",
   834 => x"10101170",
   835 => x"10101080",
   836 => x"eab40553",
   837 => x"55559d87",
   838 => x"3f80f0c4",
   839 => x"33701010",
   840 => x"80efb405",
   841 => x"9fc5710c",
   842 => x"54811151",
   843 => x"547380f0",
   844 => x"c43480d3",
   845 => x"d0527381",
   846 => x"ff06708a",
   847 => x"2980e994",
   848 => x"0552539c",
   849 => x"da3f80d3",
   850 => x"d45280f0",
   851 => x"c4337010",
   852 => x"10117010",
   853 => x"101080ea",
   854 => x"b4055356",
   855 => x"549cc03f",
   856 => x"80f0c433",
   857 => x"70101080",
   858 => x"efb405a6",
   859 => x"d8710c54",
   860 => x"81115155",
   861 => x"7480f0c4",
   862 => x"3480d3f4",
   863 => x"527481ff",
   864 => x"06708a29",
   865 => x"80e99405",
   866 => x"52539c93",
   867 => x"3f80d3fc",
   868 => x"5280f0c4",
   869 => x"33701010",
   870 => x"11701010",
   871 => x"1080eab4",
   872 => x"05535555",
   873 => x"9bf93f80",
   874 => x"f0c43370",
   875 => x"101080ef",
   876 => x"b405a78b",
   877 => x"710c5481",
   878 => x"11515473",
   879 => x"80f0c434",
   880 => x"80d49052",
   881 => x"7381ff06",
   882 => x"708a2980",
   883 => x"e9940552",
   884 => x"539bcc3f",
   885 => x"80d49852",
   886 => x"80f0c433",
   887 => x"70101011",
   888 => x"70101010",
   889 => x"80eab405",
   890 => x"5356549b",
   891 => x"b23f80f0",
   892 => x"c4337010",
   893 => x"1080efb4",
   894 => x"059eb571",
   895 => x"0c548111",
   896 => x"51557480",
   897 => x"f0c43480",
   898 => x"d4a85274",
   899 => x"81ff0670",
   900 => x"8a2980e9",
   901 => x"94055253",
   902 => x"9b853f80",
   903 => x"d4e05280",
   904 => x"f0c43370",
   905 => x"10101170",
   906 => x"10101080",
   907 => x"eab40553",
   908 => x"55559aeb",
   909 => x"3f80f0c4",
   910 => x"33701010",
   911 => x"80efb405",
   912 => x"9d9d710c",
   913 => x"54810553",
   914 => x"7280f0c4",
   915 => x"3480d2e8",
   916 => x"518d9b3f",
   917 => x"810b80f0",
   918 => x"d0348fcf",
   919 => x"3f8008ae",
   920 => x"3880f0cc",
   921 => x"0853728d",
   922 => x"3880f0d0",
   923 => x"335372ea",
   924 => x"38863d0d",
   925 => x"04722d80",
   926 => x"0b80f0cc",
   927 => x"0c80d2e8",
   928 => x"518ceb3f",
   929 => x"80f0d033",
   930 => x"5372cf38",
   931 => x"e4398fae",
   932 => x"3f800881",
   933 => x"ff0651f9",
   934 => x"d03fffbe",
   935 => x"39fc3d0d",
   936 => x"8a518cb0",
   937 => x"3f80d4b0",
   938 => x"518cc33f",
   939 => x"800b80f0",
   940 => x"c4335353",
   941 => x"72722780",
   942 => x"f3387210",
   943 => x"10107310",
   944 => x"0580e994",
   945 => x"05705254",
   946 => x"8ca43f72",
   947 => x"822b7311",
   948 => x"832b80ea",
   949 => x"b4113351",
   950 => x"53557180",
   951 => x"2eb63873",
   952 => x"519aa93f",
   953 => x"800881ff",
   954 => x"06527189",
   955 => x"269338a0",
   956 => x"518be13f",
   957 => x"81127081",
   958 => x"ff065354",
   959 => x"897227ef",
   960 => x"3880d4c8",
   961 => x"518be73f",
   962 => x"7215832b",
   963 => x"80eab405",
   964 => x"518bdb3f",
   965 => x"8a518bbc",
   966 => x"3f811370",
   967 => x"81ff0680",
   968 => x"f0c43354",
   969 => x"54557173",
   970 => x"26ff8f38",
   971 => x"8a518ba4",
   972 => x"3f863d0d",
   973 => x"04803d0d",
   974 => x"8c518b98",
   975 => x"3f823d0d",
   976 => x"04fe3d0d",
   977 => x"02930533",
   978 => x"80d4d852",
   979 => x"538b9f3f",
   980 => x"72518bbd",
   981 => x"3f80d4e4",
   982 => x"518b933f",
   983 => x"72882b80",
   984 => x"d98c0811",
   985 => x"70085353",
   986 => x"538ba63f",
   987 => x"80d4f051",
   988 => x"8afc3f80",
   989 => x"d98c0813",
   990 => x"84110852",
   991 => x"528b923f",
   992 => x"80d4fc51",
   993 => x"8ae83f80",
   994 => x"d98c0813",
   995 => x"88110852",
   996 => x"528afe3f",
   997 => x"80d58851",
   998 => x"8ad43f80",
   999 => x"d98c0813",
  1000 => x"8c110852",
  1001 => x"528aea3f",
  1002 => x"80d59451",
  1003 => x"8ac03f80",
  1004 => x"d98c0813",
  1005 => x"90110852",
  1006 => x"538ad63f",
  1007 => x"8a518a94",
  1008 => x"3f843d0d",
  1009 => x"04ff3d0d",
  1010 => x"80527151",
  1011 => x"fef33f81",
  1012 => x"127081ff",
  1013 => x"06515283",
  1014 => x"7227ef38",
  1015 => x"833d0d04",
  1016 => x"f03d0d80",
  1017 => x"0b80eff4",
  1018 => x"3380eff4",
  1019 => x"59555673",
  1020 => x"a02e0981",
  1021 => x"06963881",
  1022 => x"167081ff",
  1023 => x"0680eff4",
  1024 => x"11703353",
  1025 => x"59575473",
  1026 => x"a02eec38",
  1027 => x"80588077",
  1028 => x"33565474",
  1029 => x"742e8338",
  1030 => x"815474a0",
  1031 => x"2e83dd38",
  1032 => x"73848a38",
  1033 => x"74a02e83",
  1034 => x"d3388118",
  1035 => x"7081ff06",
  1036 => x"595a8178",
  1037 => x"26d8388a",
  1038 => x"53923dfc",
  1039 => x"05527651",
  1040 => x"9cee3f80",
  1041 => x"0881ff06",
  1042 => x"59800b80",
  1043 => x"eff43380",
  1044 => x"eff45955",
  1045 => x"5673a02e",
  1046 => x"09810696",
  1047 => x"38811670",
  1048 => x"81ff0680",
  1049 => x"eff41170",
  1050 => x"33575957",
  1051 => x"5873a02e",
  1052 => x"ec388058",
  1053 => x"80773356",
  1054 => x"5474742e",
  1055 => x"83388154",
  1056 => x"74a02e83",
  1057 => x"b8387383",
  1058 => x"e53874a0",
  1059 => x"2e83ae38",
  1060 => x"81187081",
  1061 => x"ff065955",
  1062 => x"827826d8",
  1063 => x"388a5392",
  1064 => x"3df80552",
  1065 => x"76519c88",
  1066 => x"3f80085c",
  1067 => x"800b80ef",
  1068 => x"f43380ef",
  1069 => x"f4595556",
  1070 => x"73a02e09",
  1071 => x"81069638",
  1072 => x"81167081",
  1073 => x"ff0680ef",
  1074 => x"f4117033",
  1075 => x"57525757",
  1076 => x"73a02eec",
  1077 => x"38805880",
  1078 => x"77335654",
  1079 => x"74742e83",
  1080 => x"38815474",
  1081 => x"a02e8396",
  1082 => x"387383c3",
  1083 => x"3874a02e",
  1084 => x"838c3881",
  1085 => x"187081ff",
  1086 => x"06595a83",
  1087 => x"7826d838",
  1088 => x"8a53923d",
  1089 => x"f4055276",
  1090 => x"519ba53f",
  1091 => x"80085b80",
  1092 => x"0b80eff4",
  1093 => x"3380eff4",
  1094 => x"59555673",
  1095 => x"a02e0981",
  1096 => x"06963881",
  1097 => x"167081ff",
  1098 => x"0680eff4",
  1099 => x"11703357",
  1100 => x"59575873",
  1101 => x"a02eec38",
  1102 => x"80588077",
  1103 => x"33565474",
  1104 => x"742e8338",
  1105 => x"815474a0",
  1106 => x"2e82f438",
  1107 => x"7383a138",
  1108 => x"74a02e82",
  1109 => x"ea388118",
  1110 => x"7081ff06",
  1111 => x"595a8478",
  1112 => x"26d8388a",
  1113 => x"53923df0",
  1114 => x"05527651",
  1115 => x"9ac23f80",
  1116 => x"085a800b",
  1117 => x"80eff433",
  1118 => x"80eff459",
  1119 => x"555673a0",
  1120 => x"2e098106",
  1121 => x"96388116",
  1122 => x"7081ff06",
  1123 => x"80eff411",
  1124 => x"70335759",
  1125 => x"575873a0",
  1126 => x"2eec3880",
  1127 => x"58807733",
  1128 => x"56547474",
  1129 => x"2e833881",
  1130 => x"5474a02e",
  1131 => x"82d23873",
  1132 => x"82ff3874",
  1133 => x"a02e82c8",
  1134 => x"38811870",
  1135 => x"81ff0659",
  1136 => x"54857826",
  1137 => x"d8388a53",
  1138 => x"923dec05",
  1139 => x"52765199",
  1140 => x"df3f7883",
  1141 => x"2682ea38",
  1142 => x"78828029",
  1143 => x"80d98c08",
  1144 => x"057c8412",
  1145 => x"0c7b8812",
  1146 => x"0c7a8c12",
  1147 => x"0c800890",
  1148 => x"120c5878",
  1149 => x"51faca3f",
  1150 => x"923d0d04",
  1151 => x"81167081",
  1152 => x"ff0680ef",
  1153 => x"f4117033",
  1154 => x"5c525757",
  1155 => x"78a02e09",
  1156 => x"8106fc96",
  1157 => x"38811670",
  1158 => x"81ff0680",
  1159 => x"eff41170",
  1160 => x"335c5257",
  1161 => x"5778a02e",
  1162 => x"d338fbfe",
  1163 => x"39811670",
  1164 => x"81ff0680",
  1165 => x"eff41159",
  1166 => x"5755fbd2",
  1167 => x"39811670",
  1168 => x"81ff0680",
  1169 => x"eff41170",
  1170 => x"335f5957",
  1171 => x"547ba02e",
  1172 => x"098106fc",
  1173 => x"bb388116",
  1174 => x"7081ff06",
  1175 => x"80eff411",
  1176 => x"70335f59",
  1177 => x"57547ba0",
  1178 => x"2ed338fc",
  1179 => x"a3398116",
  1180 => x"7081ff06",
  1181 => x"80eff411",
  1182 => x"59575bfb",
  1183 => x"f7398116",
  1184 => x"7081ff06",
  1185 => x"80eff411",
  1186 => x"70335759",
  1187 => x"575573a0",
  1188 => x"2e098106",
  1189 => x"fcdd3881",
  1190 => x"167081ff",
  1191 => x"0680eff4",
  1192 => x"11703357",
  1193 => x"59575573",
  1194 => x"a02ed338",
  1195 => x"fcc53981",
  1196 => x"167081ff",
  1197 => x"0680eff4",
  1198 => x"1159575b",
  1199 => x"fc993981",
  1200 => x"167081ff",
  1201 => x"0680eff4",
  1202 => x"11703357",
  1203 => x"59575573",
  1204 => x"a02e0981",
  1205 => x"06fcff38",
  1206 => x"81167081",
  1207 => x"ff0680ef",
  1208 => x"f4117033",
  1209 => x"57595755",
  1210 => x"73a02ed3",
  1211 => x"38fce739",
  1212 => x"81167081",
  1213 => x"ff0680ef",
  1214 => x"f4115257",
  1215 => x"57fcbb39",
  1216 => x"81167081",
  1217 => x"ff0680ef",
  1218 => x"f4117033",
  1219 => x"57595755",
  1220 => x"73a02e09",
  1221 => x"8106fda1",
  1222 => x"38811670",
  1223 => x"81ff0680",
  1224 => x"eff41170",
  1225 => x"33575957",
  1226 => x"5573a02e",
  1227 => x"d338fd89",
  1228 => x"39811670",
  1229 => x"81ff0680",
  1230 => x"eff41152",
  1231 => x"5757fcdd",
  1232 => x"3980d5a0",
  1233 => x"5183a73f",
  1234 => x"785183c5",
  1235 => x"3f80d5c0",
  1236 => x"51839b3f",
  1237 => x"923d0d04",
  1238 => x"fe3d0d80",
  1239 => x"0b80d98c",
  1240 => x"08545271",
  1241 => x"82802913",
  1242 => x"5181710c",
  1243 => x"81127081",
  1244 => x"ff065351",
  1245 => x"837227eb",
  1246 => x"3880d994",
  1247 => x"08841108",
  1248 => x"810a0784",
  1249 => x"120c5284",
  1250 => x"3d0d04ff",
  1251 => x"3d0d80d9",
  1252 => x"94088411",
  1253 => x"0870fe0a",
  1254 => x"0684130c",
  1255 => x"5252833d",
  1256 => x"0d04fd3d",
  1257 => x"0d80d994",
  1258 => x"08700881",
  1259 => x"0a0680e9",
  1260 => x"900c5484",
  1261 => x"e03f80e9",
  1262 => x"9008a9be",
  1263 => x"55537284",
  1264 => x"3896d054",
  1265 => x"7380f0d4",
  1266 => x"0c72802e",
  1267 => x"81ea3885",
  1268 => x"df3f80d5",
  1269 => x"e8518296",
  1270 => x"3f8c5181",
  1271 => x"f73f80d5",
  1272 => x"ec51828a",
  1273 => x"3f80e990",
  1274 => x"08802e81",
  1275 => x"a23880d6",
  1276 => x"885181fa",
  1277 => x"3f80e990",
  1278 => x"08802e81",
  1279 => x"a03880d9",
  1280 => x"8c085482",
  1281 => x"0b84150c",
  1282 => x"800b8815",
  1283 => x"0c800b8c",
  1284 => x"150c840b",
  1285 => x"90150c80",
  1286 => x"0b828415",
  1287 => x"0c810b82",
  1288 => x"88150c81",
  1289 => x"0b828c15",
  1290 => x"0c800b82",
  1291 => x"90150c81",
  1292 => x"0b828015",
  1293 => x"0c810b84",
  1294 => x"84150c82",
  1295 => x"0b848815",
  1296 => x"0c820b84",
  1297 => x"8c150c80",
  1298 => x"0b849015",
  1299 => x"0c810b84",
  1300 => x"80150c82",
  1301 => x"0b868415",
  1302 => x"0c820b86",
  1303 => x"88150c82",
  1304 => x"0b868c15",
  1305 => x"0c830b86",
  1306 => x"90150c81",
  1307 => x"0b868015",
  1308 => x"0c80d994",
  1309 => x"08841108",
  1310 => x"70810a07",
  1311 => x"84130c54",
  1312 => x"84110870",
  1313 => x"fe0a0684",
  1314 => x"130c5454",
  1315 => x"8a8f3f80",
  1316 => x"d6945180",
  1317 => x"d93f80e9",
  1318 => x"9008fee2",
  1319 => x"3880d6b8",
  1320 => x"51ec8d3f",
  1321 => x"82528351",
  1322 => x"e79d3f80",
  1323 => x"d6cc51eb",
  1324 => x"ff3fefdf",
  1325 => x"3f89e63f",
  1326 => x"e1b93ffe",
  1327 => x"9239ff3d",
  1328 => x"0d028f05",
  1329 => x"3380d9a0",
  1330 => x"0852710c",
  1331 => x"800b800c",
  1332 => x"833d0d04",
  1333 => x"ff3d0d02",
  1334 => x"8f053351",
  1335 => x"80f0d408",
  1336 => x"52712d80",
  1337 => x"0881ff06",
  1338 => x"800c833d",
  1339 => x"0d04fe3d",
  1340 => x"0d747033",
  1341 => x"53537180",
  1342 => x"2e933881",
  1343 => x"13725280",
  1344 => x"f0d40853",
  1345 => x"53712d72",
  1346 => x"335271ef",
  1347 => x"38843d0d",
  1348 => x"04f23d0d",
  1349 => x"608c3d70",
  1350 => x"5b5b5380",
  1351 => x"73565776",
  1352 => x"732480f8",
  1353 => x"38781754",
  1354 => x"8a527451",
  1355 => x"84ce3f80",
  1356 => x"08b00553",
  1357 => x"72743481",
  1358 => x"17578a52",
  1359 => x"74518497",
  1360 => x"3f800855",
  1361 => x"8008de38",
  1362 => x"8008779f",
  1363 => x"2a187081",
  1364 => x"2c5a5656",
  1365 => x"8078259e",
  1366 => x"387817ff",
  1367 => x"05557519",
  1368 => x"70335553",
  1369 => x"74337334",
  1370 => x"73753481",
  1371 => x"16ff1656",
  1372 => x"56777624",
  1373 => x"e9387619",
  1374 => x"56807634",
  1375 => x"79703354",
  1376 => x"5472802e",
  1377 => x"93388114",
  1378 => x"735280f0",
  1379 => x"d4085854",
  1380 => x"762d7333",
  1381 => x"5372ef38",
  1382 => x"903d0d04",
  1383 => x"ad7a3402",
  1384 => x"a9057330",
  1385 => x"71195656",
  1386 => x"598a5274",
  1387 => x"5183cd3f",
  1388 => x"8008b005",
  1389 => x"53727434",
  1390 => x"8117578a",
  1391 => x"52745183",
  1392 => x"963f8008",
  1393 => x"558008fe",
  1394 => x"dc38fefc",
  1395 => x"39ff3d0d",
  1396 => x"80d99808",
  1397 => x"74101075",
  1398 => x"10059412",
  1399 => x"0c52850b",
  1400 => x"98130c98",
  1401 => x"12087081",
  1402 => x"06515170",
  1403 => x"f638833d",
  1404 => x"0d04fd3d",
  1405 => x"0d80d998",
  1406 => x"0876b0ea",
  1407 => x"2994120c",
  1408 => x"54850b98",
  1409 => x"150c9814",
  1410 => x"08708106",
  1411 => x"515372f6",
  1412 => x"38853d0d",
  1413 => x"04803d0d",
  1414 => x"80d99c08",
  1415 => x"51b60b8c",
  1416 => x"120c830b",
  1417 => x"88120c82",
  1418 => x"3d0d0480",
  1419 => x"3d0d80d9",
  1420 => x"9c088411",
  1421 => x"08810680",
  1422 => x"0c51823d",
  1423 => x"0d04ff3d",
  1424 => x"0d80d99c",
  1425 => x"08528412",
  1426 => x"08708106",
  1427 => x"51517080",
  1428 => x"2ef43871",
  1429 => x"087081ff",
  1430 => x"06800c51",
  1431 => x"833d0d04",
  1432 => x"fe3d0d02",
  1433 => x"93053353",
  1434 => x"728a2e9c",
  1435 => x"3880d99c",
  1436 => x"08528412",
  1437 => x"0870892a",
  1438 => x"70810651",
  1439 => x"515170f2",
  1440 => x"3872720c",
  1441 => x"843d0d04",
  1442 => x"80d99c08",
  1443 => x"52841208",
  1444 => x"70892a70",
  1445 => x"81065151",
  1446 => x"5170f238",
  1447 => x"8d720c84",
  1448 => x"12087089",
  1449 => x"2a708106",
  1450 => x"51515170",
  1451 => x"c538d239",
  1452 => x"803d0d80",
  1453 => x"d9900851",
  1454 => x"800b8412",
  1455 => x"0c83fe80",
  1456 => x"0b88120c",
  1457 => x"800b80f0",
  1458 => x"d834800b",
  1459 => x"80f0dc34",
  1460 => x"823d0d04",
  1461 => x"fa3d0d02",
  1462 => x"a3053380",
  1463 => x"d9900880",
  1464 => x"f0d83370",
  1465 => x"81ff0670",
  1466 => x"10101180",
  1467 => x"f0dc3370",
  1468 => x"81ff0672",
  1469 => x"90291170",
  1470 => x"882b7807",
  1471 => x"770c535b",
  1472 => x"5b555559",
  1473 => x"5454738a",
  1474 => x"2e983874",
  1475 => x"80cf2e92",
  1476 => x"38738c2e",
  1477 => x"a4388116",
  1478 => x"537280f0",
  1479 => x"dc34883d",
  1480 => x"0d0471a3",
  1481 => x"26a33881",
  1482 => x"17527180",
  1483 => x"f0d83480",
  1484 => x"0b80f0dc",
  1485 => x"34883d0d",
  1486 => x"04805271",
  1487 => x"882b730c",
  1488 => x"81125297",
  1489 => x"907226f3",
  1490 => x"38800b80",
  1491 => x"f0d83480",
  1492 => x"0b80f0dc",
  1493 => x"34df398c",
  1494 => x"08028c0c",
  1495 => x"fd3d0d80",
  1496 => x"538c088c",
  1497 => x"0508528c",
  1498 => x"08880508",
  1499 => x"5182de3f",
  1500 => x"80087080",
  1501 => x"0c54853d",
  1502 => x"0d8c0c04",
  1503 => x"8c08028c",
  1504 => x"0cfd3d0d",
  1505 => x"81538c08",
  1506 => x"8c050852",
  1507 => x"8c088805",
  1508 => x"085182b9",
  1509 => x"3f800870",
  1510 => x"800c5485",
  1511 => x"3d0d8c0c",
  1512 => x"048c0802",
  1513 => x"8c0cf93d",
  1514 => x"0d800b8c",
  1515 => x"08fc050c",
  1516 => x"8c088805",
  1517 => x"088025ab",
  1518 => x"388c0888",
  1519 => x"0508308c",
  1520 => x"0888050c",
  1521 => x"800b8c08",
  1522 => x"f4050c8c",
  1523 => x"08fc0508",
  1524 => x"8838810b",
  1525 => x"8c08f405",
  1526 => x"0c8c08f4",
  1527 => x"05088c08",
  1528 => x"fc050c8c",
  1529 => x"088c0508",
  1530 => x"8025ab38",
  1531 => x"8c088c05",
  1532 => x"08308c08",
  1533 => x"8c050c80",
  1534 => x"0b8c08f0",
  1535 => x"050c8c08",
  1536 => x"fc050888",
  1537 => x"38810b8c",
  1538 => x"08f0050c",
  1539 => x"8c08f005",
  1540 => x"088c08fc",
  1541 => x"050c8053",
  1542 => x"8c088c05",
  1543 => x"08528c08",
  1544 => x"88050851",
  1545 => x"81a73f80",
  1546 => x"08708c08",
  1547 => x"f8050c54",
  1548 => x"8c08fc05",
  1549 => x"08802e8c",
  1550 => x"388c08f8",
  1551 => x"0508308c",
  1552 => x"08f8050c",
  1553 => x"8c08f805",
  1554 => x"0870800c",
  1555 => x"54893d0d",
  1556 => x"8c0c048c",
  1557 => x"08028c0c",
  1558 => x"fb3d0d80",
  1559 => x"0b8c08fc",
  1560 => x"050c8c08",
  1561 => x"88050880",
  1562 => x"2593388c",
  1563 => x"08880508",
  1564 => x"308c0888",
  1565 => x"050c810b",
  1566 => x"8c08fc05",
  1567 => x"0c8c088c",
  1568 => x"05088025",
  1569 => x"8c388c08",
  1570 => x"8c050830",
  1571 => x"8c088c05",
  1572 => x"0c81538c",
  1573 => x"088c0508",
  1574 => x"528c0888",
  1575 => x"050851ad",
  1576 => x"3f800870",
  1577 => x"8c08f805",
  1578 => x"0c548c08",
  1579 => x"fc050880",
  1580 => x"2e8c388c",
  1581 => x"08f80508",
  1582 => x"308c08f8",
  1583 => x"050c8c08",
  1584 => x"f8050870",
  1585 => x"800c5487",
  1586 => x"3d0d8c0c",
  1587 => x"048c0802",
  1588 => x"8c0cfd3d",
  1589 => x"0d810b8c",
  1590 => x"08fc050c",
  1591 => x"800b8c08",
  1592 => x"f8050c8c",
  1593 => x"088c0508",
  1594 => x"8c088805",
  1595 => x"0827ac38",
  1596 => x"8c08fc05",
  1597 => x"08802ea3",
  1598 => x"38800b8c",
  1599 => x"088c0508",
  1600 => x"2499388c",
  1601 => x"088c0508",
  1602 => x"108c088c",
  1603 => x"050c8c08",
  1604 => x"fc050810",
  1605 => x"8c08fc05",
  1606 => x"0cc9398c",
  1607 => x"08fc0508",
  1608 => x"802e80c9",
  1609 => x"388c088c",
  1610 => x"05088c08",
  1611 => x"88050826",
  1612 => x"a1388c08",
  1613 => x"8805088c",
  1614 => x"088c0508",
  1615 => x"318c0888",
  1616 => x"050c8c08",
  1617 => x"f805088c",
  1618 => x"08fc0508",
  1619 => x"078c08f8",
  1620 => x"050c8c08",
  1621 => x"fc050881",
  1622 => x"2a8c08fc",
  1623 => x"050c8c08",
  1624 => x"8c050881",
  1625 => x"2a8c088c",
  1626 => x"050cffaf",
  1627 => x"398c0890",
  1628 => x"0508802e",
  1629 => x"8f388c08",
  1630 => x"88050870",
  1631 => x"8c08f405",
  1632 => x"0c518d39",
  1633 => x"8c08f805",
  1634 => x"08708c08",
  1635 => x"f4050c51",
  1636 => x"8c08f405",
  1637 => x"08800c85",
  1638 => x"3d0d8c0c",
  1639 => x"04803d0d",
  1640 => x"865182fd",
  1641 => x"3f81519d",
  1642 => x"e43ffd3d",
  1643 => x"0d755384",
  1644 => x"d8130880",
  1645 => x"2e8a3880",
  1646 => x"5372800c",
  1647 => x"853d0d04",
  1648 => x"81805272",
  1649 => x"5189fe3f",
  1650 => x"800884d8",
  1651 => x"140cff53",
  1652 => x"8008802e",
  1653 => x"e4388008",
  1654 => x"549f5380",
  1655 => x"74708405",
  1656 => x"560cff13",
  1657 => x"53807324",
  1658 => x"ce388074",
  1659 => x"70840556",
  1660 => x"0cff1353",
  1661 => x"728025e3",
  1662 => x"38ffbc39",
  1663 => x"fd3d0d75",
  1664 => x"7755539f",
  1665 => x"74278d38",
  1666 => x"96730cff",
  1667 => x"5271800c",
  1668 => x"853d0d04",
  1669 => x"84d81308",
  1670 => x"5271802e",
  1671 => x"93387310",
  1672 => x"10127008",
  1673 => x"79720c51",
  1674 => x"5271800c",
  1675 => x"853d0d04",
  1676 => x"7251fef6",
  1677 => x"3fff5280",
  1678 => x"08d33884",
  1679 => x"d8130874",
  1680 => x"10101170",
  1681 => x"087a720c",
  1682 => x"515152dd",
  1683 => x"39f93d0d",
  1684 => x"797b5856",
  1685 => x"769f2680",
  1686 => x"e83884d8",
  1687 => x"16085473",
  1688 => x"802eaa38",
  1689 => x"76101014",
  1690 => x"70085555",
  1691 => x"73802eba",
  1692 => x"38805873",
  1693 => x"812e8f38",
  1694 => x"73ff2ea3",
  1695 => x"3880750c",
  1696 => x"7651732d",
  1697 => x"80587780",
  1698 => x"0c893d0d",
  1699 => x"047551fe",
  1700 => x"993fff58",
  1701 => x"8008ef38",
  1702 => x"84d81608",
  1703 => x"54c63996",
  1704 => x"760c810b",
  1705 => x"800c893d",
  1706 => x"0d047551",
  1707 => x"81ed3f76",
  1708 => x"53800852",
  1709 => x"755181ad",
  1710 => x"3f800880",
  1711 => x"0c893d0d",
  1712 => x"0496760c",
  1713 => x"ff0b800c",
  1714 => x"893d0d04",
  1715 => x"fc3d0d76",
  1716 => x"785653ff",
  1717 => x"54749f26",
  1718 => x"b13884d8",
  1719 => x"13085271",
  1720 => x"802eae38",
  1721 => x"74101012",
  1722 => x"70085353",
  1723 => x"81547180",
  1724 => x"2e983882",
  1725 => x"5471ff2e",
  1726 => x"91388354",
  1727 => x"71812e8a",
  1728 => x"3880730c",
  1729 => x"7451712d",
  1730 => x"80547380",
  1731 => x"0c863d0d",
  1732 => x"047251fd",
  1733 => x"953f8008",
  1734 => x"f13884d8",
  1735 => x"130852c4",
  1736 => x"39ff3d0d",
  1737 => x"735280d9",
  1738 => x"a40851fe",
  1739 => x"a03f833d",
  1740 => x"0d04fe3d",
  1741 => x"0d755374",
  1742 => x"5280d9a4",
  1743 => x"0851fdbc",
  1744 => x"3f843d0d",
  1745 => x"04803d0d",
  1746 => x"80d9a408",
  1747 => x"51fcdb3f",
  1748 => x"823d0d04",
  1749 => x"ff3d0d73",
  1750 => x"5280d9a4",
  1751 => x"0851feec",
  1752 => x"3f833d0d",
  1753 => x"04fc3d0d",
  1754 => x"800b80f0",
  1755 => x"e80c7852",
  1756 => x"7751998d",
  1757 => x"3f800854",
  1758 => x"8008ff2e",
  1759 => x"88387380",
  1760 => x"0c863d0d",
  1761 => x"0480f0e8",
  1762 => x"08557480",
  1763 => x"2ef03876",
  1764 => x"75710c53",
  1765 => x"73800c86",
  1766 => x"3d0d0498",
  1767 => x"df3f04fc",
  1768 => x"3d0d7670",
  1769 => x"79707307",
  1770 => x"83065454",
  1771 => x"54557080",
  1772 => x"c3387170",
  1773 => x"08700970",
  1774 => x"f7fbfdff",
  1775 => x"130670f8",
  1776 => x"84828180",
  1777 => x"06515153",
  1778 => x"535470a6",
  1779 => x"38841472",
  1780 => x"74708405",
  1781 => x"560c7008",
  1782 => x"700970f7",
  1783 => x"fbfdff13",
  1784 => x"0670f884",
  1785 => x"82818006",
  1786 => x"51515353",
  1787 => x"5470802e",
  1788 => x"dc387352",
  1789 => x"71708105",
  1790 => x"53335170",
  1791 => x"73708105",
  1792 => x"553470f0",
  1793 => x"3874800c",
  1794 => x"863d0d04",
  1795 => x"fd3d0d75",
  1796 => x"70718306",
  1797 => x"53555270",
  1798 => x"b8387170",
  1799 => x"087009f7",
  1800 => x"fbfdff12",
  1801 => x"0670f884",
  1802 => x"82818006",
  1803 => x"51515253",
  1804 => x"709d3884",
  1805 => x"13700870",
  1806 => x"09f7fbfd",
  1807 => x"ff120670",
  1808 => x"f8848281",
  1809 => x"80065151",
  1810 => x"52537080",
  1811 => x"2ee53872",
  1812 => x"52713351",
  1813 => x"70802e8a",
  1814 => x"38811270",
  1815 => x"33525270",
  1816 => x"f8387174",
  1817 => x"31800c85",
  1818 => x"3d0d04fa",
  1819 => x"3d0d787a",
  1820 => x"7c705455",
  1821 => x"55527280",
  1822 => x"2e80d938",
  1823 => x"71740783",
  1824 => x"06517080",
  1825 => x"2e80d438",
  1826 => x"ff135372",
  1827 => x"ff2eb138",
  1828 => x"71337433",
  1829 => x"56517471",
  1830 => x"2e098106",
  1831 => x"a9387280",
  1832 => x"2e818738",
  1833 => x"7081ff06",
  1834 => x"5170802e",
  1835 => x"80fc3881",
  1836 => x"128115ff",
  1837 => x"15555552",
  1838 => x"72ff2e09",
  1839 => x"8106d138",
  1840 => x"71337433",
  1841 => x"56517081",
  1842 => x"ff067581",
  1843 => x"ff067171",
  1844 => x"31515252",
  1845 => x"70800c88",
  1846 => x"3d0d0471",
  1847 => x"74575583",
  1848 => x"73278838",
  1849 => x"71087408",
  1850 => x"2e883874",
  1851 => x"765552ff",
  1852 => x"9739fc13",
  1853 => x"5372802e",
  1854 => x"b1387408",
  1855 => x"7009f7fb",
  1856 => x"fdff1206",
  1857 => x"70f88482",
  1858 => x"81800651",
  1859 => x"5151709a",
  1860 => x"38841584",
  1861 => x"17575583",
  1862 => x"7327d038",
  1863 => x"74087608",
  1864 => x"2ed03874",
  1865 => x"765552fe",
  1866 => x"df39800b",
  1867 => x"800c883d",
  1868 => x"0d04f33d",
  1869 => x"0d606264",
  1870 => x"725a5a5e",
  1871 => x"5e805c76",
  1872 => x"70810558",
  1873 => x"3380d6d9",
  1874 => x"11337083",
  1875 => x"2a708106",
  1876 => x"51555556",
  1877 => x"72e93875",
  1878 => x"ad2e8288",
  1879 => x"3875ab2e",
  1880 => x"82843877",
  1881 => x"30707907",
  1882 => x"80257990",
  1883 => x"32703070",
  1884 => x"72078025",
  1885 => x"73075357",
  1886 => x"57515372",
  1887 => x"802e8738",
  1888 => x"75b02e81",
  1889 => x"eb38778a",
  1890 => x"38885875",
  1891 => x"b02e8338",
  1892 => x"8a58810a",
  1893 => x"5a7b8438",
  1894 => x"fe0a5a77",
  1895 => x"527951f3",
  1896 => x"db3f8008",
  1897 => x"78537a52",
  1898 => x"5bf3ac3f",
  1899 => x"80085a80",
  1900 => x"7080d6d9",
  1901 => x"18337082",
  1902 => x"2a708106",
  1903 => x"5156565a",
  1904 => x"5572802e",
  1905 => x"80c138d0",
  1906 => x"16567578",
  1907 => x"2580d738",
  1908 => x"80792475",
  1909 => x"7b260753",
  1910 => x"72933874",
  1911 => x"7a2e80eb",
  1912 => x"387a7625",
  1913 => x"80ed3872",
  1914 => x"802e80e7",
  1915 => x"38ff7770",
  1916 => x"81055933",
  1917 => x"575980d6",
  1918 => x"d9163370",
  1919 => x"822a7081",
  1920 => x"06515454",
  1921 => x"72c13873",
  1922 => x"83065372",
  1923 => x"802e9738",
  1924 => x"738106c9",
  1925 => x"17555372",
  1926 => x"8538ffa9",
  1927 => x"16547356",
  1928 => x"777624ff",
  1929 => x"ab388079",
  1930 => x"2480f038",
  1931 => x"7b802e84",
  1932 => x"38743055",
  1933 => x"7c802e8c",
  1934 => x"38ff1753",
  1935 => x"7883387d",
  1936 => x"53727d0c",
  1937 => x"74800c8f",
  1938 => x"3d0d0481",
  1939 => x"53757b24",
  1940 => x"ff953881",
  1941 => x"75792917",
  1942 => x"78708105",
  1943 => x"5a335856",
  1944 => x"59ff9339",
  1945 => x"815c7670",
  1946 => x"81055833",
  1947 => x"56fdf439",
  1948 => x"80773354",
  1949 => x"547280f8",
  1950 => x"2eb23872",
  1951 => x"80d83270",
  1952 => x"30708025",
  1953 => x"76075151",
  1954 => x"5372802e",
  1955 => x"fdf83881",
  1956 => x"17338218",
  1957 => x"58569058",
  1958 => x"fdf83981",
  1959 => x"0a557b84",
  1960 => x"38fe0a55",
  1961 => x"7f53a273",
  1962 => x"0cff8939",
  1963 => x"8154cc39",
  1964 => x"fd3d0d77",
  1965 => x"54765375",
  1966 => x"5280d9a4",
  1967 => x"0851fcf2",
  1968 => x"3f853d0d",
  1969 => x"04f33d0d",
  1970 => x"7f618b11",
  1971 => x"70f8065c",
  1972 => x"55555e72",
  1973 => x"96268338",
  1974 => x"90598079",
  1975 => x"24747a26",
  1976 => x"07538054",
  1977 => x"72742e09",
  1978 => x"810680cb",
  1979 => x"387d518b",
  1980 => x"ca3f7883",
  1981 => x"f72680c6",
  1982 => x"3878832a",
  1983 => x"70101010",
  1984 => x"80e0e005",
  1985 => x"8c110859",
  1986 => x"595a7678",
  1987 => x"2e83b038",
  1988 => x"841708fc",
  1989 => x"06568c17",
  1990 => x"08881808",
  1991 => x"718c120c",
  1992 => x"88120c58",
  1993 => x"75178411",
  1994 => x"08810784",
  1995 => x"120c537d",
  1996 => x"518b893f",
  1997 => x"88175473",
  1998 => x"800c8f3d",
  1999 => x"0d047889",
  2000 => x"2a79832a",
  2001 => x"5b537280",
  2002 => x"2ebf3878",
  2003 => x"862ab805",
  2004 => x"5a847327",
  2005 => x"b43880db",
  2006 => x"135a9473",
  2007 => x"27ab3878",
  2008 => x"8c2a80ee",
  2009 => x"055a80d4",
  2010 => x"73279e38",
  2011 => x"788f2a80",
  2012 => x"f7055a82",
  2013 => x"d4732791",
  2014 => x"3878922a",
  2015 => x"80fc055a",
  2016 => x"8ad47327",
  2017 => x"843880fe",
  2018 => x"5a791010",
  2019 => x"1080e0e0",
  2020 => x"058c1108",
  2021 => x"58557675",
  2022 => x"2ea33884",
  2023 => x"1708fc06",
  2024 => x"707a3155",
  2025 => x"56738f24",
  2026 => x"88d53873",
  2027 => x"8025fee6",
  2028 => x"388c1708",
  2029 => x"5776752e",
  2030 => x"098106df",
  2031 => x"38811a5a",
  2032 => x"80e0f008",
  2033 => x"577680e0",
  2034 => x"e82e82c0",
  2035 => x"38841708",
  2036 => x"fc06707a",
  2037 => x"31555673",
  2038 => x"8f2481f9",
  2039 => x"3880e0e8",
  2040 => x"0b80e0f4",
  2041 => x"0c80e0e8",
  2042 => x"0b80e0f0",
  2043 => x"0c738025",
  2044 => x"feb23883",
  2045 => x"ff762783",
  2046 => x"df387589",
  2047 => x"2a76832a",
  2048 => x"55537280",
  2049 => x"2ebf3875",
  2050 => x"862ab805",
  2051 => x"54847327",
  2052 => x"b43880db",
  2053 => x"13549473",
  2054 => x"27ab3875",
  2055 => x"8c2a80ee",
  2056 => x"055480d4",
  2057 => x"73279e38",
  2058 => x"758f2a80",
  2059 => x"f7055482",
  2060 => x"d4732791",
  2061 => x"3875922a",
  2062 => x"80fc0554",
  2063 => x"8ad47327",
  2064 => x"843880fe",
  2065 => x"54731010",
  2066 => x"1080e0e0",
  2067 => x"05881108",
  2068 => x"56587478",
  2069 => x"2e86cf38",
  2070 => x"841508fc",
  2071 => x"06537573",
  2072 => x"278d3888",
  2073 => x"15085574",
  2074 => x"782e0981",
  2075 => x"06ea388c",
  2076 => x"150880e0",
  2077 => x"e00b8405",
  2078 => x"08718c1a",
  2079 => x"0c76881a",
  2080 => x"0c788813",
  2081 => x"0c788c18",
  2082 => x"0c5d5879",
  2083 => x"53807a24",
  2084 => x"83e63872",
  2085 => x"822c8171",
  2086 => x"2b5c537a",
  2087 => x"7c268198",
  2088 => x"387b7b06",
  2089 => x"537282f1",
  2090 => x"3879fc06",
  2091 => x"84055a7a",
  2092 => x"10707d06",
  2093 => x"545b7282",
  2094 => x"e038841a",
  2095 => x"5af13988",
  2096 => x"178c1108",
  2097 => x"58587678",
  2098 => x"2e098106",
  2099 => x"fcc23882",
  2100 => x"1a5afdec",
  2101 => x"39781779",
  2102 => x"81078419",
  2103 => x"0c7080e0",
  2104 => x"f40c7080",
  2105 => x"e0f00c80",
  2106 => x"e0e80b8c",
  2107 => x"120c8c11",
  2108 => x"0888120c",
  2109 => x"74810784",
  2110 => x"120c7411",
  2111 => x"75710c51",
  2112 => x"537d5187",
  2113 => x"b73f8817",
  2114 => x"54fcac39",
  2115 => x"80e0e00b",
  2116 => x"8405087a",
  2117 => x"545c7980",
  2118 => x"25fef838",
  2119 => x"82da397a",
  2120 => x"097c0670",
  2121 => x"80e0e00b",
  2122 => x"84050c5c",
  2123 => x"7a105b7a",
  2124 => x"7c268538",
  2125 => x"7a85b838",
  2126 => x"80e0e00b",
  2127 => x"88050870",
  2128 => x"841208fc",
  2129 => x"06707c31",
  2130 => x"7c72268f",
  2131 => x"72250757",
  2132 => x"575c5d55",
  2133 => x"72802e80",
  2134 => x"db38797a",
  2135 => x"1680e0d8",
  2136 => x"081b9011",
  2137 => x"5a55575b",
  2138 => x"80e0d408",
  2139 => x"ff2e8838",
  2140 => x"a08f13e0",
  2141 => x"80065776",
  2142 => x"527d5186",
  2143 => x"c03f8008",
  2144 => x"548008ff",
  2145 => x"2e903880",
  2146 => x"08762782",
  2147 => x"99387480",
  2148 => x"e0e02e82",
  2149 => x"913880e0",
  2150 => x"e00b8805",
  2151 => x"08558415",
  2152 => x"08fc0670",
  2153 => x"7a317a72",
  2154 => x"268f7225",
  2155 => x"07525553",
  2156 => x"7283e638",
  2157 => x"74798107",
  2158 => x"84170c79",
  2159 => x"167080e0",
  2160 => x"e00b8805",
  2161 => x"0c758107",
  2162 => x"84120c54",
  2163 => x"7e525785",
  2164 => x"eb3f8817",
  2165 => x"54fae039",
  2166 => x"75832a70",
  2167 => x"54548074",
  2168 => x"24819b38",
  2169 => x"72822c81",
  2170 => x"712b80e0",
  2171 => x"e4080770",
  2172 => x"80e0e00b",
  2173 => x"84050c75",
  2174 => x"10101080",
  2175 => x"e0e00588",
  2176 => x"1108585a",
  2177 => x"5d53778c",
  2178 => x"180c7488",
  2179 => x"180c7688",
  2180 => x"190c768c",
  2181 => x"160cfcf3",
  2182 => x"39797a10",
  2183 => x"101080e0",
  2184 => x"e0057057",
  2185 => x"595d8c15",
  2186 => x"08577675",
  2187 => x"2ea33884",
  2188 => x"1708fc06",
  2189 => x"707a3155",
  2190 => x"56738f24",
  2191 => x"83ca3873",
  2192 => x"80258481",
  2193 => x"388c1708",
  2194 => x"5776752e",
  2195 => x"098106df",
  2196 => x"38881581",
  2197 => x"1b708306",
  2198 => x"555b5572",
  2199 => x"c9387c83",
  2200 => x"06537280",
  2201 => x"2efdb838",
  2202 => x"ff1df819",
  2203 => x"595d8818",
  2204 => x"08782eea",
  2205 => x"38fdb539",
  2206 => x"831a53fc",
  2207 => x"96398314",
  2208 => x"70822c81",
  2209 => x"712b80e0",
  2210 => x"e4080770",
  2211 => x"80e0e00b",
  2212 => x"84050c76",
  2213 => x"10101080",
  2214 => x"e0e00588",
  2215 => x"1108595b",
  2216 => x"5e5153fe",
  2217 => x"e13980e0",
  2218 => x"a4081758",
  2219 => x"8008762e",
  2220 => x"818d3880",
  2221 => x"e0d408ff",
  2222 => x"2e83ec38",
  2223 => x"73763118",
  2224 => x"80e0a40c",
  2225 => x"73870670",
  2226 => x"57537280",
  2227 => x"2e883888",
  2228 => x"73317015",
  2229 => x"55567614",
  2230 => x"9fff06a0",
  2231 => x"80713117",
  2232 => x"70547f53",
  2233 => x"575383d5",
  2234 => x"3f800853",
  2235 => x"8008ff2e",
  2236 => x"81a03880",
  2237 => x"e0a40816",
  2238 => x"7080e0a4",
  2239 => x"0c747580",
  2240 => x"e0e00b88",
  2241 => x"050c7476",
  2242 => x"31187081",
  2243 => x"07515556",
  2244 => x"587b80e0",
  2245 => x"e02e839c",
  2246 => x"38798f26",
  2247 => x"82cb3881",
  2248 => x"0b84150c",
  2249 => x"841508fc",
  2250 => x"06707a31",
  2251 => x"7a72268f",
  2252 => x"72250752",
  2253 => x"55537280",
  2254 => x"2efcf938",
  2255 => x"80db3980",
  2256 => x"089fff06",
  2257 => x"5372feeb",
  2258 => x"387780e0",
  2259 => x"a40c80e0",
  2260 => x"e00b8805",
  2261 => x"087b1881",
  2262 => x"0784120c",
  2263 => x"5580e0d0",
  2264 => x"08782786",
  2265 => x"387780e0",
  2266 => x"d00c80e0",
  2267 => x"cc087827",
  2268 => x"fcac3877",
  2269 => x"80e0cc0c",
  2270 => x"841508fc",
  2271 => x"06707a31",
  2272 => x"7a72268f",
  2273 => x"72250752",
  2274 => x"55537280",
  2275 => x"2efca538",
  2276 => x"88398074",
  2277 => x"5456fedb",
  2278 => x"397d5182",
  2279 => x"9f3f800b",
  2280 => x"800c8f3d",
  2281 => x"0d047353",
  2282 => x"807424a9",
  2283 => x"3872822c",
  2284 => x"81712b80",
  2285 => x"e0e40807",
  2286 => x"7080e0e0",
  2287 => x"0b84050c",
  2288 => x"5d53778c",
  2289 => x"180c7488",
  2290 => x"180c7688",
  2291 => x"190c768c",
  2292 => x"160cf9b7",
  2293 => x"39831470",
  2294 => x"822c8171",
  2295 => x"2b80e0e4",
  2296 => x"08077080",
  2297 => x"e0e00b84",
  2298 => x"050c5e51",
  2299 => x"53d4397b",
  2300 => x"7b065372",
  2301 => x"fca33884",
  2302 => x"1a7b105c",
  2303 => x"5af139ff",
  2304 => x"1a811151",
  2305 => x"5af7b939",
  2306 => x"78177981",
  2307 => x"0784190c",
  2308 => x"8c180888",
  2309 => x"1908718c",
  2310 => x"120c8812",
  2311 => x"0c597080",
  2312 => x"e0f40c70",
  2313 => x"80e0f00c",
  2314 => x"80e0e80b",
  2315 => x"8c120c8c",
  2316 => x"11088812",
  2317 => x"0c748107",
  2318 => x"84120c74",
  2319 => x"1175710c",
  2320 => x"5153f9bd",
  2321 => x"39751784",
  2322 => x"11088107",
  2323 => x"84120c53",
  2324 => x"8c170888",
  2325 => x"1808718c",
  2326 => x"120c8812",
  2327 => x"0c587d51",
  2328 => x"80da3f88",
  2329 => x"1754f5cf",
  2330 => x"39728415",
  2331 => x"0cf41af8",
  2332 => x"0670841e",
  2333 => x"08810607",
  2334 => x"841e0c70",
  2335 => x"1d545b85",
  2336 => x"0b84140c",
  2337 => x"850b8814",
  2338 => x"0c8f7b27",
  2339 => x"fdcf3888",
  2340 => x"1c527d51",
  2341 => x"82903f80",
  2342 => x"e0e00b88",
  2343 => x"050880e0",
  2344 => x"a4085955",
  2345 => x"fdb73977",
  2346 => x"80e0a40c",
  2347 => x"7380e0d4",
  2348 => x"0cfc9139",
  2349 => x"7284150c",
  2350 => x"fda33904",
  2351 => x"04fd3d0d",
  2352 => x"800b80f0",
  2353 => x"e80c7651",
  2354 => x"86cc3f80",
  2355 => x"08538008",
  2356 => x"ff2e8838",
  2357 => x"72800c85",
  2358 => x"3d0d0480",
  2359 => x"f0e80854",
  2360 => x"73802ef0",
  2361 => x"38757471",
  2362 => x"0c527280",
  2363 => x"0c853d0d",
  2364 => x"04fb3d0d",
  2365 => x"77705256",
  2366 => x"c23f80e0",
  2367 => x"e00b8805",
  2368 => x"08841108",
  2369 => x"fc06707b",
  2370 => x"319fef05",
  2371 => x"e08006e0",
  2372 => x"80055656",
  2373 => x"53a08074",
  2374 => x"24943880",
  2375 => x"527551ff",
  2376 => x"9c3f80e0",
  2377 => x"e8081553",
  2378 => x"7280082e",
  2379 => x"8f387551",
  2380 => x"ff8a3f80",
  2381 => x"5372800c",
  2382 => x"873d0d04",
  2383 => x"73305275",
  2384 => x"51fefa3f",
  2385 => x"8008ff2e",
  2386 => x"a83880e0",
  2387 => x"e00b8805",
  2388 => x"08757531",
  2389 => x"81078412",
  2390 => x"0c5380e0",
  2391 => x"a4087431",
  2392 => x"80e0a40c",
  2393 => x"7551fed4",
  2394 => x"3f810b80",
  2395 => x"0c873d0d",
  2396 => x"04805275",
  2397 => x"51fec63f",
  2398 => x"80e0e00b",
  2399 => x"88050880",
  2400 => x"08713156",
  2401 => x"538f7525",
  2402 => x"ffa43880",
  2403 => x"0880e0d4",
  2404 => x"083180e0",
  2405 => x"a40c7481",
  2406 => x"0784140c",
  2407 => x"7551fe9c",
  2408 => x"3f8053ff",
  2409 => x"9039f63d",
  2410 => x"0d7c7e54",
  2411 => x"5b72802e",
  2412 => x"8283387a",
  2413 => x"51fe843f",
  2414 => x"f8138411",
  2415 => x"0870fe06",
  2416 => x"70138411",
  2417 => x"08fc065d",
  2418 => x"58595458",
  2419 => x"80e0e808",
  2420 => x"752e82de",
  2421 => x"38788416",
  2422 => x"0c807381",
  2423 => x"06545a72",
  2424 => x"7a2e81d5",
  2425 => x"38781584",
  2426 => x"11088106",
  2427 => x"515372a0",
  2428 => x"38781757",
  2429 => x"7981e638",
  2430 => x"88150853",
  2431 => x"7280e0e8",
  2432 => x"2e82f938",
  2433 => x"8c150870",
  2434 => x"8c150c73",
  2435 => x"88120c56",
  2436 => x"76810784",
  2437 => x"190c7618",
  2438 => x"77710c53",
  2439 => x"79819138",
  2440 => x"83ff7727",
  2441 => x"81c83876",
  2442 => x"892a7783",
  2443 => x"2a565372",
  2444 => x"802ebf38",
  2445 => x"76862ab8",
  2446 => x"05558473",
  2447 => x"27b43880",
  2448 => x"db135594",
  2449 => x"7327ab38",
  2450 => x"768c2a80",
  2451 => x"ee055580",
  2452 => x"d473279e",
  2453 => x"38768f2a",
  2454 => x"80f70555",
  2455 => x"82d47327",
  2456 => x"91387692",
  2457 => x"2a80fc05",
  2458 => x"558ad473",
  2459 => x"27843880",
  2460 => x"fe557410",
  2461 => x"101080e0",
  2462 => x"e0058811",
  2463 => x"08555673",
  2464 => x"762e82b3",
  2465 => x"38841408",
  2466 => x"fc065376",
  2467 => x"73278d38",
  2468 => x"88140854",
  2469 => x"73762e09",
  2470 => x"8106ea38",
  2471 => x"8c140870",
  2472 => x"8c1a0c74",
  2473 => x"881a0c78",
  2474 => x"88120c56",
  2475 => x"778c150c",
  2476 => x"7a51fc88",
  2477 => x"3f8c3d0d",
  2478 => x"04770878",
  2479 => x"71315977",
  2480 => x"05881908",
  2481 => x"54577280",
  2482 => x"e0e82e80",
  2483 => x"e0388c18",
  2484 => x"08708c15",
  2485 => x"0c738812",
  2486 => x"0c56fe89",
  2487 => x"39881508",
  2488 => x"8c160870",
  2489 => x"8c130c57",
  2490 => x"88170cfe",
  2491 => x"a3397683",
  2492 => x"2a705455",
  2493 => x"80752481",
  2494 => x"98387282",
  2495 => x"2c81712b",
  2496 => x"80e0e408",
  2497 => x"0780e0e0",
  2498 => x"0b84050c",
  2499 => x"53741010",
  2500 => x"1080e0e0",
  2501 => x"05881108",
  2502 => x"5556758c",
  2503 => x"190c7388",
  2504 => x"190c7788",
  2505 => x"170c778c",
  2506 => x"150cff84",
  2507 => x"39815afd",
  2508 => x"b4397817",
  2509 => x"73810654",
  2510 => x"57729838",
  2511 => x"77087871",
  2512 => x"31597705",
  2513 => x"8c190888",
  2514 => x"1a08718c",
  2515 => x"120c8812",
  2516 => x"0c575776",
  2517 => x"81078419",
  2518 => x"0c7780e0",
  2519 => x"e00b8805",
  2520 => x"0c80e0dc",
  2521 => x"087726fe",
  2522 => x"c73880e0",
  2523 => x"d808527a",
  2524 => x"51fafe3f",
  2525 => x"7a51fac4",
  2526 => x"3ffeba39",
  2527 => x"81788c15",
  2528 => x"0c788815",
  2529 => x"0c738c1a",
  2530 => x"0c73881a",
  2531 => x"0c5afd80",
  2532 => x"39831570",
  2533 => x"822c8171",
  2534 => x"2b80e0e4",
  2535 => x"080780e0",
  2536 => x"e00b8405",
  2537 => x"0c515374",
  2538 => x"10101080",
  2539 => x"e0e00588",
  2540 => x"11085556",
  2541 => x"fee43974",
  2542 => x"53807524",
  2543 => x"a7387282",
  2544 => x"2c81712b",
  2545 => x"80e0e408",
  2546 => x"0780e0e0",
  2547 => x"0b84050c",
  2548 => x"53758c19",
  2549 => x"0c738819",
  2550 => x"0c778817",
  2551 => x"0c778c15",
  2552 => x"0cfdcd39",
  2553 => x"83157082",
  2554 => x"2c81712b",
  2555 => x"80e0e408",
  2556 => x"0780e0e0",
  2557 => x"0b84050c",
  2558 => x"5153d639",
  2559 => x"810b800c",
  2560 => x"04803d0d",
  2561 => x"72812e89",
  2562 => x"38800b80",
  2563 => x"0c823d0d",
  2564 => x"04735180",
  2565 => x"f83ffe3d",
  2566 => x"0d80f0e0",
  2567 => x"0851708a",
  2568 => x"3880f0ec",
  2569 => x"7080f0e0",
  2570 => x"0c517075",
  2571 => x"125252ff",
  2572 => x"537087fb",
  2573 => x"80802688",
  2574 => x"387080f0",
  2575 => x"e00c7153",
  2576 => x"72800c84",
  2577 => x"3d0d04fd",
  2578 => x"3d0d800b",
  2579 => x"80d98008",
  2580 => x"54547281",
  2581 => x"2e9c3873",
  2582 => x"80f0e40c",
  2583 => x"ffb8c23f",
  2584 => x"ffb79d3f",
  2585 => x"80e8e852",
  2586 => x"8151d6b6",
  2587 => x"3f800851",
  2588 => x"a23f7280",
  2589 => x"f0e40cff",
  2590 => x"b8a73fff",
  2591 => x"b7823f80",
  2592 => x"e8e85281",
  2593 => x"51d69b3f",
  2594 => x"80085187",
  2595 => x"3f00ff39",
  2596 => x"00ff39f7",
  2597 => x"3d0d7b80",
  2598 => x"d9a40882",
  2599 => x"c811085a",
  2600 => x"545a7780",
  2601 => x"2e80da38",
  2602 => x"81881884",
  2603 => x"1908ff05",
  2604 => x"81712b59",
  2605 => x"55598074",
  2606 => x"2480ea38",
  2607 => x"807424b5",
  2608 => x"3873822b",
  2609 => x"78118805",
  2610 => x"56568180",
  2611 => x"19087706",
  2612 => x"5372802e",
  2613 => x"b6387816",
  2614 => x"70085353",
  2615 => x"79517408",
  2616 => x"53722dff",
  2617 => x"14fc17fc",
  2618 => x"1779812c",
  2619 => x"5a575754",
  2620 => x"738025d6",
  2621 => x"38770858",
  2622 => x"77ffad38",
  2623 => x"80d9a408",
  2624 => x"53bc1308",
  2625 => x"a5387951",
  2626 => x"ff833f74",
  2627 => x"0853722d",
  2628 => x"ff14fc17",
  2629 => x"fc177981",
  2630 => x"2c5a5757",
  2631 => x"54738025",
  2632 => x"ffa838d1",
  2633 => x"398057ff",
  2634 => x"93397251",
  2635 => x"bc130853",
  2636 => x"722d7951",
  2637 => x"fed73fff",
  2638 => x"3d0d80e8",
  2639 => x"f00bfc05",
  2640 => x"70085252",
  2641 => x"70ff2e91",
  2642 => x"38702dfc",
  2643 => x"12700852",
  2644 => x"5270ff2e",
  2645 => x"098106f1",
  2646 => x"38833d0d",
  2647 => x"0404ffb7",
  2648 => x"ad3f0400",
  2649 => x"00000040",
  2650 => x"3e200000",
  2651 => x"636f6d6d",
  2652 => x"616e6420",
  2653 => x"6e6f7420",
  2654 => x"666f756e",
  2655 => x"642e0a00",
  2656 => x"73657400",
  2657 => x"73657420",
  2658 => x"3c636861",
  2659 => x"6e6e656c",
  2660 => x"3e203c77",
  2661 => x"6169743e",
  2662 => x"203c6f6e",
  2663 => x"3e203c6f",
  2664 => x"66663e20",
  2665 => x"3c636f75",
  2666 => x"6e743e00",
  2667 => x"73746174",
  2668 => x"75730000",
  2669 => x"67657420",
  2670 => x"616c6c20",
  2671 => x"6368616e",
  2672 => x"6e656c20",
  2673 => x"73657474",
  2674 => x"696e6773",
  2675 => x"00000000",
  2676 => x"72756e00",
  2677 => x"67656e65",
  2678 => x"72617465",
  2679 => x"20736967",
  2680 => x"6e616c20",
  2681 => x"6f6e2061",
  2682 => x"6c6c2063",
  2683 => x"68616e6e",
  2684 => x"656c7300",
  2685 => x"73746f70",
  2686 => x"00000000",
  2687 => x"73746f70",
  2688 => x"20616c6c",
  2689 => x"20636861",
  2690 => x"6e6e656c",
  2691 => x"73000000",
  2692 => x"636c6561",
  2693 => x"72000000",
  2694 => x"636c6561",
  2695 => x"72207363",
  2696 => x"7265656e",
  2697 => x"00000000",
  2698 => x"68656c70",
  2699 => x"00000000",
  2700 => x"73757070",
  2701 => x"6f727465",
  2702 => x"6420636f",
  2703 => x"6d6d616e",
  2704 => x"64733a0a",
  2705 => x"0a000000",
  2706 => x"202d2000",
  2707 => x"30780000",
  2708 => x"0a307800",
  2709 => x"203a2000",
  2710 => x"6368616e",
  2711 => x"6e656c20",
  2712 => x"00000000",
  2713 => x"09202073",
  2714 => x"74617475",
  2715 => x"733a2000",
  2716 => x"09202020",
  2717 => x"20776169",
  2718 => x"743a2000",
  2719 => x"09202020",
  2720 => x"2020206f",
  2721 => x"6e3a2000",
  2722 => x"09202020",
  2723 => x"20206f66",
  2724 => x"663a2000",
  2725 => x"09202020",
  2726 => x"636f756e",
  2727 => x"743a2000",
  2728 => x"4572726f",
  2729 => x"723a2077",
  2730 => x"726f6e67",
  2731 => x"20636861",
  2732 => x"6e6e656c",
  2733 => x"206e756d",
  2734 => x"62657220",
  2735 => x"28000000",
  2736 => x"290a0000",
  2737 => x"68656170",
  2738 => x"20707472",
  2739 => x"3a200000",
  2740 => x"66726565",
  2741 => x"206d656d",
  2742 => x"3a200000",
  2743 => x"656e643a",
  2744 => x"20202020",
  2745 => x"20200000",
  2746 => x"0a0a0000",
  2747 => x"63656e74",
  2748 => x"72616c20",
  2749 => x"74726967",
  2750 => x"67657220",
  2751 => x"67656e65",
  2752 => x"7261746f",
  2753 => x"72200000",
  2754 => x"286f6e20",
  2755 => x"73696d29",
  2756 => x"0a000000",
  2757 => x"0a636f6d",
  2758 => x"70696c65",
  2759 => x"643a204d",
  2760 => x"61722032",
  2761 => x"38203230",
  2762 => x"31312020",
  2763 => x"31363a35",
  2764 => x"393a3134",
  2765 => x"0a000000",
  2766 => x"63656e74",
  2767 => x"72616c20",
  2768 => x"20747269",
  2769 => x"67676572",
  2770 => x"00000000",
  2771 => x"67656e65",
  2772 => x"7261746f",
  2773 => x"72000000",
  2774 => x"00202020",
  2775 => x"20202020",
  2776 => x"20202828",
  2777 => x"28282820",
  2778 => x"20202020",
  2779 => x"20202020",
  2780 => x"20202020",
  2781 => x"20202020",
  2782 => x"20881010",
  2783 => x"10101010",
  2784 => x"10101010",
  2785 => x"10101010",
  2786 => x"10040404",
  2787 => x"04040404",
  2788 => x"04040410",
  2789 => x"10101010",
  2790 => x"10104141",
  2791 => x"41414141",
  2792 => x"01010101",
  2793 => x"01010101",
  2794 => x"01010101",
  2795 => x"01010101",
  2796 => x"01010101",
  2797 => x"10101010",
  2798 => x"10104242",
  2799 => x"42424242",
  2800 => x"02020202",
  2801 => x"02020202",
  2802 => x"02020202",
  2803 => x"02020202",
  2804 => x"02020202",
  2805 => x"10101010",
  2806 => x"20000000",
  2807 => x"00000000",
  2808 => x"00000000",
  2809 => x"00000000",
  2810 => x"00000000",
  2811 => x"00000000",
  2812 => x"00000000",
  2813 => x"00000000",
  2814 => x"00000000",
  2815 => x"00000000",
  2816 => x"00000000",
  2817 => x"00000000",
  2818 => x"00000000",
  2819 => x"00000000",
  2820 => x"00000000",
  2821 => x"00000000",
  2822 => x"00000000",
  2823 => x"00000000",
  2824 => x"00000000",
  2825 => x"00000000",
  2826 => x"00000000",
  2827 => x"00000000",
  2828 => x"00000000",
  2829 => x"00000000",
  2830 => x"00000000",
  2831 => x"00000000",
  2832 => x"00000000",
  2833 => x"00000000",
  2834 => x"00000000",
  2835 => x"00000000",
  2836 => x"00000000",
  2837 => x"00000000",
  2838 => x"00000000",
  2839 => x"43000000",
  2840 => x"64756d6d",
  2841 => x"792e6578",
  2842 => x"65000000",
  2843 => x"00ffffff",
  2844 => x"ff00ffff",
  2845 => x"ffff00ff",
  2846 => x"ffffff00",
  2847 => x"00000000",
  2848 => x"00000000",
  2849 => x"00000000",
  2850 => x"00003478",
  2851 => x"80000800",
  2852 => x"80000600",
  2853 => x"80000400",
  2854 => x"80000200",
  2855 => x"80000100",
  2856 => x"80000000",
  2857 => x"00002ca8",
  2858 => x"00000000",
  2859 => x"00002f10",
  2860 => x"00002f6c",
  2861 => x"00002fc8",
  2862 => x"00000000",
  2863 => x"00000000",
  2864 => x"00000000",
  2865 => x"00000000",
  2866 => x"00000000",
  2867 => x"00000000",
  2868 => x"00000000",
  2869 => x"00000000",
  2870 => x"00000000",
  2871 => x"00002c5c",
  2872 => x"00000000",
  2873 => x"00000000",
  2874 => x"00000000",
  2875 => x"00000000",
  2876 => x"00000000",
  2877 => x"00000000",
  2878 => x"00000000",
  2879 => x"00000000",
  2880 => x"00000000",
  2881 => x"00000000",
  2882 => x"00000000",
  2883 => x"00000000",
  2884 => x"00000000",
  2885 => x"00000000",
  2886 => x"00000000",
  2887 => x"00000000",
  2888 => x"00000000",
  2889 => x"00000000",
  2890 => x"00000000",
  2891 => x"00000000",
  2892 => x"00000000",
  2893 => x"00000000",
  2894 => x"00000000",
  2895 => x"00000000",
  2896 => x"00000000",
  2897 => x"00000000",
  2898 => x"00000000",
  2899 => x"00000000",
  2900 => x"00000001",
  2901 => x"330eabcd",
  2902 => x"1234e66d",
  2903 => x"deec0005",
  2904 => x"000b0000",
  2905 => x"00000000",
  2906 => x"00000000",
  2907 => x"00000000",
  2908 => x"00000000",
  2909 => x"00000000",
  2910 => x"00000000",
  2911 => x"00000000",
  2912 => x"00000000",
  2913 => x"00000000",
  2914 => x"00000000",
  2915 => x"00000000",
  2916 => x"00000000",
  2917 => x"00000000",
  2918 => x"00000000",
  2919 => x"00000000",
  2920 => x"00000000",
  2921 => x"00000000",
  2922 => x"00000000",
  2923 => x"00000000",
  2924 => x"00000000",
  2925 => x"00000000",
  2926 => x"00000000",
  2927 => x"00000000",
  2928 => x"00000000",
  2929 => x"00000000",
  2930 => x"00000000",
  2931 => x"00000000",
  2932 => x"00000000",
  2933 => x"00000000",
  2934 => x"00000000",
  2935 => x"00000000",
  2936 => x"00000000",
  2937 => x"00000000",
  2938 => x"00000000",
  2939 => x"00000000",
  2940 => x"00000000",
  2941 => x"00000000",
  2942 => x"00000000",
  2943 => x"00000000",
  2944 => x"00000000",
  2945 => x"00000000",
  2946 => x"00000000",
  2947 => x"00000000",
  2948 => x"00000000",
  2949 => x"00000000",
  2950 => x"00000000",
  2951 => x"00000000",
  2952 => x"00000000",
  2953 => x"00000000",
  2954 => x"00000000",
  2955 => x"00000000",
  2956 => x"00000000",
  2957 => x"00000000",
  2958 => x"00000000",
  2959 => x"00000000",
  2960 => x"00000000",
  2961 => x"00000000",
  2962 => x"00000000",
  2963 => x"00000000",
  2964 => x"00000000",
  2965 => x"00000000",
  2966 => x"00000000",
  2967 => x"00000000",
  2968 => x"00000000",
  2969 => x"00000000",
  2970 => x"00000000",
  2971 => x"00000000",
  2972 => x"00000000",
  2973 => x"00000000",
  2974 => x"00000000",
  2975 => x"00000000",
  2976 => x"00000000",
  2977 => x"00000000",
  2978 => x"00000000",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00000000",
  2983 => x"00000000",
  2984 => x"00000000",
  2985 => x"00000000",
  2986 => x"00000000",
  2987 => x"00000000",
  2988 => x"00000000",
  2989 => x"00000000",
  2990 => x"00000000",
  2991 => x"00000000",
  2992 => x"00000000",
  2993 => x"00000000",
  2994 => x"00000000",
  2995 => x"00000000",
  2996 => x"00000000",
  2997 => x"00000000",
  2998 => x"00000000",
  2999 => x"00000000",
  3000 => x"00000000",
  3001 => x"00000000",
  3002 => x"00000000",
  3003 => x"00000000",
  3004 => x"00000000",
  3005 => x"00000000",
  3006 => x"00000000",
  3007 => x"00000000",
  3008 => x"00000000",
  3009 => x"00000000",
  3010 => x"00000000",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"00000000",
  3015 => x"00000000",
  3016 => x"00000000",
  3017 => x"00000000",
  3018 => x"00000000",
  3019 => x"00000000",
  3020 => x"00000000",
  3021 => x"00000000",
  3022 => x"00000000",
  3023 => x"00000000",
  3024 => x"00000000",
  3025 => x"00000000",
  3026 => x"00000000",
  3027 => x"00000000",
  3028 => x"00000000",
  3029 => x"00000000",
  3030 => x"00000000",
  3031 => x"00000000",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"00000000",
  3041 => x"00000000",
  3042 => x"00000000",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000000",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00000000",
  3050 => x"00000000",
  3051 => x"00000000",
  3052 => x"00000000",
  3053 => x"00000000",
  3054 => x"00000000",
  3055 => x"00000000",
  3056 => x"00000000",
  3057 => x"00000000",
  3058 => x"00000000",
  3059 => x"00000000",
  3060 => x"00000000",
  3061 => x"00000000",
  3062 => x"00000000",
  3063 => x"00000000",
  3064 => x"00000000",
  3065 => x"00000000",
  3066 => x"00000000",
  3067 => x"00000000",
  3068 => x"00000000",
  3069 => x"00000000",
  3070 => x"00000000",
  3071 => x"00000000",
  3072 => x"00000000",
  3073 => x"00000000",
  3074 => x"00000000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000000",
  3084 => x"00000000",
  3085 => x"00000000",
  3086 => x"00000000",
  3087 => x"00000000",
  3088 => x"00000000",
  3089 => x"00000000",
  3090 => x"00000000",
  3091 => x"00000000",
  3092 => x"00000000",
  3093 => x"ffffffff",
  3094 => x"00000000",
  3095 => x"00020000",
  3096 => x"00000000",
  3097 => x"00000000",
  3098 => x"00003060",
  3099 => x"00003060",
  3100 => x"00003068",
  3101 => x"00003068",
  3102 => x"00003070",
  3103 => x"00003070",
  3104 => x"00003078",
  3105 => x"00003078",
  3106 => x"00003080",
  3107 => x"00003080",
  3108 => x"00003088",
  3109 => x"00003088",
  3110 => x"00003090",
  3111 => x"00003090",
  3112 => x"00003098",
  3113 => x"00003098",
  3114 => x"000030a0",
  3115 => x"000030a0",
  3116 => x"000030a8",
  3117 => x"000030a8",
  3118 => x"000030b0",
  3119 => x"000030b0",
  3120 => x"000030b8",
  3121 => x"000030b8",
  3122 => x"000030c0",
  3123 => x"000030c0",
  3124 => x"000030c8",
  3125 => x"000030c8",
  3126 => x"000030d0",
  3127 => x"000030d0",
  3128 => x"000030d8",
  3129 => x"000030d8",
  3130 => x"000030e0",
  3131 => x"000030e0",
  3132 => x"000030e8",
  3133 => x"000030e8",
  3134 => x"000030f0",
  3135 => x"000030f0",
  3136 => x"000030f8",
  3137 => x"000030f8",
  3138 => x"00003100",
  3139 => x"00003100",
  3140 => x"00003108",
  3141 => x"00003108",
  3142 => x"00003110",
  3143 => x"00003110",
  3144 => x"00003118",
  3145 => x"00003118",
  3146 => x"00003120",
  3147 => x"00003120",
  3148 => x"00003128",
  3149 => x"00003128",
  3150 => x"00003130",
  3151 => x"00003130",
  3152 => x"00003138",
  3153 => x"00003138",
  3154 => x"00003140",
  3155 => x"00003140",
  3156 => x"00003148",
  3157 => x"00003148",
  3158 => x"00003150",
  3159 => x"00003150",
  3160 => x"00003158",
  3161 => x"00003158",
  3162 => x"00003160",
  3163 => x"00003160",
  3164 => x"00003168",
  3165 => x"00003168",
  3166 => x"00003170",
  3167 => x"00003170",
  3168 => x"00003178",
  3169 => x"00003178",
  3170 => x"00003180",
  3171 => x"00003180",
  3172 => x"00003188",
  3173 => x"00003188",
  3174 => x"00003190",
  3175 => x"00003190",
  3176 => x"00003198",
  3177 => x"00003198",
  3178 => x"000031a0",
  3179 => x"000031a0",
  3180 => x"000031a8",
  3181 => x"000031a8",
  3182 => x"000031b0",
  3183 => x"000031b0",
  3184 => x"000031b8",
  3185 => x"000031b8",
  3186 => x"000031c0",
  3187 => x"000031c0",
  3188 => x"000031c8",
  3189 => x"000031c8",
  3190 => x"000031d0",
  3191 => x"000031d0",
  3192 => x"000031d8",
  3193 => x"000031d8",
  3194 => x"000031e0",
  3195 => x"000031e0",
  3196 => x"000031e8",
  3197 => x"000031e8",
  3198 => x"000031f0",
  3199 => x"000031f0",
  3200 => x"000031f8",
  3201 => x"000031f8",
  3202 => x"00003200",
  3203 => x"00003200",
  3204 => x"00003208",
  3205 => x"00003208",
  3206 => x"00003210",
  3207 => x"00003210",
  3208 => x"00003218",
  3209 => x"00003218",
  3210 => x"00003220",
  3211 => x"00003220",
  3212 => x"00003228",
  3213 => x"00003228",
  3214 => x"00003230",
  3215 => x"00003230",
  3216 => x"00003238",
  3217 => x"00003238",
  3218 => x"00003240",
  3219 => x"00003240",
  3220 => x"00003248",
  3221 => x"00003248",
  3222 => x"00003250",
  3223 => x"00003250",
  3224 => x"00003258",
  3225 => x"00003258",
  3226 => x"00003260",
  3227 => x"00003260",
  3228 => x"00003268",
  3229 => x"00003268",
  3230 => x"00003270",
  3231 => x"00003270",
  3232 => x"00003278",
  3233 => x"00003278",
  3234 => x"00003280",
  3235 => x"00003280",
  3236 => x"00003288",
  3237 => x"00003288",
  3238 => x"00003290",
  3239 => x"00003290",
  3240 => x"00003298",
  3241 => x"00003298",
  3242 => x"000032a0",
  3243 => x"000032a0",
  3244 => x"000032a8",
  3245 => x"000032a8",
  3246 => x"000032b0",
  3247 => x"000032b0",
  3248 => x"000032b8",
  3249 => x"000032b8",
  3250 => x"000032c0",
  3251 => x"000032c0",
  3252 => x"000032c8",
  3253 => x"000032c8",
  3254 => x"000032d0",
  3255 => x"000032d0",
  3256 => x"000032d8",
  3257 => x"000032d8",
  3258 => x"000032e0",
  3259 => x"000032e0",
  3260 => x"000032e8",
  3261 => x"000032e8",
  3262 => x"000032f0",
  3263 => x"000032f0",
  3264 => x"000032f8",
  3265 => x"000032f8",
  3266 => x"00003300",
  3267 => x"00003300",
  3268 => x"00003308",
  3269 => x"00003308",
  3270 => x"00003310",
  3271 => x"00003310",
  3272 => x"00003318",
  3273 => x"00003318",
  3274 => x"00003320",
  3275 => x"00003320",
  3276 => x"00003328",
  3277 => x"00003328",
  3278 => x"00003330",
  3279 => x"00003330",
  3280 => x"00003338",
  3281 => x"00003338",
  3282 => x"00003340",
  3283 => x"00003340",
  3284 => x"00003348",
  3285 => x"00003348",
  3286 => x"00003350",
  3287 => x"00003350",
  3288 => x"00003358",
  3289 => x"00003358",
  3290 => x"00003360",
  3291 => x"00003360",
  3292 => x"00003368",
  3293 => x"00003368",
  3294 => x"00003370",
  3295 => x"00003370",
  3296 => x"00003378",
  3297 => x"00003378",
  3298 => x"00003380",
  3299 => x"00003380",
  3300 => x"00003388",
  3301 => x"00003388",
  3302 => x"00003390",
  3303 => x"00003390",
  3304 => x"00003398",
  3305 => x"00003398",
  3306 => x"000033a0",
  3307 => x"000033a0",
  3308 => x"000033a8",
  3309 => x"000033a8",
  3310 => x"000033b0",
  3311 => x"000033b0",
  3312 => x"000033b8",
  3313 => x"000033b8",
  3314 => x"000033c0",
  3315 => x"000033c0",
  3316 => x"000033c8",
  3317 => x"000033c8",
  3318 => x"000033d0",
  3319 => x"000033d0",
  3320 => x"000033d8",
  3321 => x"000033d8",
  3322 => x"000033e0",
  3323 => x"000033e0",
  3324 => x"000033e8",
  3325 => x"000033e8",
  3326 => x"000033f0",
  3327 => x"000033f0",
  3328 => x"000033f8",
  3329 => x"000033f8",
  3330 => x"00003400",
  3331 => x"00003400",
  3332 => x"00003408",
  3333 => x"00003408",
  3334 => x"00003410",
  3335 => x"00003410",
  3336 => x"00003418",
  3337 => x"00003418",
  3338 => x"00003420",
  3339 => x"00003420",
  3340 => x"00003428",
  3341 => x"00003428",
  3342 => x"00003430",
  3343 => x"00003430",
  3344 => x"00003438",
  3345 => x"00003438",
  3346 => x"00003440",
  3347 => x"00003440",
  3348 => x"00003448",
  3349 => x"00003448",
  3350 => x"00003450",
  3351 => x"00003450",
  3352 => x"00003458",
  3353 => x"00003458",
  3354 => x"00002c60",
  3355 => x"ffffffff",
  3356 => x"00000000",
  3357 => x"ffffffff",
  3358 => x"00000000",
  3359 => x"00000000",
	others => x"aaaaaaaa" -- mask for mem check
	--others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
