-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80c0c80c",
     3 => x"3a0b0b0b",
     4 => x"b1ff0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0bb2c42d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80c0",
   162 => x"b4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b95",
   171 => x"e62d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b97",
   179 => x"982d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80c0c40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82803fab",
   257 => x"e63f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"53510480",
   280 => x"c0c40880",
   281 => x"2ea43880",
   282 => x"c0c80882",
   283 => x"2ebd3883",
   284 => x"80800b0b",
   285 => x"0b80d0cc",
   286 => x"0c82a080",
   287 => x"0b80d0d0",
   288 => x"0c829080",
   289 => x"0b80d0d4",
   290 => x"0c04f880",
   291 => x"8080a40b",
   292 => x"0b0b80d0",
   293 => x"cc0cf880",
   294 => x"8082800b",
   295 => x"80d0d00c",
   296 => x"f8808084",
   297 => x"800b80d0",
   298 => x"d40c0480",
   299 => x"c0a8808c",
   300 => x"0b0b0b80",
   301 => x"d0cc0c80",
   302 => x"c0a88094",
   303 => x"0b80d0d0",
   304 => x"0c0b0b0b",
   305 => x"b4980b80",
   306 => x"d0d40c04",
   307 => x"ff3d0d80",
   308 => x"d0d83351",
   309 => x"70a73880",
   310 => x"c0d00870",
   311 => x"08525270",
   312 => x"802e9438",
   313 => x"841280c0",
   314 => x"d00c702d",
   315 => x"80c0d008",
   316 => x"70085252",
   317 => x"70ee3881",
   318 => x"0b80d0d8",
   319 => x"34833d0d",
   320 => x"0404803d",
   321 => x"0d0b0b80",
   322 => x"d0c80880",
   323 => x"2e8e380b",
   324 => x"0b0b0b80",
   325 => x"0b802e09",
   326 => x"81068538",
   327 => x"823d0d04",
   328 => x"0b0b80d0",
   329 => x"c8510b0b",
   330 => x"0bf5d53f",
   331 => x"823d0d04",
   332 => x"04ff3d0d",
   333 => x"028f0533",
   334 => x"70525289",
   335 => x"ab3f7151",
   336 => x"8aa13f71",
   337 => x"800c833d",
   338 => x"0d04ff3d",
   339 => x"0d028f05",
   340 => x"3380c0d8",
   341 => x"0871710c",
   342 => x"53800c83",
   343 => x"3d0d04fe",
   344 => x"3d0d800b",
   345 => x"fa808082",
   346 => x"80349b0b",
   347 => x"fa808082",
   348 => x"8134a10b",
   349 => x"fa808082",
   350 => x"823480e7",
   351 => x"0bfa8080",
   352 => x"828334ff",
   353 => x"b80bfa80",
   354 => x"80828434",
   355 => x"ffb80bfa",
   356 => x"80808285",
   357 => x"34de0bfa",
   358 => x"80808286",
   359 => x"34ffad0b",
   360 => x"fa808082",
   361 => x"8734ffbe",
   362 => x"0bfa8080",
   363 => x"828834ef",
   364 => x"0bfa8080",
   365 => x"82893480",
   366 => x"0bfa8080",
   367 => x"828a34a0",
   368 => x"0bfa8080",
   369 => x"828b3488",
   370 => x"0bfa8080",
   371 => x"828c3480",
   372 => x"0bfa8080",
   373 => x"828d3480",
   374 => x"c50bfa80",
   375 => x"80828e34",
   376 => x"800bfa80",
   377 => x"80828f34",
   378 => x"850bfa80",
   379 => x"80829034",
   380 => x"d50bfa80",
   381 => x"80829134",
   382 => x"800bfa80",
   383 => x"80829234",
   384 => x"800bfa80",
   385 => x"80829334",
   386 => x"80c00bfa",
   387 => x"80808294",
   388 => x"34800bfa",
   389 => x"80808295",
   390 => x"34ff0bfa",
   391 => x"80808296",
   392 => x"34910bfa",
   393 => x"80808297",
   394 => x"3480e20b",
   395 => x"fa808082",
   396 => x"9834950b",
   397 => x"fa808082",
   398 => x"99348a0b",
   399 => x"fa808082",
   400 => x"9a34800b",
   401 => x"fa808082",
   402 => x"9b34800b",
   403 => x"fa808082",
   404 => x"9c34820b",
   405 => x"fa808082",
   406 => x"9d348a0b",
   407 => x"fa808082",
   408 => x"9e34800b",
   409 => x"fa808082",
   410 => x"9f34800b",
   411 => x"fa808082",
   412 => x"a034810b",
   413 => x"fa808082",
   414 => x"a134930b",
   415 => x"fa808082",
   416 => x"a234ffba",
   417 => x"0bfa8080",
   418 => x"82a33493",
   419 => x"0bfa8080",
   420 => x"82a434ff",
   421 => x"ba0bfa80",
   422 => x"8082a534",
   423 => x"850bfa80",
   424 => x"8082a634",
   425 => x"c00bfa80",
   426 => x"8082a734",
   427 => x"ffb80bfa",
   428 => x"808082a8",
   429 => x"34f70bfa",
   430 => x"808082a9",
   431 => x"34fa8080",
   432 => x"82800bfa",
   433 => x"80808084",
   434 => x"0cbbe20b",
   435 => x"850a0c80",
   436 => x"c0dc0853",
   437 => x"850a0b94",
   438 => x"140c9173",
   439 => x"0c850a08",
   440 => x"708b2a70",
   441 => x"81065151",
   442 => x"5372f238",
   443 => x"b6845183",
   444 => x"d73f80c0",
   445 => x"dc087008",
   446 => x"5353a051",
   447 => x"83ed3f8a",
   448 => x"5183ab3f",
   449 => x"b6985183",
   450 => x"bf3f80c0",
   451 => x"dc088411",
   452 => x"085353a0",
   453 => x"5183d43f",
   454 => x"8a518392",
   455 => x"3fb6ac51",
   456 => x"83a63f85",
   457 => x"0a0852a0",
   458 => x"5183c03f",
   459 => x"8a5182fe",
   460 => x"3f843d0d",
   461 => x"04f73d0d",
   462 => x"80c0e008",
   463 => x"7008810a",
   464 => x"0680d0dc",
   465 => x"0c5384ee",
   466 => x"3f85873f",
   467 => x"8aca5280",
   468 => x"d0dc0884",
   469 => x"388ab152",
   470 => x"7180d0e0",
   471 => x"0c85e03f",
   472 => x"80c0d408",
   473 => x"53fac98e",
   474 => x"868c730c",
   475 => x"72087084",
   476 => x"2a810655",
   477 => x"5273f538",
   478 => x"80c0dc08",
   479 => x"53ff0b84",
   480 => x"140c9480",
   481 => x"0b88140c",
   482 => x"82d0affd",
   483 => x"fb0b8c14",
   484 => x"0c80c073",
   485 => x"0c720870",
   486 => x"862a8106",
   487 => x"555273f5",
   488 => x"38901308",
   489 => x"70832a81",
   490 => x"06555273",
   491 => x"f43881fc",
   492 => x"80810b90",
   493 => x"140c9013",
   494 => x"0870832a",
   495 => x"81065552",
   496 => x"73f43883",
   497 => x"f0820b90",
   498 => x"140c9013",
   499 => x"0870832a",
   500 => x"81065552",
   501 => x"73f43890",
   502 => x"13087096",
   503 => x"2a810655",
   504 => x"5273d338",
   505 => x"90130870",
   506 => x"832a8106",
   507 => x"555273f4",
   508 => x"3880fdc0",
   509 => x"810b9014",
   510 => x"0cbfac51",
   511 => x"81ca3f80",
   512 => x"d0dc0880",
   513 => x"2e819338",
   514 => x"bfb45181",
   515 => x"bb3fb6dc",
   516 => x"5181b53f",
   517 => x"8052fac7",
   518 => x"3f811270",
   519 => x"81ff0653",
   520 => x"53827227",
   521 => x"f138f881",
   522 => x"c08e8053",
   523 => x"a00b80c0",
   524 => x"e0085555",
   525 => x"80d0dc08",
   526 => x"802eab38",
   527 => x"7281ff06",
   528 => x"84150c72",
   529 => x"9f2a7310",
   530 => x"07537480",
   531 => x"2e9538ff",
   532 => x"157381ff",
   533 => x"0684160c",
   534 => x"739f2a74",
   535 => x"10075455",
   536 => x"74ed3888",
   537 => x"fd3f7281",
   538 => x"ff068415",
   539 => x"0c729f2a",
   540 => x"73100753",
   541 => x"80fd5182",
   542 => x"9a3f80c0",
   543 => x"e0087381",
   544 => x"ff068412",
   545 => x"0c54729f",
   546 => x"2a731007",
   547 => x"5380fd51",
   548 => x"82813f80",
   549 => x"c0e00854",
   550 => x"cd39bfc0",
   551 => x"51aa3fbf",
   552 => x"d051a53f",
   553 => x"b6dc51a0",
   554 => x"3f8052fe",
   555 => x"e939ff3d",
   556 => x"0d028f05",
   557 => x"335180d0",
   558 => x"e0085271",
   559 => x"2d800881",
   560 => x"ff06800c",
   561 => x"833d0d04",
   562 => x"fe3d0d74",
   563 => x"70335353",
   564 => x"71802e93",
   565 => x"38811372",
   566 => x"5280d0e0",
   567 => x"08535371",
   568 => x"2d723352",
   569 => x"71ef3884",
   570 => x"3d0d04f4",
   571 => x"3d0d7f02",
   572 => x"8405bb05",
   573 => x"33555788",
   574 => x"0b8c3d5b",
   575 => x"598b5380",
   576 => x"c0985279",
   577 => x"5187e83f",
   578 => x"73792e81",
   579 => x"80387856",
   580 => x"73902e80",
   581 => x"ed3802a9",
   582 => x"0558768f",
   583 => x"06547389",
   584 => x"2680c338",
   585 => x"7518b015",
   586 => x"55557375",
   587 => x"3476842a",
   588 => x"ff177081",
   589 => x"ff065855",
   590 => x"5775df38",
   591 => x"8e3d7905",
   592 => x"f6055775",
   593 => x"77347970",
   594 => x"33555573",
   595 => x"802e9338",
   596 => x"81157452",
   597 => x"80d0e008",
   598 => x"5755752d",
   599 => x"74335473",
   600 => x"ef388e3d",
   601 => x"0d047518",
   602 => x"b7155555",
   603 => x"73753476",
   604 => x"842aff17",
   605 => x"7081ff06",
   606 => x"58555775",
   607 => x"ff9c38ff",
   608 => x"bb398470",
   609 => x"575902a9",
   610 => x"0558ff8e",
   611 => x"39827057",
   612 => x"59f439fd",
   613 => x"3d0d80c0",
   614 => x"e80876b0",
   615 => x"ea299412",
   616 => x"0c54850b",
   617 => x"98150c98",
   618 => x"14087081",
   619 => x"06515372",
   620 => x"f638853d",
   621 => x"0d04803d",
   622 => x"0d80c0e8",
   623 => x"0851870b",
   624 => x"84120cb0",
   625 => x"ea0ba412",
   626 => x"0c870ba8",
   627 => x"120c823d",
   628 => x"0d04803d",
   629 => x"0d80c0ec",
   630 => x"0851b60b",
   631 => x"8c120c83",
   632 => x"0b88120c",
   633 => x"823d0d04",
   634 => x"fe3d0d02",
   635 => x"93053353",
   636 => x"728a2e9e",
   637 => x"3880c0ec",
   638 => x"08528412",
   639 => x"0870822a",
   640 => x"70810651",
   641 => x"51517080",
   642 => x"2ef03872",
   643 => x"720c843d",
   644 => x"0d0480c0",
   645 => x"ec085284",
   646 => x"12087082",
   647 => x"2a708106",
   648 => x"51515170",
   649 => x"802ef038",
   650 => x"8d720c84",
   651 => x"12087082",
   652 => x"2a708106",
   653 => x"51515170",
   654 => x"802effbe",
   655 => x"38cd3980",
   656 => x"3d0d80c0",
   657 => x"e4085180",
   658 => x"0b84120c",
   659 => x"fe800a0b",
   660 => x"88120c80",
   661 => x"0b80d0e4",
   662 => x"34800b80",
   663 => x"d0e83482",
   664 => x"3d0d04fa",
   665 => x"3d0d02a3",
   666 => x"053380c0",
   667 => x"e40880d0",
   668 => x"e4337081",
   669 => x"ff067010",
   670 => x"101180d0",
   671 => x"e8337081",
   672 => x"ff067290",
   673 => x"29117088",
   674 => x"2b780777",
   675 => x"0c535b5b",
   676 => x"55555954",
   677 => x"54738a2e",
   678 => x"98387480",
   679 => x"cf2e9238",
   680 => x"738c2ea4",
   681 => x"38811653",
   682 => x"7280d0e8",
   683 => x"34883d0d",
   684 => x"0471a326",
   685 => x"a3388117",
   686 => x"527180d0",
   687 => x"e434800b",
   688 => x"80d0e834",
   689 => x"883d0d04",
   690 => x"80527188",
   691 => x"2b730c81",
   692 => x"12529790",
   693 => x"7226f338",
   694 => x"800b80d0",
   695 => x"e434800b",
   696 => x"80d0e834",
   697 => x"df398c08",
   698 => x"028c0cf9",
   699 => x"3d0d800b",
   700 => x"8c08fc05",
   701 => x"0c8c0888",
   702 => x"05088025",
   703 => x"ab388c08",
   704 => x"88050830",
   705 => x"8c088805",
   706 => x"0c800b8c",
   707 => x"08f4050c",
   708 => x"8c08fc05",
   709 => x"08883881",
   710 => x"0b8c08f4",
   711 => x"050c8c08",
   712 => x"f405088c",
   713 => x"08fc050c",
   714 => x"8c088c05",
   715 => x"088025ab",
   716 => x"388c088c",
   717 => x"0508308c",
   718 => x"088c050c",
   719 => x"800b8c08",
   720 => x"f0050c8c",
   721 => x"08fc0508",
   722 => x"8838810b",
   723 => x"8c08f005",
   724 => x"0c8c08f0",
   725 => x"05088c08",
   726 => x"fc050c80",
   727 => x"538c088c",
   728 => x"0508528c",
   729 => x"08880508",
   730 => x"5181a73f",
   731 => x"8008708c",
   732 => x"08f8050c",
   733 => x"548c08fc",
   734 => x"0508802e",
   735 => x"8c388c08",
   736 => x"f8050830",
   737 => x"8c08f805",
   738 => x"0c8c08f8",
   739 => x"05087080",
   740 => x"0c54893d",
   741 => x"0d8c0c04",
   742 => x"8c08028c",
   743 => x"0cfb3d0d",
   744 => x"800b8c08",
   745 => x"fc050c8c",
   746 => x"08880508",
   747 => x"80259338",
   748 => x"8c088805",
   749 => x"08308c08",
   750 => x"88050c81",
   751 => x"0b8c08fc",
   752 => x"050c8c08",
   753 => x"8c050880",
   754 => x"258c388c",
   755 => x"088c0508",
   756 => x"308c088c",
   757 => x"050c8153",
   758 => x"8c088c05",
   759 => x"08528c08",
   760 => x"88050851",
   761 => x"ad3f8008",
   762 => x"708c08f8",
   763 => x"050c548c",
   764 => x"08fc0508",
   765 => x"802e8c38",
   766 => x"8c08f805",
   767 => x"08308c08",
   768 => x"f8050c8c",
   769 => x"08f80508",
   770 => x"70800c54",
   771 => x"873d0d8c",
   772 => x"0c048c08",
   773 => x"028c0cfd",
   774 => x"3d0d810b",
   775 => x"8c08fc05",
   776 => x"0c800b8c",
   777 => x"08f8050c",
   778 => x"8c088c05",
   779 => x"088c0888",
   780 => x"050827ac",
   781 => x"388c08fc",
   782 => x"0508802e",
   783 => x"a338800b",
   784 => x"8c088c05",
   785 => x"08249938",
   786 => x"8c088c05",
   787 => x"08108c08",
   788 => x"8c050c8c",
   789 => x"08fc0508",
   790 => x"108c08fc",
   791 => x"050cc939",
   792 => x"8c08fc05",
   793 => x"08802e80",
   794 => x"c9388c08",
   795 => x"8c05088c",
   796 => x"08880508",
   797 => x"26a1388c",
   798 => x"08880508",
   799 => x"8c088c05",
   800 => x"08318c08",
   801 => x"88050c8c",
   802 => x"08f80508",
   803 => x"8c08fc05",
   804 => x"08078c08",
   805 => x"f8050c8c",
   806 => x"08fc0508",
   807 => x"812a8c08",
   808 => x"fc050c8c",
   809 => x"088c0508",
   810 => x"812a8c08",
   811 => x"8c050cff",
   812 => x"af398c08",
   813 => x"90050880",
   814 => x"2e8f388c",
   815 => x"08880508",
   816 => x"708c08f4",
   817 => x"050c518d",
   818 => x"398c08f8",
   819 => x"0508708c",
   820 => x"08f4050c",
   821 => x"518c08f4",
   822 => x"0508800c",
   823 => x"853d0d8c",
   824 => x"0c04803d",
   825 => x"0d865184",
   826 => x"963f8151",
   827 => x"98d33ffc",
   828 => x"3d0d7670",
   829 => x"797b5555",
   830 => x"55558f72",
   831 => x"278c3872",
   832 => x"75078306",
   833 => x"5170802e",
   834 => x"a738ff12",
   835 => x"5271ff2e",
   836 => x"98387270",
   837 => x"81055433",
   838 => x"74708105",
   839 => x"5634ff12",
   840 => x"5271ff2e",
   841 => x"098106ea",
   842 => x"3874800c",
   843 => x"863d0d04",
   844 => x"74517270",
   845 => x"84055408",
   846 => x"71708405",
   847 => x"530c7270",
   848 => x"84055408",
   849 => x"71708405",
   850 => x"530c7270",
   851 => x"84055408",
   852 => x"71708405",
   853 => x"530c7270",
   854 => x"84055408",
   855 => x"71708405",
   856 => x"530cf012",
   857 => x"52718f26",
   858 => x"c9388372",
   859 => x"27953872",
   860 => x"70840554",
   861 => x"08717084",
   862 => x"05530cfc",
   863 => x"12527183",
   864 => x"26ed3870",
   865 => x"54ff8339",
   866 => x"fd3d0d75",
   867 => x"5384d813",
   868 => x"08802e8a",
   869 => x"38805372",
   870 => x"800c853d",
   871 => x"0d048180",
   872 => x"52725183",
   873 => x"d83f8008",
   874 => x"84d8140c",
   875 => x"ff538008",
   876 => x"802ee438",
   877 => x"8008549f",
   878 => x"53807470",
   879 => x"8405560c",
   880 => x"ff135380",
   881 => x"7324ce38",
   882 => x"80747084",
   883 => x"05560cff",
   884 => x"13537280",
   885 => x"25e338ff",
   886 => x"bc39fd3d",
   887 => x"0d757755",
   888 => x"539f7427",
   889 => x"8d389673",
   890 => x"0cff5271",
   891 => x"800c853d",
   892 => x"0d0484d8",
   893 => x"13085271",
   894 => x"802e9338",
   895 => x"73101012",
   896 => x"70087972",
   897 => x"0c515271",
   898 => x"800c853d",
   899 => x"0d047251",
   900 => x"fef63fff",
   901 => x"528008d3",
   902 => x"3884d813",
   903 => x"08741010",
   904 => x"1170087a",
   905 => x"720c5151",
   906 => x"52dd39f9",
   907 => x"3d0d797b",
   908 => x"5856769f",
   909 => x"2680e838",
   910 => x"84d81608",
   911 => x"5473802e",
   912 => x"aa387610",
   913 => x"10147008",
   914 => x"55557380",
   915 => x"2eba3880",
   916 => x"5873812e",
   917 => x"8f3873ff",
   918 => x"2ea33880",
   919 => x"750c7651",
   920 => x"732d8058",
   921 => x"77800c89",
   922 => x"3d0d0475",
   923 => x"51fe993f",
   924 => x"ff588008",
   925 => x"ef3884d8",
   926 => x"160854c6",
   927 => x"3996760c",
   928 => x"810b800c",
   929 => x"893d0d04",
   930 => x"755181ed",
   931 => x"3f765380",
   932 => x"08527551",
   933 => x"81ad3f80",
   934 => x"08800c89",
   935 => x"3d0d0496",
   936 => x"760cff0b",
   937 => x"800c893d",
   938 => x"0d04fc3d",
   939 => x"0d767856",
   940 => x"53ff5474",
   941 => x"9f26b138",
   942 => x"84d81308",
   943 => x"5271802e",
   944 => x"ae387410",
   945 => x"10127008",
   946 => x"53538154",
   947 => x"71802e98",
   948 => x"38825471",
   949 => x"ff2e9138",
   950 => x"83547181",
   951 => x"2e8a3880",
   952 => x"730c7451",
   953 => x"712d8054",
   954 => x"73800c86",
   955 => x"3d0d0472",
   956 => x"51fd953f",
   957 => x"8008f138",
   958 => x"84d81308",
   959 => x"52c439ff",
   960 => x"3d0d7352",
   961 => x"80c0f008",
   962 => x"51fea03f",
   963 => x"833d0d04",
   964 => x"fe3d0d75",
   965 => x"53745280",
   966 => x"c0f00851",
   967 => x"fdbc3f84",
   968 => x"3d0d0480",
   969 => x"3d0d80c0",
   970 => x"f00851fc",
   971 => x"db3f823d",
   972 => x"0d04ff3d",
   973 => x"0d735280",
   974 => x"c0f00851",
   975 => x"feec3f83",
   976 => x"3d0d04fc",
   977 => x"3d0d800b",
   978 => x"80d0f40c",
   979 => x"78527751",
   980 => x"92e73f80",
   981 => x"08548008",
   982 => x"ff2e8838",
   983 => x"73800c86",
   984 => x"3d0d0480",
   985 => x"d0f40855",
   986 => x"74802ef0",
   987 => x"38767571",
   988 => x"0c537380",
   989 => x"0c863d0d",
   990 => x"0492b93f",
   991 => x"04f33d0d",
   992 => x"7f618b11",
   993 => x"70f8065c",
   994 => x"55555e72",
   995 => x"96268338",
   996 => x"90598079",
   997 => x"24747a26",
   998 => x"07538054",
   999 => x"72742e09",
  1000 => x"810680cb",
  1001 => x"387d518b",
  1002 => x"ca3f7883",
  1003 => x"f72680c6",
  1004 => x"3878832a",
  1005 => x"70101010",
  1006 => x"80c8ac05",
  1007 => x"8c110859",
  1008 => x"595a7678",
  1009 => x"2e83b038",
  1010 => x"841708fc",
  1011 => x"06568c17",
  1012 => x"08881808",
  1013 => x"718c120c",
  1014 => x"88120c58",
  1015 => x"75178411",
  1016 => x"08810784",
  1017 => x"120c537d",
  1018 => x"518b893f",
  1019 => x"88175473",
  1020 => x"800c8f3d",
  1021 => x"0d047889",
  1022 => x"2a79832a",
  1023 => x"5b537280",
  1024 => x"2ebf3878",
  1025 => x"862ab805",
  1026 => x"5a847327",
  1027 => x"b43880db",
  1028 => x"135a9473",
  1029 => x"27ab3878",
  1030 => x"8c2a80ee",
  1031 => x"055a80d4",
  1032 => x"73279e38",
  1033 => x"788f2a80",
  1034 => x"f7055a82",
  1035 => x"d4732791",
  1036 => x"3878922a",
  1037 => x"80fc055a",
  1038 => x"8ad47327",
  1039 => x"843880fe",
  1040 => x"5a791010",
  1041 => x"1080c8ac",
  1042 => x"058c1108",
  1043 => x"58557675",
  1044 => x"2ea33884",
  1045 => x"1708fc06",
  1046 => x"707a3155",
  1047 => x"56738f24",
  1048 => x"88d53873",
  1049 => x"8025fee6",
  1050 => x"388c1708",
  1051 => x"5776752e",
  1052 => x"098106df",
  1053 => x"38811a5a",
  1054 => x"80c8bc08",
  1055 => x"577680c8",
  1056 => x"b42e82c0",
  1057 => x"38841708",
  1058 => x"fc06707a",
  1059 => x"31555673",
  1060 => x"8f2481f9",
  1061 => x"3880c8b4",
  1062 => x"0b80c8c0",
  1063 => x"0c80c8b4",
  1064 => x"0b80c8bc",
  1065 => x"0c738025",
  1066 => x"feb23883",
  1067 => x"ff762783",
  1068 => x"df387589",
  1069 => x"2a76832a",
  1070 => x"55537280",
  1071 => x"2ebf3875",
  1072 => x"862ab805",
  1073 => x"54847327",
  1074 => x"b43880db",
  1075 => x"13549473",
  1076 => x"27ab3875",
  1077 => x"8c2a80ee",
  1078 => x"055480d4",
  1079 => x"73279e38",
  1080 => x"758f2a80",
  1081 => x"f7055482",
  1082 => x"d4732791",
  1083 => x"3875922a",
  1084 => x"80fc0554",
  1085 => x"8ad47327",
  1086 => x"843880fe",
  1087 => x"54731010",
  1088 => x"1080c8ac",
  1089 => x"05881108",
  1090 => x"56587478",
  1091 => x"2e86cf38",
  1092 => x"841508fc",
  1093 => x"06537573",
  1094 => x"278d3888",
  1095 => x"15085574",
  1096 => x"782e0981",
  1097 => x"06ea388c",
  1098 => x"150880c8",
  1099 => x"ac0b8405",
  1100 => x"08718c1a",
  1101 => x"0c76881a",
  1102 => x"0c788813",
  1103 => x"0c788c18",
  1104 => x"0c5d5879",
  1105 => x"53807a24",
  1106 => x"83e63872",
  1107 => x"822c8171",
  1108 => x"2b5c537a",
  1109 => x"7c268198",
  1110 => x"387b7b06",
  1111 => x"537282f1",
  1112 => x"3879fc06",
  1113 => x"84055a7a",
  1114 => x"10707d06",
  1115 => x"545b7282",
  1116 => x"e038841a",
  1117 => x"5af13988",
  1118 => x"178c1108",
  1119 => x"58587678",
  1120 => x"2e098106",
  1121 => x"fcc23882",
  1122 => x"1a5afdec",
  1123 => x"39781779",
  1124 => x"81078419",
  1125 => x"0c7080c8",
  1126 => x"c00c7080",
  1127 => x"c8bc0c80",
  1128 => x"c8b40b8c",
  1129 => x"120c8c11",
  1130 => x"0888120c",
  1131 => x"74810784",
  1132 => x"120c7411",
  1133 => x"75710c51",
  1134 => x"537d5187",
  1135 => x"b73f8817",
  1136 => x"54fcac39",
  1137 => x"80c8ac0b",
  1138 => x"8405087a",
  1139 => x"545c7980",
  1140 => x"25fef838",
  1141 => x"82da397a",
  1142 => x"097c0670",
  1143 => x"80c8ac0b",
  1144 => x"84050c5c",
  1145 => x"7a105b7a",
  1146 => x"7c268538",
  1147 => x"7a85b838",
  1148 => x"80c8ac0b",
  1149 => x"88050870",
  1150 => x"841208fc",
  1151 => x"06707c31",
  1152 => x"7c72268f",
  1153 => x"72250757",
  1154 => x"575c5d55",
  1155 => x"72802e80",
  1156 => x"db38797a",
  1157 => x"1680c8a4",
  1158 => x"081b9011",
  1159 => x"5a55575b",
  1160 => x"80c8a008",
  1161 => x"ff2e8838",
  1162 => x"a08f13e0",
  1163 => x"80065776",
  1164 => x"527d5186",
  1165 => x"c03f8008",
  1166 => x"548008ff",
  1167 => x"2e903880",
  1168 => x"08762782",
  1169 => x"99387480",
  1170 => x"c8ac2e82",
  1171 => x"913880c8",
  1172 => x"ac0b8805",
  1173 => x"08558415",
  1174 => x"08fc0670",
  1175 => x"7a317a72",
  1176 => x"268f7225",
  1177 => x"07525553",
  1178 => x"7283e638",
  1179 => x"74798107",
  1180 => x"84170c79",
  1181 => x"167080c8",
  1182 => x"ac0b8805",
  1183 => x"0c758107",
  1184 => x"84120c54",
  1185 => x"7e525785",
  1186 => x"eb3f8817",
  1187 => x"54fae039",
  1188 => x"75832a70",
  1189 => x"54548074",
  1190 => x"24819b38",
  1191 => x"72822c81",
  1192 => x"712b80c8",
  1193 => x"b0080770",
  1194 => x"80c8ac0b",
  1195 => x"84050c75",
  1196 => x"10101080",
  1197 => x"c8ac0588",
  1198 => x"1108585a",
  1199 => x"5d53778c",
  1200 => x"180c7488",
  1201 => x"180c7688",
  1202 => x"190c768c",
  1203 => x"160cfcf3",
  1204 => x"39797a10",
  1205 => x"101080c8",
  1206 => x"ac057057",
  1207 => x"595d8c15",
  1208 => x"08577675",
  1209 => x"2ea33884",
  1210 => x"1708fc06",
  1211 => x"707a3155",
  1212 => x"56738f24",
  1213 => x"83ca3873",
  1214 => x"80258481",
  1215 => x"388c1708",
  1216 => x"5776752e",
  1217 => x"098106df",
  1218 => x"38881581",
  1219 => x"1b708306",
  1220 => x"555b5572",
  1221 => x"c9387c83",
  1222 => x"06537280",
  1223 => x"2efdb838",
  1224 => x"ff1df819",
  1225 => x"595d8818",
  1226 => x"08782eea",
  1227 => x"38fdb539",
  1228 => x"831a53fc",
  1229 => x"96398314",
  1230 => x"70822c81",
  1231 => x"712b80c8",
  1232 => x"b0080770",
  1233 => x"80c8ac0b",
  1234 => x"84050c76",
  1235 => x"10101080",
  1236 => x"c8ac0588",
  1237 => x"1108595b",
  1238 => x"5e5153fe",
  1239 => x"e13980c7",
  1240 => x"f0081758",
  1241 => x"8008762e",
  1242 => x"818d3880",
  1243 => x"c8a008ff",
  1244 => x"2e83ec38",
  1245 => x"73763118",
  1246 => x"80c7f00c",
  1247 => x"73870670",
  1248 => x"57537280",
  1249 => x"2e883888",
  1250 => x"73317015",
  1251 => x"55567614",
  1252 => x"9fff06a0",
  1253 => x"80713117",
  1254 => x"70547f53",
  1255 => x"575383d5",
  1256 => x"3f800853",
  1257 => x"8008ff2e",
  1258 => x"81a03880",
  1259 => x"c7f00816",
  1260 => x"7080c7f0",
  1261 => x"0c747580",
  1262 => x"c8ac0b88",
  1263 => x"050c7476",
  1264 => x"31187081",
  1265 => x"07515556",
  1266 => x"587b80c8",
  1267 => x"ac2e839c",
  1268 => x"38798f26",
  1269 => x"82cb3881",
  1270 => x"0b84150c",
  1271 => x"841508fc",
  1272 => x"06707a31",
  1273 => x"7a72268f",
  1274 => x"72250752",
  1275 => x"55537280",
  1276 => x"2efcf938",
  1277 => x"80db3980",
  1278 => x"089fff06",
  1279 => x"5372feeb",
  1280 => x"387780c7",
  1281 => x"f00c80c8",
  1282 => x"ac0b8805",
  1283 => x"087b1881",
  1284 => x"0784120c",
  1285 => x"5580c89c",
  1286 => x"08782786",
  1287 => x"387780c8",
  1288 => x"9c0c80c8",
  1289 => x"98087827",
  1290 => x"fcac3877",
  1291 => x"80c8980c",
  1292 => x"841508fc",
  1293 => x"06707a31",
  1294 => x"7a72268f",
  1295 => x"72250752",
  1296 => x"55537280",
  1297 => x"2efca538",
  1298 => x"88398074",
  1299 => x"5456fedb",
  1300 => x"397d5182",
  1301 => x"9f3f800b",
  1302 => x"800c8f3d",
  1303 => x"0d047353",
  1304 => x"807424a9",
  1305 => x"3872822c",
  1306 => x"81712b80",
  1307 => x"c8b00807",
  1308 => x"7080c8ac",
  1309 => x"0b84050c",
  1310 => x"5d53778c",
  1311 => x"180c7488",
  1312 => x"180c7688",
  1313 => x"190c768c",
  1314 => x"160cf9b7",
  1315 => x"39831470",
  1316 => x"822c8171",
  1317 => x"2b80c8b0",
  1318 => x"08077080",
  1319 => x"c8ac0b84",
  1320 => x"050c5e51",
  1321 => x"53d4397b",
  1322 => x"7b065372",
  1323 => x"fca33884",
  1324 => x"1a7b105c",
  1325 => x"5af139ff",
  1326 => x"1a811151",
  1327 => x"5af7b939",
  1328 => x"78177981",
  1329 => x"0784190c",
  1330 => x"8c180888",
  1331 => x"1908718c",
  1332 => x"120c8812",
  1333 => x"0c597080",
  1334 => x"c8c00c70",
  1335 => x"80c8bc0c",
  1336 => x"80c8b40b",
  1337 => x"8c120c8c",
  1338 => x"11088812",
  1339 => x"0c748107",
  1340 => x"84120c74",
  1341 => x"1175710c",
  1342 => x"5153f9bd",
  1343 => x"39751784",
  1344 => x"11088107",
  1345 => x"84120c53",
  1346 => x"8c170888",
  1347 => x"1808718c",
  1348 => x"120c8812",
  1349 => x"0c587d51",
  1350 => x"80da3f88",
  1351 => x"1754f5cf",
  1352 => x"39728415",
  1353 => x"0cf41af8",
  1354 => x"0670841e",
  1355 => x"08810607",
  1356 => x"841e0c70",
  1357 => x"1d545b85",
  1358 => x"0b84140c",
  1359 => x"850b8814",
  1360 => x"0c8f7b27",
  1361 => x"fdcf3888",
  1362 => x"1c527d51",
  1363 => x"82903f80",
  1364 => x"c8ac0b88",
  1365 => x"050880c7",
  1366 => x"f0085955",
  1367 => x"fdb73977",
  1368 => x"80c7f00c",
  1369 => x"7380c8a0",
  1370 => x"0cfc9139",
  1371 => x"7284150c",
  1372 => x"fda33904",
  1373 => x"04fd3d0d",
  1374 => x"800b80d0",
  1375 => x"f40c7651",
  1376 => x"86cc3f80",
  1377 => x"08538008",
  1378 => x"ff2e8838",
  1379 => x"72800c85",
  1380 => x"3d0d0480",
  1381 => x"d0f40854",
  1382 => x"73802ef0",
  1383 => x"38757471",
  1384 => x"0c527280",
  1385 => x"0c853d0d",
  1386 => x"04fb3d0d",
  1387 => x"77705256",
  1388 => x"c23f80c8",
  1389 => x"ac0b8805",
  1390 => x"08841108",
  1391 => x"fc06707b",
  1392 => x"319fef05",
  1393 => x"e08006e0",
  1394 => x"80055656",
  1395 => x"53a08074",
  1396 => x"24943880",
  1397 => x"527551ff",
  1398 => x"9c3f80c8",
  1399 => x"b4081553",
  1400 => x"7280082e",
  1401 => x"8f387551",
  1402 => x"ff8a3f80",
  1403 => x"5372800c",
  1404 => x"873d0d04",
  1405 => x"73305275",
  1406 => x"51fefa3f",
  1407 => x"8008ff2e",
  1408 => x"a83880c8",
  1409 => x"ac0b8805",
  1410 => x"08757531",
  1411 => x"81078412",
  1412 => x"0c5380c7",
  1413 => x"f0087431",
  1414 => x"80c7f00c",
  1415 => x"7551fed4",
  1416 => x"3f810b80",
  1417 => x"0c873d0d",
  1418 => x"04805275",
  1419 => x"51fec63f",
  1420 => x"80c8ac0b",
  1421 => x"88050880",
  1422 => x"08713156",
  1423 => x"538f7525",
  1424 => x"ffa43880",
  1425 => x"0880c8a0",
  1426 => x"083180c7",
  1427 => x"f00c7481",
  1428 => x"0784140c",
  1429 => x"7551fe9c",
  1430 => x"3f8053ff",
  1431 => x"9039f63d",
  1432 => x"0d7c7e54",
  1433 => x"5b72802e",
  1434 => x"8283387a",
  1435 => x"51fe843f",
  1436 => x"f8138411",
  1437 => x"0870fe06",
  1438 => x"70138411",
  1439 => x"08fc065d",
  1440 => x"58595458",
  1441 => x"80c8b408",
  1442 => x"752e82de",
  1443 => x"38788416",
  1444 => x"0c807381",
  1445 => x"06545a72",
  1446 => x"7a2e81d5",
  1447 => x"38781584",
  1448 => x"11088106",
  1449 => x"515372a0",
  1450 => x"38781757",
  1451 => x"7981e638",
  1452 => x"88150853",
  1453 => x"7280c8b4",
  1454 => x"2e82f938",
  1455 => x"8c150870",
  1456 => x"8c150c73",
  1457 => x"88120c56",
  1458 => x"76810784",
  1459 => x"190c7618",
  1460 => x"77710c53",
  1461 => x"79819138",
  1462 => x"83ff7727",
  1463 => x"81c83876",
  1464 => x"892a7783",
  1465 => x"2a565372",
  1466 => x"802ebf38",
  1467 => x"76862ab8",
  1468 => x"05558473",
  1469 => x"27b43880",
  1470 => x"db135594",
  1471 => x"7327ab38",
  1472 => x"768c2a80",
  1473 => x"ee055580",
  1474 => x"d473279e",
  1475 => x"38768f2a",
  1476 => x"80f70555",
  1477 => x"82d47327",
  1478 => x"91387692",
  1479 => x"2a80fc05",
  1480 => x"558ad473",
  1481 => x"27843880",
  1482 => x"fe557410",
  1483 => x"101080c8",
  1484 => x"ac058811",
  1485 => x"08555673",
  1486 => x"762e82b3",
  1487 => x"38841408",
  1488 => x"fc065376",
  1489 => x"73278d38",
  1490 => x"88140854",
  1491 => x"73762e09",
  1492 => x"8106ea38",
  1493 => x"8c140870",
  1494 => x"8c1a0c74",
  1495 => x"881a0c78",
  1496 => x"88120c56",
  1497 => x"778c150c",
  1498 => x"7a51fc88",
  1499 => x"3f8c3d0d",
  1500 => x"04770878",
  1501 => x"71315977",
  1502 => x"05881908",
  1503 => x"54577280",
  1504 => x"c8b42e80",
  1505 => x"e0388c18",
  1506 => x"08708c15",
  1507 => x"0c738812",
  1508 => x"0c56fe89",
  1509 => x"39881508",
  1510 => x"8c160870",
  1511 => x"8c130c57",
  1512 => x"88170cfe",
  1513 => x"a3397683",
  1514 => x"2a705455",
  1515 => x"80752481",
  1516 => x"98387282",
  1517 => x"2c81712b",
  1518 => x"80c8b008",
  1519 => x"0780c8ac",
  1520 => x"0b84050c",
  1521 => x"53741010",
  1522 => x"1080c8ac",
  1523 => x"05881108",
  1524 => x"5556758c",
  1525 => x"190c7388",
  1526 => x"190c7788",
  1527 => x"170c778c",
  1528 => x"150cff84",
  1529 => x"39815afd",
  1530 => x"b4397817",
  1531 => x"73810654",
  1532 => x"57729838",
  1533 => x"77087871",
  1534 => x"31597705",
  1535 => x"8c190888",
  1536 => x"1a08718c",
  1537 => x"120c8812",
  1538 => x"0c575776",
  1539 => x"81078419",
  1540 => x"0c7780c8",
  1541 => x"ac0b8805",
  1542 => x"0c80c8a8",
  1543 => x"087726fe",
  1544 => x"c73880c8",
  1545 => x"a408527a",
  1546 => x"51fafe3f",
  1547 => x"7a51fac4",
  1548 => x"3ffeba39",
  1549 => x"81788c15",
  1550 => x"0c788815",
  1551 => x"0c738c1a",
  1552 => x"0c73881a",
  1553 => x"0c5afd80",
  1554 => x"39831570",
  1555 => x"822c8171",
  1556 => x"2b80c8b0",
  1557 => x"080780c8",
  1558 => x"ac0b8405",
  1559 => x"0c515374",
  1560 => x"10101080",
  1561 => x"c8ac0588",
  1562 => x"11085556",
  1563 => x"fee43974",
  1564 => x"53807524",
  1565 => x"a7387282",
  1566 => x"2c81712b",
  1567 => x"80c8b008",
  1568 => x"0780c8ac",
  1569 => x"0b84050c",
  1570 => x"53758c19",
  1571 => x"0c738819",
  1572 => x"0c778817",
  1573 => x"0c778c15",
  1574 => x"0cfdcd39",
  1575 => x"83157082",
  1576 => x"2c81712b",
  1577 => x"80c8b008",
  1578 => x"0780c8ac",
  1579 => x"0b84050c",
  1580 => x"5153d639",
  1581 => x"810b800c",
  1582 => x"04803d0d",
  1583 => x"72812e89",
  1584 => x"38800b80",
  1585 => x"0c823d0d",
  1586 => x"04735180",
  1587 => x"f43ffe3d",
  1588 => x"0d80d0ec",
  1589 => x"0851708a",
  1590 => x"3880d0f8",
  1591 => x"7080d0ec",
  1592 => x"0c517075",
  1593 => x"125252ff",
  1594 => x"537087fb",
  1595 => x"80802688",
  1596 => x"387080d0",
  1597 => x"ec0c7153",
  1598 => x"72800c84",
  1599 => x"3d0d04fd",
  1600 => x"3d0d800b",
  1601 => x"80c0c808",
  1602 => x"54547281",
  1603 => x"2e9a3873",
  1604 => x"80d0f00c",
  1605 => x"d6c93fd5",
  1606 => x"e73f80d0",
  1607 => x"b4528151",
  1608 => x"dc933f80",
  1609 => x"0851a03f",
  1610 => x"7280d0f0",
  1611 => x"0cd6b03f",
  1612 => x"d5ce3f80",
  1613 => x"d0b45281",
  1614 => x"51dbfa3f",
  1615 => x"80085187",
  1616 => x"3f00ff39",
  1617 => x"00ff39f7",
  1618 => x"3d0d7b80",
  1619 => x"c0f00882",
  1620 => x"c811085a",
  1621 => x"545a7780",
  1622 => x"2e80da38",
  1623 => x"81881884",
  1624 => x"1908ff05",
  1625 => x"81712b59",
  1626 => x"55598074",
  1627 => x"2480ea38",
  1628 => x"807424b5",
  1629 => x"3873822b",
  1630 => x"78118805",
  1631 => x"56568180",
  1632 => x"19087706",
  1633 => x"5372802e",
  1634 => x"b6387816",
  1635 => x"70085353",
  1636 => x"79517408",
  1637 => x"53722dff",
  1638 => x"14fc17fc",
  1639 => x"1779812c",
  1640 => x"5a575754",
  1641 => x"738025d6",
  1642 => x"38770858",
  1643 => x"77ffad38",
  1644 => x"80c0f008",
  1645 => x"53bc1308",
  1646 => x"a5387951",
  1647 => x"ff833f74",
  1648 => x"0853722d",
  1649 => x"ff14fc17",
  1650 => x"fc177981",
  1651 => x"2c5a5757",
  1652 => x"54738025",
  1653 => x"ffa838d1",
  1654 => x"398057ff",
  1655 => x"93397251",
  1656 => x"bc130853",
  1657 => x"722d7951",
  1658 => x"fed73fff",
  1659 => x"3d0d80d0",
  1660 => x"bc0bfc05",
  1661 => x"70085252",
  1662 => x"70ff2e91",
  1663 => x"38702dfc",
  1664 => x"12700852",
  1665 => x"5270ff2e",
  1666 => x"098106f1",
  1667 => x"38833d0d",
  1668 => x"0404d5b8",
  1669 => x"3f040000",
  1670 => x"00000040",
  1671 => x"0a677265",
  1672 => x"74682072",
  1673 => x"65676973",
  1674 => x"74657273",
  1675 => x"3a000000",
  1676 => x"0a636f6e",
  1677 => x"74726f6c",
  1678 => x"3a202020",
  1679 => x"20202000",
  1680 => x"0a737461",
  1681 => x"7475733a",
  1682 => x"20202020",
  1683 => x"20202000",
  1684 => x"0a6d6163",
  1685 => x"5f6d7362",
  1686 => x"3a202020",
  1687 => x"20202000",
  1688 => x"0a6d6163",
  1689 => x"5f6c7362",
  1690 => x"3a202020",
  1691 => x"20202000",
  1692 => x"0a6d6469",
  1693 => x"6f5f636f",
  1694 => x"6e74726f",
  1695 => x"6c3a2000",
  1696 => x"0a74785f",
  1697 => x"706f696e",
  1698 => x"7465723a",
  1699 => x"20202000",
  1700 => x"0a72785f",
  1701 => x"706f696e",
  1702 => x"7465723a",
  1703 => x"20202000",
  1704 => x"0a656463",
  1705 => x"6c5f6970",
  1706 => x"3a202020",
  1707 => x"20202000",
  1708 => x"0a686173",
  1709 => x"685f6d73",
  1710 => x"623a2020",
  1711 => x"20202000",
  1712 => x"0a686173",
  1713 => x"685f6c73",
  1714 => x"623a2020",
  1715 => x"20202000",
  1716 => x"0a6d6469",
  1717 => x"6f207068",
  1718 => x"79207265",
  1719 => x"67697374",
  1720 => x"65727300",
  1721 => x"0a206d64",
  1722 => x"696f2070",
  1723 => x"68793a20",
  1724 => x"00000000",
  1725 => x"0a202072",
  1726 => x"65673a20",
  1727 => x"00000000",
  1728 => x"2d3e2000",
  1729 => x"67726574",
  1730 => x"682d3e63",
  1731 => x"6f6e7472",
  1732 => x"6f6c203a",
  1733 => x"00000000",
  1734 => x"67726574",
  1735 => x"682d3e73",
  1736 => x"74617475",
  1737 => x"7320203a",
  1738 => x"00000000",
  1739 => x"64657363",
  1740 => x"722d3e63",
  1741 => x"6f6e7472",
  1742 => x"6f6c203a",
  1743 => x"00000000",
  1744 => x"77726974",
  1745 => x"65206164",
  1746 => x"64726573",
  1747 => x"733a2000",
  1748 => x"20206c65",
  1749 => x"6e677468",
  1750 => x"3a200000",
  1751 => x"0a0a0000",
  1752 => x"72656164",
  1753 => x"20206164",
  1754 => x"64726573",
  1755 => x"733a2000",
  1756 => x"20206578",
  1757 => x"70656374",
  1758 => x"3a200000",
  1759 => x"2020676f",
  1760 => x"743a2000",
  1761 => x"20657272",
  1762 => x"6f720000",
  1763 => x"206f6b00",
  1764 => x"70686173",
  1765 => x"65207368",
  1766 => x"69667420",
  1767 => x"202d2020",
  1768 => x"76616c75",
  1769 => x"653a2000",
  1770 => x"20207374",
  1771 => x"61747573",
  1772 => x"3a200000",
  1773 => x"20202020",
  1774 => x"20000000",
  1775 => x"6f6b2020",
  1776 => x"00000000",
  1777 => x"4641494c",
  1778 => x"00000000",
  1779 => x"44445220",
  1780 => x"6d656d6f",
  1781 => x"72792069",
  1782 => x"6e666f00",
  1783 => x"0a0a6175",
  1784 => x"746f2074",
  1785 => x"5f524552",
  1786 => x"45534820",
  1787 => x"3a000000",
  1788 => x"0a636c6f",
  1789 => x"636b2065",
  1790 => x"6e61626c",
  1791 => x"6520203a",
  1792 => x"00000000",
  1793 => x"0a696e69",
  1794 => x"74616c69",
  1795 => x"7a652020",
  1796 => x"2020203a",
  1797 => x"00000000",
  1798 => x"0a636f6c",
  1799 => x"756d6e20",
  1800 => x"73697a65",
  1801 => x"2020203a",
  1802 => x"00000000",
  1803 => x"0a62616e",
  1804 => x"6b73697a",
  1805 => x"65202020",
  1806 => x"2020203a",
  1807 => x"00000000",
  1808 => x"4d627974",
  1809 => x"65000000",
  1810 => x"0a745f52",
  1811 => x"43442020",
  1812 => x"20202020",
  1813 => x"2020203a",
  1814 => x"00000000",
  1815 => x"0a745f52",
  1816 => x"46432020",
  1817 => x"20202020",
  1818 => x"2020203a",
  1819 => x"00000000",
  1820 => x"0a745f52",
  1821 => x"50202020",
  1822 => x"20202020",
  1823 => x"2020203a",
  1824 => x"00000000",
  1825 => x"0a726566",
  1826 => x"72657368",
  1827 => x"20656e2e",
  1828 => x"2020203a",
  1829 => x"00000000",
  1830 => x"0a0a4444",
  1831 => x"52206672",
  1832 => x"65717565",
  1833 => x"6e637920",
  1834 => x"3a000000",
  1835 => x"0a444452",
  1836 => x"20646174",
  1837 => x"61207769",
  1838 => x"6474683a",
  1839 => x"00000000",
  1840 => x"0a6d6f62",
  1841 => x"696c6520",
  1842 => x"73757070",
  1843 => x"6f72743a",
  1844 => x"00000000",
  1845 => x"0a0a7374",
  1846 => x"61747573",
  1847 => x"20726561",
  1848 => x"64202020",
  1849 => x"3a000000",
  1850 => x"0a0a7365",
  1851 => x"6c662072",
  1852 => x"65667265",
  1853 => x"73682020",
  1854 => x"3a000000",
  1855 => x"20353132",
  1856 => x"00000000",
  1857 => x"34303639",
  1858 => x"00000000",
  1859 => x"312f3800",
  1860 => x"20617272",
  1861 => x"61790000",
  1862 => x"0a74656d",
  1863 => x"702d636f",
  1864 => x"6d702072",
  1865 => x"6566723a",
  1866 => x"00000000",
  1867 => x"c2b04300",
  1868 => x"0a647269",
  1869 => x"76652073",
  1870 => x"7472656e",
  1871 => x"6774683a",
  1872 => x"00000000",
  1873 => x"0a706f77",
  1874 => x"65722073",
  1875 => x"6176696e",
  1876 => x"6720203a",
  1877 => x"00000000",
  1878 => x"756e6b6e",
  1879 => x"6f776e00",
  1880 => x"0a745f58",
  1881 => x"50202020",
  1882 => x"20202020",
  1883 => x"2020203a",
  1884 => x"00000000",
  1885 => x"0a745f58",
  1886 => x"53522020",
  1887 => x"20202020",
  1888 => x"2020203a",
  1889 => x"00000000",
  1890 => x"0a745f43",
  1891 => x"4b452020",
  1892 => x"20202020",
  1893 => x"2020203a",
  1894 => x"00000000",
  1895 => x"0a434153",
  1896 => x"206c6174",
  1897 => x"656e6379",
  1898 => x"2020203a",
  1899 => x"00000000",
  1900 => x"0a6d6f62",
  1901 => x"696c6520",
  1902 => x"656e6162",
  1903 => x"6c65643a",
  1904 => x"00000000",
  1905 => x"0a0a7068",
  1906 => x"7920636f",
  1907 => x"6e666967",
  1908 => x"20302020",
  1909 => x"3a000000",
  1910 => x"0a0a7068",
  1911 => x"7920636f",
  1912 => x"6e666967",
  1913 => x"20312020",
  1914 => x"3a000000",
  1915 => x"31303234",
  1916 => x"00000000",
  1917 => x"32303438",
  1918 => x"00000000",
  1919 => x"66756c6c",
  1920 => x"00000000",
  1921 => x"37300000",
  1922 => x"64656570",
  1923 => x"20706f77",
  1924 => x"65722064",
  1925 => x"6f776e00",
  1926 => x"636c6f63",
  1927 => x"6b207374",
  1928 => x"6f700000",
  1929 => x"73656c66",
  1930 => x"20726566",
  1931 => x"72657368",
  1932 => x"00000000",
  1933 => x"706f7765",
  1934 => x"7220646f",
  1935 => x"776e0000",
  1936 => x"6e6f6e65",
  1937 => x"00000000",
  1938 => x"312f3200",
  1939 => x"312f3400",
  1940 => x"312f3100",
  1941 => x"332f3400",
  1942 => x"38350000",
  1943 => x"34350000",
  1944 => x"68616c66",
  1945 => x"00000000",
  1946 => x"31350000",
  1947 => x"61646472",
  1948 => x"6573733a",
  1949 => x"20000000",
  1950 => x"20646174",
  1951 => x"613a2000",
  1952 => x"0a0a4443",
  1953 => x"4d207068",
  1954 => x"61736520",
  1955 => x"73686966",
  1956 => x"74207465",
  1957 => x"7374696e",
  1958 => x"67000000",
  1959 => x"0a696e69",
  1960 => x"7469616c",
  1961 => x"3a200000",
  1962 => x"09000000",
  1963 => x"20202020",
  1964 => x"00000000",
  1965 => x"6c6f7720",
  1966 => x"666f756e",
  1967 => x"64000000",
  1968 => x"68696768",
  1969 => x"20666f75",
  1970 => x"6e640000",
  1971 => x"0a6c6f77",
  1972 => x"3a202020",
  1973 => x"20202020",
  1974 => x"20200000",
  1975 => x"0a686967",
  1976 => x"683a2020",
  1977 => x"20202020",
  1978 => x"20200000",
  1979 => x"0a646966",
  1980 => x"663a2020",
  1981 => x"20202020",
  1982 => x"20200000",
  1983 => x"0a6d696e",
  1984 => x"5f657272",
  1985 => x"3a202020",
  1986 => x"20200000",
  1987 => x"0a6d696e",
  1988 => x"5f657272",
  1989 => x"5f706f73",
  1990 => x"3a200000",
  1991 => x"676f206d",
  1992 => x"696e5f65",
  1993 => x"72726f72",
  1994 => x"00000000",
  1995 => x"0a66696e",
  1996 => x"616c3a20",
  1997 => x"20202020",
  1998 => x"20200000",
  1999 => x"6c6f7720",
  2000 => x"4e4f5420",
  2001 => x"666f756e",
  2002 => x"64000000",
  2003 => x"68696768",
  2004 => x"204e4f54",
  2005 => x"20666f75",
  2006 => x"6e640000",
  2007 => x"676f207a",
  2008 => x"65726f00",
  2009 => x"64617461",
  2010 => x"2076616c",
  2011 => x"69640000",
  2012 => x"6c6f7720",
  2013 => x"20666f75",
  2014 => x"6e640000",
  2015 => x"0a646966",
  2016 => x"662f323a",
  2017 => x"20202020",
  2018 => x"20200000",
  2019 => x"6c6f7720",
  2020 => x"204e4f54",
  2021 => x"20666f75",
  2022 => x"6e640000",
  2023 => x"64617461",
  2024 => x"204e4f54",
  2025 => x"2076616c",
  2026 => x"69640000",
  2027 => x"74657374",
  2028 => x"2e632000",
  2029 => x"286f6e20",
  2030 => x"73696d29",
  2031 => x"0a000000",
  2032 => x"286f6e20",
  2033 => x"68617264",
  2034 => x"77617265",
  2035 => x"290a0000",
  2036 => x"636f6d70",
  2037 => x"696c6564",
  2038 => x"3a204e6f",
  2039 => x"76203236",
  2040 => x"20323031",
  2041 => x"30202031",
  2042 => x"353a3237",
  2043 => x"3a33350a",
  2044 => x"00000000",
  2045 => x"30622020",
  2046 => x"20202020",
  2047 => x"20202020",
  2048 => x"20202020",
  2049 => x"20202020",
  2050 => x"20202020",
  2051 => x"20202020",
  2052 => x"20202020",
  2053 => x"20200000",
  2054 => x"30782020",
  2055 => x"20202020",
  2056 => x"20200000",
  2057 => x"43000000",
  2058 => x"64756d6d",
  2059 => x"792e6578",
  2060 => x"65000000",
  2061 => x"00ffffff",
  2062 => x"ff00ffff",
  2063 => x"ffff00ff",
  2064 => x"ffffff00",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00002844",
  2069 => x"fff00000",
  2070 => x"80000d00",
  2071 => x"80000c00",
  2072 => x"80000800",
  2073 => x"80000600",
  2074 => x"80000200",
  2075 => x"80000100",
  2076 => x"00002074",
  2077 => x"00000000",
  2078 => x"000022dc",
  2079 => x"00002338",
  2080 => x"00002394",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00002024",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000001",
  2120 => x"330eabcd",
  2121 => x"1234e66d",
  2122 => x"deec0005",
  2123 => x"000b0000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00000000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"00000000",
  2242 => x"00000000",
  2243 => x"00000000",
  2244 => x"00000000",
  2245 => x"00000000",
  2246 => x"00000000",
  2247 => x"00000000",
  2248 => x"00000000",
  2249 => x"00000000",
  2250 => x"00000000",
  2251 => x"00000000",
  2252 => x"00000000",
  2253 => x"00000000",
  2254 => x"00000000",
  2255 => x"00000000",
  2256 => x"00000000",
  2257 => x"00000000",
  2258 => x"00000000",
  2259 => x"00000000",
  2260 => x"00000000",
  2261 => x"00000000",
  2262 => x"00000000",
  2263 => x"00000000",
  2264 => x"00000000",
  2265 => x"00000000",
  2266 => x"00000000",
  2267 => x"00000000",
  2268 => x"00000000",
  2269 => x"00000000",
  2270 => x"00000000",
  2271 => x"00000000",
  2272 => x"00000000",
  2273 => x"00000000",
  2274 => x"00000000",
  2275 => x"00000000",
  2276 => x"00000000",
  2277 => x"00000000",
  2278 => x"00000000",
  2279 => x"00000000",
  2280 => x"00000000",
  2281 => x"00000000",
  2282 => x"00000000",
  2283 => x"00000000",
  2284 => x"00000000",
  2285 => x"00000000",
  2286 => x"00000000",
  2287 => x"00000000",
  2288 => x"00000000",
  2289 => x"00000000",
  2290 => x"00000000",
  2291 => x"00000000",
  2292 => x"00000000",
  2293 => x"00000000",
  2294 => x"00000000",
  2295 => x"00000000",
  2296 => x"00000000",
  2297 => x"00000000",
  2298 => x"00000000",
  2299 => x"00000000",
  2300 => x"00000000",
  2301 => x"00000000",
  2302 => x"00000000",
  2303 => x"00000000",
  2304 => x"00000000",
  2305 => x"00000000",
  2306 => x"00000000",
  2307 => x"00000000",
  2308 => x"00000000",
  2309 => x"00000000",
  2310 => x"00000000",
  2311 => x"00000000",
  2312 => x"ffffffff",
  2313 => x"00000000",
  2314 => x"00020000",
  2315 => x"00000000",
  2316 => x"00000000",
  2317 => x"0000242c",
  2318 => x"0000242c",
  2319 => x"00002434",
  2320 => x"00002434",
  2321 => x"0000243c",
  2322 => x"0000243c",
  2323 => x"00002444",
  2324 => x"00002444",
  2325 => x"0000244c",
  2326 => x"0000244c",
  2327 => x"00002454",
  2328 => x"00002454",
  2329 => x"0000245c",
  2330 => x"0000245c",
  2331 => x"00002464",
  2332 => x"00002464",
  2333 => x"0000246c",
  2334 => x"0000246c",
  2335 => x"00002474",
  2336 => x"00002474",
  2337 => x"0000247c",
  2338 => x"0000247c",
  2339 => x"00002484",
  2340 => x"00002484",
  2341 => x"0000248c",
  2342 => x"0000248c",
  2343 => x"00002494",
  2344 => x"00002494",
  2345 => x"0000249c",
  2346 => x"0000249c",
  2347 => x"000024a4",
  2348 => x"000024a4",
  2349 => x"000024ac",
  2350 => x"000024ac",
  2351 => x"000024b4",
  2352 => x"000024b4",
  2353 => x"000024bc",
  2354 => x"000024bc",
  2355 => x"000024c4",
  2356 => x"000024c4",
  2357 => x"000024cc",
  2358 => x"000024cc",
  2359 => x"000024d4",
  2360 => x"000024d4",
  2361 => x"000024dc",
  2362 => x"000024dc",
  2363 => x"000024e4",
  2364 => x"000024e4",
  2365 => x"000024ec",
  2366 => x"000024ec",
  2367 => x"000024f4",
  2368 => x"000024f4",
  2369 => x"000024fc",
  2370 => x"000024fc",
  2371 => x"00002504",
  2372 => x"00002504",
  2373 => x"0000250c",
  2374 => x"0000250c",
  2375 => x"00002514",
  2376 => x"00002514",
  2377 => x"0000251c",
  2378 => x"0000251c",
  2379 => x"00002524",
  2380 => x"00002524",
  2381 => x"0000252c",
  2382 => x"0000252c",
  2383 => x"00002534",
  2384 => x"00002534",
  2385 => x"0000253c",
  2386 => x"0000253c",
  2387 => x"00002544",
  2388 => x"00002544",
  2389 => x"0000254c",
  2390 => x"0000254c",
  2391 => x"00002554",
  2392 => x"00002554",
  2393 => x"0000255c",
  2394 => x"0000255c",
  2395 => x"00002564",
  2396 => x"00002564",
  2397 => x"0000256c",
  2398 => x"0000256c",
  2399 => x"00002574",
  2400 => x"00002574",
  2401 => x"0000257c",
  2402 => x"0000257c",
  2403 => x"00002584",
  2404 => x"00002584",
  2405 => x"0000258c",
  2406 => x"0000258c",
  2407 => x"00002594",
  2408 => x"00002594",
  2409 => x"0000259c",
  2410 => x"0000259c",
  2411 => x"000025a4",
  2412 => x"000025a4",
  2413 => x"000025ac",
  2414 => x"000025ac",
  2415 => x"000025b4",
  2416 => x"000025b4",
  2417 => x"000025bc",
  2418 => x"000025bc",
  2419 => x"000025c4",
  2420 => x"000025c4",
  2421 => x"000025cc",
  2422 => x"000025cc",
  2423 => x"000025d4",
  2424 => x"000025d4",
  2425 => x"000025dc",
  2426 => x"000025dc",
  2427 => x"000025e4",
  2428 => x"000025e4",
  2429 => x"000025ec",
  2430 => x"000025ec",
  2431 => x"000025f4",
  2432 => x"000025f4",
  2433 => x"000025fc",
  2434 => x"000025fc",
  2435 => x"00002604",
  2436 => x"00002604",
  2437 => x"0000260c",
  2438 => x"0000260c",
  2439 => x"00002614",
  2440 => x"00002614",
  2441 => x"0000261c",
  2442 => x"0000261c",
  2443 => x"00002624",
  2444 => x"00002624",
  2445 => x"0000262c",
  2446 => x"0000262c",
  2447 => x"00002634",
  2448 => x"00002634",
  2449 => x"0000263c",
  2450 => x"0000263c",
  2451 => x"00002644",
  2452 => x"00002644",
  2453 => x"0000264c",
  2454 => x"0000264c",
  2455 => x"00002654",
  2456 => x"00002654",
  2457 => x"0000265c",
  2458 => x"0000265c",
  2459 => x"00002664",
  2460 => x"00002664",
  2461 => x"0000266c",
  2462 => x"0000266c",
  2463 => x"00002674",
  2464 => x"00002674",
  2465 => x"0000267c",
  2466 => x"0000267c",
  2467 => x"00002684",
  2468 => x"00002684",
  2469 => x"0000268c",
  2470 => x"0000268c",
  2471 => x"00002694",
  2472 => x"00002694",
  2473 => x"0000269c",
  2474 => x"0000269c",
  2475 => x"000026a4",
  2476 => x"000026a4",
  2477 => x"000026ac",
  2478 => x"000026ac",
  2479 => x"000026b4",
  2480 => x"000026b4",
  2481 => x"000026bc",
  2482 => x"000026bc",
  2483 => x"000026c4",
  2484 => x"000026c4",
  2485 => x"000026cc",
  2486 => x"000026cc",
  2487 => x"000026d4",
  2488 => x"000026d4",
  2489 => x"000026dc",
  2490 => x"000026dc",
  2491 => x"000026e4",
  2492 => x"000026e4",
  2493 => x"000026ec",
  2494 => x"000026ec",
  2495 => x"000026f4",
  2496 => x"000026f4",
  2497 => x"000026fc",
  2498 => x"000026fc",
  2499 => x"00002704",
  2500 => x"00002704",
  2501 => x"0000270c",
  2502 => x"0000270c",
  2503 => x"00002714",
  2504 => x"00002714",
  2505 => x"0000271c",
  2506 => x"0000271c",
  2507 => x"00002724",
  2508 => x"00002724",
  2509 => x"0000272c",
  2510 => x"0000272c",
  2511 => x"00002734",
  2512 => x"00002734",
  2513 => x"0000273c",
  2514 => x"0000273c",
  2515 => x"00002744",
  2516 => x"00002744",
  2517 => x"0000274c",
  2518 => x"0000274c",
  2519 => x"00002754",
  2520 => x"00002754",
  2521 => x"0000275c",
  2522 => x"0000275c",
  2523 => x"00002764",
  2524 => x"00002764",
  2525 => x"0000276c",
  2526 => x"0000276c",
  2527 => x"00002774",
  2528 => x"00002774",
  2529 => x"0000277c",
  2530 => x"0000277c",
  2531 => x"00002784",
  2532 => x"00002784",
  2533 => x"0000278c",
  2534 => x"0000278c",
  2535 => x"00002794",
  2536 => x"00002794",
  2537 => x"0000279c",
  2538 => x"0000279c",
  2539 => x"000027a4",
  2540 => x"000027a4",
  2541 => x"000027ac",
  2542 => x"000027ac",
  2543 => x"000027b4",
  2544 => x"000027b4",
  2545 => x"000027bc",
  2546 => x"000027bc",
  2547 => x"000027c4",
  2548 => x"000027c4",
  2549 => x"000027cc",
  2550 => x"000027cc",
  2551 => x"000027d4",
  2552 => x"000027d4",
  2553 => x"000027dc",
  2554 => x"000027dc",
  2555 => x"000027e4",
  2556 => x"000027e4",
  2557 => x"000027ec",
  2558 => x"000027ec",
  2559 => x"000027f4",
  2560 => x"000027f4",
  2561 => x"000027fc",
  2562 => x"000027fc",
  2563 => x"00002804",
  2564 => x"00002804",
  2565 => x"0000280c",
  2566 => x"0000280c",
  2567 => x"00002814",
  2568 => x"00002814",
  2569 => x"0000281c",
  2570 => x"0000281c",
  2571 => x"00002824",
  2572 => x"00002824",
  2573 => x"00002028",
  2574 => x"ffffffff",
  2575 => x"00000000",
  2576 => x"ffffffff",
  2577 => x"00000000",
  2578 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
