
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 15;
constant bytes : integer := 28244;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B80F3";
    when 16#00001# => romdata <= X"EA040000";
    when 16#00002# => romdata <= X"00000000";
    when 16#00003# => romdata <= X"00000000";
    when 16#00004# => romdata <= X"00000000";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"0B0B80F6";
    when 16#00009# => romdata <= X"D1040000";
    when 16#0000A# => romdata <= X"00000000";
    when 16#0000B# => romdata <= X"00000000";
    when 16#0000C# => romdata <= X"00000000";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B80F6";
    when 16#00049# => romdata <= X"83040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B80F5E6";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B81CC";
    when 16#000A2# => romdata <= X"D8738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B80";
    when 16#000A5# => romdata <= X"F5E90400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"0B0B80F6";
    when 16#000A9# => romdata <= X"B8040000";
    when 16#000AA# => romdata <= X"00000000";
    when 16#000AB# => romdata <= X"00000000";
    when 16#000AC# => romdata <= X"00000000";
    when 16#000AD# => romdata <= X"00000000";
    when 16#000AE# => romdata <= X"00000000";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"0B0B80F6";
    when 16#000B1# => romdata <= X"9F040000";
    when 16#000B2# => romdata <= X"00000000";
    when 16#000B3# => romdata <= X"00000000";
    when 16#000B4# => romdata <= X"00000000";
    when 16#000B5# => romdata <= X"00000000";
    when 16#000B6# => romdata <= X"00000000";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"81CCE80C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"FF3D0D02";
    when 16#00101# => romdata <= X"8F053370";
    when 16#00102# => romdata <= X"525280F3";
    when 16#00103# => romdata <= X"AC3F7151";
    when 16#00104# => romdata <= X"80F3F63F";
    when 16#00105# => romdata <= X"71B00C83";
    when 16#00106# => romdata <= X"3D0D04FF";
    when 16#00107# => romdata <= X"3D0D81CC";
    when 16#00108# => romdata <= X"C408B811";
    when 16#00109# => romdata <= X"08535180";
    when 16#0010A# => romdata <= X"0BB8120C";
    when 16#0010B# => romdata <= X"71B00C83";
    when 16#0010C# => romdata <= X"3D0D0480";
    when 16#0010D# => romdata <= X"0B81EFF8";
    when 16#0010E# => romdata <= X"34800BB0";
    when 16#0010F# => romdata <= X"0C04FB3D";
    when 16#00110# => romdata <= X"0D815180";
    when 16#00111# => romdata <= X"C7DD3FB0";
    when 16#00112# => romdata <= X"08538251";
    when 16#00113# => romdata <= X"80C7D43F";
    when 16#00114# => romdata <= X"B00856B0";
    when 16#00115# => romdata <= X"08833890";
    when 16#00116# => romdata <= X"5672FC06";
    when 16#00117# => romdata <= X"5575812E";
    when 16#00118# => romdata <= X"80FB3880";
    when 16#00119# => romdata <= X"54737627";
    when 16#0011A# => romdata <= X"AD387383";
    when 16#0011B# => romdata <= X"06537280";
    when 16#0011C# => romdata <= X"2EB23881";
    when 16#0011D# => romdata <= X"C0C85180";
    when 16#0011E# => romdata <= X"EE983F74";
    when 16#0011F# => romdata <= X"70840556";
    when 16#00120# => romdata <= X"0852A051";
    when 16#00121# => romdata <= X"80EEAE3F";
    when 16#00122# => romdata <= X"A05180ED";
    when 16#00123# => romdata <= X"EB3F8114";
    when 16#00124# => romdata <= X"54757426";
    when 16#00125# => romdata <= X"D5388A51";
    when 16#00126# => romdata <= X"80EDDD3F";
    when 16#00127# => romdata <= X"800BB00C";
    when 16#00128# => romdata <= X"873D0D04";
    when 16#00129# => romdata <= X"81A5B051";
    when 16#0012A# => romdata <= X"80EDE73F";
    when 16#0012B# => romdata <= X"7452A051";
    when 16#0012C# => romdata <= X"80EE823F";
    when 16#0012D# => romdata <= X"81B29C51";
    when 16#0012E# => romdata <= X"80EDD73F";
    when 16#0012F# => romdata <= X"81C0C851";
    when 16#00130# => romdata <= X"80EDCF3F";
    when 16#00131# => romdata <= X"74708405";
    when 16#00132# => romdata <= X"560852A0";
    when 16#00133# => romdata <= X"5180EDE5";
    when 16#00134# => romdata <= X"3FA05180";
    when 16#00135# => romdata <= X"EDA23F81";
    when 16#00136# => romdata <= X"1454FFB5";
    when 16#00137# => romdata <= X"3981C0C8";
    when 16#00138# => romdata <= X"5180EDAE";
    when 16#00139# => romdata <= X"3F740852";
    when 16#0013A# => romdata <= X"A05180ED";
    when 16#0013B# => romdata <= X"C83F8A51";
    when 16#0013C# => romdata <= X"80ED853F";
    when 16#0013D# => romdata <= X"800BB00C";
    when 16#0013E# => romdata <= X"873D0D04";
    when 16#0013F# => romdata <= X"FC3D0D81";
    when 16#00140# => romdata <= X"5180C69F";
    when 16#00141# => romdata <= X"3FB00852";
    when 16#00142# => romdata <= X"825180C4";
    when 16#00143# => romdata <= X"E43FB008";
    when 16#00144# => romdata <= X"81FF0672";
    when 16#00145# => romdata <= X"56538354";
    when 16#00146# => romdata <= X"72802EA2";
    when 16#00147# => romdata <= X"38735180";
    when 16#00148# => romdata <= X"C6813F81";
    when 16#00149# => romdata <= X"147081FF";
    when 16#0014A# => romdata <= X"06FF1570";
    when 16#0014B# => romdata <= X"81FF06B0";
    when 16#0014C# => romdata <= X"08797084";
    when 16#0014D# => romdata <= X"055B0C56";
    when 16#0014E# => romdata <= X"52555272";
    when 16#0014F# => romdata <= X"E03872B0";
    when 16#00150# => romdata <= X"0C863D0D";
    when 16#00151# => romdata <= X"04803D0D";
    when 16#00152# => romdata <= X"8C5180EC";
    when 16#00153# => romdata <= X"AB3F800B";
    when 16#00154# => romdata <= X"B00C823D";
    when 16#00155# => romdata <= X"0D04FB3D";
    when 16#00156# => romdata <= X"0D800B81";
    when 16#00157# => romdata <= X"A5B45256";
    when 16#00158# => romdata <= X"80ECAF3F";
    when 16#00159# => romdata <= X"75557410";
    when 16#0015A# => romdata <= X"81FE0653";
    when 16#0015B# => romdata <= X"81D05281";
    when 16#0015C# => romdata <= X"CCF00851";
    when 16#0015D# => romdata <= X"80D2D13F";
    when 16#0015E# => romdata <= X"B008982B";
    when 16#0015F# => romdata <= X"54807424";
    when 16#00160# => romdata <= X"A23881A5";
    when 16#00161# => romdata <= X"C05180EC";
    when 16#00162# => romdata <= X"893F7452";
    when 16#00163# => romdata <= X"885180EC";
    when 16#00164# => romdata <= X"A43F81A5";
    when 16#00165# => romdata <= X"CC5180EB";
    when 16#00166# => romdata <= X"F93F8116";
    when 16#00167# => romdata <= X"7083FFFF";
    when 16#00168# => romdata <= X"06575481";
    when 16#00169# => romdata <= X"157081FF";
    when 16#0016A# => romdata <= X"0670982B";
    when 16#0016B# => romdata <= X"52565473";
    when 16#0016C# => romdata <= X"8025FFB2";
    when 16#0016D# => romdata <= X"3875B00C";
    when 16#0016E# => romdata <= X"873D0D04";
    when 16#0016F# => romdata <= X"F33D0D7F";
    when 16#00170# => romdata <= X"02840580";
    when 16#00171# => romdata <= X"C3053302";
    when 16#00172# => romdata <= X"880580C6";
    when 16#00173# => romdata <= X"052281A5";
    when 16#00174# => romdata <= X"DC545B55";
    when 16#00175# => romdata <= X"5880EBBA";
    when 16#00176# => romdata <= X"3F785180";
    when 16#00177# => romdata <= X"ECFE3F81";
    when 16#00178# => romdata <= X"A5E85180";
    when 16#00179# => romdata <= X"EBAC3F73";
    when 16#0017A# => romdata <= X"52885180";
    when 16#0017B# => romdata <= X"EBC73F81";
    when 16#0017C# => romdata <= X"A6845180";
    when 16#0017D# => romdata <= X"EB9C3F80";
    when 16#0017E# => romdata <= X"57767927";
    when 16#0017F# => romdata <= X"81A13873";
    when 16#00180# => romdata <= X"108E3D5D";
    when 16#00181# => romdata <= X"5A7981FF";
    when 16#00182# => romdata <= X"06538190";
    when 16#00183# => romdata <= X"52775180";
    when 16#00184# => romdata <= X"D1B63F76";
    when 16#00185# => romdata <= X"882A5390";
    when 16#00186# => romdata <= X"52775180";
    when 16#00187# => romdata <= X"D1AA3F76";
    when 16#00188# => romdata <= X"81FF0653";
    when 16#00189# => romdata <= X"90527751";
    when 16#0018A# => romdata <= X"80D19D3F";
    when 16#0018B# => romdata <= X"811A7081";
    when 16#0018C# => romdata <= X"FF065455";
    when 16#0018D# => romdata <= X"81905277";
    when 16#0018E# => romdata <= X"5180D18C";
    when 16#0018F# => romdata <= X"3F805380";
    when 16#00190# => romdata <= X"E0527751";
    when 16#00191# => romdata <= X"80D1813F";
    when 16#00192# => romdata <= X"B008982B";
    when 16#00193# => romdata <= X"54807424";
    when 16#00194# => romdata <= X"8A388818";
    when 16#00195# => romdata <= X"087081FF";
    when 16#00196# => romdata <= X"065C567A";
    when 16#00197# => romdata <= X"81FF0681";
    when 16#00198# => romdata <= X"C0C85256";
    when 16#00199# => romdata <= X"80EAAB3F";
    when 16#0019A# => romdata <= X"75528851";
    when 16#0019B# => romdata <= X"80EAC63F";
    when 16#0019C# => romdata <= X"81AFF851";
    when 16#0019D# => romdata <= X"80EA9B3F";
    when 16#0019E# => romdata <= X"E0165480";
    when 16#0019F# => romdata <= X"DF7427B6";
    when 16#001A0# => romdata <= X"38768706";
    when 16#001A1# => romdata <= X"701D5755";
    when 16#001A2# => romdata <= X"A0763474";
    when 16#001A3# => romdata <= X"872EB938";
    when 16#001A4# => romdata <= X"81177083";
    when 16#001A5# => romdata <= X"FFFF0658";
    when 16#001A6# => romdata <= X"55787726";
    when 16#001A7# => romdata <= X"FEE73880";
    when 16#001A8# => romdata <= X"E00B8C19";
    when 16#001A9# => romdata <= X"0C8C1808";
    when 16#001AA# => romdata <= X"70812A81";
    when 16#001AB# => romdata <= X"06585A76";
    when 16#001AC# => romdata <= X"F4388F3D";
    when 16#001AD# => romdata <= X"0D047687";
    when 16#001AE# => romdata <= X"06701D55";
    when 16#001AF# => romdata <= X"55757434";
    when 16#001B0# => romdata <= X"74872E09";
    when 16#001B1# => romdata <= X"8106C938";
    when 16#001B2# => romdata <= X"7B5180E9";
    when 16#001B3# => romdata <= X"C53F8A51";
    when 16#001B4# => romdata <= X"80E9A53F";
    when 16#001B5# => romdata <= X"81177083";
    when 16#001B6# => romdata <= X"FFFF0658";
    when 16#001B7# => romdata <= X"55787726";
    when 16#001B8# => romdata <= X"FEA338FF";
    when 16#001B9# => romdata <= X"BA39FB3D";
    when 16#001BA# => romdata <= X"0D815180";
    when 16#001BB# => romdata <= X"C1833FB0";
    when 16#001BC# => romdata <= X"0881FF06";
    when 16#001BD# => romdata <= X"54825180";
    when 16#001BE# => romdata <= X"C2A93FB0";
    when 16#001BF# => romdata <= X"0881FF06";
    when 16#001C0# => romdata <= X"56835180";
    when 16#001C1# => romdata <= X"C0EB3FB0";
    when 16#001C2# => romdata <= X"0883FFFF";
    when 16#001C3# => romdata <= X"0655739C";
    when 16#001C4# => romdata <= X"3881CCF0";
    when 16#001C5# => romdata <= X"08547484";
    when 16#001C6# => romdata <= X"38818055";
    when 16#001C7# => romdata <= X"74537552";
    when 16#001C8# => romdata <= X"7351FD98";
    when 16#001C9# => romdata <= X"3F74B00C";
    when 16#001CA# => romdata <= X"873D0D04";
    when 16#001CB# => romdata <= X"81CCF408";
    when 16#001CC# => romdata <= X"54E439F8";
    when 16#001CD# => romdata <= X"3D0D02AA";
    when 16#001CE# => romdata <= X"052281CC";
    when 16#001CF# => romdata <= X"CC3381F7";
    when 16#001D0# => romdata <= X"06585876";
    when 16#001D1# => romdata <= X"81CCCC34";
    when 16#001D2# => romdata <= X"81CCF008";
    when 16#001D3# => romdata <= X"5580C053";
    when 16#001D4# => romdata <= X"81905274";
    when 16#001D5# => romdata <= X"5180CEF0";
    when 16#001D6# => romdata <= X"3F745180";
    when 16#001D7# => romdata <= X"CF9C3FB0";
    when 16#001D8# => romdata <= X"0881FF06";
    when 16#001D9# => romdata <= X"5473802E";
    when 16#001DA# => romdata <= X"84903876";
    when 16#001DB# => romdata <= X"5380D052";
    when 16#001DC# => romdata <= X"745180CE";
    when 16#001DD# => romdata <= X"D33F8059";
    when 16#001DE# => romdata <= X"8F5781CC";
    when 16#001DF# => romdata <= X"CC3381FE";
    when 16#001E0# => romdata <= X"06547381";
    when 16#001E1# => romdata <= X"CCCC3481";
    when 16#001E2# => romdata <= X"CCF00874";
    when 16#001E3# => romdata <= X"575580C0";
    when 16#001E4# => romdata <= X"53819052";
    when 16#001E5# => romdata <= X"745180CE";
    when 16#001E6# => romdata <= X"AF3F7451";
    when 16#001E7# => romdata <= X"80CEDB3F";
    when 16#001E8# => romdata <= X"B00881FF";
    when 16#001E9# => romdata <= X"06547380";
    when 16#001EA# => romdata <= X"2E83C438";
    when 16#001EB# => romdata <= X"755380D0";
    when 16#001EC# => romdata <= X"52745180";
    when 16#001ED# => romdata <= X"CE923F77";
    when 16#001EE# => romdata <= X"772C8106";
    when 16#001EF# => romdata <= X"5574802E";
    when 16#001F0# => romdata <= X"83A23881";
    when 16#001F1# => romdata <= X"CCCC3382";
    when 16#001F2# => romdata <= X"07547381";
    when 16#001F3# => romdata <= X"CCCC3481";
    when 16#001F4# => romdata <= X"CCF00874";
    when 16#001F5# => romdata <= X"575580C0";
    when 16#001F6# => romdata <= X"53819052";
    when 16#001F7# => romdata <= X"745180CD";
    when 16#001F8# => romdata <= X"E73F7451";
    when 16#001F9# => romdata <= X"80CE933F";
    when 16#001FA# => romdata <= X"B00881FF";
    when 16#001FB# => romdata <= X"06547380";
    when 16#001FC# => romdata <= X"2E82E638";
    when 16#001FD# => romdata <= X"755380D0";
    when 16#001FE# => romdata <= X"52745180";
    when 16#001FF# => romdata <= X"CDCA3F81";
    when 16#00200# => romdata <= X"CCF00855";
    when 16#00201# => romdata <= X"80C15381";
    when 16#00202# => romdata <= X"90527451";
    when 16#00203# => romdata <= X"80CDB93F";
    when 16#00204# => romdata <= X"745180CD";
    when 16#00205# => romdata <= X"E53FB008";
    when 16#00206# => romdata <= X"81FF0656";
    when 16#00207# => romdata <= X"75802E82";
    when 16#00208# => romdata <= X"8C388053";
    when 16#00209# => romdata <= X"80E05274";
    when 16#0020A# => romdata <= X"5180CD9C";
    when 16#0020B# => romdata <= X"3F745180";
    when 16#0020C# => romdata <= X"CDC83FB0";
    when 16#0020D# => romdata <= X"0881FF06";
    when 16#0020E# => romdata <= X"5473802E";
    when 16#0020F# => romdata <= X"81EF3888";
    when 16#00210# => romdata <= X"15087090";
    when 16#00211# => romdata <= X"2B70902C";
    when 16#00212# => romdata <= X"56565673";
    when 16#00213# => romdata <= X"822A8106";
    when 16#00214# => romdata <= X"5473802E";
    when 16#00215# => romdata <= X"8D388177";
    when 16#00216# => romdata <= X"2B790770";
    when 16#00217# => romdata <= X"83FFFF06";
    when 16#00218# => romdata <= X"5A5681CC";
    when 16#00219# => romdata <= X"CC338107";
    when 16#0021A# => romdata <= X"547381CC";
    when 16#0021B# => romdata <= X"CC3481CC";
    when 16#0021C# => romdata <= X"F0087457";
    when 16#0021D# => romdata <= X"5580C053";
    when 16#0021E# => romdata <= X"81905274";
    when 16#0021F# => romdata <= X"5180CCC8";
    when 16#00220# => romdata <= X"3F745180";
    when 16#00221# => romdata <= X"CCF43FB0";
    when 16#00222# => romdata <= X"0881FF06";
    when 16#00223# => romdata <= X"5473802E";
    when 16#00224# => romdata <= X"81A83875";
    when 16#00225# => romdata <= X"5380D052";
    when 16#00226# => romdata <= X"745180CC";
    when 16#00227# => romdata <= X"AB3F7681";
    when 16#00228# => romdata <= X"800A2981";
    when 16#00229# => romdata <= X"FF0A0570";
    when 16#0022A# => romdata <= X"982C5856";
    when 16#0022B# => romdata <= X"768025FD";
    when 16#0022C# => romdata <= X"C93881CC";
    when 16#0022D# => romdata <= X"CC338207";
    when 16#0022E# => romdata <= X"577681CC";
    when 16#0022F# => romdata <= X"CC3481CC";
    when 16#00230# => romdata <= X"F0085580";
    when 16#00231# => romdata <= X"C0538190";
    when 16#00232# => romdata <= X"52745180";
    when 16#00233# => romdata <= X"CBFA3F74";
    when 16#00234# => romdata <= X"5180CCA6";
    when 16#00235# => romdata <= X"3FB00881";
    when 16#00236# => romdata <= X"FF065877";
    when 16#00237# => romdata <= X"802E81B8";
    when 16#00238# => romdata <= X"38765380";
    when 16#00239# => romdata <= X"D0527451";
    when 16#0023A# => romdata <= X"80CBDD3F";
    when 16#0023B# => romdata <= X"81CCCC33";
    when 16#0023C# => romdata <= X"88075776";
    when 16#0023D# => romdata <= X"81CCCC34";
    when 16#0023E# => romdata <= X"81CCF008";
    when 16#0023F# => romdata <= X"5580C053";
    when 16#00240# => romdata <= X"81905274";
    when 16#00241# => romdata <= X"5180CBC0";
    when 16#00242# => romdata <= X"3F745180";
    when 16#00243# => romdata <= X"CBEC3FB0";
    when 16#00244# => romdata <= X"0881FF06";
    when 16#00245# => romdata <= X"5877802E";
    when 16#00246# => romdata <= X"80EF3876";
    when 16#00247# => romdata <= X"5380D052";
    when 16#00248# => romdata <= X"745180CB";
    when 16#00249# => romdata <= X"A33F78B0";
    when 16#0024A# => romdata <= X"0C8A3D0D";
    when 16#0024B# => romdata <= X"0481A688";
    when 16#0024C# => romdata <= X"5180E4DE";
    when 16#0024D# => romdata <= X"3FFF54FE";
    when 16#0024E# => romdata <= X"923981A6";
    when 16#0024F# => romdata <= X"885180E4";
    when 16#00250# => romdata <= X"D13F7681";
    when 16#00251# => romdata <= X"800A2981";
    when 16#00252# => romdata <= X"FF0A0570";
    when 16#00253# => romdata <= X"982C5856";
    when 16#00254# => romdata <= X"768025FC";
    when 16#00255# => romdata <= X"A538FEDA";
    when 16#00256# => romdata <= X"3981A688";
    when 16#00257# => romdata <= X"5180E4B2";
    when 16#00258# => romdata <= X"3FFD9C39";
    when 16#00259# => romdata <= X"81CCCC33";
    when 16#0025A# => romdata <= X"81FD0654";
    when 16#0025B# => romdata <= X"FCDC3981";
    when 16#0025C# => romdata <= X"A6885180";
    when 16#0025D# => romdata <= X"E49C3FFC";
    when 16#0025E# => romdata <= X"BE3981A6";
    when 16#0025F# => romdata <= X"885180E4";
    when 16#00260# => romdata <= X"913F8059";
    when 16#00261# => romdata <= X"8F57FBF2";
    when 16#00262# => romdata <= X"3981A688";
    when 16#00263# => romdata <= X"5180E482";
    when 16#00264# => romdata <= X"3F78B00C";
    when 16#00265# => romdata <= X"8A3D0D04";
    when 16#00266# => romdata <= X"81A68851";
    when 16#00267# => romdata <= X"80E3F33F";
    when 16#00268# => romdata <= X"FECA39FF";
    when 16#00269# => romdata <= X"3D0D8151";
    when 16#0026A# => romdata <= X"BBC73FB0";
    when 16#0026B# => romdata <= X"0881FF06";
    when 16#0026C# => romdata <= X"52818051";
    when 16#0026D# => romdata <= X"FAFD3F82";
    when 16#0026E# => romdata <= X"8051FAF7";
    when 16#0026F# => romdata <= X"3F848351";
    when 16#00270# => romdata <= X"FAF13F86";
    when 16#00271# => romdata <= X"F151FAEB";
    when 16#00272# => romdata <= X"3F71832B";
    when 16#00273# => romdata <= X"88830751";
    when 16#00274# => romdata <= X"FAE13F71";
    when 16#00275# => romdata <= X"B00C833D";
    when 16#00276# => romdata <= X"0D04FE3D";
    when 16#00277# => romdata <= X"0D029305";
    when 16#00278# => romdata <= X"33028405";
    when 16#00279# => romdata <= X"97053354";
    when 16#0027A# => romdata <= X"52717327";
    when 16#0027B# => romdata <= X"9438A051";
    when 16#0027C# => romdata <= X"80E3853F";
    when 16#0027D# => romdata <= X"81127081";
    when 16#0027E# => romdata <= X"FF065152";
    when 16#0027F# => romdata <= X"727226EE";
    when 16#00280# => romdata <= X"38843D0D";
    when 16#00281# => romdata <= X"04FE3D0D";
    when 16#00282# => romdata <= X"74708106";
    when 16#00283# => romdata <= X"53537185";
    when 16#00284# => romdata <= X"D0387281";
    when 16#00285# => romdata <= X"2A708106";
    when 16#00286# => romdata <= X"51527185";
    when 16#00287# => romdata <= X"AC387282";
    when 16#00288# => romdata <= X"2A708106";
    when 16#00289# => romdata <= X"51527185";
    when 16#0028A# => romdata <= X"88387283";
    when 16#0028B# => romdata <= X"2A708106";
    when 16#0028C# => romdata <= X"51527184";
    when 16#0028D# => romdata <= X"E4387284";
    when 16#0028E# => romdata <= X"2A708106";
    when 16#0028F# => romdata <= X"51527184";
    when 16#00290# => romdata <= X"C0387285";
    when 16#00291# => romdata <= X"2A708106";
    when 16#00292# => romdata <= X"51527184";
    when 16#00293# => romdata <= X"9C387286";
    when 16#00294# => romdata <= X"2A708106";
    when 16#00295# => romdata <= X"51527183";
    when 16#00296# => romdata <= X"F8387287";
    when 16#00297# => romdata <= X"2A708106";
    when 16#00298# => romdata <= X"51527183";
    when 16#00299# => romdata <= X"D4387288";
    when 16#0029A# => romdata <= X"2A708106";
    when 16#0029B# => romdata <= X"51527183";
    when 16#0029C# => romdata <= X"B0387289";
    when 16#0029D# => romdata <= X"2A708106";
    when 16#0029E# => romdata <= X"51527183";
    when 16#0029F# => romdata <= X"8C38728A";
    when 16#002A0# => romdata <= X"2A708106";
    when 16#002A1# => romdata <= X"51527182";
    when 16#002A2# => romdata <= X"E838728B";
    when 16#002A3# => romdata <= X"2A708106";
    when 16#002A4# => romdata <= X"51527182";
    when 16#002A5# => romdata <= X"C438728C";
    when 16#002A6# => romdata <= X"2A708106";
    when 16#002A7# => romdata <= X"51527182";
    when 16#002A8# => romdata <= X"A038728D";
    when 16#002A9# => romdata <= X"2A708106";
    when 16#002AA# => romdata <= X"51527181";
    when 16#002AB# => romdata <= X"FC38728E";
    when 16#002AC# => romdata <= X"2A708106";
    when 16#002AD# => romdata <= X"51527181";
    when 16#002AE# => romdata <= X"D838728F";
    when 16#002AF# => romdata <= X"2A708106";
    when 16#002B0# => romdata <= X"51527181";
    when 16#002B1# => romdata <= X"B4387290";
    when 16#002B2# => romdata <= X"2A708106";
    when 16#002B3# => romdata <= X"51527181";
    when 16#002B4# => romdata <= X"90387291";
    when 16#002B5# => romdata <= X"2A708106";
    when 16#002B6# => romdata <= X"51527180";
    when 16#002B7# => romdata <= X"EC387292";
    when 16#002B8# => romdata <= X"2A708106";
    when 16#002B9# => romdata <= X"51527180";
    when 16#002BA# => romdata <= X"C8387293";
    when 16#002BB# => romdata <= X"2A708106";
    when 16#002BC# => romdata <= X"515271A6";
    when 16#002BD# => romdata <= X"3872942A";
    when 16#002BE# => romdata <= X"70810651";
    when 16#002BF# => romdata <= X"52718B38";
    when 16#002C0# => romdata <= X"80732483";
    when 16#002C1# => romdata <= X"F438843D";
    when 16#002C2# => romdata <= X"0D0481A6";
    when 16#002C3# => romdata <= X"C05180E1";
    when 16#002C4# => romdata <= X"813F7280";
    when 16#002C5# => romdata <= X"25F03883";
    when 16#002C6# => romdata <= X"E03981A6";
    when 16#002C7# => romdata <= X"DC5180E0";
    when 16#002C8# => romdata <= X"F13F7294";
    when 16#002C9# => romdata <= X"2A708106";
    when 16#002CA# => romdata <= X"51527180";
    when 16#002CB# => romdata <= X"2ED238DA";
    when 16#002CC# => romdata <= X"3981A6F8";
    when 16#002CD# => romdata <= X"5180E0DA";
    when 16#002CE# => romdata <= X"3F72932A";
    when 16#002CF# => romdata <= X"70810651";
    when 16#002D0# => romdata <= X"5271802E";
    when 16#002D1# => romdata <= X"FFAF38D2";
    when 16#002D2# => romdata <= X"3981A794";
    when 16#002D3# => romdata <= X"5180E0C2";
    when 16#002D4# => romdata <= X"3F72922A";
    when 16#002D5# => romdata <= X"70810651";
    when 16#002D6# => romdata <= X"5271802E";
    when 16#002D7# => romdata <= X"FF8C38D1";
    when 16#002D8# => romdata <= X"3981A7B0";
    when 16#002D9# => romdata <= X"5180E0AA";
    when 16#002DA# => romdata <= X"3F72912A";
    when 16#002DB# => romdata <= X"70810651";
    when 16#002DC# => romdata <= X"5271802E";
    when 16#002DD# => romdata <= X"FEE838D1";
    when 16#002DE# => romdata <= X"3981A7D0";
    when 16#002DF# => romdata <= X"5180E092";
    when 16#002E0# => romdata <= X"3F72902A";
    when 16#002E1# => romdata <= X"70810651";
    when 16#002E2# => romdata <= X"5271802E";
    when 16#002E3# => romdata <= X"FEC438D1";
    when 16#002E4# => romdata <= X"3981A7F0";
    when 16#002E5# => romdata <= X"5180DFFA";
    when 16#002E6# => romdata <= X"3F728F2A";
    when 16#002E7# => romdata <= X"70810651";
    when 16#002E8# => romdata <= X"5271802E";
    when 16#002E9# => romdata <= X"FEA038D1";
    when 16#002EA# => romdata <= X"3981A890";
    when 16#002EB# => romdata <= X"5180DFE2";
    when 16#002EC# => romdata <= X"3F728E2A";
    when 16#002ED# => romdata <= X"70810651";
    when 16#002EE# => romdata <= X"5271802E";
    when 16#002EF# => romdata <= X"FDFC38D1";
    when 16#002F0# => romdata <= X"3981A8B0";
    when 16#002F1# => romdata <= X"5180DFCA";
    when 16#002F2# => romdata <= X"3F728D2A";
    when 16#002F3# => romdata <= X"70810651";
    when 16#002F4# => romdata <= X"5271802E";
    when 16#002F5# => romdata <= X"FDD838D1";
    when 16#002F6# => romdata <= X"3981A8C4";
    when 16#002F7# => romdata <= X"5180DFB2";
    when 16#002F8# => romdata <= X"3F728C2A";
    when 16#002F9# => romdata <= X"70810651";
    when 16#002FA# => romdata <= X"5271802E";
    when 16#002FB# => romdata <= X"FDB438D1";
    when 16#002FC# => romdata <= X"3981A8E4";
    when 16#002FD# => romdata <= X"5180DF9A";
    when 16#002FE# => romdata <= X"3F728B2A";
    when 16#002FF# => romdata <= X"70810651";
    when 16#00300# => romdata <= X"5271802E";
    when 16#00301# => romdata <= X"FD9038D1";
    when 16#00302# => romdata <= X"3981A98C";
    when 16#00303# => romdata <= X"5180DF82";
    when 16#00304# => romdata <= X"3F728A2A";
    when 16#00305# => romdata <= X"70810651";
    when 16#00306# => romdata <= X"5271802E";
    when 16#00307# => romdata <= X"FCEC38D1";
    when 16#00308# => romdata <= X"3981A9AC";
    when 16#00309# => romdata <= X"5180DEEA";
    when 16#0030A# => romdata <= X"3F72892A";
    when 16#0030B# => romdata <= X"70810651";
    when 16#0030C# => romdata <= X"5271802E";
    when 16#0030D# => romdata <= X"FCC838D1";
    when 16#0030E# => romdata <= X"3981A9CC";
    when 16#0030F# => romdata <= X"5180DED2";
    when 16#00310# => romdata <= X"3F72882A";
    when 16#00311# => romdata <= X"70810651";
    when 16#00312# => romdata <= X"5271802E";
    when 16#00313# => romdata <= X"FCA438D1";
    when 16#00314# => romdata <= X"3981A9F4";
    when 16#00315# => romdata <= X"5180DEBA";
    when 16#00316# => romdata <= X"3F72872A";
    when 16#00317# => romdata <= X"70810651";
    when 16#00318# => romdata <= X"5271802E";
    when 16#00319# => romdata <= X"FC8038D1";
    when 16#0031A# => romdata <= X"3981AA94";
    when 16#0031B# => romdata <= X"5180DEA2";
    when 16#0031C# => romdata <= X"3F72862A";
    when 16#0031D# => romdata <= X"70810651";
    when 16#0031E# => romdata <= X"5271802E";
    when 16#0031F# => romdata <= X"FBDC38D1";
    when 16#00320# => romdata <= X"3981AAB4";
    when 16#00321# => romdata <= X"5180DE8A";
    when 16#00322# => romdata <= X"3F72852A";
    when 16#00323# => romdata <= X"70810651";
    when 16#00324# => romdata <= X"5271802E";
    when 16#00325# => romdata <= X"FBB838D1";
    when 16#00326# => romdata <= X"3981AADC";
    when 16#00327# => romdata <= X"5180DDF2";
    when 16#00328# => romdata <= X"3F72842A";
    when 16#00329# => romdata <= X"70810651";
    when 16#0032A# => romdata <= X"5271802E";
    when 16#0032B# => romdata <= X"FB9438D1";
    when 16#0032C# => romdata <= X"3981AAFC";
    when 16#0032D# => romdata <= X"5180DDDA";
    when 16#0032E# => romdata <= X"3F72832A";
    when 16#0032F# => romdata <= X"70810651";
    when 16#00330# => romdata <= X"5271802E";
    when 16#00331# => romdata <= X"FAF038D1";
    when 16#00332# => romdata <= X"3981AB9C";
    when 16#00333# => romdata <= X"5180DDC2";
    when 16#00334# => romdata <= X"3F72822A";
    when 16#00335# => romdata <= X"70810651";
    when 16#00336# => romdata <= X"5271802E";
    when 16#00337# => romdata <= X"FACC38D1";
    when 16#00338# => romdata <= X"3981ABC4";
    when 16#00339# => romdata <= X"5180DDAA";
    when 16#0033A# => romdata <= X"3F72812A";
    when 16#0033B# => romdata <= X"70810651";
    when 16#0033C# => romdata <= X"5271802E";
    when 16#0033D# => romdata <= X"FAA838D1";
    when 16#0033E# => romdata <= X"3981ABE4";
    when 16#0033F# => romdata <= X"5180DD92";
    when 16#00340# => romdata <= X"3F843D0D";
    when 16#00341# => romdata <= X"04FD3D0D";
    when 16#00342# => romdata <= X"81ABF851";
    when 16#00343# => romdata <= X"80DD833F";
    when 16#00344# => romdata <= X"81CCFC08";
    when 16#00345# => romdata <= X"7008709E";
    when 16#00346# => romdata <= X"2A708106";
    when 16#00347# => romdata <= X"51525553";
    when 16#00348# => romdata <= X"81547283";
    when 16#00349# => romdata <= X"38725473";
    when 16#0034A# => romdata <= X"802E88C4";
    when 16#0034B# => romdata <= X"3881AC94";
    when 16#0034C# => romdata <= X"5180DCDE";
    when 16#0034D# => romdata <= X"3F81AC9C";
    when 16#0034E# => romdata <= X"5180DCD6";
    when 16#0034F# => romdata <= X"3F81CCFC";
    when 16#00350# => romdata <= X"08841108";
    when 16#00351# => romdata <= X"709D2A81";
    when 16#00352# => romdata <= X"06515553";
    when 16#00353# => romdata <= X"73802E87";
    when 16#00354# => romdata <= X"B03881AC";
    when 16#00355# => romdata <= X"B85180DC";
    when 16#00356# => romdata <= X"B93F81AC";
    when 16#00357# => romdata <= X"C45180DC";
    when 16#00358# => romdata <= X"B13F81CC";
    when 16#00359# => romdata <= X"C40880D4";
    when 16#0035A# => romdata <= X"11085254";
    when 16#0035B# => romdata <= X"80DDED3F";
    when 16#0035C# => romdata <= X"81ACE051";
    when 16#0035D# => romdata <= X"80DC9B3F";
    when 16#0035E# => romdata <= X"81CCC408";
    when 16#0035F# => romdata <= X"80D01108";
    when 16#00360# => romdata <= X"525380DD";
    when 16#00361# => romdata <= X"D73F8A51";
    when 16#00362# => romdata <= X"80DBED3F";
    when 16#00363# => romdata <= X"81ACFC51";
    when 16#00364# => romdata <= X"80DBFF3F";
    when 16#00365# => romdata <= X"81ADA051";
    when 16#00366# => romdata <= X"80DBF73F";
    when 16#00367# => romdata <= X"81ADE851";
    when 16#00368# => romdata <= X"80DBEF3F";
    when 16#00369# => romdata <= X"81AEB051";
    when 16#0036A# => romdata <= X"80DBE73F";
    when 16#0036B# => romdata <= X"81CCC408";
    when 16#0036C# => romdata <= X"70085254";
    when 16#0036D# => romdata <= X"80DDA53F";
    when 16#0036E# => romdata <= X"B00881FF";
    when 16#0036F# => romdata <= X"0653728C";
    when 16#00370# => romdata <= X"279438A0";
    when 16#00371# => romdata <= X"5180DBB0";
    when 16#00372# => romdata <= X"3F811370";
    when 16#00373# => romdata <= X"81FF0651";
    when 16#00374# => romdata <= X"538C7326";
    when 16#00375# => romdata <= X"EE3881CC";
    when 16#00376# => romdata <= X"C4088411";
    when 16#00377# => romdata <= X"08525480";
    when 16#00378# => romdata <= X"DCFA3FB0";
    when 16#00379# => romdata <= X"0881FF06";
    when 16#0037A# => romdata <= X"53728C27";
    when 16#0037B# => romdata <= X"9438A051";
    when 16#0037C# => romdata <= X"80DB853F";
    when 16#0037D# => romdata <= X"81137081";
    when 16#0037E# => romdata <= X"FF065153";
    when 16#0037F# => romdata <= X"8C7326EE";
    when 16#00380# => romdata <= X"3881CCC4";
    when 16#00381# => romdata <= X"08881108";
    when 16#00382# => romdata <= X"525480DC";
    when 16#00383# => romdata <= X"CF3FB008";
    when 16#00384# => romdata <= X"81FF0653";
    when 16#00385# => romdata <= X"728C2794";
    when 16#00386# => romdata <= X"38A05180";
    when 16#00387# => romdata <= X"DADA3F81";
    when 16#00388# => romdata <= X"137081FF";
    when 16#00389# => romdata <= X"0651538C";
    when 16#0038A# => romdata <= X"7326EE38";
    when 16#0038B# => romdata <= X"81CCC408";
    when 16#0038C# => romdata <= X"8C110852";
    when 16#0038D# => romdata <= X"5480DCA4";
    when 16#0038E# => romdata <= X"3FB00881";
    when 16#0038F# => romdata <= X"FF065372";
    when 16#00390# => romdata <= X"8C279438";
    when 16#00391# => romdata <= X"A05180DA";
    when 16#00392# => romdata <= X"AF3F8113";
    when 16#00393# => romdata <= X"7081FF06";
    when 16#00394# => romdata <= X"51538C73";
    when 16#00395# => romdata <= X"26EE3881";
    when 16#00396# => romdata <= X"AECC5180";
    when 16#00397# => romdata <= X"DAB43F81";
    when 16#00398# => romdata <= X"CCC40890";
    when 16#00399# => romdata <= X"11085254";
    when 16#0039A# => romdata <= X"80DBF13F";
    when 16#0039B# => romdata <= X"B00881FF";
    when 16#0039C# => romdata <= X"0653728C";
    when 16#0039D# => romdata <= X"279438A0";
    when 16#0039E# => romdata <= X"5180D9FC";
    when 16#0039F# => romdata <= X"3F811370";
    when 16#003A0# => romdata <= X"81FF0651";
    when 16#003A1# => romdata <= X"538C7326";
    when 16#003A2# => romdata <= X"EE3881CC";
    when 16#003A3# => romdata <= X"C4089411";
    when 16#003A4# => romdata <= X"08525480";
    when 16#003A5# => romdata <= X"DBC63FB0";
    when 16#003A6# => romdata <= X"0881FF06";
    when 16#003A7# => romdata <= X"53728C27";
    when 16#003A8# => romdata <= X"9438A051";
    when 16#003A9# => romdata <= X"80D9D13F";
    when 16#003AA# => romdata <= X"81137081";
    when 16#003AB# => romdata <= X"FF065153";
    when 16#003AC# => romdata <= X"8C7326EE";
    when 16#003AD# => romdata <= X"3881CCC4";
    when 16#003AE# => romdata <= X"08981108";
    when 16#003AF# => romdata <= X"525480DB";
    when 16#003B0# => romdata <= X"9B3FB008";
    when 16#003B1# => romdata <= X"81FF0653";
    when 16#003B2# => romdata <= X"728C2794";
    when 16#003B3# => romdata <= X"38A05180";
    when 16#003B4# => romdata <= X"D9A63F81";
    when 16#003B5# => romdata <= X"137081FF";
    when 16#003B6# => romdata <= X"0651538C";
    when 16#003B7# => romdata <= X"7326EE38";
    when 16#003B8# => romdata <= X"81CCC408";
    when 16#003B9# => romdata <= X"9C110852";
    when 16#003BA# => romdata <= X"5480DAF0";
    when 16#003BB# => romdata <= X"3FB00881";
    when 16#003BC# => romdata <= X"FF065372";
    when 16#003BD# => romdata <= X"8C279438";
    when 16#003BE# => romdata <= X"A05180D8";
    when 16#003BF# => romdata <= X"FB3F8113";
    when 16#003C0# => romdata <= X"7081FF06";
    when 16#003C1# => romdata <= X"51538C73";
    when 16#003C2# => romdata <= X"26EE3881";
    when 16#003C3# => romdata <= X"AEE85180";
    when 16#003C4# => romdata <= X"D9803F81";
    when 16#003C5# => romdata <= X"CCC40854";
    when 16#003C6# => romdata <= X"810BB015";
    when 16#003C7# => romdata <= X"0CB01408";
    when 16#003C8# => romdata <= X"53728025";
    when 16#003C9# => romdata <= X"F838A014";
    when 16#003CA# => romdata <= X"085180DA";
    when 16#003CB# => romdata <= X"AF3FB008";
    when 16#003CC# => romdata <= X"81FF0653";
    when 16#003CD# => romdata <= X"728C2794";
    when 16#003CE# => romdata <= X"38A05180";
    when 16#003CF# => romdata <= X"D8BA3F81";
    when 16#003D0# => romdata <= X"137081FF";
    when 16#003D1# => romdata <= X"0654548C";
    when 16#003D2# => romdata <= X"7326EE38";
    when 16#003D3# => romdata <= X"81CCC408";
    when 16#003D4# => romdata <= X"A4110852";
    when 16#003D5# => romdata <= X"5380DA84";
    when 16#003D6# => romdata <= X"3FB00881";
    when 16#003D7# => romdata <= X"FF065372";
    when 16#003D8# => romdata <= X"8C279438";
    when 16#003D9# => romdata <= X"A05180D8";
    when 16#003DA# => romdata <= X"8F3F8113";
    when 16#003DB# => romdata <= X"7081FF06";
    when 16#003DC# => romdata <= X"54548C73";
    when 16#003DD# => romdata <= X"26EE3881";
    when 16#003DE# => romdata <= X"CCC408A8";
    when 16#003DF# => romdata <= X"11085253";
    when 16#003E0# => romdata <= X"80D9D93F";
    when 16#003E1# => romdata <= X"B00881FF";
    when 16#003E2# => romdata <= X"0653728C";
    when 16#003E3# => romdata <= X"279438A0";
    when 16#003E4# => romdata <= X"5180D7E4";
    when 16#003E5# => romdata <= X"3F811370";
    when 16#003E6# => romdata <= X"81FF0654";
    when 16#003E7# => romdata <= X"548C7326";
    when 16#003E8# => romdata <= X"EE3881CC";
    when 16#003E9# => romdata <= X"C408AC11";
    when 16#003EA# => romdata <= X"08525380";
    when 16#003EB# => romdata <= X"D9AE3FB0";
    when 16#003EC# => romdata <= X"0881FF06";
    when 16#003ED# => romdata <= X"53728C27";
    when 16#003EE# => romdata <= X"9438A051";
    when 16#003EF# => romdata <= X"80D7B93F";
    when 16#003F0# => romdata <= X"81137081";
    when 16#003F1# => romdata <= X"FF065454";
    when 16#003F2# => romdata <= X"8C7326EE";
    when 16#003F3# => romdata <= X"3881AF84";
    when 16#003F4# => romdata <= X"5180D7BE";
    when 16#003F5# => romdata <= X"3F81CCC4";
    when 16#003F6# => romdata <= X"0880E011";
    when 16#003F7# => romdata <= X"08525380";
    when 16#003F8# => romdata <= X"D8FA3F81";
    when 16#003F9# => romdata <= X"AF985180";
    when 16#003FA# => romdata <= X"D7A83F81";
    when 16#003FB# => romdata <= X"CCC408B0";
    when 16#003FC# => romdata <= X"1108FE0A";
    when 16#003FD# => romdata <= X"06525480";
    when 16#003FE# => romdata <= X"D8E23F81";
    when 16#003FF# => romdata <= X"CCC40854";
    when 16#00400# => romdata <= X"800BB015";
    when 16#00401# => romdata <= X"0C81AFAC";
    when 16#00402# => romdata <= X"5180D786";
    when 16#00403# => romdata <= X"3F81AFC4";
    when 16#00404# => romdata <= X"5180D6FE";
    when 16#00405# => romdata <= X"3F81CCC4";
    when 16#00406# => romdata <= X"0880C011";
    when 16#00407# => romdata <= X"08525380";
    when 16#00408# => romdata <= X"D8BA3FB0";
    when 16#00409# => romdata <= X"0881FF06";
    when 16#0040A# => romdata <= X"53729827";
    when 16#0040B# => romdata <= X"9438A051";
    when 16#0040C# => romdata <= X"80D6C53F";
    when 16#0040D# => romdata <= X"81137081";
    when 16#0040E# => romdata <= X"FF065454";
    when 16#0040F# => romdata <= X"987326EE";
    when 16#00410# => romdata <= X"3881CCC4";
    when 16#00411# => romdata <= X"0880C811";
    when 16#00412# => romdata <= X"08525380";
    when 16#00413# => romdata <= X"D88E3FB0";
    when 16#00414# => romdata <= X"0881FF06";
    when 16#00415# => romdata <= X"53729827";
    when 16#00416# => romdata <= X"9438A051";
    when 16#00417# => romdata <= X"80D6993F";
    when 16#00418# => romdata <= X"81137081";
    when 16#00419# => romdata <= X"FF065454";
    when 16#0041A# => romdata <= X"987326EE";
    when 16#0041B# => romdata <= X"3881AFE0";
    when 16#0041C# => romdata <= X"5180D69E";
    when 16#0041D# => romdata <= X"3F81CCC4";
    when 16#0041E# => romdata <= X"0880C411";
    when 16#0041F# => romdata <= X"08525380";
    when 16#00420# => romdata <= X"D7DA3FB0";
    when 16#00421# => romdata <= X"0881FF06";
    when 16#00422# => romdata <= X"53729827";
    when 16#00423# => romdata <= X"9438A051";
    when 16#00424# => romdata <= X"80D5E53F";
    when 16#00425# => romdata <= X"81137081";
    when 16#00426# => romdata <= X"FF065454";
    when 16#00427# => romdata <= X"987326EE";
    when 16#00428# => romdata <= X"3881CCC4";
    when 16#00429# => romdata <= X"0880CC11";
    when 16#0042A# => romdata <= X"08525380";
    when 16#0042B# => romdata <= X"D7AE3FB0";
    when 16#0042C# => romdata <= X"0881FF06";
    when 16#0042D# => romdata <= X"53729827";
    when 16#0042E# => romdata <= X"9438A051";
    when 16#0042F# => romdata <= X"80D5B93F";
    when 16#00430# => romdata <= X"81137081";
    when 16#00431# => romdata <= X"FF065454";
    when 16#00432# => romdata <= X"987326EE";
    when 16#00433# => romdata <= X"388A5180";
    when 16#00434# => romdata <= X"D5A63F81";
    when 16#00435# => romdata <= X"CCC408B4";
    when 16#00436# => romdata <= X"110881AF";
    when 16#00437# => romdata <= X"FC535153";
    when 16#00438# => romdata <= X"80D5AF3F";
    when 16#00439# => romdata <= X"725180D6";
    when 16#0043A# => romdata <= X"F33FA051";
    when 16#0043B# => romdata <= X"80D5893F";
    when 16#0043C# => romdata <= X"72862681";
    when 16#0043D# => romdata <= X"8E387210";
    when 16#0043E# => romdata <= X"1081BCB0";
    when 16#0043F# => romdata <= X"05547308";
    when 16#00440# => romdata <= X"0481B090";
    when 16#00441# => romdata <= X"5180D58A";
    when 16#00442# => romdata <= X"3F81ACC4";
    when 16#00443# => romdata <= X"5180D582";
    when 16#00444# => romdata <= X"3F81CCC4";
    when 16#00445# => romdata <= X"0880D411";
    when 16#00446# => romdata <= X"08525480";
    when 16#00447# => romdata <= X"D6BE3F81";
    when 16#00448# => romdata <= X"ACE05180";
    when 16#00449# => romdata <= X"D4EC3F81";
    when 16#0044A# => romdata <= X"CCC40880";
    when 16#0044B# => romdata <= X"D0110852";
    when 16#0044C# => romdata <= X"5380D6A8";
    when 16#0044D# => romdata <= X"3F8A5180";
    when 16#0044E# => romdata <= X"D4BE3F81";
    when 16#0044F# => romdata <= X"ACFC5180";
    when 16#00450# => romdata <= X"D4D03F81";
    when 16#00451# => romdata <= X"ADA05180";
    when 16#00452# => romdata <= X"D4C83F81";
    when 16#00453# => romdata <= X"ADE85180";
    when 16#00454# => romdata <= X"D4C03F81";
    when 16#00455# => romdata <= X"AEB05180";
    when 16#00456# => romdata <= X"D4B83F81";
    when 16#00457# => romdata <= X"CCC40870";
    when 16#00458# => romdata <= X"08525480";
    when 16#00459# => romdata <= X"D5F63FB0";
    when 16#0045A# => romdata <= X"0881FF06";
    when 16#0045B# => romdata <= X"53F8CF39";
    when 16#0045C# => romdata <= X"81B09851";
    when 16#0045D# => romdata <= X"80D49B3F";
    when 16#0045E# => romdata <= X"F7B33981";
    when 16#0045F# => romdata <= X"B0A05180";
    when 16#00460# => romdata <= X"D4903F81";
    when 16#00461# => romdata <= X"CCC408B8";
    when 16#00462# => romdata <= X"110881B0";
    when 16#00463# => romdata <= X"AC535454";
    when 16#00464# => romdata <= X"80D3FF3F";
    when 16#00465# => romdata <= X"7252A051";
    when 16#00466# => romdata <= X"80D49A3F";
    when 16#00467# => romdata <= X"7251F0E5";
    when 16#00468# => romdata <= X"3F8A5180";
    when 16#00469# => romdata <= X"D3D23F80";
    when 16#0046A# => romdata <= X"0BB00C85";
    when 16#0046B# => romdata <= X"3D0D0481";
    when 16#0046C# => romdata <= X"B0C05180";
    when 16#0046D# => romdata <= X"D3DC3FCB";
    when 16#0046E# => romdata <= X"3981B0CC";
    when 16#0046F# => romdata <= X"5180D3D2";
    when 16#00470# => romdata <= X"3FC13981";
    when 16#00471# => romdata <= X"B0D85180";
    when 16#00472# => romdata <= X"D3C83FFF";
    when 16#00473# => romdata <= X"B63981B0";
    when 16#00474# => romdata <= X"DC5180D3";
    when 16#00475# => romdata <= X"BD3FFFAB";
    when 16#00476# => romdata <= X"3981B0E8";
    when 16#00477# => romdata <= X"5180D3B2";
    when 16#00478# => romdata <= X"3FFFA039";
    when 16#00479# => romdata <= X"81B0F451";
    when 16#0047A# => romdata <= X"80D3A73F";
    when 16#0047B# => romdata <= X"FF9539FE";
    when 16#0047C# => romdata <= X"3D0D8151";
    when 16#0047D# => romdata <= X"AAFB3FB0";
    when 16#0047E# => romdata <= X"0881FF06";
    when 16#0047F# => romdata <= X"81CCC408";
    when 16#00480# => romdata <= X"71B4120C";
    when 16#00481# => romdata <= X"53B00C84";
    when 16#00482# => romdata <= X"3D0D04FE";
    when 16#00483# => romdata <= X"3D0D880A";
    when 16#00484# => romdata <= X"53840A0B";
    when 16#00485# => romdata <= X"81CCC008";
    when 16#00486# => romdata <= X"8C110851";
    when 16#00487# => romdata <= X"52528071";
    when 16#00488# => romdata <= X"27953880";
    when 16#00489# => romdata <= X"73708405";
    when 16#0048A# => romdata <= X"550C8072";
    when 16#0048B# => romdata <= X"70840554";
    when 16#0048C# => romdata <= X"0CFF1151";
    when 16#0048D# => romdata <= X"70ED3880";
    when 16#0048E# => romdata <= X"0BB00C84";
    when 16#0048F# => romdata <= X"3D0D04FA";
    when 16#00490# => romdata <= X"3D0D880A";
    when 16#00491# => romdata <= X"57840A56";
    when 16#00492# => romdata <= X"8151AAA5";
    when 16#00493# => romdata <= X"3FB00883";
    when 16#00494# => romdata <= X"FFFF0654";
    when 16#00495# => romdata <= X"73833890";
    when 16#00496# => romdata <= X"54805574";
    when 16#00497# => romdata <= X"742781C2";
    when 16#00498# => romdata <= X"38750870";
    when 16#00499# => romdata <= X"902C5253";
    when 16#0049A# => romdata <= X"80D3F13F";
    when 16#0049B# => romdata <= X"B00881FF";
    when 16#0049C# => romdata <= X"0652718A";
    when 16#0049D# => romdata <= X"279438A0";
    when 16#0049E# => romdata <= X"5180D1FC";
    when 16#0049F# => romdata <= X"3F811270";
    when 16#004A0# => romdata <= X"81FF0651";
    when 16#004A1# => romdata <= X"528A7226";
    when 16#004A2# => romdata <= X"EE387290";
    when 16#004A3# => romdata <= X"2B70902C";
    when 16#004A4# => romdata <= X"525280D3";
    when 16#004A5# => romdata <= X"C73FB008";
    when 16#004A6# => romdata <= X"81FF0652";
    when 16#004A7# => romdata <= X"718A2794";
    when 16#004A8# => romdata <= X"38A05180";
    when 16#004A9# => romdata <= X"D1D23F81";
    when 16#004AA# => romdata <= X"127081FF";
    when 16#004AB# => romdata <= X"0653538A";
    when 16#004AC# => romdata <= X"7226EE38";
    when 16#004AD# => romdata <= X"76087090";
    when 16#004AE# => romdata <= X"2C525380";
    when 16#004AF# => romdata <= X"D39E3FB0";
    when 16#004B0# => romdata <= X"0881FF06";
    when 16#004B1# => romdata <= X"52718A27";
    when 16#004B2# => romdata <= X"9438A051";
    when 16#004B3# => romdata <= X"80D1A93F";
    when 16#004B4# => romdata <= X"81127081";
    when 16#004B5# => romdata <= X"FF065152";
    when 16#004B6# => romdata <= X"8A7226EE";
    when 16#004B7# => romdata <= X"3872902B";
    when 16#004B8# => romdata <= X"70902C52";
    when 16#004B9# => romdata <= X"5280D2F4";
    when 16#004BA# => romdata <= X"3FB00881";
    when 16#004BB# => romdata <= X"FF065271";
    when 16#004BC# => romdata <= X"8A279438";
    when 16#004BD# => romdata <= X"A05180D0";
    when 16#004BE# => romdata <= X"FF3F8112";
    when 16#004BF# => romdata <= X"7081FF06";
    when 16#004C0# => romdata <= X"53538A72";
    when 16#004C1# => romdata <= X"26EE388A";
    when 16#004C2# => romdata <= X"5180D0EC";
    when 16#004C3# => romdata <= X"3F841784";
    when 16#004C4# => romdata <= X"17811770";
    when 16#004C5# => romdata <= X"83FFFF06";
    when 16#004C6# => romdata <= X"58545757";
    when 16#004C7# => romdata <= X"737526FE";
    when 16#004C8# => romdata <= X"C03873B0";
    when 16#004C9# => romdata <= X"0C883D0D";
    when 16#004CA# => romdata <= X"04FD3D0D";
    when 16#004CB# => romdata <= X"8151A8C1";
    when 16#004CC# => romdata <= X"3FB00881";
    when 16#004CD# => romdata <= X"FF065473";
    when 16#004CE# => romdata <= X"802EA438";
    when 16#004CF# => romdata <= X"73842690";
    when 16#004D0# => romdata <= X"3881CCC0";
    when 16#004D1# => romdata <= X"0874710C";
    when 16#004D2# => romdata <= X"5373B00C";
    when 16#004D3# => romdata <= X"853D0D04";
    when 16#004D4# => romdata <= X"81CCC008";
    when 16#004D5# => romdata <= X"5380730C";
    when 16#004D6# => romdata <= X"73B00C85";
    when 16#004D7# => romdata <= X"3D0D0481";
    when 16#004D8# => romdata <= X"B2805180";
    when 16#004D9# => romdata <= X"D0AC3F81";
    when 16#004DA# => romdata <= X"B2905180";
    when 16#004DB# => romdata <= X"D0A43F81";
    when 16#004DC# => romdata <= X"CCC00870";
    when 16#004DD# => romdata <= X"08525380";
    when 16#004DE# => romdata <= X"D1E23F81";
    when 16#004DF# => romdata <= X"B2A05180";
    when 16#004E0# => romdata <= X"D0903F81";
    when 16#004E1# => romdata <= X"CCC00884";
    when 16#004E2# => romdata <= X"11085353";
    when 16#004E3# => romdata <= X"A05180D0";
    when 16#004E4# => romdata <= X"A43F81B2";
    when 16#004E5# => romdata <= X"B45180CF";
    when 16#004E6# => romdata <= X"F93F81CC";
    when 16#004E7# => romdata <= X"C0088811";
    when 16#004E8# => romdata <= X"085353A0";
    when 16#004E9# => romdata <= X"5180D08D";
    when 16#004EA# => romdata <= X"3F81B2C8";
    when 16#004EB# => romdata <= X"5180CFE2";
    when 16#004EC# => romdata <= X"3F81CCC0";
    when 16#004ED# => romdata <= X"088C1108";
    when 16#004EE# => romdata <= X"525380D1";
    when 16#004EF# => romdata <= X"9F3F8A51";
    when 16#004F0# => romdata <= X"80CFB53F";
    when 16#004F1# => romdata <= X"73B00C85";
    when 16#004F2# => romdata <= X"3D0D04BC";
    when 16#004F3# => romdata <= X"0802BC0C";
    when 16#004F4# => romdata <= X"F93D0D02";
    when 16#004F5# => romdata <= X"BC08FC05";
    when 16#004F6# => romdata <= X"0C880A0B";
    when 16#004F7# => romdata <= X"BC08F405";
    when 16#004F8# => romdata <= X"0CFC3D0D";
    when 16#004F9# => romdata <= X"823DBC08";
    when 16#004FA# => romdata <= X"F0050C81";
    when 16#004FB# => romdata <= X"51A7823F";
    when 16#004FC# => romdata <= X"B00881FF";
    when 16#004FD# => romdata <= X"06BC08F8";
    when 16#004FE# => romdata <= X"050C8251";
    when 16#004FF# => romdata <= X"A6F33FB0";
    when 16#00500# => romdata <= X"08BC08F0";
    when 16#00501# => romdata <= X"05082383";
    when 16#00502# => romdata <= X"51A6E63F";
    when 16#00503# => romdata <= X"B008BC08";
    when 16#00504# => romdata <= X"F0050882";
    when 16#00505# => romdata <= X"05238451";
    when 16#00506# => romdata <= X"A6D73FB0";
    when 16#00507# => romdata <= X"08BC08F0";
    when 16#00508# => romdata <= X"05088405";
    when 16#00509# => romdata <= X"238551A6";
    when 16#0050A# => romdata <= X"C83FB008";
    when 16#0050B# => romdata <= X"BC08F005";
    when 16#0050C# => romdata <= X"08860523";
    when 16#0050D# => romdata <= X"8651A6B9";
    when 16#0050E# => romdata <= X"3FB008BC";
    when 16#0050F# => romdata <= X"08F00508";
    when 16#00510# => romdata <= X"88052387";
    when 16#00511# => romdata <= X"51A6AA3F";
    when 16#00512# => romdata <= X"B008BC08";
    when 16#00513# => romdata <= X"F005088A";
    when 16#00514# => romdata <= X"05238851";
    when 16#00515# => romdata <= X"A69B3FB0";
    when 16#00516# => romdata <= X"08BC08F0";
    when 16#00517# => romdata <= X"05088C05";
    when 16#00518# => romdata <= X"238951A6";
    when 16#00519# => romdata <= X"8C3FB008";
    when 16#0051A# => romdata <= X"BC08F005";
    when 16#0051B# => romdata <= X"088E0523";
    when 16#0051C# => romdata <= X"800B81CC";
    when 16#0051D# => romdata <= X"C008708C";
    when 16#0051E# => romdata <= X"050851BC";
    when 16#0051F# => romdata <= X"08E4050C";
    when 16#00520# => romdata <= X"BC08EC05";
    when 16#00521# => romdata <= X"0CBC08EC";
    when 16#00522# => romdata <= X"0508BC08";
    when 16#00523# => romdata <= X"E4050827";
    when 16#00524# => romdata <= X"818F38BC";
    when 16#00525# => romdata <= X"08E40508";
    when 16#00526# => romdata <= X"BC08E805";
    when 16#00527# => romdata <= X"0CBC08F8";
    when 16#00528# => romdata <= X"0508802E";
    when 16#00529# => romdata <= X"81B638BC";
    when 16#0052A# => romdata <= X"08EC0508";
    when 16#0052B# => romdata <= X"10BC08F0";
    when 16#0052C# => romdata <= X"05080570";
    when 16#0052D# => romdata <= X"22BC08F4";
    when 16#0052E# => romdata <= X"05088205";
    when 16#0052F# => romdata <= X"2271902B";
    when 16#00530# => romdata <= X"07BC08F4";
    when 16#00531# => romdata <= X"05080CBC";
    when 16#00532# => romdata <= X"08E4050C";
    when 16#00533# => romdata <= X"BC08F805";
    when 16#00534# => romdata <= X"0CBC08EC";
    when 16#00535# => romdata <= X"05088105";
    when 16#00536# => romdata <= X"7081FF06";
    when 16#00537# => romdata <= X"BC08E405";
    when 16#00538# => romdata <= X"0CBC08F8";
    when 16#00539# => romdata <= X"050C860B";
    when 16#0053A# => romdata <= X"BC08EC05";
    when 16#0053B# => romdata <= X"08278838";
    when 16#0053C# => romdata <= X"800BBC08";
    when 16#0053D# => romdata <= X"E4050CBC";
    when 16#0053E# => romdata <= X"08E40508";
    when 16#0053F# => romdata <= X"BC08F405";
    when 16#00540# => romdata <= X"088405BC";
    when 16#00541# => romdata <= X"08E80508";
    when 16#00542# => romdata <= X"FF05BC08";
    when 16#00543# => romdata <= X"E8050CBC";
    when 16#00544# => romdata <= X"08F4050C";
    when 16#00545# => romdata <= X"BC08EC05";
    when 16#00546# => romdata <= X"0CBC08E8";
    when 16#00547# => romdata <= X"0508FF87";
    when 16#00548# => romdata <= X"38BC08FC";
    when 16#00549# => romdata <= X"05080D80";
    when 16#0054A# => romdata <= X"0BB00C89";
    when 16#0054B# => romdata <= X"3D0DBC0C";
    when 16#0054C# => romdata <= X"04BC08E4";
    when 16#0054D# => romdata <= X"0508BC08";
    when 16#0054E# => romdata <= X"F4050884";
    when 16#0054F# => romdata <= X"05BC08E8";
    when 16#00550# => romdata <= X"0508FF05";
    when 16#00551# => romdata <= X"BC08E805";
    when 16#00552# => romdata <= X"0CBC08F4";
    when 16#00553# => romdata <= X"050CBC08";
    when 16#00554# => romdata <= X"EC050CBC";
    when 16#00555# => romdata <= X"08E80508";
    when 16#00556# => romdata <= X"802EC638";
    when 16#00557# => romdata <= X"BC08EC05";
    when 16#00558# => romdata <= X"0810BC08";
    when 16#00559# => romdata <= X"F0050805";
    when 16#0055A# => romdata <= X"70227090";
    when 16#0055B# => romdata <= X"2BBC08F4";
    when 16#0055C# => romdata <= X"050808FC";
    when 16#0055D# => romdata <= X"80800671";
    when 16#0055E# => romdata <= X"902C07BC";
    when 16#0055F# => romdata <= X"08F40508";
    when 16#00560# => romdata <= X"0C52BC08";
    when 16#00561# => romdata <= X"E4050CBC";
    when 16#00562# => romdata <= X"08F8050C";
    when 16#00563# => romdata <= X"800BBC08";
    when 16#00564# => romdata <= X"E4050CBC";
    when 16#00565# => romdata <= X"08EC0508";
    when 16#00566# => romdata <= X"8626FF95";
    when 16#00567# => romdata <= X"38BC08EC";
    when 16#00568# => romdata <= X"05088105";
    when 16#00569# => romdata <= X"7081FF06";
    when 16#0056A# => romdata <= X"BC08F405";
    when 16#0056B# => romdata <= X"088405BC";
    when 16#0056C# => romdata <= X"08E80508";
    when 16#0056D# => romdata <= X"FF05BC08";
    when 16#0056E# => romdata <= X"E8050CBC";
    when 16#0056F# => romdata <= X"08F4050C";
    when 16#00570# => romdata <= X"BC08EC05";
    when 16#00571# => romdata <= X"0CBC08E4";
    when 16#00572# => romdata <= X"050CBC08";
    when 16#00573# => romdata <= X"E80508FF";
    when 16#00574# => romdata <= X"8B38FECD";
    when 16#00575# => romdata <= X"39FB3D0D";
    when 16#00576# => romdata <= X"029F0533";
    when 16#00577# => romdata <= X"79982B70";
    when 16#00578# => romdata <= X"982C5154";
    when 16#00579# => romdata <= X"55810A54";
    when 16#0057A# => romdata <= X"805672E8";
    when 16#0057B# => romdata <= X"25BD38E8";
    when 16#0057C# => romdata <= X"53751081";
    when 16#0057D# => romdata <= X"07738180";
    when 16#0057E# => romdata <= X"0A298180";
    when 16#0057F# => romdata <= X"0A057098";
    when 16#00580# => romdata <= X"2C515456";
    when 16#00581# => romdata <= X"807324E9";
    when 16#00582# => romdata <= X"38807325";
    when 16#00583# => romdata <= X"80C73873";
    when 16#00584# => romdata <= X"812A810A";
    when 16#00585# => romdata <= X"07738180";
    when 16#00586# => romdata <= X"0A2981FF";
    when 16#00587# => romdata <= X"0A057098";
    when 16#00588# => romdata <= X"2C515454";
    when 16#00589# => romdata <= X"728024E7";
    when 16#0058A# => romdata <= X"38AB3997";
    when 16#0058B# => romdata <= X"73259A38";
    when 16#0058C# => romdata <= X"9774812A";
    when 16#0058D# => romdata <= X"810A0771";
    when 16#0058E# => romdata <= X"81800A29";
    when 16#0058F# => romdata <= X"81FF0A05";
    when 16#00590# => romdata <= X"70982C51";
    when 16#00591# => romdata <= X"525553DC";
    when 16#00592# => romdata <= X"39807324";
    when 16#00593# => romdata <= X"FFA33872";
    when 16#00594# => romdata <= X"8024FFBB";
    when 16#00595# => romdata <= X"38745280";
    when 16#00596# => romdata <= X"51B1B53F";
    when 16#00597# => romdata <= X"7381FF06";
    when 16#00598# => romdata <= X"51B2B33F";
    when 16#00599# => romdata <= X"74528151";
    when 16#0059A# => romdata <= X"B1A63F73";
    when 16#0059B# => romdata <= X"882A7081";
    when 16#0059C# => romdata <= X"FF065253";
    when 16#0059D# => romdata <= X"B2A03F74";
    when 16#0059E# => romdata <= X"528251B1";
    when 16#0059F# => romdata <= X"933F7390";
    when 16#005A0# => romdata <= X"2A7081FF";
    when 16#005A1# => romdata <= X"065253B2";
    when 16#005A2# => romdata <= X"8D3F7452";
    when 16#005A3# => romdata <= X"8351B180";
    when 16#005A4# => romdata <= X"3F73982A";
    when 16#005A5# => romdata <= X"51B1FF3F";
    when 16#005A6# => romdata <= X"74528451";
    when 16#005A7# => romdata <= X"B0F23F75";
    when 16#005A8# => romdata <= X"81FF0651";
    when 16#005A9# => romdata <= X"B1F03F74";
    when 16#005AA# => romdata <= X"528551B0";
    when 16#005AB# => romdata <= X"E33F7588";
    when 16#005AC# => romdata <= X"2A7081FF";
    when 16#005AD# => romdata <= X"065253B1";
    when 16#005AE# => romdata <= X"DD3F7452";
    when 16#005AF# => romdata <= X"8651B0D0";
    when 16#005B0# => romdata <= X"3F75902A";
    when 16#005B1# => romdata <= X"7081FF06";
    when 16#005B2# => romdata <= X"5254B1CA";
    when 16#005B3# => romdata <= X"3F745287";
    when 16#005B4# => romdata <= X"51B0BD3F";
    when 16#005B5# => romdata <= X"75982A51";
    when 16#005B6# => romdata <= X"B1BC3F87";
    when 16#005B7# => romdata <= X"3D0D04F2";
    when 16#005B8# => romdata <= X"3D0D0280";
    when 16#005B9# => romdata <= X"C3053302";
    when 16#005BA# => romdata <= X"840580C7";
    when 16#005BB# => romdata <= X"05338180";
    when 16#005BC# => romdata <= X"0A712B98";
    when 16#005BD# => romdata <= X"2A81CCC0";
    when 16#005BE# => romdata <= X"088C1108";
    when 16#005BF# => romdata <= X"71084453";
    when 16#005C0# => romdata <= X"565C5557";
    when 16#005C1# => romdata <= X"80730C80";
    when 16#005C2# => romdata <= X"7071725C";
    when 16#005C3# => romdata <= X"5A5E5B80";
    when 16#005C4# => romdata <= X"56757A27";
    when 16#005C5# => romdata <= X"80D73881";
    when 16#005C6# => romdata <= X"772783CE";
    when 16#005C7# => romdata <= X"387783FF";
    when 16#005C8# => romdata <= X"FF068119";
    when 16#005C9# => romdata <= X"71101084";
    when 16#005CA# => romdata <= X"0A057930";
    when 16#005CB# => romdata <= X"7A823270";
    when 16#005CC# => romdata <= X"30728025";
    when 16#005CD# => romdata <= X"71802507";
    when 16#005CE# => romdata <= X"56585841";
    when 16#005CF# => romdata <= X"57595C7B";
    when 16#005D0# => romdata <= X"802E83D5";
    when 16#005D1# => romdata <= X"38821522";
    when 16#005D2# => romdata <= X"5372902B";
    when 16#005D3# => romdata <= X"70902C54";
    when 16#005D4# => romdata <= X"55727B25";
    when 16#005D5# => romdata <= X"8338725B";
    when 16#005D6# => romdata <= X"7C732583";
    when 16#005D7# => romdata <= X"38725D81";
    when 16#005D8# => romdata <= X"167081FF";
    when 16#005D9# => romdata <= X"06575E79";
    when 16#005DA# => romdata <= X"7626FFB1";
    when 16#005DB# => romdata <= X"38811970";
    when 16#005DC# => romdata <= X"81FF065A";
    when 16#005DD# => romdata <= X"5680E579";
    when 16#005DE# => romdata <= X"27FF9438";
    when 16#005DF# => romdata <= X"987D3590";
    when 16#005E0# => romdata <= X"2B70902C";
    when 16#005E1# => romdata <= X"7C309871";
    when 16#005E2# => romdata <= X"35902B70";
    when 16#005E3# => romdata <= X"902C5C5C";
    when 16#005E4# => romdata <= X"55565477";
    when 16#005E5# => romdata <= X"54777525";
    when 16#005E6# => romdata <= X"83387454";
    when 16#005E7# => romdata <= X"73902B70";
    when 16#005E8# => romdata <= X"902C5D55";
    when 16#005E9# => romdata <= X"7B54807C";
    when 16#005EA# => romdata <= X"2583D738";
    when 16#005EB# => romdata <= X"73902B70";
    when 16#005EC# => romdata <= X"902C5F56";
    when 16#005ED# => romdata <= X"80705D58";
    when 16#005EE# => romdata <= X"80705A56";
    when 16#005EF# => romdata <= X"757A2780";
    when 16#005F0# => romdata <= X"E4388177";
    when 16#005F1# => romdata <= X"27838C38";
    when 16#005F2# => romdata <= X"7783FFFF";
    when 16#005F3# => romdata <= X"06811971";
    when 16#005F4# => romdata <= X"1010840A";
    when 16#005F5# => romdata <= X"0579307A";
    when 16#005F6# => romdata <= X"82327030";
    when 16#005F7# => romdata <= X"72802571";
    when 16#005F8# => romdata <= X"80250753";
    when 16#005F9# => romdata <= X"51575357";
    when 16#005FA# => romdata <= X"59547380";
    when 16#005FB# => romdata <= X"2E83A438";
    when 16#005FC# => romdata <= X"82152254";
    when 16#005FD# => romdata <= X"73902B70";
    when 16#005FE# => romdata <= X"902C719F";
    when 16#005FF# => romdata <= X"2C707232";
    when 16#00600# => romdata <= X"7131799F";
    when 16#00601# => romdata <= X"2C707B32";
    when 16#00602# => romdata <= X"71315154";
    when 16#00603# => romdata <= X"51565653";
    when 16#00604# => romdata <= X"72742583";
    when 16#00605# => romdata <= X"38745681";
    when 16#00606# => romdata <= X"197081FF";
    when 16#00607# => romdata <= X"065A5579";
    when 16#00608# => romdata <= X"7926FFA4";
    when 16#00609# => romdata <= X"387D7635";
    when 16#0060A# => romdata <= X"982B7098";
    when 16#0060B# => romdata <= X"2C53547B";
    when 16#0060C# => romdata <= X"51FBA23F";
    when 16#0060D# => romdata <= X"811C7081";
    when 16#0060E# => romdata <= X"FF065D59";
    when 16#0060F# => romdata <= X"80E57C27";
    when 16#00610# => romdata <= X"FEF63881";
    when 16#00611# => romdata <= X"CCC0087F";
    when 16#00612# => romdata <= X"710C5880";
    when 16#00613# => romdata <= X"5281C19C";
    when 16#00614# => romdata <= X"51B1B33F";
    when 16#00615# => romdata <= X"81F0DC08";
    when 16#00616# => romdata <= X"80F3CA0B";
    when 16#00617# => romdata <= X"81F0DC0C";
    when 16#00618# => romdata <= X"5F805280";
    when 16#00619# => romdata <= X"51ADA93F";
    when 16#0061A# => romdata <= X"81B2D851";
    when 16#0061B# => romdata <= X"80C6A33F";
    when 16#0061C# => romdata <= X"7C5180C7";
    when 16#0061D# => romdata <= X"E73F8052";
    when 16#0061E# => romdata <= X"8751AD94";
    when 16#0061F# => romdata <= X"3F81B2E0";
    when 16#00620# => romdata <= X"5180C68E";
    when 16#00621# => romdata <= X"3F7A5180";
    when 16#00622# => romdata <= X"C7D23F80";
    when 16#00623# => romdata <= X"D2528051";
    when 16#00624# => romdata <= X"ACFE3F81";
    when 16#00625# => romdata <= X"B2E85180";
    when 16#00626# => romdata <= X"C5F83F76";
    when 16#00627# => romdata <= X"5180C7BC";
    when 16#00628# => romdata <= X"3F80C052";
    when 16#00629# => romdata <= X"8751ACE8";
    when 16#0062A# => romdata <= X"3F81B2F0";
    when 16#0062B# => romdata <= X"5180C5E2";
    when 16#0062C# => romdata <= X"3F7980E6";
    when 16#0062D# => romdata <= X"295180C7";
    when 16#0062E# => romdata <= X"A33F7E81";
    when 16#0062F# => romdata <= X"F0DC0C90";
    when 16#00630# => romdata <= X"3D0D0474";
    when 16#00631# => romdata <= X"22537290";
    when 16#00632# => romdata <= X"2B70902C";
    when 16#00633# => romdata <= X"545C727B";
    when 16#00634# => romdata <= X"25833872";
    when 16#00635# => romdata <= X"5B7C7325";
    when 16#00636# => romdata <= X"8338725D";
    when 16#00637# => romdata <= X"81167081";
    when 16#00638# => romdata <= X"FF06575E";
    when 16#00639# => romdata <= X"757A27FD";
    when 16#0063A# => romdata <= X"84387783";
    when 16#0063B# => romdata <= X"FFFF0681";
    when 16#0063C# => romdata <= X"19711010";
    when 16#0063D# => romdata <= X"880A0579";
    when 16#0063E# => romdata <= X"307A8232";
    when 16#0063F# => romdata <= X"70307280";
    when 16#00640# => romdata <= X"25718025";
    when 16#00641# => romdata <= X"07565840";
    when 16#00642# => romdata <= X"41575954";
    when 16#00643# => romdata <= X"73802EFF";
    when 16#00644# => romdata <= X"B2388215";
    when 16#00645# => romdata <= X"2253FFAE";
    when 16#00646# => romdata <= X"39742253";
    when 16#00647# => romdata <= X"FCAB3974";
    when 16#00648# => romdata <= X"22547390";
    when 16#00649# => romdata <= X"2B70902C";
    when 16#0064A# => romdata <= X"719F2C70";
    when 16#0064B# => romdata <= X"72327131";
    when 16#0064C# => romdata <= X"799F2C70";
    when 16#0064D# => romdata <= X"7B327131";
    when 16#0064E# => romdata <= X"51545156";
    when 16#0064F# => romdata <= X"56537274";
    when 16#00650# => romdata <= X"25833874";
    when 16#00651# => romdata <= X"56811970";
    when 16#00652# => romdata <= X"81FF065A";
    when 16#00653# => romdata <= X"55787A27";
    when 16#00654# => romdata <= X"FDD33877";
    when 16#00655# => romdata <= X"83FFFF06";
    when 16#00656# => romdata <= X"81197110";
    when 16#00657# => romdata <= X"10880A05";
    when 16#00658# => romdata <= X"79307A82";
    when 16#00659# => romdata <= X"32703072";
    when 16#0065A# => romdata <= X"80257180";
    when 16#0065B# => romdata <= X"25075351";
    when 16#0065C# => romdata <= X"57535759";
    when 16#0065D# => romdata <= X"5473802E";
    when 16#0065E# => romdata <= X"FFA53882";
    when 16#0065F# => romdata <= X"152254FF";
    when 16#00660# => romdata <= X"A1398170";
    when 16#00661# => romdata <= X"902B7090";
    when 16#00662# => romdata <= X"2C405754";
    when 16#00663# => romdata <= X"80705D58";
    when 16#00664# => romdata <= X"FCA63974";
    when 16#00665# => romdata <= X"2254FCDC";
    when 16#00666# => romdata <= X"39FA3D0D";
    when 16#00667# => romdata <= X"8A5180C3";
    when 16#00668# => romdata <= X"D73F97C8";
    when 16#00669# => romdata <= X"3F9A8553";
    when 16#0066A# => romdata <= X"81B2F852";
    when 16#0066B# => romdata <= X"81B38C51";
    when 16#0066C# => romdata <= X"97CD3FA3";
    when 16#0066D# => romdata <= X"EF5381B3";
    when 16#0066E# => romdata <= X"905281B3";
    when 16#0066F# => romdata <= X"B85197BF";
    when 16#00670# => romdata <= X"3FBBEA53";
    when 16#00671# => romdata <= X"81B3C052";
    when 16#00672# => romdata <= X"81B3D051";
    when 16#00673# => romdata <= X"97B13FBB";
    when 16#00674# => romdata <= X"D15381B3";
    when 16#00675# => romdata <= X"D85281B3";
    when 16#00676# => romdata <= X"F45197A3";
    when 16#00677# => romdata <= X"3FA6A953";
    when 16#00678# => romdata <= X"81B3FC52";
    when 16#00679# => romdata <= X"81B4A051";
    when 16#0067A# => romdata <= X"97953FBE";
    when 16#0067B# => romdata <= X"AD5381B4";
    when 16#0067C# => romdata <= X"A85281B4";
    when 16#0067D# => romdata <= X"C8519787";
    when 16#0067E# => romdata <= X"3FBFCB53";
    when 16#0067F# => romdata <= X"81B4CC52";
    when 16#00680# => romdata <= X"81B4F051";
    when 16#00681# => romdata <= X"96F93FBC";
    when 16#00682# => romdata <= X"815381B4";
    when 16#00683# => romdata <= X"F85281B0";
    when 16#00684# => romdata <= X"905196EB";
    when 16#00685# => romdata <= X"3FBCC253";
    when 16#00686# => romdata <= X"81B59C52";
    when 16#00687# => romdata <= X"81B5C451";
    when 16#00688# => romdata <= X"96DD3FBD";
    when 16#00689# => romdata <= X"EA5381B5";
    when 16#0068A# => romdata <= X"CC5281B5";
    when 16#0068B# => romdata <= X"EC5196CF";
    when 16#0068C# => romdata <= X"3F889B53";
    when 16#0068D# => romdata <= X"81B5F452";
    when 16#0068E# => romdata <= X"81B69051";
    when 16#0068F# => romdata <= X"96C13FA4";
    when 16#00690# => romdata <= X"BF5381B6";
    when 16#00691# => romdata <= X"985281B5";
    when 16#00692# => romdata <= X"E45196B3";
    when 16#00693# => romdata <= X"3FA48B53";
    when 16#00694# => romdata <= X"81B6B452";
    when 16#00695# => romdata <= X"81B6C851";
    when 16#00696# => romdata <= X"96A53FB9";
    when 16#00697# => romdata <= X"905381B6";
    when 16#00698# => romdata <= X"D05281B6";
    when 16#00699# => romdata <= X"EC519697";
    when 16#0069A# => romdata <= X"3FB9B653";
    when 16#0069B# => romdata <= X"81B6F452";
    when 16#0069C# => romdata <= X"81B78851";
    when 16#0069D# => romdata <= X"96893FA7";
    when 16#0069E# => romdata <= X"CB5381B7";
    when 16#0069F# => romdata <= X"905281B7";
    when 16#006A0# => romdata <= X"B45195FB";
    when 16#006A1# => romdata <= X"3F80C0A9";
    when 16#006A2# => romdata <= X"5381B7BC";
    when 16#006A3# => romdata <= X"5281B7CC";
    when 16#006A4# => romdata <= X"5195EC3F";
    when 16#006A5# => romdata <= X"80C2F453";
    when 16#006A6# => romdata <= X"81B7D052";
    when 16#006A7# => romdata <= X"81B7EC51";
    when 16#006A8# => romdata <= X"95DD3FBB";
    when 16#006A9# => romdata <= X"975381B7";
    when 16#006AA# => romdata <= X"F45281B8";
    when 16#006AB# => romdata <= X"8C5195CF";
    when 16#006AC# => romdata <= X"3F80C2FC";
    when 16#006AD# => romdata <= X"5381B894";
    when 16#006AE# => romdata <= X"5281B8A8";
    when 16#006AF# => romdata <= X"5195C03F";
    when 16#006B0# => romdata <= X"8AD65381";
    when 16#006B1# => romdata <= X"B8B05281";
    when 16#006B2# => romdata <= X"B8C45195";
    when 16#006B3# => romdata <= X"B23F8DE6";
    when 16#006B4# => romdata <= X"5381B8C8";
    when 16#006B5# => romdata <= X"5281B8F0";
    when 16#006B6# => romdata <= X"5195A43F";
    when 16#006B7# => romdata <= X"BBB35381";
    when 16#006B8# => romdata <= X"B8F85281";
    when 16#006B9# => romdata <= X"B9985195";
    when 16#006BA# => romdata <= X"963F93A3";
    when 16#006BB# => romdata <= X"5381B9A0";
    when 16#006BC# => romdata <= X"5281B9B4";
    when 16#006BD# => romdata <= X"5195883F";
    when 16#006BE# => romdata <= X"88BE5381";
    when 16#006BF# => romdata <= X"B9BC5281";
    when 16#006C0# => romdata <= X"B9C85194";
    when 16#006C1# => romdata <= X"FA3F89FC";
    when 16#006C2# => romdata <= X"5381B9CC";
    when 16#006C3# => romdata <= X"5281B9F4";
    when 16#006C4# => romdata <= X"5194EC3F";
    when 16#006C5# => romdata <= X"88BE5381";
    when 16#006C6# => romdata <= X"B9FC5281";
    when 16#006C7# => romdata <= X"B2B05194";
    when 16#006C8# => romdata <= X"DE3F8AC5";
    when 16#006C9# => romdata <= X"5381BA9C";
    when 16#006CA# => romdata <= X"5281BAAC";
    when 16#006CB# => romdata <= X"5194D03F";
    when 16#006CC# => romdata <= X"88B35381";
    when 16#006CD# => romdata <= X"A5BC5281";
    when 16#006CE# => romdata <= X"A5A05194";
    when 16#006CF# => romdata <= X"C23F80D1";
    when 16#006D0# => romdata <= X"D55381A5";
    when 16#006D1# => romdata <= X"BC5281A5";
    when 16#006D2# => romdata <= X"A85194B3";
    when 16#006D3# => romdata <= X"3F9B863F";
    when 16#006D4# => romdata <= X"94F93F81";
    when 16#006D5# => romdata <= X"0B81EFF8";
    when 16#006D6# => romdata <= X"3481DCD8";
    when 16#006D7# => romdata <= X"337081FF";
    when 16#006D8# => romdata <= X"06555573";
    when 16#006D9# => romdata <= X"B23880C4";
    when 16#006DA# => romdata <= X"9B3FB008";
    when 16#006DB# => romdata <= X"903894E9";
    when 16#006DC# => romdata <= X"3F81EFF8";
    when 16#006DD# => romdata <= X"335675E1";
    when 16#006DE# => romdata <= X"38883D0D";
    when 16#006DF# => romdata <= X"0480C497";
    when 16#006E0# => romdata <= X"3FB00881";
    when 16#006E1# => romdata <= X"FF065195";
    when 16#006E2# => romdata <= X"BE3F94CD";
    when 16#006E3# => romdata <= X"3F81EFF8";
    when 16#006E4# => romdata <= X"335675C5";
    when 16#006E5# => romdata <= X"38E33980";
    when 16#006E6# => romdata <= X"0B81DCD8";
    when 16#006E7# => romdata <= X"349BD63F";
    when 16#006E8# => romdata <= X"81CCFC08";
    when 16#006E9# => romdata <= X"70087087";
    when 16#006EA# => romdata <= X"2A810652";
    when 16#006EB# => romdata <= X"57547380";
    when 16#006EC# => romdata <= X"2E8F3876";
    when 16#006ED# => romdata <= X"802E81C5";
    when 16#006EE# => romdata <= X"38FF1770";
    when 16#006EF# => romdata <= X"81FF0658";
    when 16#006F0# => romdata <= X"5475862A";
    when 16#006F1# => romdata <= X"81065574";
    when 16#006F2# => romdata <= X"802EAA38";
    when 16#006F3# => romdata <= X"7680F738";
    when 16#006F4# => romdata <= X"81960B81";
    when 16#006F5# => romdata <= X"CCFC0884";
    when 16#006F6# => romdata <= X"110870EF";
    when 16#006F7# => romdata <= X"FF0A06AE";
    when 16#006F8# => romdata <= X"800A0784";
    when 16#006F9# => romdata <= X"130C5784";
    when 16#006FA# => romdata <= X"110870BE";
    when 16#006FB# => romdata <= X"800A0784";
    when 16#006FC# => romdata <= X"130C5755";
    when 16#006FD# => romdata <= X"5775852A";
    when 16#006FE# => romdata <= X"81065574";
    when 16#006FF# => romdata <= X"802E9638";
    when 16#00700# => romdata <= X"76BA3881";
    when 16#00701# => romdata <= X"960B81CC";
    when 16#00702# => romdata <= X"C408B811";
    when 16#00703# => romdata <= X"08575557";
    when 16#00704# => romdata <= X"800BB815";
    when 16#00705# => romdata <= X"0C75842A";
    when 16#00706# => romdata <= X"81065675";
    when 16#00707# => romdata <= X"802EFEC6";
    when 16#00708# => romdata <= X"3876802E";
    when 16#00709# => romdata <= X"AC38FF17";
    when 16#0070A# => romdata <= X"7081FF06";
    when 16#0070B# => romdata <= X"585580C2";
    when 16#0070C# => romdata <= X"D33FB008";
    when 16#0070D# => romdata <= X"802EFEB6";
    when 16#0070E# => romdata <= X"38FEC239";
    when 16#0070F# => romdata <= X"FF177081";
    when 16#00710# => romdata <= X"FF065855";
    when 16#00711# => romdata <= X"D039FF17";
    when 16#00712# => romdata <= X"7081FF06";
    when 16#00713# => romdata <= X"5854FFA5";
    when 16#00714# => romdata <= X"3981960B";
    when 16#00715# => romdata <= X"81CCFC08";
    when 16#00716# => romdata <= X"84110884";
    when 16#00717# => romdata <= X"0A078412";
    when 16#00718# => romdata <= X"0C5657A6";
    when 16#00719# => romdata <= X"CE3F8052";
    when 16#0071A# => romdata <= X"81C19C51";
    when 16#0071B# => romdata <= X"A9983F80";
    when 16#0071C# => romdata <= X"C2923FB0";
    when 16#0071D# => romdata <= X"08802EFD";
    when 16#0071E# => romdata <= X"F538FE81";
    when 16#0071F# => romdata <= X"39819676";
    when 16#00720# => romdata <= X"822A8306";
    when 16#00721# => romdata <= X"53768306";
    when 16#00722# => romdata <= X"5257F4D3";
    when 16#00723# => romdata <= X"3FFEB239";
    when 16#00724# => romdata <= X"FE3D0D81";
    when 16#00725# => romdata <= X"5195DA3F";
    when 16#00726# => romdata <= X"B00881FF";
    when 16#00727# => romdata <= X"06538251";
    when 16#00728# => romdata <= X"95CF3FB0";
    when 16#00729# => romdata <= X"0881FF06";
    when 16#0072A# => romdata <= X"527251F4";
    when 16#0072B# => romdata <= X"B23F800B";
    when 16#0072C# => romdata <= X"B00C843D";
    when 16#0072D# => romdata <= X"0D04F93D";
    when 16#0072E# => romdata <= X"0D815195";
    when 16#0072F# => romdata <= X"B43FB008";
    when 16#00730# => romdata <= X"81FF0681";
    when 16#00731# => romdata <= X"BAB45257";
    when 16#00732# => romdata <= X"BDC83F81";
    when 16#00733# => romdata <= X"BAC851BD";
    when 16#00734# => romdata <= X"C13FF880";
    when 16#00735# => romdata <= X"809A8054";
    when 16#00736# => romdata <= X"80557370";
    when 16#00737# => romdata <= X"84055508";
    when 16#00738# => romdata <= X"74708405";
    when 16#00739# => romdata <= X"56085456";
    when 16#0073A# => romdata <= X"72A03881";
    when 16#0073B# => romdata <= X"157081FF";
    when 16#0073C# => romdata <= X"06565687";
    when 16#0073D# => romdata <= X"7527E338";
    when 16#0073E# => romdata <= X"76812E80";
    when 16#0073F# => romdata <= X"D8388A51";
    when 16#00740# => romdata <= X"BCF63F76";
    when 16#00741# => romdata <= X"B00C893D";
    when 16#00742# => romdata <= X"0D048A51";
    when 16#00743# => romdata <= X"BCEA3F72";
    when 16#00744# => romdata <= X"51BEC93F";
    when 16#00745# => romdata <= X"B00881FF";
    when 16#00746# => romdata <= X"0653728C";
    when 16#00747# => romdata <= X"279338A0";
    when 16#00748# => romdata <= X"51BCD53F";
    when 16#00749# => romdata <= X"81137081";
    when 16#0074A# => romdata <= X"FF065153";
    when 16#0074B# => romdata <= X"8C7326EF";
    when 16#0074C# => romdata <= X"3881BAE0";
    when 16#0074D# => romdata <= X"51BCDB3F";
    when 16#0074E# => romdata <= X"7552A051";
    when 16#0074F# => romdata <= X"BCF73F75";
    when 16#00750# => romdata <= X"51D9C23F";
    when 16#00751# => romdata <= X"81157081";
    when 16#00752# => romdata <= X"FF065656";
    when 16#00753# => romdata <= X"877527FF";
    when 16#00754# => romdata <= X"8938FFA4";
    when 16#00755# => romdata <= X"39F88080";
    when 16#00756# => romdata <= X"9A805480";
    when 16#00757# => romdata <= X"53807470";
    when 16#00758# => romdata <= X"8405560C";
    when 16#00759# => romdata <= X"80747084";
    when 16#0075A# => romdata <= X"05560C81";
    when 16#0075B# => romdata <= X"137081FF";
    when 16#0075C# => romdata <= X"06545572";
    when 16#0075D# => romdata <= X"8726FF86";
    when 16#0075E# => romdata <= X"38807470";
    when 16#0075F# => romdata <= X"8405560C";
    when 16#00760# => romdata <= X"80747084";
    when 16#00761# => romdata <= X"05560C81";
    when 16#00762# => romdata <= X"137081FF";
    when 16#00763# => romdata <= X"06545587";
    when 16#00764# => romdata <= X"7327CA38";
    when 16#00765# => romdata <= X"FEE839FE";
    when 16#00766# => romdata <= X"3D0D8151";
    when 16#00767# => romdata <= X"93D33FB0";
    when 16#00768# => romdata <= X"0881FF06";
    when 16#00769# => romdata <= X"81CCBC08";
    when 16#0076A# => romdata <= X"7188120C";
    when 16#0076B# => romdata <= X"53B00C84";
    when 16#0076C# => romdata <= X"3D0D0480";
    when 16#0076D# => romdata <= X"3D0D8151";
    when 16#0076E# => romdata <= X"94E93FB0";
    when 16#0076F# => romdata <= X"0883FFFF";
    when 16#00770# => romdata <= X"0651D2EF";
    when 16#00771# => romdata <= X"3FB00883";
    when 16#00772# => romdata <= X"FFFF06B0";
    when 16#00773# => romdata <= X"0C823D0D";
    when 16#00774# => romdata <= X"04803D0D";
    when 16#00775# => romdata <= X"81519399";
    when 16#00776# => romdata <= X"3FB00881";
    when 16#00777# => romdata <= X"FF06519E";
    when 16#00778# => romdata <= X"A83F800B";
    when 16#00779# => romdata <= X"B00C823D";
    when 16#0077A# => romdata <= X"0D04803D";
    when 16#0077B# => romdata <= X"0D81CD88";
    when 16#0077C# => romdata <= X"0851F8BB";
    when 16#0077D# => romdata <= X"9586A171";
    when 16#0077E# => romdata <= X"0C810BB0";
    when 16#0077F# => romdata <= X"0C823D0D";
    when 16#00780# => romdata <= X"04FC3D0D";
    when 16#00781# => romdata <= X"815192E9";
    when 16#00782# => romdata <= X"3FB00881";
    when 16#00783# => romdata <= X"FF065482";
    when 16#00784# => romdata <= X"5192DE3F";
    when 16#00785# => romdata <= X"B00881FF";
    when 16#00786# => romdata <= X"0681CCFC";
    when 16#00787# => romdata <= X"08841108";
    when 16#00788# => romdata <= X"70FE8F0A";
    when 16#00789# => romdata <= X"0677982B";
    when 16#0078A# => romdata <= X"07515456";
    when 16#0078B# => romdata <= X"5372802E";
    when 16#0078C# => romdata <= X"86387181";
    when 16#0078D# => romdata <= X"0A075271";
    when 16#0078E# => romdata <= X"84160C71";
    when 16#0078F# => romdata <= X"B00C863D";
    when 16#00790# => romdata <= X"0D04FD3D";
    when 16#00791# => romdata <= X"0D81CCFC";
    when 16#00792# => romdata <= X"08841108";
    when 16#00793# => romdata <= X"55538151";
    when 16#00794# => romdata <= X"929F3FB0";
    when 16#00795# => romdata <= X"0881FF06";
    when 16#00796# => romdata <= X"74DFFFFF";
    when 16#00797# => romdata <= X"06545271";
    when 16#00798# => romdata <= X"802E8738";
    when 16#00799# => romdata <= X"73A08080";
    when 16#0079A# => romdata <= X"07538251";
    when 16#0079B# => romdata <= X"92833FB0";
    when 16#0079C# => romdata <= X"0881FF06";
    when 16#0079D# => romdata <= X"73EFFF0A";
    when 16#0079E# => romdata <= X"06555271";
    when 16#0079F# => romdata <= X"802E8738";
    when 16#007A0# => romdata <= X"7290800A";
    when 16#007A1# => romdata <= X"07548351";
    when 16#007A2# => romdata <= X"91E73FB0";
    when 16#007A3# => romdata <= X"0881FF06";
    when 16#007A4# => romdata <= X"74F7FF0A";
    when 16#007A5# => romdata <= X"06545271";
    when 16#007A6# => romdata <= X"802E8738";
    when 16#007A7# => romdata <= X"7388800A";
    when 16#007A8# => romdata <= X"07538451";
    when 16#007A9# => romdata <= X"91CB3FB0";
    when 16#007AA# => romdata <= X"0881FF06";
    when 16#007AB# => romdata <= X"73FBFF0A";
    when 16#007AC# => romdata <= X"06555271";
    when 16#007AD# => romdata <= X"802E8738";
    when 16#007AE# => romdata <= X"7284800A";
    when 16#007AF# => romdata <= X"07548551";
    when 16#007B0# => romdata <= X"91AF3FB0";
    when 16#007B1# => romdata <= X"0881FF06";
    when 16#007B2# => romdata <= X"74FDFF0A";
    when 16#007B3# => romdata <= X"06545271";
    when 16#007B4# => romdata <= X"802E8738";
    when 16#007B5# => romdata <= X"7382800A";
    when 16#007B6# => romdata <= X"075381CC";
    when 16#007B7# => romdata <= X"FC087384";
    when 16#007B8# => romdata <= X"120C5472";
    when 16#007B9# => romdata <= X"B00C853D";
    when 16#007BA# => romdata <= X"0D04FA3D";
    when 16#007BB# => romdata <= X"0D880A0B";
    when 16#007BC# => romdata <= X"81CCC008";
    when 16#007BD# => romdata <= X"8C110859";
    when 16#007BE# => romdata <= X"55568151";
    when 16#007BF# => romdata <= X"90F33FB0";
    when 16#007C0# => romdata <= X"08902B70";
    when 16#007C1# => romdata <= X"902C5653";
    when 16#007C2# => romdata <= X"80772799";
    when 16#007C3# => romdata <= X"38807754";
    when 16#007C4# => romdata <= X"547383FF";
    when 16#007C5# => romdata <= X"FF067670";
    when 16#007C6# => romdata <= X"8405580C";
    when 16#007C7# => romdata <= X"FF137515";
    when 16#007C8# => romdata <= X"555372ED";
    when 16#007C9# => romdata <= X"38800BB0";
    when 16#007CA# => romdata <= X"0C883D0D";
    when 16#007CB# => romdata <= X"04FC3D0D";
    when 16#007CC# => romdata <= X"81BAE851";
    when 16#007CD# => romdata <= X"B8DC3F81";
    when 16#007CE# => romdata <= X"CCFC0870";
    when 16#007CF# => romdata <= X"08709E2A";
    when 16#007D0# => romdata <= X"70810651";
    when 16#007D1# => romdata <= X"54545481";
    when 16#007D2# => romdata <= X"53718338";
    when 16#007D3# => romdata <= X"71537280";
    when 16#007D4# => romdata <= X"2E80D238";
    when 16#007D5# => romdata <= X"81BAF851";
    when 16#007D6# => romdata <= X"B8B83F81";
    when 16#007D7# => romdata <= X"5190923F";
    when 16#007D8# => romdata <= X"B00881FF";
    when 16#007D9# => romdata <= X"0681BAE8";
    when 16#007DA# => romdata <= X"5255B8A6";
    when 16#007DB# => romdata <= X"3F74802E";
    when 16#007DC# => romdata <= X"AB3881BB";
    when 16#007DD# => romdata <= X"8051B89A";
    when 16#007DE# => romdata <= X"3F81CCFC";
    when 16#007DF# => romdata <= X"08841108";
    when 16#007E0# => romdata <= X"70FD0A06";
    when 16#007E1# => romdata <= X"54545474";
    when 16#007E2# => romdata <= X"802E8638";
    when 16#007E3# => romdata <= X"72820A07";
    when 16#007E4# => romdata <= X"52718415";
    when 16#007E5# => romdata <= X"0C71B00C";
    when 16#007E6# => romdata <= X"863D0D04";
    when 16#007E7# => romdata <= X"81B09851";
    when 16#007E8# => romdata <= X"B7F03FCE";
    when 16#007E9# => romdata <= X"3981B098";
    when 16#007EA# => romdata <= X"51B7E73F";
    when 16#007EB# => romdata <= X"81BAF851";
    when 16#007EC# => romdata <= X"B7E03F81";
    when 16#007ED# => romdata <= X"518FBA3F";
    when 16#007EE# => romdata <= X"B00881FF";
    when 16#007EF# => romdata <= X"0681BAE8";
    when 16#007F0# => romdata <= X"5255B7CE";
    when 16#007F1# => romdata <= X"3F74FFAA";
    when 16#007F2# => romdata <= X"38D239FD";
    when 16#007F3# => romdata <= X"3D0D8151";
    when 16#007F4# => romdata <= X"8F9F3FB0";
    when 16#007F5# => romdata <= X"0881FF06";
    when 16#007F6# => romdata <= X"81BB8C52";
    when 16#007F7# => romdata <= X"54B7B33F";
    when 16#007F8# => romdata <= X"73A43881";
    when 16#007F9# => romdata <= X"B09051B7";
    when 16#007FA# => romdata <= X"A93F81CC";
    when 16#007FB# => romdata <= X"FC088411";
    when 16#007FC# => romdata <= X"0870FB0A";
    when 16#007FD# => romdata <= X"0684130C";
    when 16#007FE# => romdata <= X"53538A51";
    when 16#007FF# => romdata <= X"B6FA3F73";
    when 16#00800# => romdata <= X"B00C853D";
    when 16#00801# => romdata <= X"0D0481AC";
    when 16#00802# => romdata <= X"B851B786";
    when 16#00803# => romdata <= X"3F81CCFC";
    when 16#00804# => romdata <= X"08841108";
    when 16#00805# => romdata <= X"70840A07";
    when 16#00806# => romdata <= X"84130C53";
    when 16#00807# => romdata <= X"538A51B6";
    when 16#00808# => romdata <= X"D73F73B0";
    when 16#00809# => romdata <= X"0C853D0D";
    when 16#0080A# => romdata <= X"04FD3D0D";
    when 16#0080B# => romdata <= X"81DCD408";
    when 16#0080C# => romdata <= X"52F881C0";
    when 16#0080D# => romdata <= X"8E800B81";
    when 16#0080E# => romdata <= X"CCFC0855";
    when 16#0080F# => romdata <= X"5371802E";
    when 16#00810# => romdata <= X"80F73872";
    when 16#00811# => romdata <= X"81FF0684";
    when 16#00812# => romdata <= X"150C81CC";
    when 16#00813# => romdata <= X"B8337081";
    when 16#00814# => romdata <= X"FF065152";
    when 16#00815# => romdata <= X"71802E80";
    when 16#00816# => romdata <= X"C238729F";
    when 16#00817# => romdata <= X"2A731007";
    when 16#00818# => romdata <= X"5381DCD8";
    when 16#00819# => romdata <= X"337081FF";
    when 16#0081A# => romdata <= X"06515271";
    when 16#0081B# => romdata <= X"802ED438";
    when 16#0081C# => romdata <= X"800B81DC";
    when 16#0081D# => romdata <= X"D83491FD";
    when 16#0081E# => romdata <= X"3F81CCC8";
    when 16#0081F# => romdata <= X"33547380";
    when 16#00820# => romdata <= X"E23881CC";
    when 16#00821# => romdata <= X"FC087381";
    when 16#00822# => romdata <= X"FF068412";
    when 16#00823# => romdata <= X"0C81CCB8";
    when 16#00824# => romdata <= X"337081FF";
    when 16#00825# => romdata <= X"06515354";
    when 16#00826# => romdata <= X"71C03872";
    when 16#00827# => romdata <= X"812A739F";
    when 16#00828# => romdata <= X"2B0753FF";
    when 16#00829# => romdata <= X"BC397281";
    when 16#0082A# => romdata <= X"2A739F2B";
    when 16#0082B# => romdata <= X"075380FD";
    when 16#0082C# => romdata <= X"51B8F23F";
    when 16#0082D# => romdata <= X"81CCFC08";
    when 16#0082E# => romdata <= X"547281FF";
    when 16#0082F# => romdata <= X"0684150C";
    when 16#00830# => romdata <= X"81CCB833";
    when 16#00831# => romdata <= X"7081FF06";
    when 16#00832# => romdata <= X"53547180";
    when 16#00833# => romdata <= X"2ED83872";
    when 16#00834# => romdata <= X"9F2A7310";
    when 16#00835# => romdata <= X"075380FD";
    when 16#00836# => romdata <= X"51B8CA3F";
    when 16#00837# => romdata <= X"81CCFC08";
    when 16#00838# => romdata <= X"54D73980";
    when 16#00839# => romdata <= X"0BB00C85";
    when 16#0083A# => romdata <= X"3D0D04F7";
    when 16#0083B# => romdata <= X"3D0D853D";
    when 16#0083C# => romdata <= X"54965381";
    when 16#0083D# => romdata <= X"BBA05273";
    when 16#0083E# => romdata <= X"51BBE83F";
    when 16#0083F# => romdata <= X"9EA63F81";
    when 16#00840# => romdata <= X"518CEE3F";
    when 16#00841# => romdata <= X"80528051";
    when 16#00842# => romdata <= X"9C863F73";
    when 16#00843# => romdata <= X"53805281";
    when 16#00844# => romdata <= X"C19C51B0";
    when 16#00845# => romdata <= X"C53F8052";
    when 16#00846# => romdata <= X"81519BF4";
    when 16#00847# => romdata <= X"3F735382";
    when 16#00848# => romdata <= X"5281C19C";
    when 16#00849# => romdata <= X"51B0B33F";
    when 16#0084A# => romdata <= X"80528251";
    when 16#0084B# => romdata <= X"9BE23F73";
    when 16#0084C# => romdata <= X"53815281";
    when 16#0084D# => romdata <= X"C19C51B0";
    when 16#0084E# => romdata <= X"A13F8052";
    when 16#0084F# => romdata <= X"84519BD0";
    when 16#00850# => romdata <= X"3F735384";
    when 16#00851# => romdata <= X"5281C19C";
    when 16#00852# => romdata <= X"51B08F3F";
    when 16#00853# => romdata <= X"80528551";
    when 16#00854# => romdata <= X"9BBE3F73";
    when 16#00855# => romdata <= X"53905281";
    when 16#00856# => romdata <= X"C19C51AF";
    when 16#00857# => romdata <= X"FD3F8052";
    when 16#00858# => romdata <= X"86519BAC";
    when 16#00859# => romdata <= X"3F735383";
    when 16#0085A# => romdata <= X"5281C19C";
    when 16#0085B# => romdata <= X"51AFEB3F";
    when 16#0085C# => romdata <= X"8B3D0D04";
    when 16#0085D# => romdata <= X"FEF53F80";
    when 16#0085E# => romdata <= X"0BB00C04";
    when 16#0085F# => romdata <= X"FC3D0D81";
    when 16#00860# => romdata <= X"9FB85480";
    when 16#00861# => romdata <= X"55845274";
    when 16#00862# => romdata <= X"519B853F";
    when 16#00863# => romdata <= X"80537370";
    when 16#00864# => romdata <= X"81055533";
    when 16#00865# => romdata <= X"519BFF3F";
    when 16#00866# => romdata <= X"81137081";
    when 16#00867# => romdata <= X"FF065153";
    when 16#00868# => romdata <= X"80DC7327";
    when 16#00869# => romdata <= X"E9388115";
    when 16#0086A# => romdata <= X"7081FF06";
    when 16#0086B# => romdata <= X"56538775";
    when 16#0086C# => romdata <= X"27D33880";
    when 16#0086D# => romdata <= X"0BB00C86";
    when 16#0086E# => romdata <= X"3D0D04FD";
    when 16#0086F# => romdata <= X"3D0D81CC";
    when 16#00870# => romdata <= X"B8337081";
    when 16#00871# => romdata <= X"FF065454";
    when 16#00872# => romdata <= X"72BF26AC";
    when 16#00873# => romdata <= X"3881CCB8";
    when 16#00874# => romdata <= X"337081FF";
    when 16#00875# => romdata <= X"0681CCBC";
    when 16#00876# => romdata <= X"08528812";
    when 16#00877# => romdata <= X"0C5480E4";
    when 16#00878# => romdata <= X"5280C3BB";
    when 16#00879# => romdata <= X"518FEE3F";
    when 16#0087A# => romdata <= X"81CCB833";
    when 16#0087B# => romdata <= X"81055372";
    when 16#0087C# => romdata <= X"81CCB834";
    when 16#0087D# => romdata <= X"853D0D04";
    when 16#0087E# => romdata <= X"80E45280";
    when 16#0087F# => romdata <= X"C492518F";
    when 16#00880# => romdata <= X"D43F81CC";
    when 16#00881# => romdata <= X"B8338105";
    when 16#00882# => romdata <= X"537281CC";
    when 16#00883# => romdata <= X"B834853D";
    when 16#00884# => romdata <= X"0D04FD3D";
    when 16#00885# => romdata <= X"0D81CCB8";
    when 16#00886# => romdata <= X"337081FF";
    when 16#00887# => romdata <= X"06545472";
    when 16#00888# => romdata <= X"BF2680C9";
    when 16#00889# => romdata <= X"3881CCB8";
    when 16#0088A# => romdata <= X"337081FF";
    when 16#0088B# => romdata <= X"0681CCBC";
    when 16#0088C# => romdata <= X"08568816";
    when 16#0088D# => romdata <= X"0C5381CC";
    when 16#0088E# => romdata <= X"B8337081";
    when 16#0088F# => romdata <= X"FF065553";
    when 16#00890# => romdata <= X"73BF2E80";
    when 16#00891# => romdata <= X"D13880E4";
    when 16#00892# => romdata <= X"5280C492";
    when 16#00893# => romdata <= X"518F863F";
    when 16#00894# => romdata <= X"81CCB833";
    when 16#00895# => romdata <= X"81055372";
    when 16#00896# => romdata <= X"81CCB834";
    when 16#00897# => romdata <= X"81CCB833";
    when 16#00898# => romdata <= X"80FF0653";
    when 16#00899# => romdata <= X"7281CCB8";
    when 16#0089A# => romdata <= X"34853D0D";
    when 16#0089B# => romdata <= X"0481CCB8";
    when 16#0089C# => romdata <= X"337081FF";
    when 16#0089D# => romdata <= X"0680FF71";
    when 16#0089E# => romdata <= X"3181CCBC";
    when 16#0089F# => romdata <= X"08528812";
    when 16#008A0# => romdata <= X"0C555381";
    when 16#008A1# => romdata <= X"CCB83370";
    when 16#008A2# => romdata <= X"81FF0655";
    when 16#008A3# => romdata <= X"5373BF2E";
    when 16#008A4# => romdata <= X"098106FF";
    when 16#008A5# => romdata <= X"B13880CE";
    when 16#008A6# => romdata <= X"905280C4";
    when 16#008A7# => romdata <= X"92518EB5";
    when 16#008A8# => romdata <= X"3F81CCB8";
    when 16#008A9# => romdata <= X"33810553";
    when 16#008AA# => romdata <= X"7281CCB8";
    when 16#008AB# => romdata <= X"3481CCB8";
    when 16#008AC# => romdata <= X"3380FF06";
    when 16#008AD# => romdata <= X"537281CC";
    when 16#008AE# => romdata <= X"B834853D";
    when 16#008AF# => romdata <= X"0D04810B";
    when 16#008B0# => romdata <= X"81CCC834";
    when 16#008B1# => romdata <= X"04FE3D0D";
    when 16#008B2# => romdata <= X"81CD8008";
    when 16#008B3# => romdata <= X"98110870";
    when 16#008B4# => romdata <= X"842A7081";
    when 16#008B5# => romdata <= X"06515353";
    when 16#008B6# => romdata <= X"5370802E";
    when 16#008B7# => romdata <= X"8D3871EF";
    when 16#008B8# => romdata <= X"0698140C";
    when 16#008B9# => romdata <= X"810B81DC";
    when 16#008BA# => romdata <= X"D834843D";
    when 16#008BB# => romdata <= X"0D04FB3D";
    when 16#008BC# => romdata <= X"0D81CCFC";
    when 16#008BD# => romdata <= X"08700881";
    when 16#008BE# => romdata <= X"0A0681DC";
    when 16#008BF# => romdata <= X"D40C54B4";
    when 16#008C0# => romdata <= X"C73FB4EA";
    when 16#008C1# => romdata <= X"3F8F8B3F";
    when 16#008C2# => romdata <= X"81CD8008";
    when 16#008C3# => romdata <= X"98110888";
    when 16#008C4# => romdata <= X"0798120C";
    when 16#008C5# => romdata <= X"5481DCD4";
    when 16#008C6# => romdata <= X"0880F6E2";
    when 16#008C7# => romdata <= X"55537284";
    when 16#008C8# => romdata <= X"38888054";
    when 16#008C9# => romdata <= X"7381F0DC";
    when 16#008CA# => romdata <= X"0C72802E";
    when 16#008CB# => romdata <= X"84B03881";
    when 16#008CC# => romdata <= X"A68451B0";
    when 16#008CD# => romdata <= X"DD3F8C51";
    when 16#008CE# => romdata <= X"B0BE3F81";
    when 16#008CF# => romdata <= X"BBA051B0";
    when 16#008D0# => romdata <= X"D13F81DC";
    when 16#008D1# => romdata <= X"D408802E";
    when 16#008D2# => romdata <= X"81E83881";
    when 16#008D3# => romdata <= X"BBB851B0";
    when 16#008D4# => romdata <= X"C13F81DC";
    when 16#008D5# => romdata <= X"D4085473";
    when 16#008D6# => romdata <= X"802E82D3";
    when 16#008D7# => romdata <= X"3881CCC0";
    when 16#008D8# => romdata <= X"08548174";
    when 16#008D9# => romdata <= X"0C81CCFC";
    when 16#008DA# => romdata <= X"08841108";
    when 16#008DB# => romdata <= X"70565755";
    when 16#008DC# => romdata <= X"805373FE";
    when 16#008DD# => romdata <= X"8F0A0673";
    when 16#008DE# => romdata <= X"982B0770";
    when 16#008DF# => romdata <= X"84170C81";
    when 16#008E0# => romdata <= X"147081FF";
    when 16#008E1# => romdata <= X"06515454";
    when 16#008E2# => romdata <= X"8F7327E6";
    when 16#008E3# => romdata <= X"38758416";
    when 16#008E4# => romdata <= X"0C81CCC4";
    when 16#008E5# => romdata <= X"0854800B";
    when 16#008E6# => romdata <= X"B8150C80";
    when 16#008E7# => romdata <= X"0BF88080";
    when 16#008E8# => romdata <= X"9E800CA0";
    when 16#008E9# => romdata <= X"808D0A08";
    when 16#008EA# => romdata <= X"51B1B13F";
    when 16#008EB# => romdata <= X"8A51AFC8";
    when 16#008EC# => romdata <= X"3F825280";
    when 16#008ED# => romdata <= X"C5BE518C";
    when 16#008EE# => romdata <= X"9C3FF881";
    when 16#008EF# => romdata <= X"C08E800B";
    when 16#008F0# => romdata <= X"81CCFC08";
    when 16#008F1# => romdata <= X"565481DC";
    when 16#008F2# => romdata <= X"D408802E";
    when 16#008F3# => romdata <= X"81B73873";
    when 16#008F4# => romdata <= X"81FF0684";
    when 16#008F5# => romdata <= X"160C81CC";
    when 16#008F6# => romdata <= X"B8337081";
    when 16#008F7# => romdata <= X"FF065456";
    when 16#008F8# => romdata <= X"72802E80";
    when 16#008F9# => romdata <= X"C238739F";
    when 16#008FA# => romdata <= X"2A741007";
    when 16#008FB# => romdata <= X"5481DCD8";
    when 16#008FC# => romdata <= X"337081FF";
    when 16#008FD# => romdata <= X"06575375";
    when 16#008FE# => romdata <= X"802ED438";
    when 16#008FF# => romdata <= X"800B81DC";
    when 16#00900# => romdata <= X"D8348AF1";
    when 16#00901# => romdata <= X"3F81CCC8";
    when 16#00902# => romdata <= X"33557482";
    when 16#00903# => romdata <= X"DC3881CC";
    when 16#00904# => romdata <= X"FC087481";
    when 16#00905# => romdata <= X"FF068412";
    when 16#00906# => romdata <= X"0C81CCB8";
    when 16#00907# => romdata <= X"337081FF";
    when 16#00908# => romdata <= X"06555755";
    when 16#00909# => romdata <= X"72C03873";
    when 16#0090A# => romdata <= X"812A749F";
    when 16#0090B# => romdata <= X"2B0754FF";
    when 16#0090C# => romdata <= X"BC3981BB";
    when 16#0090D# => romdata <= X"C451AEDA";
    when 16#0090E# => romdata <= X"3F810A51";
    when 16#0090F# => romdata <= X"AED43F81";
    when 16#00910# => romdata <= X"BBD851AE";
    when 16#00911# => romdata <= X"CD3F81BC";
    when 16#00912# => romdata <= X"8051AEC6";
    when 16#00913# => romdata <= X"3FB451B0";
    when 16#00914# => romdata <= X"8B3F81BC";
    when 16#00915# => romdata <= X"9451AEBA";
    when 16#00916# => romdata <= X"3F81BC9C";
    when 16#00917# => romdata <= X"51AEB33F";
    when 16#00918# => romdata <= X"81BCA851";
    when 16#00919# => romdata <= X"AEAC3F81";
    when 16#0091A# => romdata <= X"DCD40854";
    when 16#0091B# => romdata <= X"73FDEE38";
    when 16#0091C# => romdata <= X"BE397381";
    when 16#0091D# => romdata <= X"2A749F2B";
    when 16#0091E# => romdata <= X"075480FD";
    when 16#0091F# => romdata <= X"51B1A63F";
    when 16#00920# => romdata <= X"81CCFC08";
    when 16#00921# => romdata <= X"557381FF";
    when 16#00922# => romdata <= X"0684160C";
    when 16#00923# => romdata <= X"81CCB833";
    when 16#00924# => romdata <= X"7081FF06";
    when 16#00925# => romdata <= X"56567480";
    when 16#00926# => romdata <= X"2ED83873";
    when 16#00927# => romdata <= X"9F2A7410";
    when 16#00928# => romdata <= X"075480FD";
    when 16#00929# => romdata <= X"51B0FE3F";
    when 16#0092A# => romdata <= X"81CCFC08";
    when 16#0092B# => romdata <= X"55D73981";
    when 16#0092C# => romdata <= X"CCC40874";
    when 16#0092D# => romdata <= X"B4120C56";
    when 16#0092E# => romdata <= X"818051C4";
    when 16#0092F# => romdata <= X"F63F8280";
    when 16#00930# => romdata <= X"51C4F03F";
    when 16#00931# => romdata <= X"848351C4";
    when 16#00932# => romdata <= X"EA3F86F1";
    when 16#00933# => romdata <= X"51C4E43F";
    when 16#00934# => romdata <= X"888351C4";
    when 16#00935# => romdata <= X"DE3F81CC";
    when 16#00936# => romdata <= X"FC087008";
    when 16#00937# => romdata <= X"709E2A70";
    when 16#00938# => romdata <= X"81065155";
    when 16#00939# => romdata <= X"56548155";
    when 16#0093A# => romdata <= X"72802E80";
    when 16#0093B# => romdata <= X"F7387481";
    when 16#0093C# => romdata <= X"FF068415";
    when 16#0093D# => romdata <= X"0870FD0A";
    when 16#0093E# => romdata <= X"06585653";
    when 16#0093F# => romdata <= X"72802E86";
    when 16#00940# => romdata <= X"3874820A";
    when 16#00941# => romdata <= X"07567584";
    when 16#00942# => romdata <= X"150C8414";
    when 16#00943# => romdata <= X"08BE800A";
    when 16#00944# => romdata <= X"0784150C";
    when 16#00945# => romdata <= X"84140884";
    when 16#00946# => romdata <= X"0A078415";
    when 16#00947# => romdata <= X"0C81CCC4";
    when 16#00948# => romdata <= X"0855800B";
    when 16#00949# => romdata <= X"B8160C81";
    when 16#0094A# => romdata <= X"CCC00854";
    when 16#0094B# => romdata <= X"81740C93";
    when 16#0094C# => romdata <= X"C45280C2";
    when 16#0094D# => romdata <= X"FC51899D";
    when 16#0094E# => romdata <= X"3F87E852";
    when 16#0094F# => romdata <= X"80C3BB51";
    when 16#00950# => romdata <= X"89933FE8";
    when 16#00951# => romdata <= X"D43F81CC";
    when 16#00952# => romdata <= X"C0085481";
    when 16#00953# => romdata <= X"740C81CC";
    when 16#00954# => romdata <= X"FC088411";
    when 16#00955# => romdata <= X"08705657";
    when 16#00956# => romdata <= X"558053FC";
    when 16#00957# => romdata <= X"953995C4";
    when 16#00958# => romdata <= X"3FFBCC39";
    when 16#00959# => romdata <= X"7255FF86";
    when 16#0095A# => romdata <= X"39B2EB3F";
    when 16#0095B# => romdata <= X"800B81EF";
    when 16#0095C# => romdata <= X"F034800B";
    when 16#0095D# => romdata <= X"81EFEC34";
    when 16#0095E# => romdata <= X"800B81EF";
    when 16#0095F# => romdata <= X"F40C04FC";
    when 16#00960# => romdata <= X"3D0D7652";
    when 16#00961# => romdata <= X"81EFEC33";
    when 16#00962# => romdata <= X"70101010";
    when 16#00963# => romdata <= X"71100581";
    when 16#00964# => romdata <= X"DCDC0552";
    when 16#00965# => romdata <= X"54B7DA3F";
    when 16#00966# => romdata <= X"775281EF";
    when 16#00967# => romdata <= X"EC337090";
    when 16#00968# => romdata <= X"29713170";
    when 16#00969# => romdata <= X"101081DF";
    when 16#0096A# => romdata <= X"9C055355";
    when 16#0096B# => romdata <= X"55B7C23F";
    when 16#0096C# => romdata <= X"81EFEC33";
    when 16#0096D# => romdata <= X"70101081";
    when 16#0096E# => romdata <= X"EE9C057A";
    when 16#0096F# => romdata <= X"710C5481";
    when 16#00970# => romdata <= X"05537281";
    when 16#00971# => romdata <= X"EFEC3486";
    when 16#00972# => romdata <= X"3D0D0480";
    when 16#00973# => romdata <= X"3D0D81BC";
    when 16#00974# => romdata <= X"EC51ABBE";
    when 16#00975# => romdata <= X"3F823D0D";
    when 16#00976# => romdata <= X"04FE3D0D";
    when 16#00977# => romdata <= X"81EFF408";
    when 16#00978# => romdata <= X"53728538";
    when 16#00979# => romdata <= X"843D0D04";
    when 16#0097A# => romdata <= X"722DB008";
    when 16#0097B# => romdata <= X"53800B81";
    when 16#0097C# => romdata <= X"EFF40CB0";
    when 16#0097D# => romdata <= X"088C3881";
    when 16#0097E# => romdata <= X"BCEC51AB";
    when 16#0097F# => romdata <= X"953F843D";
    when 16#00980# => romdata <= X"0D0481C0";
    when 16#00981# => romdata <= X"C851AB8A";
    when 16#00982# => romdata <= X"3F7283FF";
    when 16#00983# => romdata <= X"FF26AA38";
    when 16#00984# => romdata <= X"81FF7327";
    when 16#00985# => romdata <= X"96387252";
    when 16#00986# => romdata <= X"9051AB99";
    when 16#00987# => romdata <= X"3F8A51AA";
    when 16#00988# => romdata <= X"D73F81BC";
    when 16#00989# => romdata <= X"EC51AAEA";
    when 16#0098A# => romdata <= X"3FD43972";
    when 16#0098B# => romdata <= X"528851AB";
    when 16#0098C# => romdata <= X"843F8A51";
    when 16#0098D# => romdata <= X"AAC23FEA";
    when 16#0098E# => romdata <= X"397252A0";
    when 16#0098F# => romdata <= X"51AAF63F";
    when 16#00990# => romdata <= X"8A51AAB4";
    when 16#00991# => romdata <= X"3FDC39FA";
    when 16#00992# => romdata <= X"3D0D02A3";
    when 16#00993# => romdata <= X"05335675";
    when 16#00994# => romdata <= X"8D2E80F4";
    when 16#00995# => romdata <= X"38758832";
    when 16#00996# => romdata <= X"70307780";
    when 16#00997# => romdata <= X"FF327030";
    when 16#00998# => romdata <= X"72802571";
    when 16#00999# => romdata <= X"80250754";
    when 16#0099A# => romdata <= X"51565855";
    when 16#0099B# => romdata <= X"7495389F";
    when 16#0099C# => romdata <= X"76278C38";
    when 16#0099D# => romdata <= X"81EFF033";
    when 16#0099E# => romdata <= X"5580CE75";
    when 16#0099F# => romdata <= X"27AE3888";
    when 16#009A0# => romdata <= X"3D0D0481";
    when 16#009A1# => romdata <= X"EFF03356";
    when 16#009A2# => romdata <= X"75802EF3";
    when 16#009A3# => romdata <= X"388851A9";
    when 16#009A4# => romdata <= X"E73FA051";
    when 16#009A5# => romdata <= X"A9E23F88";
    when 16#009A6# => romdata <= X"51A9DD3F";
    when 16#009A7# => romdata <= X"81EFF033";
    when 16#009A8# => romdata <= X"FF055776";
    when 16#009A9# => romdata <= X"81EFF034";
    when 16#009AA# => romdata <= X"883D0D04";
    when 16#009AB# => romdata <= X"7551A9C8";
    when 16#009AC# => romdata <= X"3F81EFF0";
    when 16#009AD# => romdata <= X"33811155";
    when 16#009AE# => romdata <= X"577381EF";
    when 16#009AF# => romdata <= X"F0347581";
    when 16#009B0# => romdata <= X"EF9C1834";
    when 16#009B1# => romdata <= X"883D0D04";
    when 16#009B2# => romdata <= X"8A51A9AC";
    when 16#009B3# => romdata <= X"3F81EFF0";
    when 16#009B4# => romdata <= X"33811156";
    when 16#009B5# => romdata <= X"547481EF";
    when 16#009B6# => romdata <= X"F034800B";
    when 16#009B7# => romdata <= X"81EF9C15";
    when 16#009B8# => romdata <= X"34805680";
    when 16#009B9# => romdata <= X"0B81EF9C";
    when 16#009BA# => romdata <= X"17335654";
    when 16#009BB# => romdata <= X"74A02E83";
    when 16#009BC# => romdata <= X"38815474";
    when 16#009BD# => romdata <= X"802E9038";
    when 16#009BE# => romdata <= X"73802E8B";
    when 16#009BF# => romdata <= X"38811670";
    when 16#009C0# => romdata <= X"81FF0657";
    when 16#009C1# => romdata <= X"57DD3975";
    when 16#009C2# => romdata <= X"802EBF38";
    when 16#009C3# => romdata <= X"800B81EF";
    when 16#009C4# => romdata <= X"EC335555";
    when 16#009C5# => romdata <= X"747427AB";
    when 16#009C6# => romdata <= X"38735774";
    when 16#009C7# => romdata <= X"10101075";
    when 16#009C8# => romdata <= X"10057654";
    when 16#009C9# => romdata <= X"81EF9C53";
    when 16#009CA# => romdata <= X"81DCDC05";
    when 16#009CB# => romdata <= X"51B68E3F";
    when 16#009CC# => romdata <= X"B008802E";
    when 16#009CD# => romdata <= X"A6388115";
    when 16#009CE# => romdata <= X"7081FF06";
    when 16#009CF# => romdata <= X"56547675";
    when 16#009D0# => romdata <= X"26D93881";
    when 16#009D1# => romdata <= X"BCF051A8";
    when 16#009D2# => romdata <= X"C93F81BC";
    when 16#009D3# => romdata <= X"EC51A8C2";
    when 16#009D4# => romdata <= X"3F800B81";
    when 16#009D5# => romdata <= X"EFF03488";
    when 16#009D6# => romdata <= X"3D0D0474";
    when 16#009D7# => romdata <= X"101081EE";
    when 16#009D8# => romdata <= X"9C057008";
    when 16#009D9# => romdata <= X"81EFF40C";
    when 16#009DA# => romdata <= X"56800B81";
    when 16#009DB# => romdata <= X"EFF034E7";
    when 16#009DC# => romdata <= X"39F73D0D";
    when 16#009DD# => romdata <= X"02AF0533";
    when 16#009DE# => romdata <= X"59800B81";
    when 16#009DF# => romdata <= X"EF9C3381";
    when 16#009E0# => romdata <= X"EF9C5955";
    when 16#009E1# => romdata <= X"5673A02E";
    when 16#009E2# => romdata <= X"09810696";
    when 16#009E3# => romdata <= X"38811670";
    when 16#009E4# => romdata <= X"81FF0681";
    when 16#009E5# => romdata <= X"EF9C1170";
    when 16#009E6# => romdata <= X"33535957";
    when 16#009E7# => romdata <= X"5473A02E";
    when 16#009E8# => romdata <= X"EC388058";
    when 16#009E9# => romdata <= X"77792780";
    when 16#009EA# => romdata <= X"EA388077";
    when 16#009EB# => romdata <= X"33565474";
    when 16#009EC# => romdata <= X"742E8338";
    when 16#009ED# => romdata <= X"815474A0";
    when 16#009EE# => romdata <= X"2E9A3873";
    when 16#009EF# => romdata <= X"80C53874";
    when 16#009F0# => romdata <= X"A02E9138";
    when 16#009F1# => romdata <= X"81187081";
    when 16#009F2# => romdata <= X"FF065955";
    when 16#009F3# => romdata <= X"787826DA";
    when 16#009F4# => romdata <= X"3880C039";
    when 16#009F5# => romdata <= X"81167081";
    when 16#009F6# => romdata <= X"FF0681EF";
    when 16#009F7# => romdata <= X"9C117033";
    when 16#009F8# => romdata <= X"57525757";
    when 16#009F9# => romdata <= X"73A02E09";
    when 16#009FA# => romdata <= X"8106D938";
    when 16#009FB# => romdata <= X"81167081";
    when 16#009FC# => romdata <= X"FF0681EF";
    when 16#009FD# => romdata <= X"9C117033";
    when 16#009FE# => romdata <= X"57525757";
    when 16#009FF# => romdata <= X"73A02ED4";
    when 16#00A00# => romdata <= X"38C23981";
    when 16#00A01# => romdata <= X"167081FF";
    when 16#00A02# => romdata <= X"0681EF9C";
    when 16#00A03# => romdata <= X"11595755";
    when 16#00A04# => romdata <= X"FF98398A";
    when 16#00A05# => romdata <= X"538B3DFC";
    when 16#00A06# => romdata <= X"05527651";
    when 16#00A07# => romdata <= X"B8E43F8B";
    when 16#00A08# => romdata <= X"3D0D04F7";
    when 16#00A09# => romdata <= X"3D0D02AF";
    when 16#00A0A# => romdata <= X"05335980";
    when 16#00A0B# => romdata <= X"0B81EF9C";
    when 16#00A0C# => romdata <= X"3381EF9C";
    when 16#00A0D# => romdata <= X"59555673";
    when 16#00A0E# => romdata <= X"A02E0981";
    when 16#00A0F# => romdata <= X"06963881";
    when 16#00A10# => romdata <= X"167081FF";
    when 16#00A11# => romdata <= X"0681EF9C";
    when 16#00A12# => romdata <= X"11703353";
    when 16#00A13# => romdata <= X"59575473";
    when 16#00A14# => romdata <= X"A02EEC38";
    when 16#00A15# => romdata <= X"80587779";
    when 16#00A16# => romdata <= X"2780EA38";
    when 16#00A17# => romdata <= X"80773356";
    when 16#00A18# => romdata <= X"5474742E";
    when 16#00A19# => romdata <= X"83388154";
    when 16#00A1A# => romdata <= X"74A02E9A";
    when 16#00A1B# => romdata <= X"387380C5";
    when 16#00A1C# => romdata <= X"3874A02E";
    when 16#00A1D# => romdata <= X"91388118";
    when 16#00A1E# => romdata <= X"7081FF06";
    when 16#00A1F# => romdata <= X"59557878";
    when 16#00A20# => romdata <= X"26DA3880";
    when 16#00A21# => romdata <= X"C0398116";
    when 16#00A22# => romdata <= X"7081FF06";
    when 16#00A23# => romdata <= X"81EF9C11";
    when 16#00A24# => romdata <= X"70335752";
    when 16#00A25# => romdata <= X"575773A0";
    when 16#00A26# => romdata <= X"2E098106";
    when 16#00A27# => romdata <= X"D9388116";
    when 16#00A28# => romdata <= X"7081FF06";
    when 16#00A29# => romdata <= X"81EF9C11";
    when 16#00A2A# => romdata <= X"70335752";
    when 16#00A2B# => romdata <= X"575773A0";
    when 16#00A2C# => romdata <= X"2ED438C2";
    when 16#00A2D# => romdata <= X"39811670";
    when 16#00A2E# => romdata <= X"81FF0681";
    when 16#00A2F# => romdata <= X"EF9C1159";
    when 16#00A30# => romdata <= X"5755FF98";
    when 16#00A31# => romdata <= X"3990538B";
    when 16#00A32# => romdata <= X"3DFC0552";
    when 16#00A33# => romdata <= X"7651BACF";
    when 16#00A34# => romdata <= X"3F8B3D0D";
    when 16#00A35# => romdata <= X"04FC3D0D";
    when 16#00A36# => romdata <= X"8A51A59C";
    when 16#00A37# => romdata <= X"3F81BD84";
    when 16#00A38# => romdata <= X"51A5AF3F";
    when 16#00A39# => romdata <= X"800B81EF";
    when 16#00A3A# => romdata <= X"EC335353";
    when 16#00A3B# => romdata <= X"72722780";
    when 16#00A3C# => romdata <= X"F5387210";
    when 16#00A3D# => romdata <= X"10107310";
    when 16#00A3E# => romdata <= X"0581DCDC";
    when 16#00A3F# => romdata <= X"05705254";
    when 16#00A40# => romdata <= X"A5903F72";
    when 16#00A41# => romdata <= X"842B7074";
    when 16#00A42# => romdata <= X"31822B81";
    when 16#00A43# => romdata <= X"DF9C1133";
    when 16#00A44# => romdata <= X"51535571";
    when 16#00A45# => romdata <= X"802EB738";
    when 16#00A46# => romdata <= X"7351B1C2";
    when 16#00A47# => romdata <= X"3FB00881";
    when 16#00A48# => romdata <= X"FF065271";
    when 16#00A49# => romdata <= X"89269338";
    when 16#00A4A# => romdata <= X"A051A4CC";
    when 16#00A4B# => romdata <= X"3F811270";
    when 16#00A4C# => romdata <= X"81FF0653";
    when 16#00A4D# => romdata <= X"54897227";
    when 16#00A4E# => romdata <= X"EF3881BD";
    when 16#00A4F# => romdata <= X"9C51A4D2";
    when 16#00A50# => romdata <= X"3F747331";
    when 16#00A51# => romdata <= X"822B81DF";
    when 16#00A52# => romdata <= X"9C0551A4";
    when 16#00A53# => romdata <= X"C53F8A51";
    when 16#00A54# => romdata <= X"A4A63F81";
    when 16#00A55# => romdata <= X"137081FF";
    when 16#00A56# => romdata <= X"0681EFEC";
    when 16#00A57# => romdata <= X"33545455";
    when 16#00A58# => romdata <= X"717326FF";
    when 16#00A59# => romdata <= X"8D388A51";
    when 16#00A5A# => romdata <= X"A48E3F81";
    when 16#00A5B# => romdata <= X"EFEC33B0";
    when 16#00A5C# => romdata <= X"0C863D0D";
    when 16#00A5D# => romdata <= X"04FE3D0D";
    when 16#00A5E# => romdata <= X"81F0CC22";
    when 16#00A5F# => romdata <= X"FF055170";
    when 16#00A60# => romdata <= X"81F0CC23";
    when 16#00A61# => romdata <= X"7083FFFF";
    when 16#00A62# => romdata <= X"06517080";
    when 16#00A63# => romdata <= X"C43881F0";
    when 16#00A64# => romdata <= X"D0335170";
    when 16#00A65# => romdata <= X"81FF2EB9";
    when 16#00A66# => romdata <= X"38701010";
    when 16#00A67# => romdata <= X"1081EFFC";
    when 16#00A68# => romdata <= X"05527133";
    when 16#00A69# => romdata <= X"81F0D034";
    when 16#00A6A# => romdata <= X"FE723481";
    when 16#00A6B# => romdata <= X"F0D03370";
    when 16#00A6C# => romdata <= X"10101081";
    when 16#00A6D# => romdata <= X"EFFC0552";
    when 16#00A6E# => romdata <= X"53821122";
    when 16#00A6F# => romdata <= X"81F0CC23";
    when 16#00A70# => romdata <= X"84120853";
    when 16#00A71# => romdata <= X"722D81F0";
    when 16#00A72# => romdata <= X"CC225170";
    when 16#00A73# => romdata <= X"802EFFBE";
    when 16#00A74# => romdata <= X"38843D0D";
    when 16#00A75# => romdata <= X"04F93D0D";
    when 16#00A76# => romdata <= X"02AA0522";
    when 16#00A77# => romdata <= X"56805574";
    when 16#00A78# => romdata <= X"10101081";
    when 16#00A79# => romdata <= X"EFFC0570";
    when 16#00A7A# => romdata <= X"33525270";
    when 16#00A7B# => romdata <= X"81FE2E99";
    when 16#00A7C# => romdata <= X"38811570";
    when 16#00A7D# => romdata <= X"81FF0656";
    when 16#00A7E# => romdata <= X"52748A2E";
    when 16#00A7F# => romdata <= X"098106DF";
    when 16#00A80# => romdata <= X"38810BB0";
    when 16#00A81# => romdata <= X"0C893D0D";
    when 16#00A82# => romdata <= X"0481F0D0";
    when 16#00A83# => romdata <= X"337081FF";
    when 16#00A84# => romdata <= X"0681F0CC";
    when 16#00A85# => romdata <= X"22535458";
    when 16#00A86# => romdata <= X"7281FF2E";
    when 16#00A87# => romdata <= X"B0387283";
    when 16#00A88# => romdata <= X"2B547076";
    when 16#00A89# => romdata <= X"2780DE38";
    when 16#00A8A# => romdata <= X"75713170";
    when 16#00A8B# => romdata <= X"83FFFF06";
    when 16#00A8C# => romdata <= X"7481EFFC";
    when 16#00A8D# => romdata <= X"17337083";
    when 16#00A8E# => romdata <= X"2B81EFFE";
    when 16#00A8F# => romdata <= X"11225658";
    when 16#00A90# => romdata <= X"56525757";
    when 16#00A91# => romdata <= X"7281FF2E";
    when 16#00A92# => romdata <= X"098106D6";
    when 16#00A93# => romdata <= X"38727234";
    when 16#00A94# => romdata <= X"75821323";
    when 16#00A95# => romdata <= X"7984130C";
    when 16#00A96# => romdata <= X"7781FF06";
    when 16#00A97# => romdata <= X"5473732E";
    when 16#00A98# => romdata <= X"96387610";
    when 16#00A99# => romdata <= X"101081EF";
    when 16#00A9A# => romdata <= X"FC055374";
    when 16#00A9B# => romdata <= X"73348051";
    when 16#00A9C# => romdata <= X"70B00C89";
    when 16#00A9D# => romdata <= X"3D0D0474";
    when 16#00A9E# => romdata <= X"81F0D034";
    when 16#00A9F# => romdata <= X"7581F0CC";
    when 16#00AA0# => romdata <= X"238051EC";
    when 16#00AA1# => romdata <= X"39707631";
    when 16#00AA2# => romdata <= X"517081EF";
    when 16#00AA3# => romdata <= X"FE1523FF";
    when 16#00AA4# => romdata <= X"BC39FF3D";
    when 16#00AA5# => romdata <= X"0D8A5271";
    when 16#00AA6# => romdata <= X"10101081";
    when 16#00AA7# => romdata <= X"EFF40551";
    when 16#00AA8# => romdata <= X"FE7134FF";
    when 16#00AA9# => romdata <= X"127081FF";
    when 16#00AAA# => romdata <= X"06535171";
    when 16#00AAB# => romdata <= X"EA38FF0B";
    when 16#00AAC# => romdata <= X"81F0D034";
    when 16#00AAD# => romdata <= X"833D0D04";
    when 16#00AAE# => romdata <= X"FE3D0D02";
    when 16#00AAF# => romdata <= X"93053302";
    when 16#00AB0# => romdata <= X"84059705";
    when 16#00AB1# => romdata <= X"33545271";
    when 16#00AB2# => romdata <= X"812E9238";
    when 16#00AB3# => romdata <= X"7180D52E";
    when 16#00AB4# => romdata <= X"BB3881BD";
    when 16#00AB5# => romdata <= X"A051A1BA";
    when 16#00AB6# => romdata <= X"3F843D0D";
    when 16#00AB7# => romdata <= X"0481BDAC";
    when 16#00AB8# => romdata <= X"51A1AF3F";
    when 16#00AB9# => romdata <= X"72912E81";
    when 16#00ABA# => romdata <= X"F6387291";
    when 16#00ABB# => romdata <= X"24B53872";
    when 16#00ABC# => romdata <= X"8C2E81F6";
    when 16#00ABD# => romdata <= X"38728C24";
    when 16#00ABE# => romdata <= X"80E33872";
    when 16#00ABF# => romdata <= X"862E81D4";
    when 16#00AC0# => romdata <= X"3881BDB8";
    when 16#00AC1# => romdata <= X"51A18B3F";
    when 16#00AC2# => romdata <= X"843D0D04";
    when 16#00AC3# => romdata <= X"81BDC851";
    when 16#00AC4# => romdata <= X"A1803F72";
    when 16#00AC5# => romdata <= X"8926EA38";
    when 16#00AC6# => romdata <= X"72101081";
    when 16#00AC7# => romdata <= X"C0F40552";
    when 16#00AC8# => romdata <= X"71080472";
    when 16#00AC9# => romdata <= X"A82E81CD";
    when 16#00ACA# => romdata <= X"38A87325";
    when 16#00ACB# => romdata <= X"9C387280";
    when 16#00ACC# => romdata <= X"C52E81CC";
    when 16#00ACD# => romdata <= X"387280E1";
    when 16#00ACE# => romdata <= X"2E098106";
    when 16#00ACF# => romdata <= X"C43881BD";
    when 16#00AD0# => romdata <= X"D451A0CE";
    when 16#00AD1# => romdata <= X"3F843D0D";
    when 16#00AD2# => romdata <= X"04729A2E";
    when 16#00AD3# => romdata <= X"098106FF";
    when 16#00AD4# => romdata <= X"B03881BD";
    when 16#00AD5# => romdata <= X"E451A0BA";
    when 16#00AD6# => romdata <= X"3F843D0D";
    when 16#00AD7# => romdata <= X"04728F2E";
    when 16#00AD8# => romdata <= X"098106FF";
    when 16#00AD9# => romdata <= X"9C3881BE";
    when 16#00ADA# => romdata <= X"8051A0A6";
    when 16#00ADB# => romdata <= X"3F843D0D";
    when 16#00ADC# => romdata <= X"0481BE9C";
    when 16#00ADD# => romdata <= X"51A09B3F";
    when 16#00ADE# => romdata <= X"843D0D04";
    when 16#00ADF# => romdata <= X"81BBA051";
    when 16#00AE0# => romdata <= X"A0903F84";
    when 16#00AE1# => romdata <= X"3D0D0481";
    when 16#00AE2# => romdata <= X"BEB451A0";
    when 16#00AE3# => romdata <= X"853F843D";
    when 16#00AE4# => romdata <= X"0D0481BE";
    when 16#00AE5# => romdata <= X"C8519FFA";
    when 16#00AE6# => romdata <= X"3F843D0D";
    when 16#00AE7# => romdata <= X"0481BED8";
    when 16#00AE8# => romdata <= X"519FEF3F";
    when 16#00AE9# => romdata <= X"843D0D04";
    when 16#00AEA# => romdata <= X"81BEEC51";
    when 16#00AEB# => romdata <= X"9FE43F84";
    when 16#00AEC# => romdata <= X"3D0D0481";
    when 16#00AED# => romdata <= X"BF88519F";
    when 16#00AEE# => romdata <= X"D93F843D";
    when 16#00AEF# => romdata <= X"0D0481BF";
    when 16#00AF0# => romdata <= X"A0519FCE";
    when 16#00AF1# => romdata <= X"3F843D0D";
    when 16#00AF2# => romdata <= X"0481BFB4";
    when 16#00AF3# => romdata <= X"519FC33F";
    when 16#00AF4# => romdata <= X"843D0D04";
    when 16#00AF5# => romdata <= X"81BFC451";
    when 16#00AF6# => romdata <= X"9FB83F84";
    when 16#00AF7# => romdata <= X"3D0D0481";
    when 16#00AF8# => romdata <= X"BFD4519F";
    when 16#00AF9# => romdata <= X"AD3F843D";
    when 16#00AFA# => romdata <= X"0D0481BF";
    when 16#00AFB# => romdata <= X"E8519FA2";
    when 16#00AFC# => romdata <= X"3F843D0D";
    when 16#00AFD# => romdata <= X"0481BFF8";
    when 16#00AFE# => romdata <= X"519F973F";
    when 16#00AFF# => romdata <= X"843D0D04";
    when 16#00B00# => romdata <= X"81C09851";
    when 16#00B01# => romdata <= X"9F8C3F84";
    when 16#00B02# => romdata <= X"3D0D04F7";
    when 16#00B03# => romdata <= X"3D0D02B3";
    when 16#00B04# => romdata <= X"05337C70";
    when 16#00B05# => romdata <= X"08C08080";
    when 16#00B06# => romdata <= X"0659545A";
    when 16#00B07# => romdata <= X"80567583";
    when 16#00B08# => romdata <= X"2B7707BF";
    when 16#00B09# => romdata <= X"E0800770";
    when 16#00B0A# => romdata <= X"70840552";
    when 16#00B0B# => romdata <= X"0871088C";
    when 16#00B0C# => romdata <= X"2ABFFE80";
    when 16#00B0D# => romdata <= X"06790771";
    when 16#00B0E# => romdata <= X"982A728C";
    when 16#00B0F# => romdata <= X"2A9FFF06";
    when 16#00B10# => romdata <= X"73852A70";
    when 16#00B11# => romdata <= X"8F06759F";
    when 16#00B12# => romdata <= X"06565158";
    when 16#00B13# => romdata <= X"5D585255";
    when 16#00B14# => romdata <= X"58748D38";
    when 16#00B15# => romdata <= X"8116568F";
    when 16#00B16# => romdata <= X"7627C338";
    when 16#00B17# => romdata <= X"8B3D0D04";
    when 16#00B18# => romdata <= X"81C0B051";
    when 16#00B19# => romdata <= X"9EAC3F75";
    when 16#00B1A# => romdata <= X"519FF13F";
    when 16#00B1B# => romdata <= X"8452B008";
    when 16#00B1C# => romdata <= X"51FFBAE6";
    when 16#00B1D# => romdata <= X"3F81C0BC";
    when 16#00B1E# => romdata <= X"519E973F";
    when 16#00B1F# => romdata <= X"74528851";
    when 16#00B20# => romdata <= X"9EB33F84";
    when 16#00B21# => romdata <= X"52B00851";
    when 16#00B22# => romdata <= X"FFBACF3F";
    when 16#00B23# => romdata <= X"81C0C451";
    when 16#00B24# => romdata <= X"9E803F78";
    when 16#00B25# => romdata <= X"5290519E";
    when 16#00B26# => romdata <= X"9C3F8652";
    when 16#00B27# => romdata <= X"B00851FF";
    when 16#00B28# => romdata <= X"BAB83F81";
    when 16#00B29# => romdata <= X"C0CC519D";
    when 16#00B2A# => romdata <= X"E93F7251";
    when 16#00B2B# => romdata <= X"9FAE3F84";
    when 16#00B2C# => romdata <= X"52B00851";
    when 16#00B2D# => romdata <= X"FFBAA33F";
    when 16#00B2E# => romdata <= X"81C0D451";
    when 16#00B2F# => romdata <= X"9DD43F73";
    when 16#00B30# => romdata <= X"519F993F";
    when 16#00B31# => romdata <= X"8452B008";
    when 16#00B32# => romdata <= X"51FFBA8E";
    when 16#00B33# => romdata <= X"3F81C0DC";
    when 16#00B34# => romdata <= X"519DBF3F";
    when 16#00B35# => romdata <= X"7752A051";
    when 16#00B36# => romdata <= X"9DDB3F8A";
    when 16#00B37# => romdata <= X"52B00851";
    when 16#00B38# => romdata <= X"FFB9F73F";
    when 16#00B39# => romdata <= X"7992388A";
    when 16#00B3A# => romdata <= X"519D8D3F";
    when 16#00B3B# => romdata <= X"8116568F";
    when 16#00B3C# => romdata <= X"7627FEAA";
    when 16#00B3D# => romdata <= X"38FEE539";
    when 16#00B3E# => romdata <= X"7881FF06";
    when 16#00B3F# => romdata <= X"527451FB";
    when 16#00B40# => romdata <= X"B73F8A51";
    when 16#00B41# => romdata <= X"9CF23FE4";
    when 16#00B42# => romdata <= X"39F83D0D";
    when 16#00B43# => romdata <= X"02AB0533";
    when 16#00B44# => romdata <= X"59805675";
    when 16#00B45# => romdata <= X"852BE090";
    when 16#00B46# => romdata <= X"11E08012";
    when 16#00B47# => romdata <= X"0870982A";
    when 16#00B48# => romdata <= X"718C2A9F";
    when 16#00B49# => romdata <= X"FF067285";
    when 16#00B4A# => romdata <= X"2A708F06";
    when 16#00B4B# => romdata <= X"749F0655";
    when 16#00B4C# => romdata <= X"51585B53";
    when 16#00B4D# => romdata <= X"56595574";
    when 16#00B4E# => romdata <= X"802E81A7";
    when 16#00B4F# => romdata <= X"3875BF26";
    when 16#00B50# => romdata <= X"81AF3881";
    when 16#00B51# => romdata <= X"C0E4519C";
    when 16#00B52# => romdata <= X"C93F7551";
    when 16#00B53# => romdata <= X"9E8E3F86";
    when 16#00B54# => romdata <= X"52B00851";
    when 16#00B55# => romdata <= X"FFB9833F";
    when 16#00B56# => romdata <= X"81C0BC51";
    when 16#00B57# => romdata <= X"9CB43F74";
    when 16#00B58# => romdata <= X"5288519C";
    when 16#00B59# => romdata <= X"D03F8452";
    when 16#00B5A# => romdata <= X"B00851FF";
    when 16#00B5B# => romdata <= X"B8EC3F81";
    when 16#00B5C# => romdata <= X"C0C4519C";
    when 16#00B5D# => romdata <= X"9D3F7652";
    when 16#00B5E# => romdata <= X"90519CB9";
    when 16#00B5F# => romdata <= X"3F8652B0";
    when 16#00B60# => romdata <= X"0851FFB8";
    when 16#00B61# => romdata <= X"D53F81C0";
    when 16#00B62# => romdata <= X"CC519C86";
    when 16#00B63# => romdata <= X"3F72519D";
    when 16#00B64# => romdata <= X"CB3F8452";
    when 16#00B65# => romdata <= X"B00851FF";
    when 16#00B66# => romdata <= X"B8C03F81";
    when 16#00B67# => romdata <= X"C0D4519B";
    when 16#00B68# => romdata <= X"F13F7351";
    when 16#00B69# => romdata <= X"9DB63F84";
    when 16#00B6A# => romdata <= X"52B00851";
    when 16#00B6B# => romdata <= X"FFB8AB3F";
    when 16#00B6C# => romdata <= X"81C0DC51";
    when 16#00B6D# => romdata <= X"9BDC3F77";
    when 16#00B6E# => romdata <= X"08C08080";
    when 16#00B6F# => romdata <= X"0652A051";
    when 16#00B70# => romdata <= X"9BF33F8A";
    when 16#00B71# => romdata <= X"52B00851";
    when 16#00B72# => romdata <= X"FFB88F3F";
    when 16#00B73# => romdata <= X"7881B238";
    when 16#00B74# => romdata <= X"8A519BA4";
    when 16#00B75# => romdata <= X"3F805374";
    when 16#00B76# => romdata <= X"812E81DF";
    when 16#00B77# => romdata <= X"3876862E";
    when 16#00B78# => romdata <= X"81BB3881";
    when 16#00B79# => romdata <= X"165680FF";
    when 16#00B7A# => romdata <= X"7627FEA7";
    when 16#00B7B# => romdata <= X"388A3D0D";
    when 16#00B7C# => romdata <= X"0481C0EC";
    when 16#00B7D# => romdata <= X"519B9B3F";
    when 16#00B7E# => romdata <= X"C016519C";
    when 16#00B7F# => romdata <= X"DF3F8652";
    when 16#00B80# => romdata <= X"B00851FF";
    when 16#00B81# => romdata <= X"B7D43F81";
    when 16#00B82# => romdata <= X"C0BC519B";
    when 16#00B83# => romdata <= X"853F7452";
    when 16#00B84# => romdata <= X"88519BA1";
    when 16#00B85# => romdata <= X"3F8452B0";
    when 16#00B86# => romdata <= X"0851FFB7";
    when 16#00B87# => romdata <= X"BD3F81C0";
    when 16#00B88# => romdata <= X"C4519AEE";
    when 16#00B89# => romdata <= X"3F765290";
    when 16#00B8A# => romdata <= X"519B8A3F";
    when 16#00B8B# => romdata <= X"8652B008";
    when 16#00B8C# => romdata <= X"51FFB7A6";
    when 16#00B8D# => romdata <= X"3F81C0CC";
    when 16#00B8E# => romdata <= X"519AD73F";
    when 16#00B8F# => romdata <= X"72519C9C";
    when 16#00B90# => romdata <= X"3F8452B0";
    when 16#00B91# => romdata <= X"0851FFB7";
    when 16#00B92# => romdata <= X"913F81C0";
    when 16#00B93# => romdata <= X"D4519AC2";
    when 16#00B94# => romdata <= X"3F73519C";
    when 16#00B95# => romdata <= X"873F8452";
    when 16#00B96# => romdata <= X"B00851FF";
    when 16#00B97# => romdata <= X"B6FC3F81";
    when 16#00B98# => romdata <= X"C0DC519A";
    when 16#00B99# => romdata <= X"AD3F7708";
    when 16#00B9A# => romdata <= X"C0808006";
    when 16#00B9B# => romdata <= X"52A0519A";
    when 16#00B9C# => romdata <= X"C43F8A52";
    when 16#00B9D# => romdata <= X"B00851FF";
    when 16#00B9E# => romdata <= X"B6E03F78";
    when 16#00B9F# => romdata <= X"802EFED0";
    when 16#00BA0# => romdata <= X"387681FF";
    when 16#00BA1# => romdata <= X"06527451";
    when 16#00BA2# => romdata <= X"F8AE3F8A";
    when 16#00BA3# => romdata <= X"5199E93F";
    when 16#00BA4# => romdata <= X"80537481";
    when 16#00BA5# => romdata <= X"2E098106";
    when 16#00BA6# => romdata <= X"FEC3389F";
    when 16#00BA7# => romdata <= X"39728106";
    when 16#00BA8# => romdata <= X"5776802E";
    when 16#00BA9# => romdata <= X"FEBD3878";
    when 16#00BAA# => romdata <= X"527751FA";
    when 16#00BAB# => romdata <= X"DE3F8116";
    when 16#00BAC# => romdata <= X"5680FF76";
    when 16#00BAD# => romdata <= X"27FCDC38";
    when 16#00BAE# => romdata <= X"FEB33974";
    when 16#00BAF# => romdata <= X"5376862E";
    when 16#00BB0# => romdata <= X"098106FE";
    when 16#00BB1# => romdata <= X"9E38D639";
    when 16#00BB2# => romdata <= X"FE3D0D74";
    when 16#00BB3# => romdata <= X"02840597";
    when 16#00BB4# => romdata <= X"05330288";
    when 16#00BB5# => romdata <= X"059B0533";
    when 16#00BB6# => romdata <= X"88130C8C";
    when 16#00BB7# => romdata <= X"120C538C";
    when 16#00BB8# => romdata <= X"13087081";
    when 16#00BB9# => romdata <= X"2A810651";
    when 16#00BBA# => romdata <= X"5271F438";
    when 16#00BBB# => romdata <= X"8C130870";
    when 16#00BBC# => romdata <= X"81FF06B0";
    when 16#00BBD# => romdata <= X"0C51843D";
    when 16#00BBE# => romdata <= X"0D04803D";
    when 16#00BBF# => romdata <= X"0D728C11";
    when 16#00BC0# => romdata <= X"0870872A";
    when 16#00BC1# => romdata <= X"81328106";
    when 16#00BC2# => romdata <= X"B00C5151";
    when 16#00BC3# => romdata <= X"823D0D04";
    when 16#00BC4# => romdata <= X"FD3D0D02";
    when 16#00BC5# => romdata <= X"97053302";
    when 16#00BC6# => romdata <= X"84059B05";
    when 16#00BC7# => romdata <= X"337181B0";
    when 16#00BC8# => romdata <= X"0781BF06";
    when 16#00BC9# => romdata <= X"535454F8";
    when 16#00BCA# => romdata <= X"80809880";
    when 16#00BCB# => romdata <= X"71710C73";
    when 16#00BCC# => romdata <= X"842A9007";
    when 16#00BCD# => romdata <= X"710C738F";
    when 16#00BCE# => romdata <= X"06710C52";
    when 16#00BCF# => romdata <= X"7281CCD0";
    when 16#00BD0# => romdata <= X"347381CC";
    when 16#00BD1# => romdata <= X"D434853D";
    when 16#00BD2# => romdata <= X"0D04FD3D";
    when 16#00BD3# => romdata <= X"0D029705";
    when 16#00BD4# => romdata <= X"3381CCD4";
    when 16#00BD5# => romdata <= X"33547305";
    when 16#00BD6# => romdata <= X"87060284";
    when 16#00BD7# => romdata <= X"059A0522";
    when 16#00BD8# => romdata <= X"81CCD033";
    when 16#00BD9# => romdata <= X"54730570";
    when 16#00BDA# => romdata <= X"81FF0672";
    when 16#00BDB# => romdata <= X"81B00754";
    when 16#00BDC# => romdata <= X"515454F8";
    when 16#00BDD# => romdata <= X"80809880";
    when 16#00BDE# => romdata <= X"71710C73";
    when 16#00BDF# => romdata <= X"842A9007";
    when 16#00BE0# => romdata <= X"710C738F";
    when 16#00BE1# => romdata <= X"06710C52";
    when 16#00BE2# => romdata <= X"7281CCD0";
    when 16#00BE3# => romdata <= X"347381CC";
    when 16#00BE4# => romdata <= X"D434853D";
    when 16#00BE5# => romdata <= X"0D04FF3D";
    when 16#00BE6# => romdata <= X"0D028F05";
    when 16#00BE7# => romdata <= X"33F88080";
    when 16#00BE8# => romdata <= X"98840C81";
    when 16#00BE9# => romdata <= X"CCD03381";
    when 16#00BEA# => romdata <= X"05517081";
    when 16#00BEB# => romdata <= X"CCD03483";
    when 16#00BEC# => romdata <= X"3D0D04FF";
    when 16#00BED# => romdata <= X"3D0D8052";
    when 16#00BEE# => romdata <= X"7181B007";
    when 16#00BEF# => romdata <= X"81BF06F8";
    when 16#00BF0# => romdata <= X"80809880";
    when 16#00BF1# => romdata <= X"0C900BF8";
    when 16#00BF2# => romdata <= X"80809880";
    when 16#00BF3# => romdata <= X"0C800BF8";
    when 16#00BF4# => romdata <= X"80809880";
    when 16#00BF5# => romdata <= X"0C805180";
    when 16#00BF6# => romdata <= X"0BF88080";
    when 16#00BF7# => romdata <= X"98840C81";
    when 16#00BF8# => romdata <= X"117081FF";
    when 16#00BF9# => romdata <= X"06515180";
    when 16#00BFA# => romdata <= X"E57127EB";
    when 16#00BFB# => romdata <= X"38811270";
    when 16#00BFC# => romdata <= X"81FF0653";
    when 16#00BFD# => romdata <= X"51877227";
    when 16#00BFE# => romdata <= X"FFBE3881";
    when 16#00BFF# => romdata <= X"B00BF880";
    when 16#00C00# => romdata <= X"8098800C";
    when 16#00C01# => romdata <= X"900BF880";
    when 16#00C02# => romdata <= X"8098800C";
    when 16#00C03# => romdata <= X"800BF880";
    when 16#00C04# => romdata <= X"8098800C";
    when 16#00C05# => romdata <= X"800B81CC";
    when 16#00C06# => romdata <= X"D034800B";
    when 16#00C07# => romdata <= X"81CCD434";
    when 16#00C08# => romdata <= X"833D0D04";
    when 16#00C09# => romdata <= X"FF3D0D80";
    when 16#00C0A# => romdata <= X"C00BF880";
    when 16#00C0B# => romdata <= X"8098800C";
    when 16#00C0C# => romdata <= X"81A10BF8";
    when 16#00C0D# => romdata <= X"80809880";
    when 16#00C0E# => romdata <= X"0C81C00B";
    when 16#00C0F# => romdata <= X"F8808098";
    when 16#00C10# => romdata <= X"800C81A4";
    when 16#00C11# => romdata <= X"0BF88080";
    when 16#00C12# => romdata <= X"98800C81";
    when 16#00C13# => romdata <= X"A60BF880";
    when 16#00C14# => romdata <= X"8098800C";
    when 16#00C15# => romdata <= X"81A20BF8";
    when 16#00C16# => romdata <= X"80809880";
    when 16#00C17# => romdata <= X"0CAF0BF8";
    when 16#00C18# => romdata <= X"80809880";
    when 16#00C19# => romdata <= X"0CA50BF8";
    when 16#00C1A# => romdata <= X"80809880";
    when 16#00C1B# => romdata <= X"0C81810B";
    when 16#00C1C# => romdata <= X"F8808098";
    when 16#00C1D# => romdata <= X"800C9D0B";
    when 16#00C1E# => romdata <= X"F8808098";
    when 16#00C1F# => romdata <= X"800C81FA";
    when 16#00C20# => romdata <= X"0BF88080";
    when 16#00C21# => romdata <= X"98800C80";
    when 16#00C22# => romdata <= X"0BF88080";
    when 16#00C23# => romdata <= X"98800C80";
    when 16#00C24# => romdata <= X"527181B0";
    when 16#00C25# => romdata <= X"0781BF06";
    when 16#00C26# => romdata <= X"F8808098";
    when 16#00C27# => romdata <= X"800C900B";
    when 16#00C28# => romdata <= X"F8808098";
    when 16#00C29# => romdata <= X"800C800B";
    when 16#00C2A# => romdata <= X"F8808098";
    when 16#00C2B# => romdata <= X"800C8051";
    when 16#00C2C# => romdata <= X"800BF880";
    when 16#00C2D# => romdata <= X"8098840C";
    when 16#00C2E# => romdata <= X"81117081";
    when 16#00C2F# => romdata <= X"FF065151";
    when 16#00C30# => romdata <= X"80E57127";
    when 16#00C31# => romdata <= X"EB388112";
    when 16#00C32# => romdata <= X"7081FF06";
    when 16#00C33# => romdata <= X"53518772";
    when 16#00C34# => romdata <= X"27FFBE38";
    when 16#00C35# => romdata <= X"81B00BF8";
    when 16#00C36# => romdata <= X"80809880";
    when 16#00C37# => romdata <= X"0C900BF8";
    when 16#00C38# => romdata <= X"80809880";
    when 16#00C39# => romdata <= X"0C800BF8";
    when 16#00C3A# => romdata <= X"80809880";
    when 16#00C3B# => romdata <= X"0C800B81";
    when 16#00C3C# => romdata <= X"CCD03480";
    when 16#00C3D# => romdata <= X"0B81CCD4";
    when 16#00C3E# => romdata <= X"3481AF0B";
    when 16#00C3F# => romdata <= X"F8808098";
    when 16#00C40# => romdata <= X"800C833D";
    when 16#00C41# => romdata <= X"0D04803D";
    when 16#00C42# => romdata <= X"0D028F05";
    when 16#00C43# => romdata <= X"337381F0";
    when 16#00C44# => romdata <= X"D40C5170";
    when 16#00C45# => romdata <= X"81F0D834";
    when 16#00C46# => romdata <= X"823D0D04";
    when 16#00C47# => romdata <= X"EE3D0D64";
    when 16#00C48# => romdata <= X"02840580";
    when 16#00C49# => romdata <= X"D7053302";
    when 16#00C4A# => romdata <= X"880580DB";
    when 16#00C4B# => romdata <= X"05335957";
    when 16#00C4C# => romdata <= X"59807681";
    when 16#00C4D# => romdata <= X"0677812A";
    when 16#00C4E# => romdata <= X"81067883";
    when 16#00C4F# => romdata <= X"2B818006";
    when 16#00C50# => romdata <= X"79822A81";
    when 16#00C51# => romdata <= X"06575E41";
    when 16#00C52# => romdata <= X"5F5D81FF";
    when 16#00C53# => romdata <= X"42727D2E";
    when 16#00C54# => romdata <= X"09810683";
    when 16#00C55# => romdata <= X"387C4276";
    when 16#00C56# => romdata <= X"8A2E83B9";
    when 16#00C57# => romdata <= X"38881908";
    when 16#00C58# => romdata <= X"5574802E";
    when 16#00C59# => romdata <= X"83A43885";
    when 16#00C5A# => romdata <= X"19335AFF";
    when 16#00C5B# => romdata <= X"53767A26";
    when 16#00C5C# => romdata <= X"8E388419";
    when 16#00C5D# => romdata <= X"33547377";
    when 16#00C5E# => romdata <= X"26853876";
    when 16#00C5F# => romdata <= X"74315374";
    when 16#00C60# => romdata <= X"13703354";
    when 16#00C61# => romdata <= X"587281FF";
    when 16#00C62# => romdata <= X"06831A33";
    when 16#00C63# => romdata <= X"70982B81";
    when 16#00C64# => romdata <= X"FF0A119B";
    when 16#00C65# => romdata <= X"2A81055B";
    when 16#00C66# => romdata <= X"45424081";
    when 16#00C67# => romdata <= X"53748338";
    when 16#00C68# => romdata <= X"74537281";
    when 16#00C69# => romdata <= X"FF064380";
    when 16#00C6A# => romdata <= X"7A81FF06";
    when 16#00C6B# => romdata <= X"545CFF54";
    when 16#00C6C# => romdata <= X"7673268B";
    when 16#00C6D# => romdata <= X"38841933";
    when 16#00C6E# => romdata <= X"53767327";
    when 16#00C6F# => romdata <= X"83F43873";
    when 16#00C70# => romdata <= X"7481FF06";
    when 16#00C71# => romdata <= X"5553805A";
    when 16#00C72# => romdata <= X"797324AB";
    when 16#00C73# => romdata <= X"38747A2E";
    when 16#00C74# => romdata <= X"09810682";
    when 16#00C75# => romdata <= X"E1386098";
    when 16#00C76# => romdata <= X"2B81FF0A";
    when 16#00C77# => romdata <= X"119B2A82";
    when 16#00C78# => romdata <= X"1B337171";
    when 16#00C79# => romdata <= X"29117081";
    when 16#00C7A# => romdata <= X"FF067871";
    when 16#00C7B# => romdata <= X"298C1F08";
    when 16#00C7C# => romdata <= X"0552455D";
    when 16#00C7D# => romdata <= X"575D537F";
    when 16#00C7E# => romdata <= X"63057081";
    when 16#00C7F# => romdata <= X"FF067061";
    when 16#00C80# => romdata <= X"2B7081FF";
    when 16#00C81# => romdata <= X"067B622B";
    when 16#00C82# => romdata <= X"7081FF06";
    when 16#00C83# => romdata <= X"7B832A81";
    when 16#00C84# => romdata <= X"065F5358";
    when 16#00C85# => romdata <= X"525E4255";
    when 16#00C86# => romdata <= X"78802E8F";
    when 16#00C87# => romdata <= X"3881CCD0";
    when 16#00C88# => romdata <= X"33610556";
    when 16#00C89# => romdata <= X"7580E624";
    when 16#00C8A# => romdata <= X"83C5387F";
    when 16#00C8B# => romdata <= X"78296130";
    when 16#00C8C# => romdata <= X"41577C7E";
    when 16#00C8D# => romdata <= X"2C982B70";
    when 16#00C8E# => romdata <= X"982C5555";
    when 16#00C8F# => romdata <= X"73772581";
    when 16#00C90# => romdata <= X"8238FF1C";
    when 16#00C91# => romdata <= X"7D81065A";
    when 16#00C92# => romdata <= X"537C732E";
    when 16#00C93# => romdata <= X"83C4387E";
    when 16#00C94# => romdata <= X"86A63861";
    when 16#00C95# => romdata <= X"84EB387D";
    when 16#00C96# => romdata <= X"802E82A4";
    when 16#00C97# => romdata <= X"38791470";
    when 16#00C98# => romdata <= X"33705854";
    when 16#00C99# => romdata <= X"55805578";
    when 16#00C9A# => romdata <= X"752E8538";
    when 16#00C9B# => romdata <= X"72842A56";
    when 16#00C9C# => romdata <= X"75832A70";
    when 16#00C9D# => romdata <= X"81065153";
    when 16#00C9E# => romdata <= X"72802E84";
    when 16#00C9F# => romdata <= X"3881C055";
    when 16#00CA0# => romdata <= X"75822A70";
    when 16#00CA1# => romdata <= X"81065153";
    when 16#00CA2# => romdata <= X"72802E85";
    when 16#00CA3# => romdata <= X"3874B007";
    when 16#00CA4# => romdata <= X"5575812A";
    when 16#00CA5# => romdata <= X"70810651";
    when 16#00CA6# => romdata <= X"5372802E";
    when 16#00CA7# => romdata <= X"8538748C";
    when 16#00CA8# => romdata <= X"07557581";
    when 16#00CA9# => romdata <= X"06537280";
    when 16#00CAA# => romdata <= X"2E853874";
    when 16#00CAB# => romdata <= X"83075574";
    when 16#00CAC# => romdata <= X"51F9E33F";
    when 16#00CAD# => romdata <= X"7714982B";
    when 16#00CAE# => romdata <= X"70982C55";
    when 16#00CAF# => romdata <= X"56767424";
    when 16#00CB0# => romdata <= X"FF9B3862";
    when 16#00CB1# => romdata <= X"802E9538";
    when 16#00CB2# => romdata <= X"61FF1D54";
    when 16#00CB3# => romdata <= X"547C732E";
    when 16#00CB4# => romdata <= X"81FB3873";
    when 16#00CB5# => romdata <= X"51F9BF3F";
    when 16#00CB6# => romdata <= X"7E81EA38";
    when 16#00CB7# => romdata <= X"7F528151";
    when 16#00CB8# => romdata <= X"F8E83F81";
    when 16#00CB9# => romdata <= X"1D7081FF";
    when 16#00CBA# => romdata <= X"065E547B";
    when 16#00CBB# => romdata <= X"7D26FEC2";
    when 16#00CBC# => romdata <= X"3860527B";
    when 16#00CBD# => romdata <= X"3070982B";
    when 16#00CBE# => romdata <= X"70982C53";
    when 16#00CBF# => romdata <= X"585BF8CA";
    when 16#00CC0# => romdata <= X"3F605372";
    when 16#00CC1# => romdata <= X"B00C943D";
    when 16#00CC2# => romdata <= X"0D048219";
    when 16#00CC3# => romdata <= X"33851A33";
    when 16#00CC4# => romdata <= X"5B53FCF1";
    when 16#00CC5# => romdata <= X"3981CCD4";
    when 16#00CC6# => romdata <= X"33537287";
    when 16#00CC7# => romdata <= X"26819A38";
    when 16#00CC8# => romdata <= X"81135680";
    when 16#00CC9# => romdata <= X"527581FF";
    when 16#00CCA# => romdata <= X"0651F7E4";
    when 16#00CCB# => romdata <= X"3F805372";
    when 16#00CCC# => romdata <= X"B00C943D";
    when 16#00CCD# => romdata <= X"0D047380";
    when 16#00CCE# => romdata <= X"2EAF38FF";
    when 16#00CCF# => romdata <= X"147081FF";
    when 16#00CD0# => romdata <= X"06555A73";
    when 16#00CD1# => romdata <= X"81FF2EA1";
    when 16#00CD2# => romdata <= X"38747081";
    when 16#00CD3# => romdata <= X"0556337C";
    when 16#00CD4# => romdata <= X"057083FF";
    when 16#00CD5# => romdata <= X"FF06FF16";
    when 16#00CD6# => romdata <= X"7081FF06";
    when 16#00CD7# => romdata <= X"575C5D53";
    when 16#00CD8# => romdata <= X"7381FF2E";
    when 16#00CD9# => romdata <= X"098106E1";
    when 16#00CDA# => romdata <= X"3860982B";
    when 16#00CDB# => romdata <= X"81FF0A11";
    when 16#00CDC# => romdata <= X"9B2A707E";
    when 16#00CDD# => romdata <= X"291E8C1C";
    when 16#00CDE# => romdata <= X"08055C42";
    when 16#00CDF# => romdata <= X"55FCF839";
    when 16#00CE0# => romdata <= X"79147033";
    when 16#00CE1# => romdata <= X"5259F88E";
    when 16#00CE2# => romdata <= X"3F771498";
    when 16#00CE3# => romdata <= X"2B70982C";
    when 16#00CE4# => romdata <= X"55567377";
    when 16#00CE5# => romdata <= X"25FEAC38";
    when 16#00CE6# => romdata <= X"79147033";
    when 16#00CE7# => romdata <= X"5259F7F6";
    when 16#00CE8# => romdata <= X"3F771498";
    when 16#00CE9# => romdata <= X"2B70982C";
    when 16#00CEA# => romdata <= X"55567674";
    when 16#00CEB# => romdata <= X"24D238FE";
    when 16#00CEC# => romdata <= X"92397673";
    when 16#00CED# => romdata <= X"3154FC87";
    when 16#00CEE# => romdata <= X"39805280";
    when 16#00CEF# => romdata <= X"51F6D13F";
    when 16#00CF0# => romdata <= X"8053FEEB";
    when 16#00CF1# => romdata <= X"397351F7";
    when 16#00CF2# => romdata <= X"CD3FFE90";
    when 16#00CF3# => romdata <= X"39617B32";
    when 16#00CF4# => romdata <= X"7081FF06";
    when 16#00CF5# => romdata <= X"55557D80";
    when 16#00CF6# => romdata <= X"2EFDF838";
    when 16#00CF7# => romdata <= X"7A812A74";
    when 16#00CF8# => romdata <= X"32705254";
    when 16#00CF9# => romdata <= X"F7B03F7E";
    when 16#00CFA# => romdata <= X"802EFDF0";
    when 16#00CFB# => romdata <= X"38D73981";
    when 16#00CFC# => romdata <= X"CCD4337C";
    when 16#00CFD# => romdata <= X"05538052";
    when 16#00CFE# => romdata <= X"7281FF06";
    when 16#00CFF# => romdata <= X"51F6913F";
    when 16#00D00# => romdata <= X"805376A0";
    when 16#00D01# => romdata <= X"2EFDFC38";
    when 16#00D02# => romdata <= X"7F782961";
    when 16#00D03# => romdata <= X"304157FC";
    when 16#00D04# => romdata <= X"A1397E87";
    when 16#00D05# => romdata <= X"AD386185";
    when 16#00D06# => romdata <= X"EB387D80";
    when 16#00D07# => romdata <= X"2E80EC38";
    when 16#00D08# => romdata <= X"79147033";
    when 16#00D09# => romdata <= X"7C077052";
    when 16#00D0A# => romdata <= X"54568055";
    when 16#00D0B# => romdata <= X"78752E85";
    when 16#00D0C# => romdata <= X"3872842A";
    when 16#00D0D# => romdata <= X"5675832A";
    when 16#00D0E# => romdata <= X"70810651";
    when 16#00D0F# => romdata <= X"5372802E";
    when 16#00D10# => romdata <= X"843881C0";
    when 16#00D11# => romdata <= X"5575822A";
    when 16#00D12# => romdata <= X"70810651";
    when 16#00D13# => romdata <= X"5372802E";
    when 16#00D14# => romdata <= X"853874B0";
    when 16#00D15# => romdata <= X"07557581";
    when 16#00D16# => romdata <= X"2A708106";
    when 16#00D17# => romdata <= X"51537280";
    when 16#00D18# => romdata <= X"2E853874";
    when 16#00D19# => romdata <= X"8C075575";
    when 16#00D1A# => romdata <= X"81065372";
    when 16#00D1B# => romdata <= X"802E8538";
    when 16#00D1C# => romdata <= X"74830755";
    when 16#00D1D# => romdata <= X"7451F69E";
    when 16#00D1E# => romdata <= X"3F771498";
    when 16#00D1F# => romdata <= X"2B70982C";
    when 16#00D20# => romdata <= X"55537674";
    when 16#00D21# => romdata <= X"24FF9938";
    when 16#00D22# => romdata <= X"FCB93979";
    when 16#00D23# => romdata <= X"1470337C";
    when 16#00D24# => romdata <= X"075256F6";
    when 16#00D25# => romdata <= X"813F7714";
    when 16#00D26# => romdata <= X"982B7098";
    when 16#00D27# => romdata <= X"2C555973";
    when 16#00D28# => romdata <= X"7725FC9F";
    when 16#00D29# => romdata <= X"38791470";
    when 16#00D2A# => romdata <= X"337C0752";
    when 16#00D2B# => romdata <= X"56F5E73F";
    when 16#00D2C# => romdata <= X"7714982B";
    when 16#00D2D# => romdata <= X"70982C55";
    when 16#00D2E# => romdata <= X"59767424";
    when 16#00D2F# => romdata <= X"CE38FC83";
    when 16#00D30# => romdata <= X"397D802E";
    when 16#00D31# => romdata <= X"80F03879";
    when 16#00D32# => romdata <= X"14703370";
    when 16#00D33# => romdata <= X"58545580";
    when 16#00D34# => romdata <= X"5578752E";
    when 16#00D35# => romdata <= X"85387284";
    when 16#00D36# => romdata <= X"2A567583";
    when 16#00D37# => romdata <= X"2A708106";
    when 16#00D38# => romdata <= X"51537280";
    when 16#00D39# => romdata <= X"2E843881";
    when 16#00D3A# => romdata <= X"C0557582";
    when 16#00D3B# => romdata <= X"2A708106";
    when 16#00D3C# => romdata <= X"51537280";
    when 16#00D3D# => romdata <= X"2E853874";
    when 16#00D3E# => romdata <= X"B0075575";
    when 16#00D3F# => romdata <= X"812A7081";
    when 16#00D40# => romdata <= X"06515372";
    when 16#00D41# => romdata <= X"802E8538";
    when 16#00D42# => romdata <= X"748C0755";
    when 16#00D43# => romdata <= X"75810653";
    when 16#00D44# => romdata <= X"72802E85";
    when 16#00D45# => romdata <= X"38748307";
    when 16#00D46# => romdata <= X"55740970";
    when 16#00D47# => romdata <= X"81FF0652";
    when 16#00D48# => romdata <= X"53F4F33F";
    when 16#00D49# => romdata <= X"7714982B";
    when 16#00D4A# => romdata <= X"70982C55";
    when 16#00D4B# => romdata <= X"56767424";
    when 16#00D4C# => romdata <= X"FF9538FB";
    when 16#00D4D# => romdata <= X"8E397914";
    when 16#00D4E# => romdata <= X"70337009";
    when 16#00D4F# => romdata <= X"7081FF06";
    when 16#00D50# => romdata <= X"54585455";
    when 16#00D51# => romdata <= X"F4D03F77";
    when 16#00D52# => romdata <= X"14982B70";
    when 16#00D53# => romdata <= X"982C5559";
    when 16#00D54# => romdata <= X"737725FA";
    when 16#00D55# => romdata <= X"EE387914";
    when 16#00D56# => romdata <= X"70337009";
    when 16#00D57# => romdata <= X"7081FF06";
    when 16#00D58# => romdata <= X"54585455";
    when 16#00D59# => romdata <= X"F4B03F77";
    when 16#00D5A# => romdata <= X"14982B70";
    when 16#00D5B# => romdata <= X"982C5559";
    when 16#00D5C# => romdata <= X"767424C2";
    when 16#00D5D# => romdata <= X"38FACC39";
    when 16#00D5E# => romdata <= X"61802E81";
    when 16#00D5F# => romdata <= X"CE387D80";
    when 16#00D60# => romdata <= X"2E80F738";
    when 16#00D61# => romdata <= X"79147033";
    when 16#00D62# => romdata <= X"70585455";
    when 16#00D63# => romdata <= X"80557875";
    when 16#00D64# => romdata <= X"2E853872";
    when 16#00D65# => romdata <= X"842A5675";
    when 16#00D66# => romdata <= X"832A7081";
    when 16#00D67# => romdata <= X"06515372";
    when 16#00D68# => romdata <= X"802E8438";
    when 16#00D69# => romdata <= X"81C05575";
    when 16#00D6A# => romdata <= X"822A7081";
    when 16#00D6B# => romdata <= X"06515372";
    when 16#00D6C# => romdata <= X"802E8538";
    when 16#00D6D# => romdata <= X"74B00755";
    when 16#00D6E# => romdata <= X"75812A70";
    when 16#00D6F# => romdata <= X"81065153";
    when 16#00D70# => romdata <= X"72802E85";
    when 16#00D71# => romdata <= X"38748C07";
    when 16#00D72# => romdata <= X"55758106";
    when 16#00D73# => romdata <= X"5372802E";
    when 16#00D74# => romdata <= X"85387483";
    when 16#00D75# => romdata <= X"07557409";
    when 16#00D76# => romdata <= X"7081FF06";
    when 16#00D77# => romdata <= X"70535753";
    when 16#00D78# => romdata <= X"F3B43F75";
    when 16#00D79# => romdata <= X"51F3AF3F";
    when 16#00D7A# => romdata <= X"7714982B";
    when 16#00D7B# => romdata <= X"70982C55";
    when 16#00D7C# => romdata <= X"55767424";
    when 16#00D7D# => romdata <= X"FF8E38F9";
    when 16#00D7E# => romdata <= X"CA397914";
    when 16#00D7F# => romdata <= X"70337009";
    when 16#00D80# => romdata <= X"7081FF06";
    when 16#00D81# => romdata <= X"70555955";
    when 16#00D82# => romdata <= X"5659F38A";
    when 16#00D83# => romdata <= X"3F7551F3";
    when 16#00D84# => romdata <= X"853F7714";
    when 16#00D85# => romdata <= X"982B7098";
    when 16#00D86# => romdata <= X"2C555973";
    when 16#00D87# => romdata <= X"7725F9A3";
    when 16#00D88# => romdata <= X"38791470";
    when 16#00D89# => romdata <= X"33700970";
    when 16#00D8A# => romdata <= X"81FF0670";
    when 16#00D8B# => romdata <= X"55595556";
    when 16#00D8C# => romdata <= X"59F2E33F";
    when 16#00D8D# => romdata <= X"7551F2DE";
    when 16#00D8E# => romdata <= X"3F771498";
    when 16#00D8F# => romdata <= X"2B70982C";
    when 16#00D90# => romdata <= X"55597674";
    when 16#00D91# => romdata <= X"24FFB338";
    when 16#00D92# => romdata <= X"F8F9397D";
    when 16#00D93# => romdata <= X"802E80F4";
    when 16#00D94# => romdata <= X"38791470";
    when 16#00D95# => romdata <= X"33705854";
    when 16#00D96# => romdata <= X"55805578";
    when 16#00D97# => romdata <= X"752E8538";
    when 16#00D98# => romdata <= X"72842A56";
    when 16#00D99# => romdata <= X"75832A70";
    when 16#00D9A# => romdata <= X"81065153";
    when 16#00D9B# => romdata <= X"72802E84";
    when 16#00D9C# => romdata <= X"3881C055";
    when 16#00D9D# => romdata <= X"75822A70";
    when 16#00D9E# => romdata <= X"81065153";
    when 16#00D9F# => romdata <= X"72802E85";
    when 16#00DA0# => romdata <= X"3874B007";
    when 16#00DA1# => romdata <= X"5575812A";
    when 16#00DA2# => romdata <= X"70810651";
    when 16#00DA3# => romdata <= X"5372802E";
    when 16#00DA4# => romdata <= X"8538748C";
    when 16#00DA5# => romdata <= X"07557581";
    when 16#00DA6# => romdata <= X"06537280";
    when 16#00DA7# => romdata <= X"2E853874";
    when 16#00DA8# => romdata <= X"83075574";
    when 16#00DA9# => romdata <= X"81FF0670";
    when 16#00DAA# => romdata <= X"5256F1EA";
    when 16#00DAB# => romdata <= X"3F7551F1";
    when 16#00DAC# => romdata <= X"E53F7714";
    when 16#00DAD# => romdata <= X"982B7098";
    when 16#00DAE# => romdata <= X"2C555576";
    when 16#00DAF# => romdata <= X"7424FF91";
    when 16#00DB0# => romdata <= X"38F88039";
    when 16#00DB1# => romdata <= X"79147033";
    when 16#00DB2# => romdata <= X"70535753";
    when 16#00DB3# => romdata <= X"F1C83F75";
    when 16#00DB4# => romdata <= X"51F1C33F";
    when 16#00DB5# => romdata <= X"7714982B";
    when 16#00DB6# => romdata <= X"70982C55";
    when 16#00DB7# => romdata <= X"59737725";
    when 16#00DB8# => romdata <= X"F7E13879";
    when 16#00DB9# => romdata <= X"14703370";
    when 16#00DBA# => romdata <= X"535753F1";
    when 16#00DBB# => romdata <= X"A93F7551";
    when 16#00DBC# => romdata <= X"F1A43F77";
    when 16#00DBD# => romdata <= X"14982B70";
    when 16#00DBE# => romdata <= X"982C5559";
    when 16#00DBF# => romdata <= X"767424C4";
    when 16#00DC0# => romdata <= X"38F7C039";
    when 16#00DC1# => romdata <= X"7D802E80";
    when 16#00DC2# => romdata <= X"F2387914";
    when 16#00DC3# => romdata <= X"70337C07";
    when 16#00DC4# => romdata <= X"70525456";
    when 16#00DC5# => romdata <= X"80557875";
    when 16#00DC6# => romdata <= X"2E853872";
    when 16#00DC7# => romdata <= X"842A5675";
    when 16#00DC8# => romdata <= X"832A7081";
    when 16#00DC9# => romdata <= X"06515372";
    when 16#00DCA# => romdata <= X"802E8438";
    when 16#00DCB# => romdata <= X"81C05575";
    when 16#00DCC# => romdata <= X"822A7081";
    when 16#00DCD# => romdata <= X"06515372";
    when 16#00DCE# => romdata <= X"802E8538";
    when 16#00DCF# => romdata <= X"74B00755";
    when 16#00DD0# => romdata <= X"75812A70";
    when 16#00DD1# => romdata <= X"81065153";
    when 16#00DD2# => romdata <= X"72802E85";
    when 16#00DD3# => romdata <= X"38748C07";
    when 16#00DD4# => romdata <= X"55758106";
    when 16#00DD5# => romdata <= X"5372802E";
    when 16#00DD6# => romdata <= X"85387483";
    when 16#00DD7# => romdata <= X"07557409";
    when 16#00DD8# => romdata <= X"7081FF06";
    when 16#00DD9# => romdata <= X"5256F0AE";
    when 16#00DDA# => romdata <= X"3F771498";
    when 16#00DDB# => romdata <= X"2B70982C";
    when 16#00DDC# => romdata <= X"55537674";
    when 16#00DDD# => romdata <= X"24FF9338";
    when 16#00DDE# => romdata <= X"F6C93979";
    when 16#00DDF# => romdata <= X"1470337C";
    when 16#00DE0# => romdata <= X"07700970";
    when 16#00DE1# => romdata <= X"81FF0654";
    when 16#00DE2# => romdata <= X"555659F0";
    when 16#00DE3# => romdata <= X"893F7714";
    when 16#00DE4# => romdata <= X"982B7098";
    when 16#00DE5# => romdata <= X"2C555973";
    when 16#00DE6# => romdata <= X"7725F6A7";
    when 16#00DE7# => romdata <= X"38791470";
    when 16#00DE8# => romdata <= X"337C0770";
    when 16#00DE9# => romdata <= X"097081FF";
    when 16#00DEA# => romdata <= X"06545556";
    when 16#00DEB# => romdata <= X"59EFE73F";
    when 16#00DEC# => romdata <= X"7714982B";
    when 16#00DED# => romdata <= X"70982C55";
    when 16#00DEE# => romdata <= X"59767424";
    when 16#00DEF# => romdata <= X"FFBD38F6";
    when 16#00DF0# => romdata <= X"82396180";
    when 16#00DF1# => romdata <= X"2E81D438";
    when 16#00DF2# => romdata <= X"7D802E80";
    when 16#00DF3# => romdata <= X"F9387914";
    when 16#00DF4# => romdata <= X"70337C07";
    when 16#00DF5# => romdata <= X"70525456";
    when 16#00DF6# => romdata <= X"80557875";
    when 16#00DF7# => romdata <= X"2E853872";
    when 16#00DF8# => romdata <= X"842A5675";
    when 16#00DF9# => romdata <= X"832A7081";
    when 16#00DFA# => romdata <= X"06515372";
    when 16#00DFB# => romdata <= X"802E8438";
    when 16#00DFC# => romdata <= X"81C05575";
    when 16#00DFD# => romdata <= X"822A7081";
    when 16#00DFE# => romdata <= X"06515372";
    when 16#00DFF# => romdata <= X"802E8538";
    when 16#00E00# => romdata <= X"74B00755";
    when 16#00E01# => romdata <= X"75812A70";
    when 16#00E02# => romdata <= X"81065153";
    when 16#00E03# => romdata <= X"72802E85";
    when 16#00E04# => romdata <= X"38748C07";
    when 16#00E05# => romdata <= X"55758106";
    when 16#00E06# => romdata <= X"5372802E";
    when 16#00E07# => romdata <= X"85387483";
    when 16#00E08# => romdata <= X"07557409";
    when 16#00E09# => romdata <= X"7081FF06";
    when 16#00E0A# => romdata <= X"70535456";
    when 16#00E0B# => romdata <= X"EEE83F72";
    when 16#00E0C# => romdata <= X"51EEE33F";
    when 16#00E0D# => romdata <= X"7714982B";
    when 16#00E0E# => romdata <= X"70982C55";
    when 16#00E0F# => romdata <= X"56767424";
    when 16#00E10# => romdata <= X"FF8C38F4";
    when 16#00E11# => romdata <= X"FE397914";
    when 16#00E12# => romdata <= X"70337C07";
    when 16#00E13# => romdata <= X"70097081";
    when 16#00E14# => romdata <= X"FF067055";
    when 16#00E15# => romdata <= X"53575753";
    when 16#00E16# => romdata <= X"EEBC3F72";
    when 16#00E17# => romdata <= X"51EEB73F";
    when 16#00E18# => romdata <= X"7714982B";
    when 16#00E19# => romdata <= X"70982C55";
    when 16#00E1A# => romdata <= X"59737725";
    when 16#00E1B# => romdata <= X"F4D53879";
    when 16#00E1C# => romdata <= X"1470337C";
    when 16#00E1D# => romdata <= X"07700970";
    when 16#00E1E# => romdata <= X"81FF0670";
    when 16#00E1F# => romdata <= X"55535757";
    when 16#00E20# => romdata <= X"53EE933F";
    when 16#00E21# => romdata <= X"7251EE8E";
    when 16#00E22# => romdata <= X"3F771498";
    when 16#00E23# => romdata <= X"2B70982C";
    when 16#00E24# => romdata <= X"55597674";
    when 16#00E25# => romdata <= X"24FFAF38";
    when 16#00E26# => romdata <= X"F4A9397D";
    when 16#00E27# => romdata <= X"802E80F6";
    when 16#00E28# => romdata <= X"38791470";
    when 16#00E29# => romdata <= X"337C0770";
    when 16#00E2A# => romdata <= X"52545680";
    when 16#00E2B# => romdata <= X"5578752E";
    when 16#00E2C# => romdata <= X"85387284";
    when 16#00E2D# => romdata <= X"2A567583";
    when 16#00E2E# => romdata <= X"2A708106";
    when 16#00E2F# => romdata <= X"51537280";
    when 16#00E30# => romdata <= X"2E843881";
    when 16#00E31# => romdata <= X"C0557582";
    when 16#00E32# => romdata <= X"2A708106";
    when 16#00E33# => romdata <= X"51537280";
    when 16#00E34# => romdata <= X"2E853874";
    when 16#00E35# => romdata <= X"B0075575";
    when 16#00E36# => romdata <= X"812A7081";
    when 16#00E37# => romdata <= X"06515372";
    when 16#00E38# => romdata <= X"802E8538";
    when 16#00E39# => romdata <= X"748C0755";
    when 16#00E3A# => romdata <= X"75810653";
    when 16#00E3B# => romdata <= X"72802E85";
    when 16#00E3C# => romdata <= X"38748307";
    when 16#00E3D# => romdata <= X"557481FF";
    when 16#00E3E# => romdata <= X"06705256";
    when 16#00E3F# => romdata <= X"ED983F75";
    when 16#00E40# => romdata <= X"51ED933F";
    when 16#00E41# => romdata <= X"7714982B";
    when 16#00E42# => romdata <= X"70982C55";
    when 16#00E43# => romdata <= X"53767424";
    when 16#00E44# => romdata <= X"FF8F38F3";
    when 16#00E45# => romdata <= X"AE397914";
    when 16#00E46# => romdata <= X"70337C07";
    when 16#00E47# => romdata <= X"70535456";
    when 16#00E48# => romdata <= X"ECF43F72";
    when 16#00E49# => romdata <= X"51ECEF3F";
    when 16#00E4A# => romdata <= X"7714982B";
    when 16#00E4B# => romdata <= X"70982C55";
    when 16#00E4C# => romdata <= X"59737725";
    when 16#00E4D# => romdata <= X"F38D3879";
    when 16#00E4E# => romdata <= X"1470337C";
    when 16#00E4F# => romdata <= X"07705354";
    when 16#00E50# => romdata <= X"56ECD33F";
    when 16#00E51# => romdata <= X"7251ECCE";
    when 16#00E52# => romdata <= X"3F771498";
    when 16#00E53# => romdata <= X"2B70982C";
    when 16#00E54# => romdata <= X"55597674";
    when 16#00E55# => romdata <= X"24C038F2";
    when 16#00E56# => romdata <= X"EA39F83D";
    when 16#00E57# => romdata <= X"0D7A7D02";
    when 16#00E58# => romdata <= X"8805AF05";
    when 16#00E59# => romdata <= X"335A5559";
    when 16#00E5A# => romdata <= X"80747081";
    when 16#00E5B# => romdata <= X"05563375";
    when 16#00E5C# => romdata <= X"58565774";
    when 16#00E5D# => romdata <= X"772E0981";
    when 16#00E5E# => romdata <= X"06883876";
    when 16#00E5F# => romdata <= X"B00C8A3D";
    when 16#00E60# => romdata <= X"0D047453";
    when 16#00E61# => romdata <= X"77527851";
    when 16#00E62# => romdata <= X"EF923FB0";
    when 16#00E63# => romdata <= X"0881FF06";
    when 16#00E64# => romdata <= X"77057083";
    when 16#00E65# => romdata <= X"FFFF0677";
    when 16#00E66# => romdata <= X"70810559";
    when 16#00E67# => romdata <= X"33525855";
    when 16#00E68# => romdata <= X"74802ED7";
    when 16#00E69# => romdata <= X"38745377";
    when 16#00E6A# => romdata <= X"527851EE";
    when 16#00E6B# => romdata <= X"EF3FB008";
    when 16#00E6C# => romdata <= X"81FF0677";
    when 16#00E6D# => romdata <= X"057083FF";
    when 16#00E6E# => romdata <= X"FF067770";
    when 16#00E6F# => romdata <= X"81055933";
    when 16#00E70# => romdata <= X"52585574";
    when 16#00E71# => romdata <= X"FFBC38FF";
    when 16#00E72# => romdata <= X"B239FE3D";
    when 16#00E73# => romdata <= X"0D029305";
    when 16#00E74# => romdata <= X"335381F0";
    when 16#00E75# => romdata <= X"D8335281";
    when 16#00E76# => romdata <= X"F0D40851";
    when 16#00E77# => romdata <= X"EEBE3FB0";
    when 16#00E78# => romdata <= X"0881FF06";
    when 16#00E79# => romdata <= X"B00C843D";
    when 16#00E7A# => romdata <= X"0D04D282";
    when 16#00E7B# => romdata <= X"3F04FB3D";
    when 16#00E7C# => romdata <= X"0D777955";
    when 16#00E7D# => romdata <= X"55805675";
    when 16#00E7E# => romdata <= X"7524AB38";
    when 16#00E7F# => romdata <= X"8074249D";
    when 16#00E80# => romdata <= X"38805373";
    when 16#00E81# => romdata <= X"52745180";
    when 16#00E82# => romdata <= X"E13FB008";
    when 16#00E83# => romdata <= X"5475802E";
    when 16#00E84# => romdata <= X"8538B008";
    when 16#00E85# => romdata <= X"305473B0";
    when 16#00E86# => romdata <= X"0C873D0D";
    when 16#00E87# => romdata <= X"04733076";
    when 16#00E88# => romdata <= X"81325754";
    when 16#00E89# => romdata <= X"DC397430";
    when 16#00E8A# => romdata <= X"55815673";
    when 16#00E8B# => romdata <= X"8025D238";
    when 16#00E8C# => romdata <= X"EC39FA3D";
    when 16#00E8D# => romdata <= X"0D787A57";
    when 16#00E8E# => romdata <= X"55805776";
    when 16#00E8F# => romdata <= X"7524A438";
    when 16#00E90# => romdata <= X"759F2C54";
    when 16#00E91# => romdata <= X"81537574";
    when 16#00E92# => romdata <= X"32743152";
    when 16#00E93# => romdata <= X"74519B3F";
    when 16#00E94# => romdata <= X"B0085476";
    when 16#00E95# => romdata <= X"802E8538";
    when 16#00E96# => romdata <= X"B0083054";
    when 16#00E97# => romdata <= X"73B00C88";
    when 16#00E98# => romdata <= X"3D0D0474";
    when 16#00E99# => romdata <= X"30558157";
    when 16#00E9A# => romdata <= X"D739FC3D";
    when 16#00E9B# => romdata <= X"0D767853";
    when 16#00E9C# => romdata <= X"54815380";
    when 16#00E9D# => romdata <= X"74732652";
    when 16#00E9E# => romdata <= X"5572802E";
    when 16#00E9F# => romdata <= X"98387080";
    when 16#00EA0# => romdata <= X"2EA93880";
    when 16#00EA1# => romdata <= X"7224A438";
    when 16#00EA2# => romdata <= X"71107310";
    when 16#00EA3# => romdata <= X"75722653";
    when 16#00EA4# => romdata <= X"545272EA";
    when 16#00EA5# => romdata <= X"38735178";
    when 16#00EA6# => romdata <= X"83387451";
    when 16#00EA7# => romdata <= X"70B00C86";
    when 16#00EA8# => romdata <= X"3D0D0472";
    when 16#00EA9# => romdata <= X"812A7281";
    when 16#00EAA# => romdata <= X"2A535372";
    when 16#00EAB# => romdata <= X"802EE638";
    when 16#00EAC# => romdata <= X"717426EF";
    when 16#00EAD# => romdata <= X"38737231";
    when 16#00EAE# => romdata <= X"75740774";
    when 16#00EAF# => romdata <= X"812A7481";
    when 16#00EB0# => romdata <= X"2A555556";
    when 16#00EB1# => romdata <= X"54E53910";
    when 16#00EB2# => romdata <= X"10101010";
    when 16#00EB3# => romdata <= X"10101010";
    when 16#00EB4# => romdata <= X"10101010";
    when 16#00EB5# => romdata <= X"10101010";
    when 16#00EB6# => romdata <= X"10101010";
    when 16#00EB7# => romdata <= X"10101010";
    when 16#00EB8# => romdata <= X"10101010";
    when 16#00EB9# => romdata <= X"10105351";
    when 16#00EBA# => romdata <= X"047381FF";
    when 16#00EBB# => romdata <= X"06738306";
    when 16#00EBC# => romdata <= X"09810583";
    when 16#00EBD# => romdata <= X"05101010";
    when 16#00EBE# => romdata <= X"2B0772FC";
    when 16#00EBF# => romdata <= X"060C5151";
    when 16#00EC0# => romdata <= X"043C0472";
    when 16#00EC1# => romdata <= X"72807281";
    when 16#00EC2# => romdata <= X"06FF0509";
    when 16#00EC3# => romdata <= X"72060571";
    when 16#00EC4# => romdata <= X"1052720A";
    when 16#00EC5# => romdata <= X"100A5372";
    when 16#00EC6# => romdata <= X"ED385151";
    when 16#00EC7# => romdata <= X"535104B0";
    when 16#00EC8# => romdata <= X"08B408B8";
    when 16#00EC9# => romdata <= X"08757580";
    when 16#00ECA# => romdata <= X"F4B22D50";
    when 16#00ECB# => romdata <= X"50B00856";
    when 16#00ECC# => romdata <= X"B80CB40C";
    when 16#00ECD# => romdata <= X"B00C5104";
    when 16#00ECE# => romdata <= X"B008B408";
    when 16#00ECF# => romdata <= X"B8087575";
    when 16#00ED0# => romdata <= X"80F3EE2D";
    when 16#00ED1# => romdata <= X"5050B008";
    when 16#00ED2# => romdata <= X"56B80CB4";
    when 16#00ED3# => romdata <= X"0CB00C51";
    when 16#00ED4# => romdata <= X"04B008B4";
    when 16#00ED5# => romdata <= X"08B80880";
    when 16#00ED6# => romdata <= X"C5C52DB8";
    when 16#00ED7# => romdata <= X"0CB40CB0";
    when 16#00ED8# => romdata <= X"0C04FF3D";
    when 16#00ED9# => romdata <= X"0D028F05";
    when 16#00EDA# => romdata <= X"3381CD8C";
    when 16#00EDB# => romdata <= X"0852710C";
    when 16#00EDC# => romdata <= X"800BB00C";
    when 16#00EDD# => romdata <= X"833D0D04";
    when 16#00EDE# => romdata <= X"FF3D0D02";
    when 16#00EDF# => romdata <= X"8F053351";
    when 16#00EE0# => romdata <= X"81F0DC08";
    when 16#00EE1# => romdata <= X"52712DB0";
    when 16#00EE2# => romdata <= X"0881FF06";
    when 16#00EE3# => romdata <= X"B00C833D";
    when 16#00EE4# => romdata <= X"0D04FE3D";
    when 16#00EE5# => romdata <= X"0D747033";
    when 16#00EE6# => romdata <= X"53537180";
    when 16#00EE7# => romdata <= X"2E933881";
    when 16#00EE8# => romdata <= X"13725281";
    when 16#00EE9# => romdata <= X"F0DC0853";
    when 16#00EEA# => romdata <= X"53712D72";
    when 16#00EEB# => romdata <= X"335271EF";
    when 16#00EEC# => romdata <= X"38843D0D";
    when 16#00EED# => romdata <= X"04F43D0D";
    when 16#00EEE# => romdata <= X"7F028405";
    when 16#00EEF# => romdata <= X"BB053355";
    when 16#00EF0# => romdata <= X"57880B8C";
    when 16#00EF1# => romdata <= X"3D5B5989";
    when 16#00EF2# => romdata <= X"5381CAA4";
    when 16#00EF3# => romdata <= X"52795186";
    when 16#00EF4# => romdata <= X"923F7379";
    when 16#00EF5# => romdata <= X"2E80FF38";
    when 16#00EF6# => romdata <= X"78567390";
    when 16#00EF7# => romdata <= X"2E80EC38";
    when 16#00EF8# => romdata <= X"02A70558";
    when 16#00EF9# => romdata <= X"768F0654";
    when 16#00EFA# => romdata <= X"73892680";
    when 16#00EFB# => romdata <= X"C2387518";
    when 16#00EFC# => romdata <= X"B0155555";
    when 16#00EFD# => romdata <= X"73753476";
    when 16#00EFE# => romdata <= X"842AFF17";
    when 16#00EFF# => romdata <= X"7081FF06";
    when 16#00F00# => romdata <= X"58555775";
    when 16#00F01# => romdata <= X"DF38781A";
    when 16#00F02# => romdata <= X"55757534";
    when 16#00F03# => romdata <= X"79703355";
    when 16#00F04# => romdata <= X"5573802E";
    when 16#00F05# => romdata <= X"93388115";
    when 16#00F06# => romdata <= X"745281F0";
    when 16#00F07# => romdata <= X"DC085755";
    when 16#00F08# => romdata <= X"752D7433";
    when 16#00F09# => romdata <= X"5473EF38";
    when 16#00F0A# => romdata <= X"78B00C8E";
    when 16#00F0B# => romdata <= X"3D0D0475";
    when 16#00F0C# => romdata <= X"18B71555";
    when 16#00F0D# => romdata <= X"55737534";
    when 16#00F0E# => romdata <= X"76842AFF";
    when 16#00F0F# => romdata <= X"177081FF";
    when 16#00F10# => romdata <= X"06585557";
    when 16#00F11# => romdata <= X"75FF9D38";
    when 16#00F12# => romdata <= X"FFBC3984";
    when 16#00F13# => romdata <= X"70575902";
    when 16#00F14# => romdata <= X"A70558FF";
    when 16#00F15# => romdata <= X"8F398270";
    when 16#00F16# => romdata <= X"5759F439";
    when 16#00F17# => romdata <= X"F13D0D61";
    when 16#00F18# => romdata <= X"8D3D705B";
    when 16#00F19# => romdata <= X"5C5A807A";
    when 16#00F1A# => romdata <= X"5657767A";
    when 16#00F1B# => romdata <= X"24818538";
    when 16#00F1C# => romdata <= X"7817548A";
    when 16#00F1D# => romdata <= X"52745184";
    when 16#00F1E# => romdata <= X"B83FB008";
    when 16#00F1F# => romdata <= X"B0055372";
    when 16#00F20# => romdata <= X"74348117";
    when 16#00F21# => romdata <= X"578A5274";
    when 16#00F22# => romdata <= X"5184813F";
    when 16#00F23# => romdata <= X"B00855B0";
    when 16#00F24# => romdata <= X"08DE38B0";
    when 16#00F25# => romdata <= X"08779F2A";
    when 16#00F26# => romdata <= X"1870812C";
    when 16#00F27# => romdata <= X"5A565680";
    when 16#00F28# => romdata <= X"78259E38";
    when 16#00F29# => romdata <= X"7817FF05";
    when 16#00F2A# => romdata <= X"55751970";
    when 16#00F2B# => romdata <= X"33555374";
    when 16#00F2C# => romdata <= X"33733473";
    when 16#00F2D# => romdata <= X"75348116";
    when 16#00F2E# => romdata <= X"FF165656";
    when 16#00F2F# => romdata <= X"777624E9";
    when 16#00F30# => romdata <= X"38761958";
    when 16#00F31# => romdata <= X"80783480";
    when 16#00F32# => romdata <= X"7A241770";
    when 16#00F33# => romdata <= X"81FF067C";
    when 16#00F34# => romdata <= X"70335657";
    when 16#00F35# => romdata <= X"55567280";
    when 16#00F36# => romdata <= X"2E933881";
    when 16#00F37# => romdata <= X"15735281";
    when 16#00F38# => romdata <= X"F0DC0858";
    when 16#00F39# => romdata <= X"55762D74";
    when 16#00F3A# => romdata <= X"335372EF";
    when 16#00F3B# => romdata <= X"3873B00C";
    when 16#00F3C# => romdata <= X"913D0D04";
    when 16#00F3D# => romdata <= X"AD7B3402";
    when 16#00F3E# => romdata <= X"AD057A30";
    when 16#00F3F# => romdata <= X"71195656";
    when 16#00F40# => romdata <= X"598A5274";
    when 16#00F41# => romdata <= X"5183AA3F";
    when 16#00F42# => romdata <= X"B008B005";
    when 16#00F43# => romdata <= X"53727434";
    when 16#00F44# => romdata <= X"8117578A";
    when 16#00F45# => romdata <= X"52745182";
    when 16#00F46# => romdata <= X"F33FB008";
    when 16#00F47# => romdata <= X"55B008FE";
    when 16#00F48# => romdata <= X"CF38FEEF";
    when 16#00F49# => romdata <= X"39FD3D0D";
    when 16#00F4A# => romdata <= X"81CD8008";
    when 16#00F4B# => romdata <= X"76B2E429";
    when 16#00F4C# => romdata <= X"94120C54";
    when 16#00F4D# => romdata <= X"850B9815";
    when 16#00F4E# => romdata <= X"0C981408";
    when 16#00F4F# => romdata <= X"70810651";
    when 16#00F50# => romdata <= X"5372F638";
    when 16#00F51# => romdata <= X"853D0D04";
    when 16#00F52# => romdata <= X"803D0D81";
    when 16#00F53# => romdata <= X"CD800851";
    when 16#00F54# => romdata <= X"870B8412";
    when 16#00F55# => romdata <= X"0CFF0BA4";
    when 16#00F56# => romdata <= X"120CA70B";
    when 16#00F57# => romdata <= X"A8120CB2";
    when 16#00F58# => romdata <= X"E40B9412";
    when 16#00F59# => romdata <= X"0C870B98";
    when 16#00F5A# => romdata <= X"120C823D";
    when 16#00F5B# => romdata <= X"0D04803D";
    when 16#00F5C# => romdata <= X"0D81CD84";
    when 16#00F5D# => romdata <= X"0851B80B";
    when 16#00F5E# => romdata <= X"8C120C83";
    when 16#00F5F# => romdata <= X"0B88120C";
    when 16#00F60# => romdata <= X"823D0D04";
    when 16#00F61# => romdata <= X"803D0D81";
    when 16#00F62# => romdata <= X"CD840884";
    when 16#00F63# => romdata <= X"11088106";
    when 16#00F64# => romdata <= X"B00C5182";
    when 16#00F65# => romdata <= X"3D0D04FF";
    when 16#00F66# => romdata <= X"3D0D81CD";
    when 16#00F67# => romdata <= X"84085284";
    when 16#00F68# => romdata <= X"12087081";
    when 16#00F69# => romdata <= X"06515170";
    when 16#00F6A# => romdata <= X"802EF438";
    when 16#00F6B# => romdata <= X"71087081";
    when 16#00F6C# => romdata <= X"FF06B00C";
    when 16#00F6D# => romdata <= X"51833D0D";
    when 16#00F6E# => romdata <= X"04FE3D0D";
    when 16#00F6F# => romdata <= X"02930533";
    when 16#00F70# => romdata <= X"53728A2E";
    when 16#00F71# => romdata <= X"9C3881CD";
    when 16#00F72# => romdata <= X"84085284";
    when 16#00F73# => romdata <= X"12087089";
    when 16#00F74# => romdata <= X"2A708106";
    when 16#00F75# => romdata <= X"51515170";
    when 16#00F76# => romdata <= X"F2387272";
    when 16#00F77# => romdata <= X"0C843D0D";
    when 16#00F78# => romdata <= X"0481CD84";
    when 16#00F79# => romdata <= X"08528412";
    when 16#00F7A# => romdata <= X"0870892A";
    when 16#00F7B# => romdata <= X"70810651";
    when 16#00F7C# => romdata <= X"515170F2";
    when 16#00F7D# => romdata <= X"388D720C";
    when 16#00F7E# => romdata <= X"84120870";
    when 16#00F7F# => romdata <= X"892A7081";
    when 16#00F80# => romdata <= X"06515151";
    when 16#00F81# => romdata <= X"70C538D2";
    when 16#00F82# => romdata <= X"39FA3D0D";
    when 16#00F83# => romdata <= X"02A30533";
    when 16#00F84# => romdata <= X"81CCF808";
    when 16#00F85# => romdata <= X"81F0E033";
    when 16#00F86# => romdata <= X"7081FF06";
    when 16#00F87# => romdata <= X"70101011";
    when 16#00F88# => romdata <= X"81F0E433";
    when 16#00F89# => romdata <= X"7081FF06";
    when 16#00F8A# => romdata <= X"72902911";
    when 16#00F8B# => romdata <= X"70882B78";
    when 16#00F8C# => romdata <= X"07770C53";
    when 16#00F8D# => romdata <= X"5B5B5555";
    when 16#00F8E# => romdata <= X"59545473";
    when 16#00F8F# => romdata <= X"8A2E9838";
    when 16#00F90# => romdata <= X"7480CF2E";
    when 16#00F91# => romdata <= X"9238738C";
    when 16#00F92# => romdata <= X"2EA43881";
    when 16#00F93# => romdata <= X"16537281";
    when 16#00F94# => romdata <= X"F0E43488";
    when 16#00F95# => romdata <= X"3D0D0471";
    when 16#00F96# => romdata <= X"A326A338";
    when 16#00F97# => romdata <= X"81175271";
    when 16#00F98# => romdata <= X"81F0E034";
    when 16#00F99# => romdata <= X"800B81F0";
    when 16#00F9A# => romdata <= X"E434883D";
    when 16#00F9B# => romdata <= X"0D048052";
    when 16#00F9C# => romdata <= X"71882B73";
    when 16#00F9D# => romdata <= X"0C811252";
    when 16#00F9E# => romdata <= X"97907226";
    when 16#00F9F# => romdata <= X"F338800B";
    when 16#00FA0# => romdata <= X"81F0E034";
    when 16#00FA1# => romdata <= X"800B81F0";
    when 16#00FA2# => romdata <= X"E434DF39";
    when 16#00FA3# => romdata <= X"BC0802BC";
    when 16#00FA4# => romdata <= X"0CFD3D0D";
    when 16#00FA5# => romdata <= X"8053BC08";
    when 16#00FA6# => romdata <= X"8C050852";
    when 16#00FA7# => romdata <= X"BC088805";
    when 16#00FA8# => romdata <= X"0851F7C6";
    when 16#00FA9# => romdata <= X"3FB00870";
    when 16#00FAA# => romdata <= X"B00C5485";
    when 16#00FAB# => romdata <= X"3D0DBC0C";
    when 16#00FAC# => romdata <= X"04BC0802";
    when 16#00FAD# => romdata <= X"BC0CFD3D";
    when 16#00FAE# => romdata <= X"0D8153BC";
    when 16#00FAF# => romdata <= X"088C0508";
    when 16#00FB0# => romdata <= X"52BC0888";
    when 16#00FB1# => romdata <= X"050851F7";
    when 16#00FB2# => romdata <= X"A13FB008";
    when 16#00FB3# => romdata <= X"70B00C54";
    when 16#00FB4# => romdata <= X"853D0DBC";
    when 16#00FB5# => romdata <= X"0C04803D";
    when 16#00FB6# => romdata <= X"0D865184";
    when 16#00FB7# => romdata <= X"963F8151";
    when 16#00FB8# => romdata <= X"A1D33FFC";
    when 16#00FB9# => romdata <= X"3D0D7670";
    when 16#00FBA# => romdata <= X"797B5555";
    when 16#00FBB# => romdata <= X"55558F72";
    when 16#00FBC# => romdata <= X"278C3872";
    when 16#00FBD# => romdata <= X"75078306";
    when 16#00FBE# => romdata <= X"5170802E";
    when 16#00FBF# => romdata <= X"A738FF12";
    when 16#00FC0# => romdata <= X"5271FF2E";
    when 16#00FC1# => romdata <= X"98387270";
    when 16#00FC2# => romdata <= X"81055433";
    when 16#00FC3# => romdata <= X"74708105";
    when 16#00FC4# => romdata <= X"5634FF12";
    when 16#00FC5# => romdata <= X"5271FF2E";
    when 16#00FC6# => romdata <= X"098106EA";
    when 16#00FC7# => romdata <= X"3874B00C";
    when 16#00FC8# => romdata <= X"863D0D04";
    when 16#00FC9# => romdata <= X"74517270";
    when 16#00FCA# => romdata <= X"84055408";
    when 16#00FCB# => romdata <= X"71708405";
    when 16#00FCC# => romdata <= X"530C7270";
    when 16#00FCD# => romdata <= X"84055408";
    when 16#00FCE# => romdata <= X"71708405";
    when 16#00FCF# => romdata <= X"530C7270";
    when 16#00FD0# => romdata <= X"84055408";
    when 16#00FD1# => romdata <= X"71708405";
    when 16#00FD2# => romdata <= X"530C7270";
    when 16#00FD3# => romdata <= X"84055408";
    when 16#00FD4# => romdata <= X"71708405";
    when 16#00FD5# => romdata <= X"530CF012";
    when 16#00FD6# => romdata <= X"52718F26";
    when 16#00FD7# => romdata <= X"C9388372";
    when 16#00FD8# => romdata <= X"27953872";
    when 16#00FD9# => romdata <= X"70840554";
    when 16#00FDA# => romdata <= X"08717084";
    when 16#00FDB# => romdata <= X"05530CFC";
    when 16#00FDC# => romdata <= X"12527183";
    when 16#00FDD# => romdata <= X"26ED3870";
    when 16#00FDE# => romdata <= X"54FF8339";
    when 16#00FDF# => romdata <= X"FD3D0D75";
    when 16#00FE0# => romdata <= X"5384D813";
    when 16#00FE1# => romdata <= X"08802E8A";
    when 16#00FE2# => romdata <= X"38805372";
    when 16#00FE3# => romdata <= X"B00C853D";
    when 16#00FE4# => romdata <= X"0D048180";
    when 16#00FE5# => romdata <= X"5272518D";
    when 16#00FE6# => romdata <= X"9B3FB008";
    when 16#00FE7# => romdata <= X"84D8140C";
    when 16#00FE8# => romdata <= X"FF53B008";
    when 16#00FE9# => romdata <= X"802EE438";
    when 16#00FEA# => romdata <= X"B008549F";
    when 16#00FEB# => romdata <= X"53807470";
    when 16#00FEC# => romdata <= X"8405560C";
    when 16#00FED# => romdata <= X"FF135380";
    when 16#00FEE# => romdata <= X"7324CE38";
    when 16#00FEF# => romdata <= X"80747084";
    when 16#00FF0# => romdata <= X"05560CFF";
    when 16#00FF1# => romdata <= X"13537280";
    when 16#00FF2# => romdata <= X"25E338FF";
    when 16#00FF3# => romdata <= X"BC39FD3D";
    when 16#00FF4# => romdata <= X"0D757755";
    when 16#00FF5# => romdata <= X"539F7427";
    when 16#00FF6# => romdata <= X"8D389673";
    when 16#00FF7# => romdata <= X"0CFF5271";
    when 16#00FF8# => romdata <= X"B00C853D";
    when 16#00FF9# => romdata <= X"0D0484D8";
    when 16#00FFA# => romdata <= X"13085271";
    when 16#00FFB# => romdata <= X"802E9338";
    when 16#00FFC# => romdata <= X"73101012";
    when 16#00FFD# => romdata <= X"70087972";
    when 16#00FFE# => romdata <= X"0C515271";
    when 16#00FFF# => romdata <= X"B00C853D";
    when 16#01000# => romdata <= X"0D047251";
    when 16#01001# => romdata <= X"FEF63FFF";
    when 16#01002# => romdata <= X"52B008D3";
    when 16#01003# => romdata <= X"3884D813";
    when 16#01004# => romdata <= X"08741010";
    when 16#01005# => romdata <= X"1170087A";
    when 16#01006# => romdata <= X"720C5151";
    when 16#01007# => romdata <= X"52DD39F9";
    when 16#01008# => romdata <= X"3D0D797B";
    when 16#01009# => romdata <= X"5856769F";
    when 16#0100A# => romdata <= X"2680E838";
    when 16#0100B# => romdata <= X"84D81608";
    when 16#0100C# => romdata <= X"5473802E";
    when 16#0100D# => romdata <= X"AA387610";
    when 16#0100E# => romdata <= X"10147008";
    when 16#0100F# => romdata <= X"55557380";
    when 16#01010# => romdata <= X"2EBA3880";
    when 16#01011# => romdata <= X"5873812E";
    when 16#01012# => romdata <= X"8F3873FF";
    when 16#01013# => romdata <= X"2EA33880";
    when 16#01014# => romdata <= X"750C7651";
    when 16#01015# => romdata <= X"732D8058";
    when 16#01016# => romdata <= X"77B00C89";
    when 16#01017# => romdata <= X"3D0D0475";
    when 16#01018# => romdata <= X"51FE993F";
    when 16#01019# => romdata <= X"FF58B008";
    when 16#0101A# => romdata <= X"EF3884D8";
    when 16#0101B# => romdata <= X"160854C6";
    when 16#0101C# => romdata <= X"3996760C";
    when 16#0101D# => romdata <= X"810BB00C";
    when 16#0101E# => romdata <= X"893D0D04";
    when 16#0101F# => romdata <= X"755181ED";
    when 16#01020# => romdata <= X"3F7653B0";
    when 16#01021# => romdata <= X"08527551";
    when 16#01022# => romdata <= X"81AD3FB0";
    when 16#01023# => romdata <= X"08B00C89";
    when 16#01024# => romdata <= X"3D0D0496";
    when 16#01025# => romdata <= X"760CFF0B";
    when 16#01026# => romdata <= X"B00C893D";
    when 16#01027# => romdata <= X"0D04FC3D";
    when 16#01028# => romdata <= X"0D767856";
    when 16#01029# => romdata <= X"53FF5474";
    when 16#0102A# => romdata <= X"9F26B138";
    when 16#0102B# => romdata <= X"84D81308";
    when 16#0102C# => romdata <= X"5271802E";
    when 16#0102D# => romdata <= X"AE387410";
    when 16#0102E# => romdata <= X"10127008";
    when 16#0102F# => romdata <= X"53538154";
    when 16#01030# => romdata <= X"71802E98";
    when 16#01031# => romdata <= X"38825471";
    when 16#01032# => romdata <= X"FF2E9138";
    when 16#01033# => romdata <= X"83547181";
    when 16#01034# => romdata <= X"2E8A3880";
    when 16#01035# => romdata <= X"730C7451";
    when 16#01036# => romdata <= X"712D8054";
    when 16#01037# => romdata <= X"73B00C86";
    when 16#01038# => romdata <= X"3D0D0472";
    when 16#01039# => romdata <= X"51FD953F";
    when 16#0103A# => romdata <= X"B008F138";
    when 16#0103B# => romdata <= X"84D81308";
    when 16#0103C# => romdata <= X"52C439FF";
    when 16#0103D# => romdata <= X"3D0D7352";
    when 16#0103E# => romdata <= X"81CD9008";
    when 16#0103F# => romdata <= X"51FEA03F";
    when 16#01040# => romdata <= X"833D0D04";
    when 16#01041# => romdata <= X"FE3D0D75";
    when 16#01042# => romdata <= X"53745281";
    when 16#01043# => romdata <= X"CD900851";
    when 16#01044# => romdata <= X"FDBC3F84";
    when 16#01045# => romdata <= X"3D0D0480";
    when 16#01046# => romdata <= X"3D0D81CD";
    when 16#01047# => romdata <= X"900851FC";
    when 16#01048# => romdata <= X"DB3F823D";
    when 16#01049# => romdata <= X"0D04FF3D";
    when 16#0104A# => romdata <= X"0D735281";
    when 16#0104B# => romdata <= X"CD900851";
    when 16#0104C# => romdata <= X"FEEC3F83";
    when 16#0104D# => romdata <= X"3D0D04FC";
    when 16#0104E# => romdata <= X"3D0D800B";
    when 16#0104F# => romdata <= X"81F0EC0C";
    when 16#01050# => romdata <= X"78527751";
    when 16#01051# => romdata <= X"9CAA3FB0";
    when 16#01052# => romdata <= X"0854B008";
    when 16#01053# => romdata <= X"FF2E8838";
    when 16#01054# => romdata <= X"73B00C86";
    when 16#01055# => romdata <= X"3D0D0481";
    when 16#01056# => romdata <= X"F0EC0855";
    when 16#01057# => romdata <= X"74802EF0";
    when 16#01058# => romdata <= X"38767571";
    when 16#01059# => romdata <= X"0C5373B0";
    when 16#0105A# => romdata <= X"0C863D0D";
    when 16#0105B# => romdata <= X"049BFC3F";
    when 16#0105C# => romdata <= X"04FC3D0D";
    when 16#0105D# => romdata <= X"76707970";
    when 16#0105E# => romdata <= X"73078306";
    when 16#0105F# => romdata <= X"54545455";
    when 16#01060# => romdata <= X"7080C338";
    when 16#01061# => romdata <= X"71700870";
    when 16#01062# => romdata <= X"0970F7FB";
    when 16#01063# => romdata <= X"FDFF1306";
    when 16#01064# => romdata <= X"70F88482";
    when 16#01065# => romdata <= X"81800651";
    when 16#01066# => romdata <= X"51535354";
    when 16#01067# => romdata <= X"70A63884";
    when 16#01068# => romdata <= X"14727470";
    when 16#01069# => romdata <= X"8405560C";
    when 16#0106A# => romdata <= X"70087009";
    when 16#0106B# => romdata <= X"70F7FBFD";
    when 16#0106C# => romdata <= X"FF130670";
    when 16#0106D# => romdata <= X"F8848281";
    when 16#0106E# => romdata <= X"80065151";
    when 16#0106F# => romdata <= X"53535470";
    when 16#01070# => romdata <= X"802EDC38";
    when 16#01071# => romdata <= X"73527170";
    when 16#01072# => romdata <= X"81055333";
    when 16#01073# => romdata <= X"51707370";
    when 16#01074# => romdata <= X"81055534";
    when 16#01075# => romdata <= X"70F03874";
    when 16#01076# => romdata <= X"B00C863D";
    when 16#01077# => romdata <= X"0D04FD3D";
    when 16#01078# => romdata <= X"0D757071";
    when 16#01079# => romdata <= X"83065355";
    when 16#0107A# => romdata <= X"5270B838";
    when 16#0107B# => romdata <= X"71700870";
    when 16#0107C# => romdata <= X"09F7FBFD";
    when 16#0107D# => romdata <= X"FF120670";
    when 16#0107E# => romdata <= X"F8848281";
    when 16#0107F# => romdata <= X"80065151";
    when 16#01080# => romdata <= X"5253709D";
    when 16#01081# => romdata <= X"38841370";
    when 16#01082# => romdata <= X"087009F7";
    when 16#01083# => romdata <= X"FBFDFF12";
    when 16#01084# => romdata <= X"0670F884";
    when 16#01085# => romdata <= X"82818006";
    when 16#01086# => romdata <= X"51515253";
    when 16#01087# => romdata <= X"70802EE5";
    when 16#01088# => romdata <= X"38725271";
    when 16#01089# => romdata <= X"33517080";
    when 16#0108A# => romdata <= X"2E8A3881";
    when 16#0108B# => romdata <= X"12703352";
    when 16#0108C# => romdata <= X"5270F838";
    when 16#0108D# => romdata <= X"717431B0";
    when 16#0108E# => romdata <= X"0C853D0D";
    when 16#0108F# => romdata <= X"04FA3D0D";
    when 16#01090# => romdata <= X"787A7C70";
    when 16#01091# => romdata <= X"54555552";
    when 16#01092# => romdata <= X"72802E80";
    when 16#01093# => romdata <= X"D9387174";
    when 16#01094# => romdata <= X"07830651";
    when 16#01095# => romdata <= X"70802E80";
    when 16#01096# => romdata <= X"D438FF13";
    when 16#01097# => romdata <= X"5372FF2E";
    when 16#01098# => romdata <= X"B1387133";
    when 16#01099# => romdata <= X"74335651";
    when 16#0109A# => romdata <= X"74712E09";
    when 16#0109B# => romdata <= X"8106A938";
    when 16#0109C# => romdata <= X"72802E81";
    when 16#0109D# => romdata <= X"87387081";
    when 16#0109E# => romdata <= X"FF065170";
    when 16#0109F# => romdata <= X"802E80FC";
    when 16#010A0# => romdata <= X"38811281";
    when 16#010A1# => romdata <= X"15FF1555";
    when 16#010A2# => romdata <= X"555272FF";
    when 16#010A3# => romdata <= X"2E098106";
    when 16#010A4# => romdata <= X"D1387133";
    when 16#010A5# => romdata <= X"74335651";
    when 16#010A6# => romdata <= X"7081FF06";
    when 16#010A7# => romdata <= X"7581FF06";
    when 16#010A8# => romdata <= X"71713151";
    when 16#010A9# => romdata <= X"525270B0";
    when 16#010AA# => romdata <= X"0C883D0D";
    when 16#010AB# => romdata <= X"04717457";
    when 16#010AC# => romdata <= X"55837327";
    when 16#010AD# => romdata <= X"88387108";
    when 16#010AE# => romdata <= X"74082E88";
    when 16#010AF# => romdata <= X"38747655";
    when 16#010B0# => romdata <= X"52FF9739";
    when 16#010B1# => romdata <= X"FC135372";
    when 16#010B2# => romdata <= X"802EB138";
    when 16#010B3# => romdata <= X"74087009";
    when 16#010B4# => romdata <= X"F7FBFDFF";
    when 16#010B5# => romdata <= X"120670F8";
    when 16#010B6# => romdata <= X"84828180";
    when 16#010B7# => romdata <= X"06515151";
    when 16#010B8# => romdata <= X"709A3884";
    when 16#010B9# => romdata <= X"15841757";
    when 16#010BA# => romdata <= X"55837327";
    when 16#010BB# => romdata <= X"D0387408";
    when 16#010BC# => romdata <= X"76082ED0";
    when 16#010BD# => romdata <= X"38747655";
    when 16#010BE# => romdata <= X"52FEDF39";
    when 16#010BF# => romdata <= X"800BB00C";
    when 16#010C0# => romdata <= X"883D0D04";
    when 16#010C1# => romdata <= X"F33D0D60";
    when 16#010C2# => romdata <= X"6264725A";
    when 16#010C3# => romdata <= X"5A5E5E80";
    when 16#010C4# => romdata <= X"5C767081";
    when 16#010C5# => romdata <= X"05583381";
    when 16#010C6# => romdata <= X"CAB11133";
    when 16#010C7# => romdata <= X"70832A70";
    when 16#010C8# => romdata <= X"81065155";
    when 16#010C9# => romdata <= X"555672E9";
    when 16#010CA# => romdata <= X"3875AD2E";
    when 16#010CB# => romdata <= X"82883875";
    when 16#010CC# => romdata <= X"AB2E8284";
    when 16#010CD# => romdata <= X"38773070";
    when 16#010CE# => romdata <= X"79078025";
    when 16#010CF# => romdata <= X"79903270";
    when 16#010D0# => romdata <= X"30707207";
    when 16#010D1# => romdata <= X"80257307";
    when 16#010D2# => romdata <= X"53575751";
    when 16#010D3# => romdata <= X"5372802E";
    when 16#010D4# => romdata <= X"873875B0";
    when 16#010D5# => romdata <= X"2E81EB38";
    when 16#010D6# => romdata <= X"778A3888";
    when 16#010D7# => romdata <= X"5875B02E";
    when 16#010D8# => romdata <= X"83388A58";
    when 16#010D9# => romdata <= X"810A5A7B";
    when 16#010DA# => romdata <= X"8438FE0A";
    when 16#010DB# => romdata <= X"5A775279";
    when 16#010DC# => romdata <= X"51F6BE3F";
    when 16#010DD# => romdata <= X"B0087853";
    when 16#010DE# => romdata <= X"7A525BF6";
    when 16#010DF# => romdata <= X"8F3FB008";
    when 16#010E0# => romdata <= X"5A807081";
    when 16#010E1# => romdata <= X"CAB11833";
    when 16#010E2# => romdata <= X"70822A70";
    when 16#010E3# => romdata <= X"81065156";
    when 16#010E4# => romdata <= X"565A5572";
    when 16#010E5# => romdata <= X"802E80C1";
    when 16#010E6# => romdata <= X"38D01656";
    when 16#010E7# => romdata <= X"75782580";
    when 16#010E8# => romdata <= X"D7388079";
    when 16#010E9# => romdata <= X"24757B26";
    when 16#010EA# => romdata <= X"07537293";
    when 16#010EB# => romdata <= X"38747A2E";
    when 16#010EC# => romdata <= X"80EB387A";
    when 16#010ED# => romdata <= X"762580ED";
    when 16#010EE# => romdata <= X"3872802E";
    when 16#010EF# => romdata <= X"80E738FF";
    when 16#010F0# => romdata <= X"77708105";
    when 16#010F1# => romdata <= X"59335759";
    when 16#010F2# => romdata <= X"81CAB116";
    when 16#010F3# => romdata <= X"3370822A";
    when 16#010F4# => romdata <= X"70810651";
    when 16#010F5# => romdata <= X"545472C1";
    when 16#010F6# => romdata <= X"38738306";
    when 16#010F7# => romdata <= X"5372802E";
    when 16#010F8# => romdata <= X"97387381";
    when 16#010F9# => romdata <= X"06C91755";
    when 16#010FA# => romdata <= X"53728538";
    when 16#010FB# => romdata <= X"FFA91654";
    when 16#010FC# => romdata <= X"73567776";
    when 16#010FD# => romdata <= X"24FFAB38";
    when 16#010FE# => romdata <= X"80792480";
    when 16#010FF# => romdata <= X"F0387B80";
    when 16#01100# => romdata <= X"2E843874";
    when 16#01101# => romdata <= X"30557C80";
    when 16#01102# => romdata <= X"2E8C38FF";
    when 16#01103# => romdata <= X"17537883";
    when 16#01104# => romdata <= X"387D5372";
    when 16#01105# => romdata <= X"7D0C74B0";
    when 16#01106# => romdata <= X"0C8F3D0D";
    when 16#01107# => romdata <= X"04815375";
    when 16#01108# => romdata <= X"7B24FF95";
    when 16#01109# => romdata <= X"38817579";
    when 16#0110A# => romdata <= X"29177870";
    when 16#0110B# => romdata <= X"81055A33";
    when 16#0110C# => romdata <= X"585659FF";
    when 16#0110D# => romdata <= X"9339815C";
    when 16#0110E# => romdata <= X"76708105";
    when 16#0110F# => romdata <= X"583356FD";
    when 16#01110# => romdata <= X"F4398077";
    when 16#01111# => romdata <= X"33545472";
    when 16#01112# => romdata <= X"80F82EB2";
    when 16#01113# => romdata <= X"387280D8";
    when 16#01114# => romdata <= X"32703070";
    when 16#01115# => romdata <= X"80257607";
    when 16#01116# => romdata <= X"51515372";
    when 16#01117# => romdata <= X"802EFDF8";
    when 16#01118# => romdata <= X"38811733";
    when 16#01119# => romdata <= X"82185856";
    when 16#0111A# => romdata <= X"9058FDF8";
    when 16#0111B# => romdata <= X"39810A55";
    when 16#0111C# => romdata <= X"7B8438FE";
    when 16#0111D# => romdata <= X"0A557F53";
    when 16#0111E# => romdata <= X"A2730CFF";
    when 16#0111F# => romdata <= X"89398154";
    when 16#01120# => romdata <= X"CC39FD3D";
    when 16#01121# => romdata <= X"0D775476";
    when 16#01122# => romdata <= X"53755281";
    when 16#01123# => romdata <= X"CD900851";
    when 16#01124# => romdata <= X"FCF23F85";
    when 16#01125# => romdata <= X"3D0D04F3";
    when 16#01126# => romdata <= X"3D0D6062";
    when 16#01127# => romdata <= X"64725A5A";
    when 16#01128# => romdata <= X"5D5D805E";
    when 16#01129# => romdata <= X"76708105";
    when 16#0112A# => romdata <= X"583381CA";
    when 16#0112B# => romdata <= X"B1113370";
    when 16#0112C# => romdata <= X"832A7081";
    when 16#0112D# => romdata <= X"06515555";
    when 16#0112E# => romdata <= X"5672E938";
    when 16#0112F# => romdata <= X"75AD2E81";
    when 16#01130# => romdata <= X"FF3875AB";
    when 16#01131# => romdata <= X"2E81FB38";
    when 16#01132# => romdata <= X"77307079";
    when 16#01133# => romdata <= X"07802579";
    when 16#01134# => romdata <= X"90327030";
    when 16#01135# => romdata <= X"70720780";
    when 16#01136# => romdata <= X"25730753";
    when 16#01137# => romdata <= X"57575153";
    when 16#01138# => romdata <= X"72802E87";
    when 16#01139# => romdata <= X"3875B02E";
    when 16#0113A# => romdata <= X"81E23877";
    when 16#0113B# => romdata <= X"8A388858";
    when 16#0113C# => romdata <= X"75B02E83";
    when 16#0113D# => romdata <= X"388A5877";
    when 16#0113E# => romdata <= X"52FF51F3";
    when 16#0113F# => romdata <= X"8F3FB008";
    when 16#01140# => romdata <= X"78535AFF";
    when 16#01141# => romdata <= X"51F3AA3F";
    when 16#01142# => romdata <= X"B0085B80";
    when 16#01143# => romdata <= X"705A5581";
    when 16#01144# => romdata <= X"CAB11633";
    when 16#01145# => romdata <= X"70822A70";
    when 16#01146# => romdata <= X"81065154";
    when 16#01147# => romdata <= X"5472802E";
    when 16#01148# => romdata <= X"80C138D0";
    when 16#01149# => romdata <= X"16567578";
    when 16#0114A# => romdata <= X"2580D738";
    when 16#0114B# => romdata <= X"80792475";
    when 16#0114C# => romdata <= X"7B260753";
    when 16#0114D# => romdata <= X"72933874";
    when 16#0114E# => romdata <= X"7A2E80EB";
    when 16#0114F# => romdata <= X"387A7625";
    when 16#01150# => romdata <= X"80ED3872";
    when 16#01151# => romdata <= X"802E80E7";
    when 16#01152# => romdata <= X"38FF7770";
    when 16#01153# => romdata <= X"81055933";
    when 16#01154# => romdata <= X"575981CA";
    when 16#01155# => romdata <= X"B1163370";
    when 16#01156# => romdata <= X"822A7081";
    when 16#01157# => romdata <= X"06515454";
    when 16#01158# => romdata <= X"72C13873";
    when 16#01159# => romdata <= X"83065372";
    when 16#0115A# => romdata <= X"802E9738";
    when 16#0115B# => romdata <= X"738106C9";
    when 16#0115C# => romdata <= X"17555372";
    when 16#0115D# => romdata <= X"8538FFA9";
    when 16#0115E# => romdata <= X"16547356";
    when 16#0115F# => romdata <= X"777624FF";
    when 16#01160# => romdata <= X"AB388079";
    when 16#01161# => romdata <= X"24818938";
    when 16#01162# => romdata <= X"7D802E84";
    when 16#01163# => romdata <= X"38743055";
    when 16#01164# => romdata <= X"7B802E8C";
    when 16#01165# => romdata <= X"38FF1753";
    when 16#01166# => romdata <= X"7883387C";
    when 16#01167# => romdata <= X"53727C0C";
    when 16#01168# => romdata <= X"74B00C8F";
    when 16#01169# => romdata <= X"3D0D0481";
    when 16#0116A# => romdata <= X"53757B24";
    when 16#0116B# => romdata <= X"FF953881";
    when 16#0116C# => romdata <= X"75792917";
    when 16#0116D# => romdata <= X"78708105";
    when 16#0116E# => romdata <= X"5A335856";
    when 16#0116F# => romdata <= X"59FF9339";
    when 16#01170# => romdata <= X"815E7670";
    when 16#01171# => romdata <= X"81055833";
    when 16#01172# => romdata <= X"56FDFD39";
    when 16#01173# => romdata <= X"80773354";
    when 16#01174# => romdata <= X"547280F8";
    when 16#01175# => romdata <= X"2E80C338";
    when 16#01176# => romdata <= X"7280D832";
    when 16#01177# => romdata <= X"70307080";
    when 16#01178# => romdata <= X"25760751";
    when 16#01179# => romdata <= X"51537280";
    when 16#0117A# => romdata <= X"2EFE8038";
    when 16#0117B# => romdata <= X"81173382";
    when 16#0117C# => romdata <= X"18585690";
    when 16#0117D# => romdata <= X"705358FF";
    when 16#0117E# => romdata <= X"51F1913F";
    when 16#0117F# => romdata <= X"B0087853";
    when 16#01180# => romdata <= X"5AFF51F1";
    when 16#01181# => romdata <= X"AC3FB008";
    when 16#01182# => romdata <= X"5B80705A";
    when 16#01183# => romdata <= X"55FE8039";
    when 16#01184# => romdata <= X"FF605455";
    when 16#01185# => romdata <= X"A2730CFE";
    when 16#01186# => romdata <= X"F7398154";
    when 16#01187# => romdata <= X"FFBA39FD";
    when 16#01188# => romdata <= X"3D0D7754";
    when 16#01189# => romdata <= X"76537552";
    when 16#0118A# => romdata <= X"81CD9008";
    when 16#0118B# => romdata <= X"51FCE83F";
    when 16#0118C# => romdata <= X"853D0D04";
    when 16#0118D# => romdata <= X"F33D0D7F";
    when 16#0118E# => romdata <= X"618B1170";
    when 16#0118F# => romdata <= X"F8065C55";
    when 16#01190# => romdata <= X"555E7296";
    when 16#01191# => romdata <= X"26833890";
    when 16#01192# => romdata <= X"59807924";
    when 16#01193# => romdata <= X"747A2607";
    when 16#01194# => romdata <= X"53805472";
    when 16#01195# => romdata <= X"742E0981";
    when 16#01196# => romdata <= X"0680CB38";
    when 16#01197# => romdata <= X"7D518BCA";
    when 16#01198# => romdata <= X"3F7883F7";
    when 16#01199# => romdata <= X"2680C638";
    when 16#0119A# => romdata <= X"78832A70";
    when 16#0119B# => romdata <= X"10101081";
    when 16#0119C# => romdata <= X"D4CC058C";
    when 16#0119D# => romdata <= X"11085959";
    when 16#0119E# => romdata <= X"5A76782E";
    when 16#0119F# => romdata <= X"83B03884";
    when 16#011A0# => romdata <= X"1708FC06";
    when 16#011A1# => romdata <= X"568C1708";
    when 16#011A2# => romdata <= X"88180871";
    when 16#011A3# => romdata <= X"8C120C88";
    when 16#011A4# => romdata <= X"120C5875";
    when 16#011A5# => romdata <= X"17841108";
    when 16#011A6# => romdata <= X"81078412";
    when 16#011A7# => romdata <= X"0C537D51";
    when 16#011A8# => romdata <= X"8B893F88";
    when 16#011A9# => romdata <= X"175473B0";
    when 16#011AA# => romdata <= X"0C8F3D0D";
    when 16#011AB# => romdata <= X"0478892A";
    when 16#011AC# => romdata <= X"79832A5B";
    when 16#011AD# => romdata <= X"5372802E";
    when 16#011AE# => romdata <= X"BF387886";
    when 16#011AF# => romdata <= X"2AB8055A";
    when 16#011B0# => romdata <= X"847327B4";
    when 16#011B1# => romdata <= X"3880DB13";
    when 16#011B2# => romdata <= X"5A947327";
    when 16#011B3# => romdata <= X"AB38788C";
    when 16#011B4# => romdata <= X"2A80EE05";
    when 16#011B5# => romdata <= X"5A80D473";
    when 16#011B6# => romdata <= X"279E3878";
    when 16#011B7# => romdata <= X"8F2A80F7";
    when 16#011B8# => romdata <= X"055A82D4";
    when 16#011B9# => romdata <= X"73279138";
    when 16#011BA# => romdata <= X"78922A80";
    when 16#011BB# => romdata <= X"FC055A8A";
    when 16#011BC# => romdata <= X"D4732784";
    when 16#011BD# => romdata <= X"3880FE5A";
    when 16#011BE# => romdata <= X"79101010";
    when 16#011BF# => romdata <= X"81D4CC05";
    when 16#011C0# => romdata <= X"8C110858";
    when 16#011C1# => romdata <= X"5576752E";
    when 16#011C2# => romdata <= X"A3388417";
    when 16#011C3# => romdata <= X"08FC0670";
    when 16#011C4# => romdata <= X"7A315556";
    when 16#011C5# => romdata <= X"738F2488";
    when 16#011C6# => romdata <= X"D5387380";
    when 16#011C7# => romdata <= X"25FEE638";
    when 16#011C8# => romdata <= X"8C170857";
    when 16#011C9# => romdata <= X"76752E09";
    when 16#011CA# => romdata <= X"8106DF38";
    when 16#011CB# => romdata <= X"811A5A81";
    when 16#011CC# => romdata <= X"D4DC0857";
    when 16#011CD# => romdata <= X"7681D4D4";
    when 16#011CE# => romdata <= X"2E82C038";
    when 16#011CF# => romdata <= X"841708FC";
    when 16#011D0# => romdata <= X"06707A31";
    when 16#011D1# => romdata <= X"5556738F";
    when 16#011D2# => romdata <= X"2481F938";
    when 16#011D3# => romdata <= X"81D4D40B";
    when 16#011D4# => romdata <= X"81D4E00C";
    when 16#011D5# => romdata <= X"81D4D40B";
    when 16#011D6# => romdata <= X"81D4DC0C";
    when 16#011D7# => romdata <= X"738025FE";
    when 16#011D8# => romdata <= X"B23883FF";
    when 16#011D9# => romdata <= X"762783DF";
    when 16#011DA# => romdata <= X"3875892A";
    when 16#011DB# => romdata <= X"76832A55";
    when 16#011DC# => romdata <= X"5372802E";
    when 16#011DD# => romdata <= X"BF387586";
    when 16#011DE# => romdata <= X"2AB80554";
    when 16#011DF# => romdata <= X"847327B4";
    when 16#011E0# => romdata <= X"3880DB13";
    when 16#011E1# => romdata <= X"54947327";
    when 16#011E2# => romdata <= X"AB38758C";
    when 16#011E3# => romdata <= X"2A80EE05";
    when 16#011E4# => romdata <= X"5480D473";
    when 16#011E5# => romdata <= X"279E3875";
    when 16#011E6# => romdata <= X"8F2A80F7";
    when 16#011E7# => romdata <= X"055482D4";
    when 16#011E8# => romdata <= X"73279138";
    when 16#011E9# => romdata <= X"75922A80";
    when 16#011EA# => romdata <= X"FC05548A";
    when 16#011EB# => romdata <= X"D4732784";
    when 16#011EC# => romdata <= X"3880FE54";
    when 16#011ED# => romdata <= X"73101010";
    when 16#011EE# => romdata <= X"81D4CC05";
    when 16#011EF# => romdata <= X"88110856";
    when 16#011F0# => romdata <= X"5874782E";
    when 16#011F1# => romdata <= X"86CF3884";
    when 16#011F2# => romdata <= X"1508FC06";
    when 16#011F3# => romdata <= X"53757327";
    when 16#011F4# => romdata <= X"8D388815";
    when 16#011F5# => romdata <= X"08557478";
    when 16#011F6# => romdata <= X"2E098106";
    when 16#011F7# => romdata <= X"EA388C15";
    when 16#011F8# => romdata <= X"0881D4CC";
    when 16#011F9# => romdata <= X"0B840508";
    when 16#011FA# => romdata <= X"718C1A0C";
    when 16#011FB# => romdata <= X"76881A0C";
    when 16#011FC# => romdata <= X"7888130C";
    when 16#011FD# => romdata <= X"788C180C";
    when 16#011FE# => romdata <= X"5D587953";
    when 16#011FF# => romdata <= X"807A2483";
    when 16#01200# => romdata <= X"E6387282";
    when 16#01201# => romdata <= X"2C81712B";
    when 16#01202# => romdata <= X"5C537A7C";
    when 16#01203# => romdata <= X"26819838";
    when 16#01204# => romdata <= X"7B7B0653";
    when 16#01205# => romdata <= X"7282F138";
    when 16#01206# => romdata <= X"79FC0684";
    when 16#01207# => romdata <= X"055A7A10";
    when 16#01208# => romdata <= X"707D0654";
    when 16#01209# => romdata <= X"5B7282E0";
    when 16#0120A# => romdata <= X"38841A5A";
    when 16#0120B# => romdata <= X"F1398817";
    when 16#0120C# => romdata <= X"8C110858";
    when 16#0120D# => romdata <= X"5876782E";
    when 16#0120E# => romdata <= X"098106FC";
    when 16#0120F# => romdata <= X"C238821A";
    when 16#01210# => romdata <= X"5AFDEC39";
    when 16#01211# => romdata <= X"78177981";
    when 16#01212# => romdata <= X"0784190C";
    when 16#01213# => romdata <= X"7081D4E0";
    when 16#01214# => romdata <= X"0C7081D4";
    when 16#01215# => romdata <= X"DC0C81D4";
    when 16#01216# => romdata <= X"D40B8C12";
    when 16#01217# => romdata <= X"0C8C1108";
    when 16#01218# => romdata <= X"88120C74";
    when 16#01219# => romdata <= X"81078412";
    when 16#0121A# => romdata <= X"0C741175";
    when 16#0121B# => romdata <= X"710C5153";
    when 16#0121C# => romdata <= X"7D5187B7";
    when 16#0121D# => romdata <= X"3F881754";
    when 16#0121E# => romdata <= X"FCAC3981";
    when 16#0121F# => romdata <= X"D4CC0B84";
    when 16#01220# => romdata <= X"05087A54";
    when 16#01221# => romdata <= X"5C798025";
    when 16#01222# => romdata <= X"FEF83882";
    when 16#01223# => romdata <= X"DA397A09";
    when 16#01224# => romdata <= X"7C067081";
    when 16#01225# => romdata <= X"D4CC0B84";
    when 16#01226# => romdata <= X"050C5C7A";
    when 16#01227# => romdata <= X"105B7A7C";
    when 16#01228# => romdata <= X"2685387A";
    when 16#01229# => romdata <= X"85B83881";
    when 16#0122A# => romdata <= X"D4CC0B88";
    when 16#0122B# => romdata <= X"05087084";
    when 16#0122C# => romdata <= X"1208FC06";
    when 16#0122D# => romdata <= X"707C317C";
    when 16#0122E# => romdata <= X"72268F72";
    when 16#0122F# => romdata <= X"25075757";
    when 16#01230# => romdata <= X"5C5D5572";
    when 16#01231# => romdata <= X"802E80DB";
    when 16#01232# => romdata <= X"38797A16";
    when 16#01233# => romdata <= X"81D4C408";
    when 16#01234# => romdata <= X"1B90115A";
    when 16#01235# => romdata <= X"55575B81";
    when 16#01236# => romdata <= X"D4C008FF";
    when 16#01237# => romdata <= X"2E8838A0";
    when 16#01238# => romdata <= X"8F13E080";
    when 16#01239# => romdata <= X"06577652";
    when 16#0123A# => romdata <= X"7D5186C0";
    when 16#0123B# => romdata <= X"3FB00854";
    when 16#0123C# => romdata <= X"B008FF2E";
    when 16#0123D# => romdata <= X"9038B008";
    when 16#0123E# => romdata <= X"76278299";
    when 16#0123F# => romdata <= X"387481D4";
    when 16#01240# => romdata <= X"CC2E8291";
    when 16#01241# => romdata <= X"3881D4CC";
    when 16#01242# => romdata <= X"0B880508";
    when 16#01243# => romdata <= X"55841508";
    when 16#01244# => romdata <= X"FC06707A";
    when 16#01245# => romdata <= X"317A7226";
    when 16#01246# => romdata <= X"8F722507";
    when 16#01247# => romdata <= X"52555372";
    when 16#01248# => romdata <= X"83E63874";
    when 16#01249# => romdata <= X"79810784";
    when 16#0124A# => romdata <= X"170C7916";
    when 16#0124B# => romdata <= X"7081D4CC";
    when 16#0124C# => romdata <= X"0B88050C";
    when 16#0124D# => romdata <= X"75810784";
    when 16#0124E# => romdata <= X"120C547E";
    when 16#0124F# => romdata <= X"525785EB";
    when 16#01250# => romdata <= X"3F881754";
    when 16#01251# => romdata <= X"FAE03975";
    when 16#01252# => romdata <= X"832A7054";
    when 16#01253# => romdata <= X"54807424";
    when 16#01254# => romdata <= X"819B3872";
    when 16#01255# => romdata <= X"822C8171";
    when 16#01256# => romdata <= X"2B81D4D0";
    when 16#01257# => romdata <= X"08077081";
    when 16#01258# => romdata <= X"D4CC0B84";
    when 16#01259# => romdata <= X"050C7510";
    when 16#0125A# => romdata <= X"101081D4";
    when 16#0125B# => romdata <= X"CC058811";
    when 16#0125C# => romdata <= X"08585A5D";
    when 16#0125D# => romdata <= X"53778C18";
    when 16#0125E# => romdata <= X"0C748818";
    when 16#0125F# => romdata <= X"0C768819";
    when 16#01260# => romdata <= X"0C768C16";
    when 16#01261# => romdata <= X"0CFCF339";
    when 16#01262# => romdata <= X"797A1010";
    when 16#01263# => romdata <= X"1081D4CC";
    when 16#01264# => romdata <= X"05705759";
    when 16#01265# => romdata <= X"5D8C1508";
    when 16#01266# => romdata <= X"5776752E";
    when 16#01267# => romdata <= X"A3388417";
    when 16#01268# => romdata <= X"08FC0670";
    when 16#01269# => romdata <= X"7A315556";
    when 16#0126A# => romdata <= X"738F2483";
    when 16#0126B# => romdata <= X"CA387380";
    when 16#0126C# => romdata <= X"25848138";
    when 16#0126D# => romdata <= X"8C170857";
    when 16#0126E# => romdata <= X"76752E09";
    when 16#0126F# => romdata <= X"8106DF38";
    when 16#01270# => romdata <= X"8815811B";
    when 16#01271# => romdata <= X"70830655";
    when 16#01272# => romdata <= X"5B5572C9";
    when 16#01273# => romdata <= X"387C8306";
    when 16#01274# => romdata <= X"5372802E";
    when 16#01275# => romdata <= X"FDB838FF";
    when 16#01276# => romdata <= X"1DF81959";
    when 16#01277# => romdata <= X"5D881808";
    when 16#01278# => romdata <= X"782EEA38";
    when 16#01279# => romdata <= X"FDB53983";
    when 16#0127A# => romdata <= X"1A53FC96";
    when 16#0127B# => romdata <= X"39831470";
    when 16#0127C# => romdata <= X"822C8171";
    when 16#0127D# => romdata <= X"2B81D4D0";
    when 16#0127E# => romdata <= X"08077081";
    when 16#0127F# => romdata <= X"D4CC0B84";
    when 16#01280# => romdata <= X"050C7610";
    when 16#01281# => romdata <= X"101081D4";
    when 16#01282# => romdata <= X"CC058811";
    when 16#01283# => romdata <= X"08595B5E";
    when 16#01284# => romdata <= X"5153FEE1";
    when 16#01285# => romdata <= X"3981D490";
    when 16#01286# => romdata <= X"081758B0";
    when 16#01287# => romdata <= X"08762E81";
    when 16#01288# => romdata <= X"8D3881D4";
    when 16#01289# => romdata <= X"C008FF2E";
    when 16#0128A# => romdata <= X"83EC3873";
    when 16#0128B# => romdata <= X"76311881";
    when 16#0128C# => romdata <= X"D4900C73";
    when 16#0128D# => romdata <= X"87067057";
    when 16#0128E# => romdata <= X"5372802E";
    when 16#0128F# => romdata <= X"88388873";
    when 16#01290# => romdata <= X"31701555";
    when 16#01291# => romdata <= X"5676149F";
    when 16#01292# => romdata <= X"FF06A080";
    when 16#01293# => romdata <= X"71311770";
    when 16#01294# => romdata <= X"547F5357";
    when 16#01295# => romdata <= X"5383D53F";
    when 16#01296# => romdata <= X"B00853B0";
    when 16#01297# => romdata <= X"08FF2E81";
    when 16#01298# => romdata <= X"A03881D4";
    when 16#01299# => romdata <= X"90081670";
    when 16#0129A# => romdata <= X"81D4900C";
    when 16#0129B# => romdata <= X"747581D4";
    when 16#0129C# => romdata <= X"CC0B8805";
    when 16#0129D# => romdata <= X"0C747631";
    when 16#0129E# => romdata <= X"18708107";
    when 16#0129F# => romdata <= X"51555658";
    when 16#012A0# => romdata <= X"7B81D4CC";
    when 16#012A1# => romdata <= X"2E839C38";
    when 16#012A2# => romdata <= X"798F2682";
    when 16#012A3# => romdata <= X"CB38810B";
    when 16#012A4# => romdata <= X"84150C84";
    when 16#012A5# => romdata <= X"1508FC06";
    when 16#012A6# => romdata <= X"707A317A";
    when 16#012A7# => romdata <= X"72268F72";
    when 16#012A8# => romdata <= X"25075255";
    when 16#012A9# => romdata <= X"5372802E";
    when 16#012AA# => romdata <= X"FCF93880";
    when 16#012AB# => romdata <= X"DB39B008";
    when 16#012AC# => romdata <= X"9FFF0653";
    when 16#012AD# => romdata <= X"72FEEB38";
    when 16#012AE# => romdata <= X"7781D490";
    when 16#012AF# => romdata <= X"0C81D4CC";
    when 16#012B0# => romdata <= X"0B880508";
    when 16#012B1# => romdata <= X"7B188107";
    when 16#012B2# => romdata <= X"84120C55";
    when 16#012B3# => romdata <= X"81D4BC08";
    when 16#012B4# => romdata <= X"78278638";
    when 16#012B5# => romdata <= X"7781D4BC";
    when 16#012B6# => romdata <= X"0C81D4B8";
    when 16#012B7# => romdata <= X"087827FC";
    when 16#012B8# => romdata <= X"AC387781";
    when 16#012B9# => romdata <= X"D4B80C84";
    when 16#012BA# => romdata <= X"1508FC06";
    when 16#012BB# => romdata <= X"707A317A";
    when 16#012BC# => romdata <= X"72268F72";
    when 16#012BD# => romdata <= X"25075255";
    when 16#012BE# => romdata <= X"5372802E";
    when 16#012BF# => romdata <= X"FCA53888";
    when 16#012C0# => romdata <= X"39807454";
    when 16#012C1# => romdata <= X"56FEDB39";
    when 16#012C2# => romdata <= X"7D51829F";
    when 16#012C3# => romdata <= X"3F800BB0";
    when 16#012C4# => romdata <= X"0C8F3D0D";
    when 16#012C5# => romdata <= X"04735380";
    when 16#012C6# => romdata <= X"7424A938";
    when 16#012C7# => romdata <= X"72822C81";
    when 16#012C8# => romdata <= X"712B81D4";
    when 16#012C9# => romdata <= X"D0080770";
    when 16#012CA# => romdata <= X"81D4CC0B";
    when 16#012CB# => romdata <= X"84050C5D";
    when 16#012CC# => romdata <= X"53778C18";
    when 16#012CD# => romdata <= X"0C748818";
    when 16#012CE# => romdata <= X"0C768819";
    when 16#012CF# => romdata <= X"0C768C16";
    when 16#012D0# => romdata <= X"0CF9B739";
    when 16#012D1# => romdata <= X"83147082";
    when 16#012D2# => romdata <= X"2C81712B";
    when 16#012D3# => romdata <= X"81D4D008";
    when 16#012D4# => romdata <= X"077081D4";
    when 16#012D5# => romdata <= X"CC0B8405";
    when 16#012D6# => romdata <= X"0C5E5153";
    when 16#012D7# => romdata <= X"D4397B7B";
    when 16#012D8# => romdata <= X"065372FC";
    when 16#012D9# => romdata <= X"A338841A";
    when 16#012DA# => romdata <= X"7B105C5A";
    when 16#012DB# => romdata <= X"F139FF1A";
    when 16#012DC# => romdata <= X"8111515A";
    when 16#012DD# => romdata <= X"F7B93978";
    when 16#012DE# => romdata <= X"17798107";
    when 16#012DF# => romdata <= X"84190C8C";
    when 16#012E0# => romdata <= X"18088819";
    when 16#012E1# => romdata <= X"08718C12";
    when 16#012E2# => romdata <= X"0C88120C";
    when 16#012E3# => romdata <= X"597081D4";
    when 16#012E4# => romdata <= X"E00C7081";
    when 16#012E5# => romdata <= X"D4DC0C81";
    when 16#012E6# => romdata <= X"D4D40B8C";
    when 16#012E7# => romdata <= X"120C8C11";
    when 16#012E8# => romdata <= X"0888120C";
    when 16#012E9# => romdata <= X"74810784";
    when 16#012EA# => romdata <= X"120C7411";
    when 16#012EB# => romdata <= X"75710C51";
    when 16#012EC# => romdata <= X"53F9BD39";
    when 16#012ED# => romdata <= X"75178411";
    when 16#012EE# => romdata <= X"08810784";
    when 16#012EF# => romdata <= X"120C538C";
    when 16#012F0# => romdata <= X"17088818";
    when 16#012F1# => romdata <= X"08718C12";
    when 16#012F2# => romdata <= X"0C88120C";
    when 16#012F3# => romdata <= X"587D5180";
    when 16#012F4# => romdata <= X"DA3F8817";
    when 16#012F5# => romdata <= X"54F5CF39";
    when 16#012F6# => romdata <= X"7284150C";
    when 16#012F7# => romdata <= X"F41AF806";
    when 16#012F8# => romdata <= X"70841E08";
    when 16#012F9# => romdata <= X"81060784";
    when 16#012FA# => romdata <= X"1E0C701D";
    when 16#012FB# => romdata <= X"545B850B";
    when 16#012FC# => romdata <= X"84140C85";
    when 16#012FD# => romdata <= X"0B88140C";
    when 16#012FE# => romdata <= X"8F7B27FD";
    when 16#012FF# => romdata <= X"CF38881C";
    when 16#01300# => romdata <= X"527D5182";
    when 16#01301# => romdata <= X"903F81D4";
    when 16#01302# => romdata <= X"CC0B8805";
    when 16#01303# => romdata <= X"0881D490";
    when 16#01304# => romdata <= X"085955FD";
    when 16#01305# => romdata <= X"B7397781";
    when 16#01306# => romdata <= X"D4900C73";
    when 16#01307# => romdata <= X"81D4C00C";
    when 16#01308# => romdata <= X"FC913972";
    when 16#01309# => romdata <= X"84150CFD";
    when 16#0130A# => romdata <= X"A3390404";
    when 16#0130B# => romdata <= X"FD3D0D80";
    when 16#0130C# => romdata <= X"0B81F0EC";
    when 16#0130D# => romdata <= X"0C765186";
    when 16#0130E# => romdata <= X"CB3FB008";
    when 16#0130F# => romdata <= X"53B008FF";
    when 16#01310# => romdata <= X"2E883872";
    when 16#01311# => romdata <= X"B00C853D";
    when 16#01312# => romdata <= X"0D0481F0";
    when 16#01313# => romdata <= X"EC085473";
    when 16#01314# => romdata <= X"802EF038";
    when 16#01315# => romdata <= X"7574710C";
    when 16#01316# => romdata <= X"5272B00C";
    when 16#01317# => romdata <= X"853D0D04";
    when 16#01318# => romdata <= X"FB3D0D77";
    when 16#01319# => romdata <= X"705256C2";
    when 16#0131A# => romdata <= X"3F81D4CC";
    when 16#0131B# => romdata <= X"0B880508";
    when 16#0131C# => romdata <= X"841108FC";
    when 16#0131D# => romdata <= X"06707B31";
    when 16#0131E# => romdata <= X"9FEF05E0";
    when 16#0131F# => romdata <= X"8006E080";
    when 16#01320# => romdata <= X"05565653";
    when 16#01321# => romdata <= X"A0807424";
    when 16#01322# => romdata <= X"94388052";
    when 16#01323# => romdata <= X"7551FF9C";
    when 16#01324# => romdata <= X"3F81D4D4";
    when 16#01325# => romdata <= X"08155372";
    when 16#01326# => romdata <= X"B0082E8F";
    when 16#01327# => romdata <= X"387551FF";
    when 16#01328# => romdata <= X"8A3F8053";
    when 16#01329# => romdata <= X"72B00C87";
    when 16#0132A# => romdata <= X"3D0D0473";
    when 16#0132B# => romdata <= X"30527551";
    when 16#0132C# => romdata <= X"FEFA3FB0";
    when 16#0132D# => romdata <= X"08FF2EA8";
    when 16#0132E# => romdata <= X"3881D4CC";
    when 16#0132F# => romdata <= X"0B880508";
    when 16#01330# => romdata <= X"75753181";
    when 16#01331# => romdata <= X"0784120C";
    when 16#01332# => romdata <= X"5381D490";
    when 16#01333# => romdata <= X"08743181";
    when 16#01334# => romdata <= X"D4900C75";
    when 16#01335# => romdata <= X"51FED43F";
    when 16#01336# => romdata <= X"810BB00C";
    when 16#01337# => romdata <= X"873D0D04";
    when 16#01338# => romdata <= X"80527551";
    when 16#01339# => romdata <= X"FEC63F81";
    when 16#0133A# => romdata <= X"D4CC0B88";
    when 16#0133B# => romdata <= X"0508B008";
    when 16#0133C# => romdata <= X"71315653";
    when 16#0133D# => romdata <= X"8F7525FF";
    when 16#0133E# => romdata <= X"A438B008";
    when 16#0133F# => romdata <= X"81D4C008";
    when 16#01340# => romdata <= X"3181D490";
    when 16#01341# => romdata <= X"0C748107";
    when 16#01342# => romdata <= X"84140C75";
    when 16#01343# => romdata <= X"51FE9C3F";
    when 16#01344# => romdata <= X"8053FF90";
    when 16#01345# => romdata <= X"39F63D0D";
    when 16#01346# => romdata <= X"7C7E545B";
    when 16#01347# => romdata <= X"72802E82";
    when 16#01348# => romdata <= X"83387A51";
    when 16#01349# => romdata <= X"FE843FF8";
    when 16#0134A# => romdata <= X"13841108";
    when 16#0134B# => romdata <= X"70FE0670";
    when 16#0134C# => romdata <= X"13841108";
    when 16#0134D# => romdata <= X"FC065D58";
    when 16#0134E# => romdata <= X"59545881";
    when 16#0134F# => romdata <= X"D4D40875";
    when 16#01350# => romdata <= X"2E82DE38";
    when 16#01351# => romdata <= X"7884160C";
    when 16#01352# => romdata <= X"80738106";
    when 16#01353# => romdata <= X"545A727A";
    when 16#01354# => romdata <= X"2E81D538";
    when 16#01355# => romdata <= X"78158411";
    when 16#01356# => romdata <= X"08810651";
    when 16#01357# => romdata <= X"5372A038";
    when 16#01358# => romdata <= X"78175779";
    when 16#01359# => romdata <= X"81E63888";
    when 16#0135A# => romdata <= X"15085372";
    when 16#0135B# => romdata <= X"81D4D42E";
    when 16#0135C# => romdata <= X"82F9388C";
    when 16#0135D# => romdata <= X"1508708C";
    when 16#0135E# => romdata <= X"150C7388";
    when 16#0135F# => romdata <= X"120C5676";
    when 16#01360# => romdata <= X"81078419";
    when 16#01361# => romdata <= X"0C761877";
    when 16#01362# => romdata <= X"710C5379";
    when 16#01363# => romdata <= X"81913883";
    when 16#01364# => romdata <= X"FF772781";
    when 16#01365# => romdata <= X"C8387689";
    when 16#01366# => romdata <= X"2A77832A";
    when 16#01367# => romdata <= X"56537280";
    when 16#01368# => romdata <= X"2EBF3876";
    when 16#01369# => romdata <= X"862AB805";
    when 16#0136A# => romdata <= X"55847327";
    when 16#0136B# => romdata <= X"B43880DB";
    when 16#0136C# => romdata <= X"13559473";
    when 16#0136D# => romdata <= X"27AB3876";
    when 16#0136E# => romdata <= X"8C2A80EE";
    when 16#0136F# => romdata <= X"055580D4";
    when 16#01370# => romdata <= X"73279E38";
    when 16#01371# => romdata <= X"768F2A80";
    when 16#01372# => romdata <= X"F7055582";
    when 16#01373# => romdata <= X"D4732791";
    when 16#01374# => romdata <= X"3876922A";
    when 16#01375# => romdata <= X"80FC0555";
    when 16#01376# => romdata <= X"8AD47327";
    when 16#01377# => romdata <= X"843880FE";
    when 16#01378# => romdata <= X"55741010";
    when 16#01379# => romdata <= X"1081D4CC";
    when 16#0137A# => romdata <= X"05881108";
    when 16#0137B# => romdata <= X"55567376";
    when 16#0137C# => romdata <= X"2E82B338";
    when 16#0137D# => romdata <= X"841408FC";
    when 16#0137E# => romdata <= X"06537673";
    when 16#0137F# => romdata <= X"278D3888";
    when 16#01380# => romdata <= X"14085473";
    when 16#01381# => romdata <= X"762E0981";
    when 16#01382# => romdata <= X"06EA388C";
    when 16#01383# => romdata <= X"1408708C";
    when 16#01384# => romdata <= X"1A0C7488";
    when 16#01385# => romdata <= X"1A0C7888";
    when 16#01386# => romdata <= X"120C5677";
    when 16#01387# => romdata <= X"8C150C7A";
    when 16#01388# => romdata <= X"51FC883F";
    when 16#01389# => romdata <= X"8C3D0D04";
    when 16#0138A# => romdata <= X"77087871";
    when 16#0138B# => romdata <= X"31597705";
    when 16#0138C# => romdata <= X"88190854";
    when 16#0138D# => romdata <= X"577281D4";
    when 16#0138E# => romdata <= X"D42E80E0";
    when 16#0138F# => romdata <= X"388C1808";
    when 16#01390# => romdata <= X"708C150C";
    when 16#01391# => romdata <= X"7388120C";
    when 16#01392# => romdata <= X"56FE8939";
    when 16#01393# => romdata <= X"8815088C";
    when 16#01394# => romdata <= X"1608708C";
    when 16#01395# => romdata <= X"130C5788";
    when 16#01396# => romdata <= X"170CFEA3";
    when 16#01397# => romdata <= X"3976832A";
    when 16#01398# => romdata <= X"70545580";
    when 16#01399# => romdata <= X"75248198";
    when 16#0139A# => romdata <= X"3872822C";
    when 16#0139B# => romdata <= X"81712B81";
    when 16#0139C# => romdata <= X"D4D00807";
    when 16#0139D# => romdata <= X"81D4CC0B";
    when 16#0139E# => romdata <= X"84050C53";
    when 16#0139F# => romdata <= X"74101010";
    when 16#013A0# => romdata <= X"81D4CC05";
    when 16#013A1# => romdata <= X"88110855";
    when 16#013A2# => romdata <= X"56758C19";
    when 16#013A3# => romdata <= X"0C738819";
    when 16#013A4# => romdata <= X"0C778817";
    when 16#013A5# => romdata <= X"0C778C15";
    when 16#013A6# => romdata <= X"0CFF8439";
    when 16#013A7# => romdata <= X"815AFDB4";
    when 16#013A8# => romdata <= X"39781773";
    when 16#013A9# => romdata <= X"81065457";
    when 16#013AA# => romdata <= X"72983877";
    when 16#013AB# => romdata <= X"08787131";
    when 16#013AC# => romdata <= X"5977058C";
    when 16#013AD# => romdata <= X"1908881A";
    when 16#013AE# => romdata <= X"08718C12";
    when 16#013AF# => romdata <= X"0C88120C";
    when 16#013B0# => romdata <= X"57577681";
    when 16#013B1# => romdata <= X"0784190C";
    when 16#013B2# => romdata <= X"7781D4CC";
    when 16#013B3# => romdata <= X"0B88050C";
    when 16#013B4# => romdata <= X"81D4C808";
    when 16#013B5# => romdata <= X"7726FEC7";
    when 16#013B6# => romdata <= X"3881D4C4";
    when 16#013B7# => romdata <= X"08527A51";
    when 16#013B8# => romdata <= X"FAFE3F7A";
    when 16#013B9# => romdata <= X"51FAC43F";
    when 16#013BA# => romdata <= X"FEBA3981";
    when 16#013BB# => romdata <= X"788C150C";
    when 16#013BC# => romdata <= X"7888150C";
    when 16#013BD# => romdata <= X"738C1A0C";
    when 16#013BE# => romdata <= X"73881A0C";
    when 16#013BF# => romdata <= X"5AFD8039";
    when 16#013C0# => romdata <= X"83157082";
    when 16#013C1# => romdata <= X"2C81712B";
    when 16#013C2# => romdata <= X"81D4D008";
    when 16#013C3# => romdata <= X"0781D4CC";
    when 16#013C4# => romdata <= X"0B84050C";
    when 16#013C5# => romdata <= X"51537410";
    when 16#013C6# => romdata <= X"101081D4";
    when 16#013C7# => romdata <= X"CC058811";
    when 16#013C8# => romdata <= X"085556FE";
    when 16#013C9# => romdata <= X"E4397453";
    when 16#013CA# => romdata <= X"807524A7";
    when 16#013CB# => romdata <= X"3872822C";
    when 16#013CC# => romdata <= X"81712B81";
    when 16#013CD# => romdata <= X"D4D00807";
    when 16#013CE# => romdata <= X"81D4CC0B";
    when 16#013CF# => romdata <= X"84050C53";
    when 16#013D0# => romdata <= X"758C190C";
    when 16#013D1# => romdata <= X"7388190C";
    when 16#013D2# => romdata <= X"7788170C";
    when 16#013D3# => romdata <= X"778C150C";
    when 16#013D4# => romdata <= X"FDCD3983";
    when 16#013D5# => romdata <= X"1570822C";
    when 16#013D6# => romdata <= X"81712B81";
    when 16#013D7# => romdata <= X"D4D00807";
    when 16#013D8# => romdata <= X"81D4CC0B";
    when 16#013D9# => romdata <= X"84050C51";
    when 16#013DA# => romdata <= X"53D63981";
    when 16#013DB# => romdata <= X"0BB00C04";
    when 16#013DC# => romdata <= X"803D0D72";
    when 16#013DD# => romdata <= X"812E8938";
    when 16#013DE# => romdata <= X"800BB00C";
    when 16#013DF# => romdata <= X"823D0D04";
    when 16#013E0# => romdata <= X"7351B23F";
    when 16#013E1# => romdata <= X"FE3D0D81";
    when 16#013E2# => romdata <= X"F0E80851";
    when 16#013E3# => romdata <= X"708A3881";
    when 16#013E4# => romdata <= X"F0F07081";
    when 16#013E5# => romdata <= X"F0E80C51";
    when 16#013E6# => romdata <= X"70751252";
    when 16#013E7# => romdata <= X"52FF5370";
    when 16#013E8# => romdata <= X"87FB8080";
    when 16#013E9# => romdata <= X"26883870";
    when 16#013EA# => romdata <= X"81F0E80C";
    when 16#013EB# => romdata <= X"715372B0";
    when 16#013EC# => romdata <= X"0C843D0D";
    when 16#013ED# => romdata <= X"0400FF39";
    when 16#013EE# => romdata <= X"00000000";
    when 16#013EF# => romdata <= X"00000000";
    when 16#013F0# => romdata <= X"00000000";
    when 16#013F1# => romdata <= X"00000000";
    when 16#013F2# => romdata <= X"00CAC5CA";
    when 16#013F3# => romdata <= X"C5C0C0C0";
    when 16#013F4# => romdata <= X"C0C0C0C0";
    when 16#013F5# => romdata <= X"C0C0C0CF";
    when 16#013F6# => romdata <= X"CFCFCF00";
    when 16#013F7# => romdata <= X"00000F0F";
    when 16#013F8# => romdata <= X"0F0F8F8F";
    when 16#013F9# => romdata <= X"CFCFCFCF";
    when 16#013FA# => romdata <= X"CFCF4F0F";
    when 16#013FB# => romdata <= X"0F0F0000";
    when 16#013FC# => romdata <= X"CFCFCFCF";
    when 16#013FD# => romdata <= X"0F0F0F0F";
    when 16#013FE# => romdata <= X"0F0F0F0F";
    when 16#013FF# => romdata <= X"0F0FFEFE";
    when 16#01400# => romdata <= X"FEFC0000";
    when 16#01401# => romdata <= X"CFCFCFCF";
    when 16#01402# => romdata <= X"CFCFCFCF";
    when 16#01403# => romdata <= X"CFCFCFCF";
    when 16#01404# => romdata <= X"CFFFFF7E";
    when 16#01405# => romdata <= X"7E000000";
    when 16#01406# => romdata <= X"00000000";
    when 16#01407# => romdata <= X"00000000";
    when 16#01408# => romdata <= X"00000000";
    when 16#01409# => romdata <= X"00003F3F";
    when 16#0140A# => romdata <= X"3F3F0101";
    when 16#0140B# => romdata <= X"01010101";
    when 16#0140C# => romdata <= X"01010101";
    when 16#0140D# => romdata <= X"3F3F3F3F";
    when 16#0140E# => romdata <= X"0000383C";
    when 16#0140F# => romdata <= X"3E3E3F3F";
    when 16#01410# => romdata <= X"3F3B3B39";
    when 16#01411# => romdata <= X"39383838";
    when 16#01412# => romdata <= X"38383800";
    when 16#01413# => romdata <= X"003F3F3F";
    when 16#01414# => romdata <= X"3F383838";
    when 16#01415# => romdata <= X"38383838";
    when 16#01416# => romdata <= X"38383C3F";
    when 16#01417# => romdata <= X"3F1F0F00";
    when 16#01418# => romdata <= X"003F3F3F";
    when 16#01419# => romdata <= X"3F030303";
    when 16#0141A# => romdata <= X"03030303";
    when 16#0141B# => romdata <= X"03033F3F";
    when 16#0141C# => romdata <= X"3F3E0000";
    when 16#0141D# => romdata <= X"00000000";
    when 16#0141E# => romdata <= X"00000000";
    when 16#0141F# => romdata <= X"00000000";
    when 16#01420# => romdata <= X"00000000";
    when 16#01421# => romdata <= X"00000000";
    when 16#01422# => romdata <= X"00000000";
    when 16#01423# => romdata <= X"00000000";
    when 16#01424# => romdata <= X"00000000";
    when 16#01425# => romdata <= X"00000000";
    when 16#01426# => romdata <= X"00000000";
    when 16#01427# => romdata <= X"00000000";
    when 16#01428# => romdata <= X"00000000";
    when 16#01429# => romdata <= X"00000000";
    when 16#0142A# => romdata <= X"00000000";
    when 16#0142B# => romdata <= X"00000000";
    when 16#0142C# => romdata <= X"00000000";
    when 16#0142D# => romdata <= X"00000000";
    when 16#0142E# => romdata <= X"00000000";
    when 16#0142F# => romdata <= X"00000000";
    when 16#01430# => romdata <= X"00000000";
    when 16#01431# => romdata <= X"00000000";
    when 16#01432# => romdata <= X"00000000";
    when 16#01433# => romdata <= X"00000000";
    when 16#01434# => romdata <= X"00000000";
    when 16#01435# => romdata <= X"8080C0C0";
    when 16#01436# => romdata <= X"E0E06000";
    when 16#01437# => romdata <= X"00000000";
    when 16#01438# => romdata <= X"00000000";
    when 16#01439# => romdata <= X"00000000";
    when 16#0143A# => romdata <= X"00000000";
    when 16#0143B# => romdata <= X"00000000";
    when 16#0143C# => romdata <= X"00000000";
    when 16#0143D# => romdata <= X"00000000";
    when 16#0143E# => romdata <= X"00000000";
    when 16#0143F# => romdata <= X"00000000";
    when 16#01440# => romdata <= X"00000000";
    when 16#01441# => romdata <= X"00000000";
    when 16#01442# => romdata <= X"00000000";
    when 16#01443# => romdata <= X"00000000";
    when 16#01444# => romdata <= X"00000000";
    when 16#01445# => romdata <= X"00000000";
    when 16#01446# => romdata <= X"00000000";
    when 16#01447# => romdata <= X"00000000";
    when 16#01448# => romdata <= X"00000000";
    when 16#01449# => romdata <= X"00000000";
    when 16#0144A# => romdata <= X"00000000";
    when 16#0144B# => romdata <= X"806098EE";
    when 16#0144C# => romdata <= X"77BBDDEC";
    when 16#0144D# => romdata <= X"EE6E0200";
    when 16#0144E# => romdata <= X"00000000";
    when 16#0144F# => romdata <= X"00E08080";
    when 16#01450# => romdata <= X"E00000E0";
    when 16#01451# => romdata <= X"A0A00000";
    when 16#01452# => romdata <= X"E0000000";
    when 16#01453# => romdata <= X"00E0C000";
    when 16#01454# => romdata <= X"C0E00000";
    when 16#01455# => romdata <= X"E08080E0";
    when 16#01456# => romdata <= X"0000C020";
    when 16#01457# => romdata <= X"20C00000";
    when 16#01458# => romdata <= X"E0000000";
    when 16#01459# => romdata <= X"20E02000";
    when 16#0145A# => romdata <= X"0020A060";
    when 16#0145B# => romdata <= X"20000000";
    when 16#0145C# => romdata <= X"00000000";
    when 16#0145D# => romdata <= X"00000000";
    when 16#0145E# => romdata <= X"00000000";
    when 16#0145F# => romdata <= X"00000000";
    when 16#01460# => romdata <= X"00000000";
    when 16#01461# => romdata <= X"00000000";
    when 16#01462# => romdata <= X"00030007";
    when 16#01463# => romdata <= X"00070701";
    when 16#01464# => romdata <= X"00000000";
    when 16#01465# => romdata <= X"00000000";
    when 16#01466# => romdata <= X"00000300";
    when 16#01467# => romdata <= X"C0030000";
    when 16#01468# => romdata <= X"034242C0";
    when 16#01469# => romdata <= X"00C34242";
    when 16#0146A# => romdata <= X"0000C380";
    when 16#0146B# => romdata <= X"01C00340";
    when 16#0146C# => romdata <= X"C04300C0";
    when 16#0146D# => romdata <= X"43408001";
    when 16#0146E# => romdata <= X"C20201C0";
    when 16#0146F# => romdata <= X"00C38202";
    when 16#01470# => romdata <= X"80C00300";
    when 16#01471# => romdata <= X"00C04342";
    when 16#01472# => romdata <= X"8202C040";
    when 16#01473# => romdata <= X"40800000";
    when 16#01474# => romdata <= X"C0404000";
    when 16#01475# => romdata <= X"80404000";
    when 16#01476# => romdata <= X"00C04040";
    when 16#01477# => romdata <= X"8000C040";
    when 16#01478# => romdata <= X"4000C080";
    when 16#01479# => romdata <= X"00C00000";
    when 16#0147A# => romdata <= X"00000000";
    when 16#0147B# => romdata <= X"00000000";
    when 16#0147C# => romdata <= X"00000000";
    when 16#0147D# => romdata <= X"00000000";
    when 16#0147E# => romdata <= X"00FF0000";
    when 16#0147F# => romdata <= X"0000C645";
    when 16#01480# => romdata <= X"44800785";
    when 16#01481# => romdata <= X"45408007";
    when 16#01482# => romdata <= X"80424700";
    when 16#01483# => romdata <= X"80474000";
    when 16#01484# => romdata <= X"07C14344";
    when 16#01485# => romdata <= X"00C38404";
    when 16#01486# => romdata <= X"C30007C1";
    when 16#01487# => romdata <= X"42418700";
    when 16#01488# => romdata <= X"80404784";
    when 16#01489# => romdata <= X"04C34047";
    when 16#0148A# => romdata <= X"8101C640";
    when 16#0148B# => romdata <= X"40070505";
    when 16#0148C# => romdata <= X"00040502";
    when 16#0148D# => romdata <= X"00000704";
    when 16#0148E# => romdata <= X"04030007";
    when 16#0148F# => romdata <= X"05050007";
    when 16#01490# => romdata <= X"00020700";
    when 16#01491# => romdata <= X"00000000";
    when 16#01492# => romdata <= X"00000000";
    when 16#01493# => romdata <= X"00000000";
    when 16#01494# => romdata <= X"00000000";
    when 16#01495# => romdata <= X"0000FF00";
    when 16#01496# => romdata <= X"00000007";
    when 16#01497# => romdata <= X"01030500";
    when 16#01498# => romdata <= X"03040403";
    when 16#01499# => romdata <= X"00040502";
    when 16#0149A# => romdata <= X"00040502";
    when 16#0149B# => romdata <= X"00000705";
    when 16#0149C# => romdata <= X"05000700";
    when 16#0149D# => romdata <= X"02070000";
    when 16#0149E# => romdata <= X"07040403";
    when 16#0149F# => romdata <= X"00030404";
    when 16#014A0# => romdata <= X"03000701";
    when 16#014A1# => romdata <= X"03050007";
    when 16#014A2# => romdata <= X"01010000";
    when 16#014A3# => romdata <= X"00000000";
    when 16#014A4# => romdata <= X"00000000";
    when 16#014A5# => romdata <= X"00000000";
    when 16#014A6# => romdata <= X"00000000";
    when 16#014A7# => romdata <= X"00000000";
    when 16#014A8# => romdata <= X"71756974";
    when 16#014A9# => romdata <= X"00000000";
    when 16#014AA# => romdata <= X"68656C70";
    when 16#014AB# => romdata <= X"00000000";
    when 16#014AC# => romdata <= X"0A307800";
    when 16#014AD# => romdata <= X"69326320";
    when 16#014AE# => romdata <= X"464D430A";
    when 16#014AF# => romdata <= X"00000000";
    when 16#014B0# => romdata <= X"61646472";
    when 16#014B1# => romdata <= X"6573733A";
    when 16#014B2# => romdata <= X"20307800";
    when 16#014B3# => romdata <= X"2020202D";
    when 16#014B4# => romdata <= X"2D3E2020";
    when 16#014B5# => romdata <= X"2041434B";
    when 16#014B6# => romdata <= X"0A000000";
    when 16#014B7# => romdata <= X"72656164";
    when 16#014B8# => romdata <= X"20646174";
    when 16#014B9# => romdata <= X"61202800";
    when 16#014BA# => romdata <= X"20627974";
    when 16#014BB# => romdata <= X"65732920";
    when 16#014BC# => romdata <= X"66726F6D";
    when 16#014BD# => romdata <= X"20493243";
    when 16#014BE# => romdata <= X"2D616464";
    when 16#014BF# => romdata <= X"72657373";
    when 16#014C0# => romdata <= X"20307800";
    when 16#014C1# => romdata <= X"0A0A0000";
    when 16#014C2# => romdata <= X"6E6F6163";
    when 16#014C3# => romdata <= X"6B200000";
    when 16#014C4# => romdata <= X"6368726F";
    when 16#014C5# => romdata <= X"6E74656C";
    when 16#014C6# => romdata <= X"20726567";
    when 16#014C7# => romdata <= X"20307800";
    when 16#014C8# => romdata <= X"3A203078";
    when 16#014C9# => romdata <= X"00000000";
    when 16#014CA# => romdata <= X"206E6163";
    when 16#014CB# => romdata <= X"6B000000";
    when 16#014CC# => romdata <= X"6572726F";
    when 16#014CD# => romdata <= X"7220286E";
    when 16#014CE# => romdata <= X"61636B29";
    when 16#014CF# => romdata <= X"0A000000";
    when 16#014D0# => romdata <= X"0A202063";
    when 16#014D1# => romdata <= X"68616E6E";
    when 16#014D2# => romdata <= X"656C2033";
    when 16#014D3# => romdata <= X"20696E70";
    when 16#014D4# => romdata <= X"7574206F";
    when 16#014D5# => romdata <= X"76657266";
    when 16#014D6# => romdata <= X"6C6F7700";
    when 16#014D7# => romdata <= X"0A202063";
    when 16#014D8# => romdata <= X"68616E6E";
    when 16#014D9# => romdata <= X"656C2032";
    when 16#014DA# => romdata <= X"20696E70";
    when 16#014DB# => romdata <= X"7574206F";
    when 16#014DC# => romdata <= X"76657266";
    when 16#014DD# => romdata <= X"6C6F7700";
    when 16#014DE# => romdata <= X"0A202063";
    when 16#014DF# => romdata <= X"68616E6E";
    when 16#014E0# => romdata <= X"656C2031";
    when 16#014E1# => romdata <= X"20696E70";
    when 16#014E2# => romdata <= X"7574206F";
    when 16#014E3# => romdata <= X"76657266";
    when 16#014E4# => romdata <= X"6C6F7700";
    when 16#014E5# => romdata <= X"0A202063";
    when 16#014E6# => romdata <= X"68616E6E";
    when 16#014E7# => romdata <= X"656C2030";
    when 16#014E8# => romdata <= X"20696E70";
    when 16#014E9# => romdata <= X"7574206F";
    when 16#014EA# => romdata <= X"76657266";
    when 16#014EB# => romdata <= X"6C6F7700";
    when 16#014EC# => romdata <= X"0A202063";
    when 16#014ED# => romdata <= X"68616E6E";
    when 16#014EE# => romdata <= X"656C2033";
    when 16#014EF# => romdata <= X"20717561";
    when 16#014F0# => romdata <= X"6473756D";
    when 16#014F1# => romdata <= X"206F7665";
    when 16#014F2# => romdata <= X"72666C6F";
    when 16#014F3# => romdata <= X"77000000";
    when 16#014F4# => romdata <= X"0A202063";
    when 16#014F5# => romdata <= X"68616E6E";
    when 16#014F6# => romdata <= X"656C2032";
    when 16#014F7# => romdata <= X"20717561";
    when 16#014F8# => romdata <= X"6473756D";
    when 16#014F9# => romdata <= X"206F7665";
    when 16#014FA# => romdata <= X"72666C6F";
    when 16#014FB# => romdata <= X"77000000";
    when 16#014FC# => romdata <= X"0A202063";
    when 16#014FD# => romdata <= X"68616E6E";
    when 16#014FE# => romdata <= X"656C2031";
    when 16#014FF# => romdata <= X"20717561";
    when 16#01500# => romdata <= X"6473756D";
    when 16#01501# => romdata <= X"206F7665";
    when 16#01502# => romdata <= X"72666C6F";
    when 16#01503# => romdata <= X"77000000";
    when 16#01504# => romdata <= X"0A202063";
    when 16#01505# => romdata <= X"68616E6E";
    when 16#01506# => romdata <= X"656C2030";
    when 16#01507# => romdata <= X"20717561";
    when 16#01508# => romdata <= X"6473756D";
    when 16#01509# => romdata <= X"206F7665";
    when 16#0150A# => romdata <= X"72666C6F";
    when 16#0150B# => romdata <= X"77000000";
    when 16#0150C# => romdata <= X"0A202073";
    when 16#0150D# => romdata <= X"756D2076";
    when 16#0150E# => romdata <= X"616C7565";
    when 16#0150F# => romdata <= X"20637574";
    when 16#01510# => romdata <= X"74656400";
    when 16#01511# => romdata <= X"0A202063";
    when 16#01512# => romdata <= X"68616E6E";
    when 16#01513# => romdata <= X"656C2033";
    when 16#01514# => romdata <= X"20646976";
    when 16#01515# => romdata <= X"6964656E";
    when 16#01516# => romdata <= X"64206375";
    when 16#01517# => romdata <= X"74746564";
    when 16#01518# => romdata <= X"00000000";
    when 16#01519# => romdata <= X"0A202063";
    when 16#0151A# => romdata <= X"68616E6E";
    when 16#0151B# => romdata <= X"656C2033";
    when 16#0151C# => romdata <= X"206E6F69";
    when 16#0151D# => romdata <= X"73652063";
    when 16#0151E# => romdata <= X"6F6D7065";
    when 16#0151F# => romdata <= X"6E736174";
    when 16#01520# => romdata <= X"696F6E20";
    when 16#01521# => romdata <= X"746F2062";
    when 16#01522# => romdata <= X"69670000";
    when 16#01523# => romdata <= X"0A202063";
    when 16#01524# => romdata <= X"68616E6E";
    when 16#01525# => romdata <= X"656C2033";
    when 16#01526# => romdata <= X"206E6F69";
    when 16#01527# => romdata <= X"73652076";
    when 16#01528# => romdata <= X"616C7565";
    when 16#01529# => romdata <= X"20637574";
    when 16#0152A# => romdata <= X"74656400";
    when 16#0152B# => romdata <= X"0A202063";
    when 16#0152C# => romdata <= X"68616E6E";
    when 16#0152D# => romdata <= X"656C2032";
    when 16#0152E# => romdata <= X"20646976";
    when 16#0152F# => romdata <= X"6964656E";
    when 16#01530# => romdata <= X"64206375";
    when 16#01531# => romdata <= X"74746564";
    when 16#01532# => romdata <= X"00000000";
    when 16#01533# => romdata <= X"0A202063";
    when 16#01534# => romdata <= X"68616E6E";
    when 16#01535# => romdata <= X"656C2032";
    when 16#01536# => romdata <= X"206E6F69";
    when 16#01537# => romdata <= X"73652063";
    when 16#01538# => romdata <= X"6F6D7065";
    when 16#01539# => romdata <= X"6E736174";
    when 16#0153A# => romdata <= X"696F6E20";
    when 16#0153B# => romdata <= X"746F2062";
    when 16#0153C# => romdata <= X"69670000";
    when 16#0153D# => romdata <= X"0A202063";
    when 16#0153E# => romdata <= X"68616E6E";
    when 16#0153F# => romdata <= X"656C2032";
    when 16#01540# => romdata <= X"206E6F69";
    when 16#01541# => romdata <= X"73652076";
    when 16#01542# => romdata <= X"616C7565";
    when 16#01543# => romdata <= X"20637574";
    when 16#01544# => romdata <= X"74656400";
    when 16#01545# => romdata <= X"0A202063";
    when 16#01546# => romdata <= X"68616E6E";
    when 16#01547# => romdata <= X"656C2031";
    when 16#01548# => romdata <= X"20646976";
    when 16#01549# => romdata <= X"6964656E";
    when 16#0154A# => romdata <= X"64206375";
    when 16#0154B# => romdata <= X"74746564";
    when 16#0154C# => romdata <= X"00000000";
    when 16#0154D# => romdata <= X"0A202063";
    when 16#0154E# => romdata <= X"68616E6E";
    when 16#0154F# => romdata <= X"656C2031";
    when 16#01550# => romdata <= X"206E6F69";
    when 16#01551# => romdata <= X"73652063";
    when 16#01552# => romdata <= X"6F6D7065";
    when 16#01553# => romdata <= X"6E736174";
    when 16#01554# => romdata <= X"696F6E20";
    when 16#01555# => romdata <= X"746F2062";
    when 16#01556# => romdata <= X"69670000";
    when 16#01557# => romdata <= X"0A202063";
    when 16#01558# => romdata <= X"68616E6E";
    when 16#01559# => romdata <= X"656C2031";
    when 16#0155A# => romdata <= X"206E6F69";
    when 16#0155B# => romdata <= X"73652076";
    when 16#0155C# => romdata <= X"616C7565";
    when 16#0155D# => romdata <= X"20637574";
    when 16#0155E# => romdata <= X"74656400";
    when 16#0155F# => romdata <= X"0A202063";
    when 16#01560# => romdata <= X"68616E6E";
    when 16#01561# => romdata <= X"656C2030";
    when 16#01562# => romdata <= X"20646976";
    when 16#01563# => romdata <= X"6964656E";
    when 16#01564# => romdata <= X"64206375";
    when 16#01565# => romdata <= X"74746564";
    when 16#01566# => romdata <= X"00000000";
    when 16#01567# => romdata <= X"0A202063";
    when 16#01568# => romdata <= X"68616E6E";
    when 16#01569# => romdata <= X"656C2030";
    when 16#0156A# => romdata <= X"206E6F69";
    when 16#0156B# => romdata <= X"73652063";
    when 16#0156C# => romdata <= X"6F6D7065";
    when 16#0156D# => romdata <= X"6E736174";
    when 16#0156E# => romdata <= X"696F6E20";
    when 16#0156F# => romdata <= X"746F2062";
    when 16#01570# => romdata <= X"69670000";
    when 16#01571# => romdata <= X"0A202063";
    when 16#01572# => romdata <= X"68616E6E";
    when 16#01573# => romdata <= X"656C2030";
    when 16#01574# => romdata <= X"206E6F69";
    when 16#01575# => romdata <= X"73652076";
    when 16#01576# => romdata <= X"616C7565";
    when 16#01577# => romdata <= X"20637574";
    when 16#01578# => romdata <= X"74656400";
    when 16#01579# => romdata <= X"0A202073";
    when 16#0157A# => romdata <= X"6F667477";
    when 16#0157B# => romdata <= X"61726520";
    when 16#0157C# => romdata <= X"6572726F";
    when 16#0157D# => romdata <= X"72000000";
    when 16#0157E# => romdata <= X"0A657874";
    when 16#0157F# => romdata <= X"65726E61";
    when 16#01580# => romdata <= X"6C20636C";
    when 16#01581# => romdata <= X"6F636B20";
    when 16#01582# => romdata <= X"20202020";
    when 16#01583# => romdata <= X"2020203A";
    when 16#01584# => romdata <= X"20000000";
    when 16#01585# => romdata <= X"61637469";
    when 16#01586# => romdata <= X"76650000";
    when 16#01587# => romdata <= X"0A6D6963";
    when 16#01588# => romdata <= X"726F7075";
    when 16#01589# => romdata <= X"6C736520";
    when 16#0158A# => romdata <= X"736F7572";
    when 16#0158B# => romdata <= X"63652020";
    when 16#0158C# => romdata <= X"2020203A";
    when 16#0158D# => romdata <= X"20000000";
    when 16#0158E# => romdata <= X"65787465";
    when 16#0158F# => romdata <= X"726E616C";
    when 16#01590# => romdata <= X"00000000";
    when 16#01591# => romdata <= X"0A6D6963";
    when 16#01592# => romdata <= X"726F7075";
    when 16#01593# => romdata <= X"6C736520";
    when 16#01594# => romdata <= X"6576656E";
    when 16#01595# => romdata <= X"74206C69";
    when 16#01596# => romdata <= X"6D69743A";
    when 16#01597# => romdata <= X"20000000";
    when 16#01598# => romdata <= X"0A6D6561";
    when 16#01599# => romdata <= X"73757265";
    when 16#0159A# => romdata <= X"6D656E74";
    when 16#0159B# => romdata <= X"206C656E";
    when 16#0159C# => romdata <= X"67746820";
    when 16#0159D# => romdata <= X"2020203A";
    when 16#0159E# => romdata <= X"20000000";
    when 16#0159F# => romdata <= X"0A626561";
    when 16#015A0# => romdata <= X"6D20706F";
    when 16#015A1# => romdata <= X"73697469";
    when 16#015A2# => romdata <= X"6F6E206D";
    when 16#015A3# => romdata <= X"6F6E6974";
    when 16#015A4# => romdata <= X"6F722072";
    when 16#015A5# => romdata <= X"65676973";
    when 16#015A6# => romdata <= X"74657273";
    when 16#015A7# => romdata <= X"00000000";
    when 16#015A8# => romdata <= X"0A202020";
    when 16#015A9# => romdata <= X"20202020";
    when 16#015AA# => romdata <= X"20202020";
    when 16#015AB# => romdata <= X"20202020";
    when 16#015AC# => romdata <= X"20202020";
    when 16#015AD# => romdata <= X"20202020";
    when 16#015AE# => romdata <= X"20636861";
    when 16#015AF# => romdata <= X"6E6E656C";
    when 16#015B0# => romdata <= X"20302020";
    when 16#015B1# => romdata <= X"20636861";
    when 16#015B2# => romdata <= X"6E6E656C";
    when 16#015B3# => romdata <= X"20312020";
    when 16#015B4# => romdata <= X"20636861";
    when 16#015B5# => romdata <= X"6E6E656C";
    when 16#015B6# => romdata <= X"20322020";
    when 16#015B7# => romdata <= X"20636861";
    when 16#015B8# => romdata <= X"6E6E656C";
    when 16#015B9# => romdata <= X"20330000";
    when 16#015BA# => romdata <= X"0A202020";
    when 16#015BB# => romdata <= X"20202020";
    when 16#015BC# => romdata <= X"20202020";
    when 16#015BD# => romdata <= X"20202020";
    when 16#015BE# => romdata <= X"20202020";
    when 16#015BF# => romdata <= X"20202020";
    when 16#015C0# => romdata <= X"202D2D2D";
    when 16#015C1# => romdata <= X"2D20686F";
    when 16#015C2# => romdata <= X"72697A6F";
    when 16#015C3# => romdata <= X"6E74616C";
    when 16#015C4# => romdata <= X"202D2D2D";
    when 16#015C5# => romdata <= X"2D2D2020";
    when 16#015C6# => romdata <= X"202D2D2D";
    when 16#015C7# => romdata <= X"2D2D2D20";
    when 16#015C8# => romdata <= X"76657274";
    when 16#015C9# => romdata <= X"6963616C";
    when 16#015CA# => romdata <= X"202D2D2D";
    when 16#015CB# => romdata <= X"2D2D0000";
    when 16#015CC# => romdata <= X"0A736361";
    when 16#015CD# => romdata <= X"6C657220";
    when 16#015CE# => romdata <= X"76616C75";
    when 16#015CF# => romdata <= X"65732020";
    when 16#015D0# => romdata <= X"20202020";
    when 16#015D1# => romdata <= X"20202020";
    when 16#015D2# => romdata <= X"20000000";
    when 16#015D3# => romdata <= X"0A6E6F69";
    when 16#015D4# => romdata <= X"73652063";
    when 16#015D5# => romdata <= X"6F6D7065";
    when 16#015D6# => romdata <= X"6E736174";
    when 16#015D7# => romdata <= X"696F6E20";
    when 16#015D8# => romdata <= X"20202020";
    when 16#015D9# => romdata <= X"20000000";
    when 16#015DA# => romdata <= X"0A6D6561";
    when 16#015DB# => romdata <= X"73757265";
    when 16#015DC# => romdata <= X"6D656E74";
    when 16#015DD# => romdata <= X"20202020";
    when 16#015DE# => romdata <= X"20202020";
    when 16#015DF# => romdata <= X"20202020";
    when 16#015E0# => romdata <= X"20000000";
    when 16#015E1# => romdata <= X"0A73616D";
    when 16#015E2# => romdata <= X"706C6573";
    when 16#015E3# => romdata <= X"20286469";
    when 16#015E4# => romdata <= X"7629203A";
    when 16#015E5# => romdata <= X"20000000";
    when 16#015E6# => romdata <= X"0A73756D";
    when 16#015E7# => romdata <= X"20636861";
    when 16#015E8# => romdata <= X"6E6E656C";
    when 16#015E9# => romdata <= X"2020203A";
    when 16#015EA# => romdata <= X"20000000";
    when 16#015EB# => romdata <= X"0A0A706F";
    when 16#015EC# => romdata <= X"73697469";
    when 16#015ED# => romdata <= X"6F6E2063";
    when 16#015EE# => romdata <= X"6F6D7075";
    when 16#015EF# => romdata <= X"74617469";
    when 16#015F0# => romdata <= X"6F6E0000";
    when 16#015F1# => romdata <= X"0A202073";
    when 16#015F2# => romdata <= X"63616C65";
    when 16#015F3# => romdata <= X"72207661";
    when 16#015F4# => romdata <= X"6C756573";
    when 16#015F5# => romdata <= X"20202020";
    when 16#015F6# => romdata <= X"20202020";
    when 16#015F7# => romdata <= X"20000000";
    when 16#015F8# => romdata <= X"0A20206F";
    when 16#015F9# => romdata <= X"66667365";
    when 16#015FA# => romdata <= X"74202020";
    when 16#015FB# => romdata <= X"20202020";
    when 16#015FC# => romdata <= X"20202020";
    when 16#015FD# => romdata <= X"20202020";
    when 16#015FE# => romdata <= X"20000000";
    when 16#015FF# => romdata <= X"0A6F7574";
    when 16#01600# => romdata <= X"70757420";
    when 16#01601# => romdata <= X"73656C65";
    when 16#01602# => romdata <= X"6374203A";
    when 16#01603# => romdata <= X"20000000";
    when 16#01604# => romdata <= X"74657374";
    when 16#01605# => romdata <= X"67656E00";
    when 16#01606# => romdata <= X"4E4F5420";
    when 16#01607# => romdata <= X"00000000";
    when 16#01608# => romdata <= X"6368616E";
    when 16#01609# => romdata <= X"6E656C20";
    when 16#0160A# => romdata <= X"30000000";
    when 16#0160B# => romdata <= X"0A63616C";
    when 16#0160C# => romdata <= X"63207374";
    when 16#0160D# => romdata <= X"61746520";
    when 16#0160E# => romdata <= X"2020203A";
    when 16#0160F# => romdata <= X"20307800";
    when 16#01610# => romdata <= X"76657274";
    when 16#01611# => romdata <= X"6963616C";
    when 16#01612# => romdata <= X"00000000";
    when 16#01613# => romdata <= X"686F7269";
    when 16#01614# => romdata <= X"7A6F6E74";
    when 16#01615# => romdata <= X"616C0000";
    when 16#01616# => romdata <= X"73756D00";
    when 16#01617# => romdata <= X"6368616E";
    when 16#01618# => romdata <= X"6E656C20";
    when 16#01619# => romdata <= X"33000000";
    when 16#0161A# => romdata <= X"6368616E";
    when 16#0161B# => romdata <= X"6E656C20";
    when 16#0161C# => romdata <= X"32000000";
    when 16#0161D# => romdata <= X"6368616E";
    when 16#0161E# => romdata <= X"6E656C20";
    when 16#0161F# => romdata <= X"31000000";
    when 16#01620# => romdata <= X"786D6F64";
    when 16#01621# => romdata <= X"656D2074";
    when 16#01622# => romdata <= X"72616E73";
    when 16#01623# => romdata <= X"6D69742E";
    when 16#01624# => romdata <= X"2E2E0A00";
    when 16#01625# => romdata <= X"20627974";
    when 16#01626# => romdata <= X"65732074";
    when 16#01627# => romdata <= X"72616E73";
    when 16#01628# => romdata <= X"6D697474";
    when 16#01629# => romdata <= X"65640A00";
    when 16#0162A# => romdata <= X"63616E63";
    when 16#0162B# => romdata <= X"656C0A00";
    when 16#0162C# => romdata <= X"72657472";
    when 16#0162D# => romdata <= X"79206F75";
    when 16#0162E# => romdata <= X"740A0000";
    when 16#0162F# => romdata <= X"786D6F64";
    when 16#01630# => romdata <= X"656D2072";
    when 16#01631# => romdata <= X"65636569";
    when 16#01632# => romdata <= X"76652E2E";
    when 16#01633# => romdata <= X"2E0A0000";
    when 16#01634# => romdata <= X"20627974";
    when 16#01635# => romdata <= X"65732072";
    when 16#01636# => romdata <= X"65636569";
    when 16#01637# => romdata <= X"7665640A";
    when 16#01638# => romdata <= X"00000000";
    when 16#01639# => romdata <= X"72782062";
    when 16#0163A# => romdata <= X"75666665";
    when 16#0163B# => romdata <= X"72206675";
    when 16#0163C# => romdata <= X"6C6C0A00";
    when 16#0163D# => romdata <= X"74696D65";
    when 16#0163E# => romdata <= X"206F7574";
    when 16#0163F# => romdata <= X"0A000000";
    when 16#01640# => romdata <= X"64656275";
    when 16#01641# => romdata <= X"67207265";
    when 16#01642# => romdata <= X"67697374";
    when 16#01643# => romdata <= X"65727300";
    when 16#01644# => romdata <= X"0A6D6F64";
    when 16#01645# => romdata <= X"65202020";
    when 16#01646# => romdata <= X"20202020";
    when 16#01647# => romdata <= X"203A2000";
    when 16#01648# => romdata <= X"0A616464";
    when 16#01649# => romdata <= X"72657373";
    when 16#0164A# => romdata <= X"20302020";
    when 16#0164B# => romdata <= X"203A2030";
    when 16#0164C# => romdata <= X"78000000";
    when 16#0164D# => romdata <= X"0A616464";
    when 16#0164E# => romdata <= X"72657373";
    when 16#0164F# => romdata <= X"20312020";
    when 16#01650# => romdata <= X"203A2030";
    when 16#01651# => romdata <= X"78000000";
    when 16#01652# => romdata <= X"0A627566";
    when 16#01653# => romdata <= X"66657220";
    when 16#01654# => romdata <= X"73697A65";
    when 16#01655# => romdata <= X"203A2000";
    when 16#01656# => romdata <= X"6D61783A";
    when 16#01657# => romdata <= X"20000000";
    when 16#01658# => romdata <= X"6D696E3A";
    when 16#01659# => romdata <= X"20000000";
    when 16#0165A# => romdata <= X"63683A20";
    when 16#0165B# => romdata <= X"00000000";
    when 16#0165C# => romdata <= X"73706C3A";
    when 16#0165D# => romdata <= X"20000000";
    when 16#0165E# => romdata <= X"73686F77";
    when 16#0165F# => romdata <= X"2042504D";
    when 16#01660# => romdata <= X"20726567";
    when 16#01661# => romdata <= X"69737465";
    when 16#01662# => romdata <= X"72730000";
    when 16#01663# => romdata <= X"62706D00";
    when 16#01664# => romdata <= X"73656C65";
    when 16#01665# => romdata <= X"6374206F";
    when 16#01666# => romdata <= X"75747075";
    when 16#01667# => romdata <= X"74206368";
    when 16#01668# => romdata <= X"616E6E65";
    when 16#01669# => romdata <= X"6C202830";
    when 16#0166A# => romdata <= X"2E2E3320";
    when 16#0166B# => romdata <= X"73756D20";
    when 16#0166C# => romdata <= X"68207629";
    when 16#0166D# => romdata <= X"00000000";
    when 16#0166E# => romdata <= X"73656C65";
    when 16#0166F# => romdata <= X"63740000";
    when 16#01670# => romdata <= X"73797374";
    when 16#01671# => romdata <= X"656D2072";
    when 16#01672# => romdata <= X"65736574";
    when 16#01673# => romdata <= X"00000000";
    when 16#01674# => romdata <= X"72657365";
    when 16#01675# => romdata <= X"74000000";
    when 16#01676# => romdata <= X"73686F77";
    when 16#01677# => romdata <= X"20737973";
    when 16#01678# => romdata <= X"74656D20";
    when 16#01679# => romdata <= X"696E666F";
    when 16#0167A# => romdata <= X"203C7665";
    when 16#0167B# => romdata <= X"72626F73";
    when 16#0167C# => romdata <= X"653E0000";
    when 16#0167D# => romdata <= X"73797369";
    when 16#0167E# => romdata <= X"6E666F00";
    when 16#0167F# => romdata <= X"73686F77";
    when 16#01680# => romdata <= X"2F736574";
    when 16#01681# => romdata <= X"20646562";
    when 16#01682# => romdata <= X"75672072";
    when 16#01683# => romdata <= X"65676973";
    when 16#01684# => romdata <= X"74657273";
    when 16#01685# => romdata <= X"203C7365";
    when 16#01686# => romdata <= X"74206D6F";
    when 16#01687# => romdata <= X"64653E00";
    when 16#01688# => romdata <= X"64656275";
    when 16#01689# => romdata <= X"67000000";
    when 16#0168A# => romdata <= X"636C6B20";
    when 16#0168B# => romdata <= X"736F7572";
    when 16#0168C# => romdata <= X"63653A20";
    when 16#0168D# => romdata <= X"2030203D";
    when 16#0168E# => romdata <= X"20696E74";
    when 16#0168F# => romdata <= X"2C203120";
    when 16#01690# => romdata <= X"3D206578";
    when 16#01691# => romdata <= X"74000000";
    when 16#01692# => romdata <= X"636C6B00";
    when 16#01693# => romdata <= X"6D696372";
    when 16#01694# => romdata <= X"6F70756C";
    when 16#01695# => romdata <= X"73652073";
    when 16#01696# => romdata <= X"6F757263";
    when 16#01697# => romdata <= X"653A2030";
    when 16#01698# => romdata <= X"203D2069";
    when 16#01699# => romdata <= X"6E742C20";
    when 16#0169A# => romdata <= X"31203D20";
    when 16#0169B# => romdata <= X"65787400";
    when 16#0169C# => romdata <= X"6D696372";
    when 16#0169D# => romdata <= X"6F000000";
    when 16#0169E# => romdata <= X"74657374";
    when 16#0169F# => romdata <= X"67656E65";
    when 16#016A0# => romdata <= X"7261746F";
    when 16#016A1# => romdata <= X"72203C73";
    when 16#016A2# => romdata <= X"63616C65";
    when 16#016A3# => romdata <= X"723E203C";
    when 16#016A4# => romdata <= X"72657374";
    when 16#016A5# => romdata <= X"6172743E";
    when 16#016A6# => romdata <= X"00000000";
    when 16#016A7# => romdata <= X"3C6D7574";
    when 16#016A8# => romdata <= X"655F6E3E";
    when 16#016A9# => romdata <= X"203C7273";
    when 16#016AA# => romdata <= X"745F6E3E";
    when 16#016AB# => romdata <= X"203C6270";
    when 16#016AC# => romdata <= X"625F6E3E";
    when 16#016AD# => romdata <= X"203C6F73";
    when 16#016AE# => romdata <= X"72313E20";
    when 16#016AF# => romdata <= X"3C6F7372";
    when 16#016B0# => romdata <= X"323E0000";
    when 16#016B1# => romdata <= X"64616363";
    when 16#016B2# => romdata <= X"6F6E6600";
    when 16#016B3# => romdata <= X"3C6D756C";
    when 16#016B4# => romdata <= X"7469706C";
    when 16#016B5# => romdata <= X"6965723E";
    when 16#016B6# => romdata <= X"20696E69";
    when 16#016B7# => romdata <= X"7469616C";
    when 16#016B8# => romdata <= X"697A6520";
    when 16#016B9# => romdata <= X"62756666";
    when 16#016BA# => romdata <= X"65720000";
    when 16#016BB# => romdata <= X"64616374";
    when 16#016BC# => romdata <= X"65737400";
    when 16#016BD# => romdata <= X"72657365";
    when 16#016BE# => romdata <= X"74206361";
    when 16#016BF# => romdata <= X"6C63756C";
    when 16#016C0# => romdata <= X"6174696F";
    when 16#016C1# => romdata <= X"6E206572";
    when 16#016C2# => romdata <= X"726F7273";
    when 16#016C3# => romdata <= X"00000000";
    when 16#016C4# => romdata <= X"63616C63";
    when 16#016C5# => romdata <= X"72657300";
    when 16#016C6# => romdata <= X"73686F77";
    when 16#016C7# => romdata <= X"20646562";
    when 16#016C8# => romdata <= X"75672062";
    when 16#016C9# => romdata <= X"75666665";
    when 16#016CA# => romdata <= X"72203C6C";
    when 16#016CB# => romdata <= X"656E6774";
    when 16#016CC# => romdata <= X"683E0000";
    when 16#016CD# => romdata <= X"636C6561";
    when 16#016CE# => romdata <= X"72206465";
    when 16#016CF# => romdata <= X"62756720";
    when 16#016D0# => romdata <= X"62756666";
    when 16#016D1# => romdata <= X"65720000";
    when 16#016D2# => romdata <= X"62636C65";
    when 16#016D3# => romdata <= X"61720000";
    when 16#016D4# => romdata <= X"62756666";
    when 16#016D5# => romdata <= X"6572206F";
    when 16#016D6# => romdata <= X"6E204C43";
    when 16#016D7# => romdata <= X"44203C63";
    when 16#016D8# => romdata <= X"683E203C";
    when 16#016D9# => romdata <= X"636F6D62";
    when 16#016DA# => romdata <= X"3E000000";
    when 16#016DB# => romdata <= X"73636F70";
    when 16#016DC# => romdata <= X"65000000";
    when 16#016DD# => romdata <= X"64656275";
    when 16#016DE# => romdata <= X"67207472";
    when 16#016DF# => romdata <= X"61636520";
    when 16#016E0# => romdata <= X"3C636C65";
    when 16#016E1# => romdata <= X"61723E00";
    when 16#016E2# => romdata <= X"74726163";
    when 16#016E3# => romdata <= X"65000000";
    when 16#016E4# => romdata <= X"73657475";
    when 16#016E5# => romdata <= X"70206368";
    when 16#016E6# => romdata <= X"616E6E65";
    when 16#016E7# => romdata <= X"6C207465";
    when 16#016E8# => romdata <= X"7374203C";
    when 16#016E9# => romdata <= X"63683E20";
    when 16#016EA# => romdata <= X"3C76616C";
    when 16#016EB# => romdata <= X"302E2E37";
    when 16#016EC# => romdata <= X"3E000000";
    when 16#016ED# => romdata <= X"63687465";
    when 16#016EE# => romdata <= X"73740000";
    when 16#016EF# => romdata <= X"72756E6E";
    when 16#016F0# => romdata <= X"696E6720";
    when 16#016F1# => romdata <= X"6C696768";
    when 16#016F2# => romdata <= X"74000000";
    when 16#016F3# => romdata <= X"72756E00";
    when 16#016F4# => romdata <= X"72756E20";
    when 16#016F5# => romdata <= X"64697370";
    when 16#016F6# => romdata <= X"6C617920";
    when 16#016F7# => romdata <= X"74657374";
    when 16#016F8# => romdata <= X"2066756E";
    when 16#016F9# => romdata <= X"6374696F";
    when 16#016FA# => romdata <= X"6E000000";
    when 16#016FB# => romdata <= X"64697370";
    when 16#016FC# => romdata <= X"6C617900";
    when 16#016FD# => romdata <= X"73657420";
    when 16#016FE# => romdata <= X"6261636B";
    when 16#016FF# => romdata <= X"6C696768";
    when 16#01700# => romdata <= X"74203C30";
    when 16#01701# => romdata <= X"2E2E3331";
    when 16#01702# => romdata <= X"3E000000";
    when 16#01703# => romdata <= X"6261636B";
    when 16#01704# => romdata <= X"00000000";
    when 16#01705# => romdata <= X"73686F77";
    when 16#01706# => romdata <= X"206C6F67";
    when 16#01707# => romdata <= X"6F206F6E";
    when 16#01708# => romdata <= X"20676C63";
    when 16#01709# => romdata <= X"64000000";
    when 16#0170A# => romdata <= X"6C6F676F";
    when 16#0170B# => romdata <= X"00000000";
    when 16#0170C# => romdata <= X"63686563";
    when 16#0170D# => romdata <= X"6B204932";
    when 16#0170E# => romdata <= X"43206164";
    when 16#0170F# => romdata <= X"64726573";
    when 16#01710# => romdata <= X"73000000";
    when 16#01711# => romdata <= X"69326300";
    when 16#01712# => romdata <= X"72656164";
    when 16#01713# => romdata <= X"20454550";
    when 16#01714# => romdata <= X"524F4D20";
    when 16#01715# => romdata <= X"3C627573";
    when 16#01716# => romdata <= X"3E203C69";
    when 16#01717# => romdata <= X"32635F61";
    when 16#01718# => romdata <= X"6464723E";
    when 16#01719# => romdata <= X"203C6C65";
    when 16#0171A# => romdata <= X"6E677468";
    when 16#0171B# => romdata <= X"3E000000";
    when 16#0171C# => romdata <= X"65657072";
    when 16#0171D# => romdata <= X"6F6D0000";
    when 16#0171E# => romdata <= X"41444320";
    when 16#0171F# => romdata <= X"72656769";
    when 16#01720# => romdata <= X"73746572";
    when 16#01721# => romdata <= X"20747261";
    when 16#01722# => romdata <= X"6E736665";
    when 16#01723# => romdata <= X"72203C76";
    when 16#01724# => romdata <= X"616C7565";
    when 16#01725# => romdata <= X"3E000000";
    when 16#01726# => romdata <= X"61747261";
    when 16#01727# => romdata <= X"6E730000";
    when 16#01728# => romdata <= X"696E6974";
    when 16#01729# => romdata <= X"20414443";
    when 16#0172A# => romdata <= X"20726567";
    when 16#0172B# => romdata <= X"69737465";
    when 16#0172C# => romdata <= X"72730000";
    when 16#0172D# => romdata <= X"61696E69";
    when 16#0172E# => romdata <= X"74000000";
    when 16#0172F# => romdata <= X"616C6961";
    when 16#01730# => romdata <= X"7320666F";
    when 16#01731# => romdata <= X"72207800";
    when 16#01732# => romdata <= X"6D656D00";
    when 16#01733# => romdata <= X"77726974";
    when 16#01734# => romdata <= X"6520776F";
    when 16#01735# => romdata <= X"7264203C";
    when 16#01736# => romdata <= X"61646472";
    when 16#01737# => romdata <= X"3E203C6C";
    when 16#01738# => romdata <= X"656E6774";
    when 16#01739# => romdata <= X"683E203C";
    when 16#0173A# => romdata <= X"76616C75";
    when 16#0173B# => romdata <= X"65287329";
    when 16#0173C# => romdata <= X"3E000000";
    when 16#0173D# => romdata <= X"776D656D";
    when 16#0173E# => romdata <= X"00000000";
    when 16#0173F# => romdata <= X"6558616D";
    when 16#01740# => romdata <= X"696E6520";
    when 16#01741# => romdata <= X"6D656D6F";
    when 16#01742# => romdata <= X"7279203C";
    when 16#01743# => romdata <= X"61646472";
    when 16#01744# => romdata <= X"3E203C6C";
    when 16#01745# => romdata <= X"656E6774";
    when 16#01746# => romdata <= X"683E0000";
    when 16#01747# => romdata <= X"636C6561";
    when 16#01748# => romdata <= X"72207363";
    when 16#01749# => romdata <= X"7265656E";
    when 16#0174A# => romdata <= X"00000000";
    when 16#0174B# => romdata <= X"636C6561";
    when 16#0174C# => romdata <= X"72000000";
    when 16#0174D# => romdata <= X"0A646562";
    when 16#0174E# => romdata <= X"75672074";
    when 16#0174F# => romdata <= X"72616365";
    when 16#01750# => romdata <= X"206D656D";
    when 16#01751# => romdata <= X"6F727900";
    when 16#01752# => romdata <= X"0A74696D";
    when 16#01753# => romdata <= X"65207374";
    when 16#01754# => romdata <= X"616D7020";
    when 16#01755# => romdata <= X"20202073";
    when 16#01756# => romdata <= X"74617465";
    when 16#01757# => romdata <= X"00000000";
    when 16#01758# => romdata <= X"20203078";
    when 16#01759# => romdata <= X"00000000";
    when 16#0175A# => romdata <= X"65787465";
    when 16#0175B# => romdata <= X"726E616C";
    when 16#0175C# => romdata <= X"20636C6F";
    when 16#0175D# => romdata <= X"636B2000";
    when 16#0175E# => romdata <= X"61637469";
    when 16#0175F# => romdata <= X"76650A00";
    when 16#01760# => romdata <= X"73656C65";
    when 16#01761# => romdata <= X"63746564";
    when 16#01762# => romdata <= X"0A000000";
    when 16#01763# => romdata <= X"6D696372";
    when 16#01764# => romdata <= X"6F70756C";
    when 16#01765# => romdata <= X"73652073";
    when 16#01766# => romdata <= X"6F757263";
    when 16#01767# => romdata <= X"653A2000";
    when 16#01768# => romdata <= X"6265616D";
    when 16#01769# => romdata <= X"20706F73";
    when 16#0176A# => romdata <= X"6974696F";
    when 16#0176B# => romdata <= X"6E206D6F";
    when 16#0176C# => romdata <= X"6E69746F";
    when 16#0176D# => romdata <= X"72000000";
    when 16#0176E# => romdata <= X"20286F6E";
    when 16#0176F# => romdata <= X"2073696D";
    when 16#01770# => romdata <= X"290A0000";
    when 16#01771# => romdata <= X"0A485720";
    when 16#01772# => romdata <= X"73796E74";
    when 16#01773# => romdata <= X"68657369";
    when 16#01774# => romdata <= X"7A65643A";
    when 16#01775# => romdata <= X"20000000";
    when 16#01776# => romdata <= X"0A535720";
    when 16#01777# => romdata <= X"636F6D70";
    when 16#01778# => romdata <= X"696C6564";
    when 16#01779# => romdata <= X"2020203A";
    when 16#0177A# => romdata <= X"20417567";
    when 16#0177B# => romdata <= X"20313820";
    when 16#0177C# => romdata <= X"32303131";
    when 16#0177D# => romdata <= X"20203131";
    when 16#0177E# => romdata <= X"3A32323A";
    when 16#0177F# => romdata <= X"35300000";
    when 16#01780# => romdata <= X"0A737973";
    when 16#01781# => romdata <= X"74656D20";
    when 16#01782# => romdata <= X"636C6F63";
    when 16#01783# => romdata <= X"6B20203A";
    when 16#01784# => romdata <= X"20000000";
    when 16#01785# => romdata <= X"204D487A";
    when 16#01786# => romdata <= X"0A000000";
    when 16#01787# => romdata <= X"44454255";
    when 16#01788# => romdata <= X"47204D4F";
    when 16#01789# => romdata <= X"44450000";
    when 16#0178A# => romdata <= X"204F4E0A";
    when 16#0178B# => romdata <= X"00000000";
    when 16#0178C# => romdata <= X"0000117B";
    when 16#0178D# => romdata <= X"000011E4";
    when 16#0178E# => romdata <= X"000011D9";
    when 16#0178F# => romdata <= X"000011CE";
    when 16#01790# => romdata <= X"000011C3";
    when 16#01791# => romdata <= X"000011B9";
    when 16#01792# => romdata <= X"000011AF";
    when 16#01793# => romdata <= X"000002C2";
    when 16#01794# => romdata <= X"FC1902C4";
    when 16#01795# => romdata <= X"FFFEFD3F";
    when 16#01796# => romdata <= X"03E7FD3B";
    when 16#01797# => romdata <= X"0000485D";
    when 16#01798# => romdata <= X"999B4888";
    when 16#01799# => romdata <= X"FFC4B7CE";
    when 16#0179A# => romdata <= X"6665B74E";
    when 16#0179B# => romdata <= X"3E200000";
    when 16#0179C# => romdata <= X"636F6D6D";
    when 16#0179D# => romdata <= X"616E6420";
    when 16#0179E# => romdata <= X"6E6F7420";
    when 16#0179F# => romdata <= X"666F756E";
    when 16#017A0# => romdata <= X"642E0A00";
    when 16#017A1# => romdata <= X"73757070";
    when 16#017A2# => romdata <= X"6F727465";
    when 16#017A3# => romdata <= X"6420636F";
    when 16#017A4# => romdata <= X"6D6D616E";
    when 16#017A5# => romdata <= X"64733A0A";
    when 16#017A6# => romdata <= X"0A000000";
    when 16#017A7# => romdata <= X"202D2000";
    when 16#017A8# => romdata <= X"76656E64";
    when 16#017A9# => romdata <= X"6F723F20";
    when 16#017AA# => romdata <= X"20000000";
    when 16#017AB# => romdata <= X"67616973";
    when 16#017AC# => romdata <= X"6C657220";
    when 16#017AD# => romdata <= X"20000000";
    when 16#017AE# => romdata <= X"756E6B6E";
    when 16#017AF# => romdata <= X"6F776E20";
    when 16#017B0# => romdata <= X"64657669";
    when 16#017B1# => romdata <= X"63650000";
    when 16#017B2# => romdata <= X"485A4452";
    when 16#017B3# => romdata <= X"20202020";
    when 16#017B4# => romdata <= X"20000000";
    when 16#017B5# => romdata <= X"56474120";
    when 16#017B6# => romdata <= X"636F6E74";
    when 16#017B7# => romdata <= X"726F6C6C";
    when 16#017B8# => romdata <= X"65720000";
    when 16#017B9# => romdata <= X"47656E65";
    when 16#017BA# => romdata <= X"72616C20";
    when 16#017BB# => romdata <= X"50757270";
    when 16#017BC# => romdata <= X"6F736520";
    when 16#017BD# => romdata <= X"492F4F20";
    when 16#017BE# => romdata <= X"706F7274";
    when 16#017BF# => romdata <= X"00000000";
    when 16#017C0# => romdata <= X"4475616C";
    when 16#017C1# => romdata <= X"2D706F72";
    when 16#017C2# => romdata <= X"74204148";
    when 16#017C3# => romdata <= X"42205352";
    when 16#017C4# => romdata <= X"414D206D";
    when 16#017C5# => romdata <= X"6F64756C";
    when 16#017C6# => romdata <= X"65000000";
    when 16#017C7# => romdata <= X"64656275";
    when 16#017C8# => romdata <= X"67206275";
    when 16#017C9# => romdata <= X"66666572";
    when 16#017CA# => romdata <= X"20636F6E";
    when 16#017CB# => romdata <= X"74726F6C";
    when 16#017CC# => romdata <= X"00000000";
    when 16#017CD# => romdata <= X"74726967";
    when 16#017CE# => romdata <= X"67657220";
    when 16#017CF# => romdata <= X"67656E65";
    when 16#017D0# => romdata <= X"7261746F";
    when 16#017D1# => romdata <= X"72000000";
    when 16#017D2# => romdata <= X"64656275";
    when 16#017D3# => romdata <= X"6720636F";
    when 16#017D4# => romdata <= X"6E736F6C";
    when 16#017D5# => romdata <= X"65000000";
    when 16#017D6# => romdata <= X"64656275";
    when 16#017D7# => romdata <= X"67207472";
    when 16#017D8# => romdata <= X"61636572";
    when 16#017D9# => romdata <= X"206D656D";
    when 16#017DA# => romdata <= X"6F727900";
    when 16#017DB# => romdata <= X"4541444F";
    when 16#017DC# => romdata <= X"47533130";
    when 16#017DD# => romdata <= X"32206469";
    when 16#017DE# => romdata <= X"73706C61";
    when 16#017DF# => romdata <= X"79206472";
    when 16#017E0# => romdata <= X"69766572";
    when 16#017E1# => romdata <= X"00000000";
    when 16#017E2# => romdata <= X"44434D20";
    when 16#017E3# => romdata <= X"70686173";
    when 16#017E4# => romdata <= X"65207368";
    when 16#017E5# => romdata <= X"69667420";
    when 16#017E6# => romdata <= X"636F6E74";
    when 16#017E7# => romdata <= X"726F6C00";
    when 16#017E8# => romdata <= X"5A505520";
    when 16#017E9# => romdata <= X"4D656D6F";
    when 16#017EA# => romdata <= X"72792077";
    when 16#017EB# => romdata <= X"72617070";
    when 16#017EC# => romdata <= X"65720000";
    when 16#017ED# => romdata <= X"5A505520";
    when 16#017EE# => romdata <= X"41484220";
    when 16#017EF# => romdata <= X"57726170";
    when 16#017F0# => romdata <= X"70657200";
    when 16#017F1# => romdata <= X"4148422F";
    when 16#017F2# => romdata <= X"41504220";
    when 16#017F3# => romdata <= X"42726964";
    when 16#017F4# => romdata <= X"67650000";
    when 16#017F5# => romdata <= X"4D6F6475";
    when 16#017F6# => romdata <= X"6C617220";
    when 16#017F7# => romdata <= X"54696D65";
    when 16#017F8# => romdata <= X"7220556E";
    when 16#017F9# => romdata <= X"69740000";
    when 16#017FA# => romdata <= X"47656E65";
    when 16#017FB# => romdata <= X"72696320";
    when 16#017FC# => romdata <= X"55415254";
    when 16#017FD# => romdata <= X"00000000";
    when 16#017FE# => romdata <= X"414D4241";
    when 16#017FF# => romdata <= X"20577261";
    when 16#01800# => romdata <= X"70706572";
    when 16#01801# => romdata <= X"20666F72";
    when 16#01802# => romdata <= X"204F4320";
    when 16#01803# => romdata <= X"4932432D";
    when 16#01804# => romdata <= X"6D617374";
    when 16#01805# => romdata <= X"65720000";
    when 16#01806# => romdata <= X"53504920";
    when 16#01807# => romdata <= X"4D656D6F";
    when 16#01808# => romdata <= X"72792043";
    when 16#01809# => romdata <= X"6F6E7472";
    when 16#0180A# => romdata <= X"6F6C6C65";
    when 16#0180B# => romdata <= X"72000000";
    when 16#0180C# => romdata <= X"20206170";
    when 16#0180D# => romdata <= X"62736C76";
    when 16#0180E# => romdata <= X"00000000";
    when 16#0180F# => romdata <= X"76656E64";
    when 16#01810# => romdata <= X"20307800";
    when 16#01811# => romdata <= X"64657620";
    when 16#01812# => romdata <= X"30780000";
    when 16#01813# => romdata <= X"76657220";
    when 16#01814# => romdata <= X"00000000";
    when 16#01815# => romdata <= X"69727120";
    when 16#01816# => romdata <= X"00000000";
    when 16#01817# => romdata <= X"61646472";
    when 16#01818# => romdata <= X"20307800";
    when 16#01819# => romdata <= X"6168626D";
    when 16#0181A# => romdata <= X"73740000";
    when 16#0181B# => romdata <= X"61686273";
    when 16#0181C# => romdata <= X"6C760000";
    when 16#0181D# => romdata <= X"00002B01";
    when 16#0181E# => romdata <= X"00002BC9";
    when 16#0181F# => romdata <= X"00002BBE";
    when 16#01820# => romdata <= X"00002BB3";
    when 16#01821# => romdata <= X"00002B92";
    when 16#01822# => romdata <= X"00002B87";
    when 16#01823# => romdata <= X"00002B7C";
    when 16#01824# => romdata <= X"00002B71";
    when 16#01825# => romdata <= X"00002BA8";
    when 16#01826# => romdata <= X"00002B9D";
    when 16#01827# => romdata <= X"04580808";
    when 16#01828# => romdata <= X"20FF0000";
    when 16#01829# => romdata <= X"000060AC";
    when 16#0182A# => romdata <= X"0000618C";
    when 16#0182B# => romdata <= X"02010305";
    when 16#0182C# => romdata <= X"05070501";
    when 16#0182D# => romdata <= X"03030505";
    when 16#0182E# => romdata <= X"02030104";
    when 16#0182F# => romdata <= X"05050505";
    when 16#01830# => romdata <= X"05050505";
    when 16#01831# => romdata <= X"05050101";
    when 16#01832# => romdata <= X"04050404";
    when 16#01833# => romdata <= X"07050505";
    when 16#01834# => romdata <= X"05050505";
    when 16#01835# => romdata <= X"05030405";
    when 16#01836# => romdata <= X"05050505";
    when 16#01837# => romdata <= X"05050505";
    when 16#01838# => romdata <= X"05050505";
    when 16#01839# => romdata <= X"05050503";
    when 16#0183A# => romdata <= X"04030505";
    when 16#0183B# => romdata <= X"02050504";
    when 16#0183C# => romdata <= X"05050405";
    when 16#0183D# => romdata <= X"04010204";
    when 16#0183E# => romdata <= X"02050404";
    when 16#0183F# => romdata <= X"05050404";
    when 16#01840# => romdata <= X"04040507";
    when 16#01841# => romdata <= X"05040404";
    when 16#01842# => romdata <= X"02040500";
    when 16#01843# => romdata <= X"04050200";
    when 16#01844# => romdata <= X"04080303";
    when 16#01845# => romdata <= X"04090003";
    when 16#01846# => romdata <= X"06000000";
    when 16#01847# => romdata <= X"00020204";
    when 16#01848# => romdata <= X"04040400";
    when 16#01849# => romdata <= X"04060003";
    when 16#0184A# => romdata <= X"05000000";
    when 16#0184B# => romdata <= X"00000404";
    when 16#0184C# => romdata <= X"05050204";
    when 16#0184D# => romdata <= X"05060305";
    when 16#0184E# => romdata <= X"04030705";
    when 16#0184F# => romdata <= X"04050303";
    when 16#01850# => romdata <= X"02040502";
    when 16#01851# => romdata <= X"03020405";
    when 16#01852# => romdata <= X"06060604";
    when 16#01853# => romdata <= X"05050505";
    when 16#01854# => romdata <= X"05050504";
    when 16#01855# => romdata <= X"04040404";
    when 16#01856# => romdata <= X"03030303";
    when 16#01857# => romdata <= X"05050505";
    when 16#01858# => romdata <= X"05050505";
    when 16#01859# => romdata <= X"05040404";
    when 16#0185A# => romdata <= X"04050404";
    when 16#0185B# => romdata <= X"04040404";
    when 16#0185C# => romdata <= X"04040503";
    when 16#0185D# => romdata <= X"04040404";
    when 16#0185E# => romdata <= X"02020303";
    when 16#0185F# => romdata <= X"04040404";
    when 16#01860# => romdata <= X"04040405";
    when 16#01861# => romdata <= X"04040404";
    when 16#01862# => romdata <= X"04030303";
    when 16#01863# => romdata <= X"00005F07";
    when 16#01864# => romdata <= X"0007741C";
    when 16#01865# => romdata <= X"771C172E";
    when 16#01866# => romdata <= X"6A3E2B3A";
    when 16#01867# => romdata <= X"06493608";
    when 16#01868# => romdata <= X"36493036";
    when 16#01869# => romdata <= X"49597648";
    when 16#0186A# => romdata <= X"073C4281";
    when 16#0186B# => romdata <= X"81423C0A";
    when 16#0186C# => romdata <= X"041F040A";
    when 16#0186D# => romdata <= X"08083E08";
    when 16#0186E# => romdata <= X"08806008";
    when 16#0186F# => romdata <= X"080840C0";
    when 16#01870# => romdata <= X"300C033E";
    when 16#01871# => romdata <= X"4141413E";
    when 16#01872# => romdata <= X"44427F40";
    when 16#01873# => romdata <= X"40466151";
    when 16#01874# => romdata <= X"49462241";
    when 16#01875# => romdata <= X"49493618";
    when 16#01876# => romdata <= X"14127F10";
    when 16#01877# => romdata <= X"27454545";
    when 16#01878# => romdata <= X"393E4949";
    when 16#01879# => romdata <= X"49300101";
    when 16#0187A# => romdata <= X"710D0336";
    when 16#0187B# => romdata <= X"49494936";
    when 16#0187C# => romdata <= X"06494929";
    when 16#0187D# => romdata <= X"1E36D008";
    when 16#0187E# => romdata <= X"14224114";
    when 16#0187F# => romdata <= X"14141414";
    when 16#01880# => romdata <= X"41221408";
    when 16#01881# => romdata <= X"02510906";
    when 16#01882# => romdata <= X"3C4299A5";
    when 16#01883# => romdata <= X"BD421C7C";
    when 16#01884# => romdata <= X"1211127C";
    when 16#01885# => romdata <= X"7F494949";
    when 16#01886# => romdata <= X"363E4141";
    when 16#01887# => romdata <= X"41227F41";
    when 16#01888# => romdata <= X"41413E7F";
    when 16#01889# => romdata <= X"49494941";
    when 16#0188A# => romdata <= X"7F090909";
    when 16#0188B# => romdata <= X"013E4149";
    when 16#0188C# => romdata <= X"497A7F08";
    when 16#0188D# => romdata <= X"08087F41";
    when 16#0188E# => romdata <= X"7F414041";
    when 16#0188F# => romdata <= X"413F7F08";
    when 16#01890# => romdata <= X"1422417F";
    when 16#01891# => romdata <= X"40404040";
    when 16#01892# => romdata <= X"7F060C06";
    when 16#01893# => romdata <= X"7F7F0608";
    when 16#01894# => romdata <= X"307F3E41";
    when 16#01895# => romdata <= X"41413E7F";
    when 16#01896# => romdata <= X"09090906";
    when 16#01897# => romdata <= X"3E4161C1";
    when 16#01898# => romdata <= X"BE7F0919";
    when 16#01899# => romdata <= X"29462649";
    when 16#0189A# => romdata <= X"49493201";
    when 16#0189B# => romdata <= X"017F0101";
    when 16#0189C# => romdata <= X"3F404040";
    when 16#0189D# => romdata <= X"3F073840";
    when 16#0189E# => romdata <= X"38071F60";
    when 16#0189F# => romdata <= X"1F601F63";
    when 16#018A0# => romdata <= X"14081463";
    when 16#018A1# => romdata <= X"01067806";
    when 16#018A2# => romdata <= X"01615149";
    when 16#018A3# => romdata <= X"45437F41";
    when 16#018A4# => romdata <= X"41030C30";
    when 16#018A5# => romdata <= X"C041417F";
    when 16#018A6# => romdata <= X"04020102";
    when 16#018A7# => romdata <= X"04808080";
    when 16#018A8# => romdata <= X"80800102";
    when 16#018A9# => romdata <= X"20545454";
    when 16#018AA# => romdata <= X"787F4444";
    when 16#018AB# => romdata <= X"44383844";
    when 16#018AC# => romdata <= X"44443844";
    when 16#018AD# => romdata <= X"44447F38";
    when 16#018AE# => romdata <= X"54545458";
    when 16#018AF# => romdata <= X"087E0901";
    when 16#018B0# => romdata <= X"18A4A4A4";
    when 16#018B1# => romdata <= X"787F0404";
    when 16#018B2# => romdata <= X"787D807D";
    when 16#018B3# => romdata <= X"7F102844";
    when 16#018B4# => romdata <= X"3F407C04";
    when 16#018B5# => romdata <= X"7804787C";
    when 16#018B6# => romdata <= X"04047838";
    when 16#018B7# => romdata <= X"444438FC";
    when 16#018B8# => romdata <= X"24242418";
    when 16#018B9# => romdata <= X"18242424";
    when 16#018BA# => romdata <= X"FC7C0804";
    when 16#018BB# => romdata <= X"04485454";
    when 16#018BC# => romdata <= X"24043F44";
    when 16#018BD# => romdata <= X"403C4040";
    when 16#018BE# => romdata <= X"7C1C2040";
    when 16#018BF# => romdata <= X"201C1C60";
    when 16#018C0# => romdata <= X"601C6060";
    when 16#018C1# => romdata <= X"1C442810";
    when 16#018C2# => romdata <= X"28449CA0";
    when 16#018C3# => romdata <= X"601C6454";
    when 16#018C4# => romdata <= X"544C187E";
    when 16#018C5# => romdata <= X"8181FFFF";
    when 16#018C6# => romdata <= X"81817E18";
    when 16#018C7# => romdata <= X"18040810";
    when 16#018C8# => romdata <= X"0C143E55";
    when 16#018C9# => romdata <= X"55FF8181";
    when 16#018CA# => romdata <= X"81FF8060";
    when 16#018CB# => romdata <= X"80608060";
    when 16#018CC# => romdata <= X"60600060";
    when 16#018CD# => romdata <= X"60006060";
    when 16#018CE# => romdata <= X"047F0414";
    when 16#018CF# => romdata <= X"7F140201";
    when 16#018D0# => romdata <= X"01024629";
    when 16#018D1# => romdata <= X"1608344A";
    when 16#018D2# => romdata <= X"31483000";
    when 16#018D3# => romdata <= X"18243E41";
    when 16#018D4# => romdata <= X"227F4941";
    when 16#018D5# => romdata <= X"03040403";
    when 16#018D6# => romdata <= X"03040304";
    when 16#018D7# => romdata <= X"04030403";
    when 16#018D8# => romdata <= X"183C3C18";
    when 16#018D9# => romdata <= X"08080808";
    when 16#018DA# => romdata <= X"03010203";
    when 16#018DB# => romdata <= X"020E020E";
    when 16#018DC# => romdata <= X"060E0048";
    when 16#018DD# => romdata <= X"30384438";
    when 16#018DE# => romdata <= X"54483844";
    when 16#018DF# => romdata <= X"FE44487E";
    when 16#018E0# => romdata <= X"49014438";
    when 16#018E1# => romdata <= X"28384403";
    when 16#018E2# => romdata <= X"147C1403";
    when 16#018E3# => romdata <= X"E7E74E55";
    when 16#018E4# => romdata <= X"55390101";
    when 16#018E5# => romdata <= X"0001011C";
    when 16#018E6# => romdata <= X"2A555522";
    when 16#018E7# => romdata <= X"1C1D151E";
    when 16#018E8# => romdata <= X"18240018";
    when 16#018E9# => romdata <= X"24080808";
    when 16#018EA# => romdata <= X"18080808";
    when 16#018EB# => romdata <= X"3C42BD95";
    when 16#018EC# => romdata <= X"A9423C01";
    when 16#018ED# => romdata <= X"01010101";
    when 16#018EE# => romdata <= X"06090906";
    when 16#018EF# => romdata <= X"44445F44";
    when 16#018F0# => romdata <= X"44191512";
    when 16#018F1# => romdata <= X"15150A02";
    when 16#018F2# => romdata <= X"01FC2020";
    when 16#018F3# => romdata <= X"1C0E7F01";
    when 16#018F4# => romdata <= X"7F011818";
    when 16#018F5# => romdata <= X"00804002";
    when 16#018F6# => romdata <= X"1F060909";
    when 16#018F7# => romdata <= X"06241800";
    when 16#018F8# => romdata <= X"2418824F";
    when 16#018F9# => romdata <= X"304C62F1";
    when 16#018FA# => romdata <= X"824F300C";
    when 16#018FB# => romdata <= X"D2B1955F";
    when 16#018FC# => romdata <= X"304C62F1";
    when 16#018FD# => romdata <= X"30484520";
    when 16#018FE# => romdata <= X"60392E38";
    when 16#018FF# => romdata <= X"6060382E";
    when 16#01900# => romdata <= X"3960701D";
    when 16#01901# => romdata <= X"131D7072";
    when 16#01902# => romdata <= X"1D121E71";
    when 16#01903# => romdata <= X"701D121D";
    when 16#01904# => romdata <= X"70603B25";
    when 16#01905# => romdata <= X"3B607E11";
    when 16#01906# => romdata <= X"7F49411E";
    when 16#01907# => romdata <= X"2161927C";
    when 16#01908# => romdata <= X"5556447C";
    when 16#01909# => romdata <= X"5655447C";
    when 16#0190A# => romdata <= X"5655467D";
    when 16#0190B# => romdata <= X"54544545";
    when 16#0190C# => romdata <= X"7E44447E";
    when 16#0190D# => romdata <= X"45467D46";
    when 16#0190E# => romdata <= X"457C4508";
    when 16#0190F# => romdata <= X"7F49413E";
    when 16#01910# => romdata <= X"7E091222";
    when 16#01911# => romdata <= X"7D384546";
    when 16#01912# => romdata <= X"44383844";
    when 16#01913# => romdata <= X"46453838";
    when 16#01914# => romdata <= X"46454638";
    when 16#01915# => romdata <= X"3A454546";
    when 16#01916# => romdata <= X"39384544";
    when 16#01917# => romdata <= X"45382214";
    when 16#01918# => romdata <= X"081422BC";
    when 16#01919# => romdata <= X"625A463D";
    when 16#0191A# => romdata <= X"3C41423C";
    when 16#0191B# => romdata <= X"3C42413C";
    when 16#0191C# => romdata <= X"3C42413E";
    when 16#0191D# => romdata <= X"3D40403D";
    when 16#0191E# => romdata <= X"0608F209";
    when 16#0191F# => romdata <= X"067F2222";
    when 16#01920# => romdata <= X"1CFE0989";
    when 16#01921# => romdata <= X"76205556";
    when 16#01922# => romdata <= X"78205655";
    when 16#01923# => romdata <= X"78225555";
    when 16#01924# => romdata <= X"7A235556";
    when 16#01925# => romdata <= X"7B205554";
    when 16#01926# => romdata <= X"79275557";
    when 16#01927# => romdata <= X"78205438";
    when 16#01928# => romdata <= X"54483844";
    when 16#01929# => romdata <= X"C4385556";
    when 16#0192A# => romdata <= X"58385655";
    when 16#0192B# => romdata <= X"583A5555";
    when 16#0192C# => romdata <= X"5A395454";
    when 16#0192D# => romdata <= X"59017A7A";
    when 16#0192E# => romdata <= X"01027902";
    when 16#0192F# => romdata <= X"02780260";
    when 16#01930# => romdata <= X"91927C7B";
    when 16#01931# => romdata <= X"090A7338";
    when 16#01932# => romdata <= X"45463838";
    when 16#01933# => romdata <= X"4645383A";
    when 16#01934# => romdata <= X"45453A3B";
    when 16#01935# => romdata <= X"45463B39";
    when 16#01936# => romdata <= X"44443908";
    when 16#01937# => romdata <= X"082A0808";
    when 16#01938# => romdata <= X"B8644C3A";
    when 16#01939# => romdata <= X"3C41427C";
    when 16#0193A# => romdata <= X"3C42417C";
    when 16#0193B# => romdata <= X"3A41417A";
    when 16#0193C# => romdata <= X"3D40407D";
    when 16#0193D# => romdata <= X"986219FF";
    when 16#0193E# => romdata <= X"423C9A60";
    when 16#0193F# => romdata <= X"1A000000";
    when 16#01940# => romdata <= X"30622020";
    when 16#01941# => romdata <= X"20202020";
    when 16#01942# => romdata <= X"20202020";
    when 16#01943# => romdata <= X"20202020";
    when 16#01944# => romdata <= X"20202020";
    when 16#01945# => romdata <= X"20202020";
    when 16#01946# => romdata <= X"20202020";
    when 16#01947# => romdata <= X"20202020";
    when 16#01948# => romdata <= X"20200000";
    when 16#01949# => romdata <= X"20202020";
    when 16#0194A# => romdata <= X"20202020";
    when 16#0194B# => romdata <= X"00000000";
    when 16#0194C# => romdata <= X"00202020";
    when 16#0194D# => romdata <= X"20202020";
    when 16#0194E# => romdata <= X"20202828";
    when 16#0194F# => romdata <= X"28282820";
    when 16#01950# => romdata <= X"20202020";
    when 16#01951# => romdata <= X"20202020";
    when 16#01952# => romdata <= X"20202020";
    when 16#01953# => romdata <= X"20202020";
    when 16#01954# => romdata <= X"20881010";
    when 16#01955# => romdata <= X"10101010";
    when 16#01956# => romdata <= X"10101010";
    when 16#01957# => romdata <= X"10101010";
    when 16#01958# => romdata <= X"10040404";
    when 16#01959# => romdata <= X"04040404";
    when 16#0195A# => romdata <= X"04040410";
    when 16#0195B# => romdata <= X"10101010";
    when 16#0195C# => romdata <= X"10104141";
    when 16#0195D# => romdata <= X"41414141";
    when 16#0195E# => romdata <= X"01010101";
    when 16#0195F# => romdata <= X"01010101";
    when 16#01960# => romdata <= X"01010101";
    when 16#01961# => romdata <= X"01010101";
    when 16#01962# => romdata <= X"01010101";
    when 16#01963# => romdata <= X"10101010";
    when 16#01964# => romdata <= X"10104242";
    when 16#01965# => romdata <= X"42424242";
    when 16#01966# => romdata <= X"02020202";
    when 16#01967# => romdata <= X"02020202";
    when 16#01968# => romdata <= X"02020202";
    when 16#01969# => romdata <= X"02020202";
    when 16#0196A# => romdata <= X"02020202";
    when 16#0196B# => romdata <= X"10101010";
    when 16#0196C# => romdata <= X"20000000";
    when 16#0196D# => romdata <= X"00000000";
    when 16#0196E# => romdata <= X"00000000";
    when 16#0196F# => romdata <= X"00000000";
    when 16#01970# => romdata <= X"00000000";
    when 16#01971# => romdata <= X"00000000";
    when 16#01972# => romdata <= X"00000000";
    when 16#01973# => romdata <= X"00000000";
    when 16#01974# => romdata <= X"00000000";
    when 16#01975# => romdata <= X"00000000";
    when 16#01976# => romdata <= X"00000000";
    when 16#01977# => romdata <= X"00000000";
    when 16#01978# => romdata <= X"00000000";
    when 16#01979# => romdata <= X"00000000";
    when 16#0197A# => romdata <= X"00000000";
    when 16#0197B# => romdata <= X"00000000";
    when 16#0197C# => romdata <= X"00000000";
    when 16#0197D# => romdata <= X"00000000";
    when 16#0197E# => romdata <= X"00000000";
    when 16#0197F# => romdata <= X"00000000";
    when 16#01980# => romdata <= X"00000000";
    when 16#01981# => romdata <= X"00000000";
    when 16#01982# => romdata <= X"00000000";
    when 16#01983# => romdata <= X"00000000";
    when 16#01984# => romdata <= X"00000000";
    when 16#01985# => romdata <= X"00000000";
    when 16#01986# => romdata <= X"00000000";
    when 16#01987# => romdata <= X"00000000";
    when 16#01988# => romdata <= X"00000000";
    when 16#01989# => romdata <= X"00000000";
    when 16#0198A# => romdata <= X"00000000";
    when 16#0198B# => romdata <= X"00000000";
    when 16#0198C# => romdata <= X"00000000";
    when 16#0198D# => romdata <= X"43000000";
    when 16#0198E# => romdata <= X"00000000";
    when 16#0198F# => romdata <= X"80000C00";
    when 16#01990# => romdata <= X"80000B00";
    when 16#01991# => romdata <= X"80000800";
    when 16#01992# => romdata <= X"00000000";
    when 16#01993# => romdata <= X"FF000000";
    when 16#01994# => romdata <= X"00000000";
    when 16#01995# => romdata <= X"00000000";
    when 16#01996# => romdata <= X"00FFFFFF";
    when 16#01997# => romdata <= X"FF00FFFF";
    when 16#01998# => romdata <= X"FFFF00FF";
    when 16#01999# => romdata <= X"FFFFFF00";
    when 16#0199A# => romdata <= X"00000000";
    when 16#0199B# => romdata <= X"00000000";
    when 16#0199C# => romdata <= X"80000A00";
    when 16#0199D# => romdata <= X"80000700";
    when 16#0199E# => romdata <= X"80000600";
    when 16#0199F# => romdata <= X"80000400";
    when 16#019A0# => romdata <= X"80000200";
    when 16#019A1# => romdata <= X"80000100";
    when 16#019A2# => romdata <= X"80000004";
    when 16#019A3# => romdata <= X"80000000";
    when 16#019A4# => romdata <= X"00006694";
    when 16#019A5# => romdata <= X"00000000";
    when 16#019A6# => romdata <= X"000068FC";
    when 16#019A7# => romdata <= X"00006958";
    when 16#019A8# => romdata <= X"000069B4";
    when 16#019A9# => romdata <= X"00000000";
    when 16#019AA# => romdata <= X"00000000";
    when 16#019AB# => romdata <= X"00000000";
    when 16#019AC# => romdata <= X"00000000";
    when 16#019AD# => romdata <= X"00000000";
    when 16#019AE# => romdata <= X"00000000";
    when 16#019AF# => romdata <= X"00000000";
    when 16#019B0# => romdata <= X"00000000";
    when 16#019B1# => romdata <= X"00000000";
    when 16#019B2# => romdata <= X"00006634";
    when 16#019B3# => romdata <= X"00000000";
    when 16#019B4# => romdata <= X"00000000";
    when 16#019B5# => romdata <= X"00000000";
    when 16#019B6# => romdata <= X"00000000";
    when 16#019B7# => romdata <= X"00000000";
    when 16#019B8# => romdata <= X"00000000";
    when 16#019B9# => romdata <= X"00000000";
    when 16#019BA# => romdata <= X"00000000";
    when 16#019BB# => romdata <= X"00000000";
    when 16#019BC# => romdata <= X"00000000";
    when 16#019BD# => romdata <= X"00000000";
    when 16#019BE# => romdata <= X"00000000";
    when 16#019BF# => romdata <= X"00000000";
    when 16#019C0# => romdata <= X"00000000";
    when 16#019C1# => romdata <= X"00000000";
    when 16#019C2# => romdata <= X"00000000";
    when 16#019C3# => romdata <= X"00000000";
    when 16#019C4# => romdata <= X"00000000";
    when 16#019C5# => romdata <= X"00000000";
    when 16#019C6# => romdata <= X"00000000";
    when 16#019C7# => romdata <= X"00000000";
    when 16#019C8# => romdata <= X"00000000";
    when 16#019C9# => romdata <= X"00000000";
    when 16#019CA# => romdata <= X"00000000";
    when 16#019CB# => romdata <= X"00000000";
    when 16#019CC# => romdata <= X"00000000";
    when 16#019CD# => romdata <= X"00000000";
    when 16#019CE# => romdata <= X"00000000";
    when 16#019CF# => romdata <= X"00000001";
    when 16#019D0# => romdata <= X"330EABCD";
    when 16#019D1# => romdata <= X"1234E66D";
    when 16#019D2# => romdata <= X"DEEC0005";
    when 16#019D3# => romdata <= X"000B0000";
    when 16#019D4# => romdata <= X"00000000";
    when 16#019D5# => romdata <= X"00000000";
    when 16#019D6# => romdata <= X"00000000";
    when 16#019D7# => romdata <= X"00000000";
    when 16#019D8# => romdata <= X"00000000";
    when 16#019D9# => romdata <= X"00000000";
    when 16#019DA# => romdata <= X"00000000";
    when 16#019DB# => romdata <= X"00000000";
    when 16#019DC# => romdata <= X"00000000";
    when 16#019DD# => romdata <= X"00000000";
    when 16#019DE# => romdata <= X"00000000";
    when 16#019DF# => romdata <= X"00000000";
    when 16#019E0# => romdata <= X"00000000";
    when 16#019E1# => romdata <= X"00000000";
    when 16#019E2# => romdata <= X"00000000";
    when 16#019E3# => romdata <= X"00000000";
    when 16#019E4# => romdata <= X"00000000";
    when 16#019E5# => romdata <= X"00000000";
    when 16#019E6# => romdata <= X"00000000";
    when 16#019E7# => romdata <= X"00000000";
    when 16#019E8# => romdata <= X"00000000";
    when 16#019E9# => romdata <= X"00000000";
    when 16#019EA# => romdata <= X"00000000";
    when 16#019EB# => romdata <= X"00000000";
    when 16#019EC# => romdata <= X"00000000";
    when 16#019ED# => romdata <= X"00000000";
    when 16#019EE# => romdata <= X"00000000";
    when 16#019EF# => romdata <= X"00000000";
    when 16#019F0# => romdata <= X"00000000";
    when 16#019F1# => romdata <= X"00000000";
    when 16#019F2# => romdata <= X"00000000";
    when 16#019F3# => romdata <= X"00000000";
    when 16#019F4# => romdata <= X"00000000";
    when 16#019F5# => romdata <= X"00000000";
    when 16#019F6# => romdata <= X"00000000";
    when 16#019F7# => romdata <= X"00000000";
    when 16#019F8# => romdata <= X"00000000";
    when 16#019F9# => romdata <= X"00000000";
    when 16#019FA# => romdata <= X"00000000";
    when 16#019FB# => romdata <= X"00000000";
    when 16#019FC# => romdata <= X"00000000";
    when 16#019FD# => romdata <= X"00000000";
    when 16#019FE# => romdata <= X"00000000";
    when 16#019FF# => romdata <= X"00000000";
    when 16#01A00# => romdata <= X"00000000";
    when 16#01A01# => romdata <= X"00000000";
    when 16#01A02# => romdata <= X"00000000";
    when 16#01A03# => romdata <= X"00000000";
    when 16#01A04# => romdata <= X"00000000";
    when 16#01A05# => romdata <= X"00000000";
    when 16#01A06# => romdata <= X"00000000";
    when 16#01A07# => romdata <= X"00000000";
    when 16#01A08# => romdata <= X"00000000";
    when 16#01A09# => romdata <= X"00000000";
    when 16#01A0A# => romdata <= X"00000000";
    when 16#01A0B# => romdata <= X"00000000";
    when 16#01A0C# => romdata <= X"00000000";
    when 16#01A0D# => romdata <= X"00000000";
    when 16#01A0E# => romdata <= X"00000000";
    when 16#01A0F# => romdata <= X"00000000";
    when 16#01A10# => romdata <= X"00000000";
    when 16#01A11# => romdata <= X"00000000";
    when 16#01A12# => romdata <= X"00000000";
    when 16#01A13# => romdata <= X"00000000";
    when 16#01A14# => romdata <= X"00000000";
    when 16#01A15# => romdata <= X"00000000";
    when 16#01A16# => romdata <= X"00000000";
    when 16#01A17# => romdata <= X"00000000";
    when 16#01A18# => romdata <= X"00000000";
    when 16#01A19# => romdata <= X"00000000";
    when 16#01A1A# => romdata <= X"00000000";
    when 16#01A1B# => romdata <= X"00000000";
    when 16#01A1C# => romdata <= X"00000000";
    when 16#01A1D# => romdata <= X"00000000";
    when 16#01A1E# => romdata <= X"00000000";
    when 16#01A1F# => romdata <= X"00000000";
    when 16#01A20# => romdata <= X"00000000";
    when 16#01A21# => romdata <= X"00000000";
    when 16#01A22# => romdata <= X"00000000";
    when 16#01A23# => romdata <= X"00000000";
    when 16#01A24# => romdata <= X"00000000";
    when 16#01A25# => romdata <= X"00000000";
    when 16#01A26# => romdata <= X"00000000";
    when 16#01A27# => romdata <= X"00000000";
    when 16#01A28# => romdata <= X"00000000";
    when 16#01A29# => romdata <= X"00000000";
    when 16#01A2A# => romdata <= X"00000000";
    when 16#01A2B# => romdata <= X"00000000";
    when 16#01A2C# => romdata <= X"00000000";
    when 16#01A2D# => romdata <= X"00000000";
    when 16#01A2E# => romdata <= X"00000000";
    when 16#01A2F# => romdata <= X"00000000";
    when 16#01A30# => romdata <= X"00000000";
    when 16#01A31# => romdata <= X"00000000";
    when 16#01A32# => romdata <= X"00000000";
    when 16#01A33# => romdata <= X"00000000";
    when 16#01A34# => romdata <= X"00000000";
    when 16#01A35# => romdata <= X"00000000";
    when 16#01A36# => romdata <= X"00000000";
    when 16#01A37# => romdata <= X"00000000";
    when 16#01A38# => romdata <= X"00000000";
    when 16#01A39# => romdata <= X"00000000";
    when 16#01A3A# => romdata <= X"00000000";
    when 16#01A3B# => romdata <= X"00000000";
    when 16#01A3C# => romdata <= X"00000000";
    when 16#01A3D# => romdata <= X"00000000";
    when 16#01A3E# => romdata <= X"00000000";
    when 16#01A3F# => romdata <= X"00000000";
    when 16#01A40# => romdata <= X"00000000";
    when 16#01A41# => romdata <= X"00000000";
    when 16#01A42# => romdata <= X"00000000";
    when 16#01A43# => romdata <= X"00000000";
    when 16#01A44# => romdata <= X"00000000";
    when 16#01A45# => romdata <= X"00000000";
    when 16#01A46# => romdata <= X"00000000";
    when 16#01A47# => romdata <= X"00000000";
    when 16#01A48# => romdata <= X"00000000";
    when 16#01A49# => romdata <= X"00000000";
    when 16#01A4A# => romdata <= X"00000000";
    when 16#01A4B# => romdata <= X"00000000";
    when 16#01A4C# => romdata <= X"00000000";
    when 16#01A4D# => romdata <= X"00000000";
    when 16#01A4E# => romdata <= X"00000000";
    when 16#01A4F# => romdata <= X"00000000";
    when 16#01A50# => romdata <= X"00000000";
    when 16#01A51# => romdata <= X"00000000";
    when 16#01A52# => romdata <= X"00000000";
    when 16#01A53# => romdata <= X"00000000";
    when 16#01A54# => romdata <= X"00000000";
    when 16#01A55# => romdata <= X"00000000";
    when 16#01A56# => romdata <= X"00000000";
    when 16#01A57# => romdata <= X"00000000";
    when 16#01A58# => romdata <= X"00000000";
    when 16#01A59# => romdata <= X"00000000";
    when 16#01A5A# => romdata <= X"00000000";
    when 16#01A5B# => romdata <= X"00000000";
    when 16#01A5C# => romdata <= X"00000000";
    when 16#01A5D# => romdata <= X"00000000";
    when 16#01A5E# => romdata <= X"00000000";
    when 16#01A5F# => romdata <= X"00000000";
    when 16#01A60# => romdata <= X"00000000";
    when 16#01A61# => romdata <= X"00000000";
    when 16#01A62# => romdata <= X"00000000";
    when 16#01A63# => romdata <= X"00000000";
    when 16#01A64# => romdata <= X"00000000";
    when 16#01A65# => romdata <= X"00000000";
    when 16#01A66# => romdata <= X"00000000";
    when 16#01A67# => romdata <= X"00000000";
    when 16#01A68# => romdata <= X"00000000";
    when 16#01A69# => romdata <= X"00000000";
    when 16#01A6A# => romdata <= X"00000000";
    when 16#01A6B# => romdata <= X"00000000";
    when 16#01A6C# => romdata <= X"00000000";
    when 16#01A6D# => romdata <= X"00000000";
    when 16#01A6E# => romdata <= X"00000000";
    when 16#01A6F# => romdata <= X"00000000";
    when 16#01A70# => romdata <= X"00000000";
    when 16#01A71# => romdata <= X"00000000";
    when 16#01A72# => romdata <= X"00000000";
    when 16#01A73# => romdata <= X"00000000";
    when 16#01A74# => romdata <= X"00000000";
    when 16#01A75# => romdata <= X"00000000";
    when 16#01A76# => romdata <= X"00000000";
    when 16#01A77# => romdata <= X"00000000";
    when 16#01A78# => romdata <= X"00000000";
    when 16#01A79# => romdata <= X"00000000";
    when 16#01A7A# => romdata <= X"00000000";
    when 16#01A7B# => romdata <= X"00000000";
    when 16#01A7C# => romdata <= X"00000000";
    when 16#01A7D# => romdata <= X"00000000";
    when 16#01A7E# => romdata <= X"00000000";
    when 16#01A7F# => romdata <= X"00000000";
    when 16#01A80# => romdata <= X"00000000";
    when 16#01A81# => romdata <= X"00000000";
    when 16#01A82# => romdata <= X"00000000";
    when 16#01A83# => romdata <= X"00000000";
    when 16#01A84# => romdata <= X"00000000";
    when 16#01A85# => romdata <= X"00000000";
    when 16#01A86# => romdata <= X"00000000";
    when 16#01A87# => romdata <= X"00000000";
    when 16#01A88# => romdata <= X"00000000";
    when 16#01A89# => romdata <= X"00000000";
    when 16#01A8A# => romdata <= X"00000000";
    when 16#01A8B# => romdata <= X"00000000";
    when 16#01A8C# => romdata <= X"00000000";
    when 16#01A8D# => romdata <= X"00000000";
    when 16#01A8E# => romdata <= X"00000000";
    when 16#01A8F# => romdata <= X"00000000";
    when 16#01A90# => romdata <= X"FFFFFFFF";
    when 16#01A91# => romdata <= X"00000000";
    when 16#01A92# => romdata <= X"00020000";
    when 16#01A93# => romdata <= X"00000000";
    when 16#01A94# => romdata <= X"00000000";
    when 16#01A95# => romdata <= X"00006A4C";
    when 16#01A96# => romdata <= X"00006A4C";
    when 16#01A97# => romdata <= X"00006A54";
    when 16#01A98# => romdata <= X"00006A54";
    when 16#01A99# => romdata <= X"00006A5C";
    when 16#01A9A# => romdata <= X"00006A5C";
    when 16#01A9B# => romdata <= X"00006A64";
    when 16#01A9C# => romdata <= X"00006A64";
    when 16#01A9D# => romdata <= X"00006A6C";
    when 16#01A9E# => romdata <= X"00006A6C";
    when 16#01A9F# => romdata <= X"00006A74";
    when 16#01AA0# => romdata <= X"00006A74";
    when 16#01AA1# => romdata <= X"00006A7C";
    when 16#01AA2# => romdata <= X"00006A7C";
    when 16#01AA3# => romdata <= X"00006A84";
    when 16#01AA4# => romdata <= X"00006A84";
    when 16#01AA5# => romdata <= X"00006A8C";
    when 16#01AA6# => romdata <= X"00006A8C";
    when 16#01AA7# => romdata <= X"00006A94";
    when 16#01AA8# => romdata <= X"00006A94";
    when 16#01AA9# => romdata <= X"00006A9C";
    when 16#01AAA# => romdata <= X"00006A9C";
    when 16#01AAB# => romdata <= X"00006AA4";
    when 16#01AAC# => romdata <= X"00006AA4";
    when 16#01AAD# => romdata <= X"00006AAC";
    when 16#01AAE# => romdata <= X"00006AAC";
    when 16#01AAF# => romdata <= X"00006AB4";
    when 16#01AB0# => romdata <= X"00006AB4";
    when 16#01AB1# => romdata <= X"00006ABC";
    when 16#01AB2# => romdata <= X"00006ABC";
    when 16#01AB3# => romdata <= X"00006AC4";
    when 16#01AB4# => romdata <= X"00006AC4";
    when 16#01AB5# => romdata <= X"00006ACC";
    when 16#01AB6# => romdata <= X"00006ACC";
    when 16#01AB7# => romdata <= X"00006AD4";
    when 16#01AB8# => romdata <= X"00006AD4";
    when 16#01AB9# => romdata <= X"00006ADC";
    when 16#01ABA# => romdata <= X"00006ADC";
    when 16#01ABB# => romdata <= X"00006AE4";
    when 16#01ABC# => romdata <= X"00006AE4";
    when 16#01ABD# => romdata <= X"00006AEC";
    when 16#01ABE# => romdata <= X"00006AEC";
    when 16#01ABF# => romdata <= X"00006AF4";
    when 16#01AC0# => romdata <= X"00006AF4";
    when 16#01AC1# => romdata <= X"00006AFC";
    when 16#01AC2# => romdata <= X"00006AFC";
    when 16#01AC3# => romdata <= X"00006B04";
    when 16#01AC4# => romdata <= X"00006B04";
    when 16#01AC5# => romdata <= X"00006B0C";
    when 16#01AC6# => romdata <= X"00006B0C";
    when 16#01AC7# => romdata <= X"00006B14";
    when 16#01AC8# => romdata <= X"00006B14";
    when 16#01AC9# => romdata <= X"00006B1C";
    when 16#01ACA# => romdata <= X"00006B1C";
    when 16#01ACB# => romdata <= X"00006B24";
    when 16#01ACC# => romdata <= X"00006B24";
    when 16#01ACD# => romdata <= X"00006B2C";
    when 16#01ACE# => romdata <= X"00006B2C";
    when 16#01ACF# => romdata <= X"00006B34";
    when 16#01AD0# => romdata <= X"00006B34";
    when 16#01AD1# => romdata <= X"00006B3C";
    when 16#01AD2# => romdata <= X"00006B3C";
    when 16#01AD3# => romdata <= X"00006B44";
    when 16#01AD4# => romdata <= X"00006B44";
    when 16#01AD5# => romdata <= X"00006B4C";
    when 16#01AD6# => romdata <= X"00006B4C";
    when 16#01AD7# => romdata <= X"00006B54";
    when 16#01AD8# => romdata <= X"00006B54";
    when 16#01AD9# => romdata <= X"00006B5C";
    when 16#01ADA# => romdata <= X"00006B5C";
    when 16#01ADB# => romdata <= X"00006B64";
    when 16#01ADC# => romdata <= X"00006B64";
    when 16#01ADD# => romdata <= X"00006B6C";
    when 16#01ADE# => romdata <= X"00006B6C";
    when 16#01ADF# => romdata <= X"00006B74";
    when 16#01AE0# => romdata <= X"00006B74";
    when 16#01AE1# => romdata <= X"00006B7C";
    when 16#01AE2# => romdata <= X"00006B7C";
    when 16#01AE3# => romdata <= X"00006B84";
    when 16#01AE4# => romdata <= X"00006B84";
    when 16#01AE5# => romdata <= X"00006B8C";
    when 16#01AE6# => romdata <= X"00006B8C";
    when 16#01AE7# => romdata <= X"00006B94";
    when 16#01AE8# => romdata <= X"00006B94";
    when 16#01AE9# => romdata <= X"00006B9C";
    when 16#01AEA# => romdata <= X"00006B9C";
    when 16#01AEB# => romdata <= X"00006BA4";
    when 16#01AEC# => romdata <= X"00006BA4";
    when 16#01AED# => romdata <= X"00006BAC";
    when 16#01AEE# => romdata <= X"00006BAC";
    when 16#01AEF# => romdata <= X"00006BB4";
    when 16#01AF0# => romdata <= X"00006BB4";
    when 16#01AF1# => romdata <= X"00006BBC";
    when 16#01AF2# => romdata <= X"00006BBC";
    when 16#01AF3# => romdata <= X"00006BC4";
    when 16#01AF4# => romdata <= X"00006BC4";
    when 16#01AF5# => romdata <= X"00006BCC";
    when 16#01AF6# => romdata <= X"00006BCC";
    when 16#01AF7# => romdata <= X"00006BD4";
    when 16#01AF8# => romdata <= X"00006BD4";
    when 16#01AF9# => romdata <= X"00006BDC";
    when 16#01AFA# => romdata <= X"00006BDC";
    when 16#01AFB# => romdata <= X"00006BE4";
    when 16#01AFC# => romdata <= X"00006BE4";
    when 16#01AFD# => romdata <= X"00006BEC";
    when 16#01AFE# => romdata <= X"00006BEC";
    when 16#01AFF# => romdata <= X"00006BF4";
    when 16#01B00# => romdata <= X"00006BF4";
    when 16#01B01# => romdata <= X"00006BFC";
    when 16#01B02# => romdata <= X"00006BFC";
    when 16#01B03# => romdata <= X"00006C04";
    when 16#01B04# => romdata <= X"00006C04";
    when 16#01B05# => romdata <= X"00006C0C";
    when 16#01B06# => romdata <= X"00006C0C";
    when 16#01B07# => romdata <= X"00006C14";
    when 16#01B08# => romdata <= X"00006C14";
    when 16#01B09# => romdata <= X"00006C1C";
    when 16#01B0A# => romdata <= X"00006C1C";
    when 16#01B0B# => romdata <= X"00006C24";
    when 16#01B0C# => romdata <= X"00006C24";
    when 16#01B0D# => romdata <= X"00006C2C";
    when 16#01B0E# => romdata <= X"00006C2C";
    when 16#01B0F# => romdata <= X"00006C34";
    when 16#01B10# => romdata <= X"00006C34";
    when 16#01B11# => romdata <= X"00006C3C";
    when 16#01B12# => romdata <= X"00006C3C";
    when 16#01B13# => romdata <= X"00006C44";
    when 16#01B14# => romdata <= X"00006C44";
    when 16#01B15# => romdata <= X"00006C4C";
    when 16#01B16# => romdata <= X"00006C4C";
    when 16#01B17# => romdata <= X"00006C54";
    when 16#01B18# => romdata <= X"00006C54";
    when 16#01B19# => romdata <= X"00006C5C";
    when 16#01B1A# => romdata <= X"00006C5C";
    when 16#01B1B# => romdata <= X"00006C64";
    when 16#01B1C# => romdata <= X"00006C64";
    when 16#01B1D# => romdata <= X"00006C6C";
    when 16#01B1E# => romdata <= X"00006C6C";
    when 16#01B1F# => romdata <= X"00006C74";
    when 16#01B20# => romdata <= X"00006C74";
    when 16#01B21# => romdata <= X"00006C7C";
    when 16#01B22# => romdata <= X"00006C7C";
    when 16#01B23# => romdata <= X"00006C84";
    when 16#01B24# => romdata <= X"00006C84";
    when 16#01B25# => romdata <= X"00006C8C";
    when 16#01B26# => romdata <= X"00006C8C";
    when 16#01B27# => romdata <= X"00006C94";
    when 16#01B28# => romdata <= X"00006C94";
    when 16#01B29# => romdata <= X"00006C9C";
    when 16#01B2A# => romdata <= X"00006C9C";
    when 16#01B2B# => romdata <= X"00006CA4";
    when 16#01B2C# => romdata <= X"00006CA4";
    when 16#01B2D# => romdata <= X"00006CAC";
    when 16#01B2E# => romdata <= X"00006CAC";
    when 16#01B2F# => romdata <= X"00006CB4";
    when 16#01B30# => romdata <= X"00006CB4";
    when 16#01B31# => romdata <= X"00006CBC";
    when 16#01B32# => romdata <= X"00006CBC";
    when 16#01B33# => romdata <= X"00006CC4";
    when 16#01B34# => romdata <= X"00006CC4";
    when 16#01B35# => romdata <= X"00006CCC";
    when 16#01B36# => romdata <= X"00006CCC";
    when 16#01B37# => romdata <= X"00006CD4";
    when 16#01B38# => romdata <= X"00006CD4";
    when 16#01B39# => romdata <= X"00006CDC";
    when 16#01B3A# => romdata <= X"00006CDC";
    when 16#01B3B# => romdata <= X"00006CE4";
    when 16#01B3C# => romdata <= X"00006CE4";
    when 16#01B3D# => romdata <= X"00006CEC";
    when 16#01B3E# => romdata <= X"00006CEC";
    when 16#01B3F# => romdata <= X"00006CF4";
    when 16#01B40# => romdata <= X"00006CF4";
    when 16#01B41# => romdata <= X"00006CFC";
    when 16#01B42# => romdata <= X"00006CFC";
    when 16#01B43# => romdata <= X"00006D04";
    when 16#01B44# => romdata <= X"00006D04";
    when 16#01B45# => romdata <= X"00006D0C";
    when 16#01B46# => romdata <= X"00006D0C";
    when 16#01B47# => romdata <= X"00006D14";
    when 16#01B48# => romdata <= X"00006D14";
    when 16#01B49# => romdata <= X"00006D1C";
    when 16#01B4A# => romdata <= X"00006D1C";
    when 16#01B4B# => romdata <= X"00006D24";
    when 16#01B4C# => romdata <= X"00006D24";
    when 16#01B4D# => romdata <= X"00006D2C";
    when 16#01B4E# => romdata <= X"00006D2C";
    when 16#01B4F# => romdata <= X"00006D34";
    when 16#01B50# => romdata <= X"00006D34";
    when 16#01B51# => romdata <= X"00006D3C";
    when 16#01B52# => romdata <= X"00006D3C";
    when 16#01B53# => romdata <= X"00006D44";
    when 16#01B54# => romdata <= X"00006D44";
    when 16#01B55# => romdata <= X"00006D4C";
    when 16#01B56# => romdata <= X"00006D4C";
    when 16#01B57# => romdata <= X"00006D54";
    when 16#01B58# => romdata <= X"00006D54";
    when 16#01B59# => romdata <= X"00006D5C";
    when 16#01B5A# => romdata <= X"00006D5C";
    when 16#01B5B# => romdata <= X"00006D64";
    when 16#01B5C# => romdata <= X"00006D64";
    when 16#01B5D# => romdata <= X"00006D6C";
    when 16#01B5E# => romdata <= X"00006D6C";
    when 16#01B5F# => romdata <= X"00006D74";
    when 16#01B60# => romdata <= X"00006D74";
    when 16#01B61# => romdata <= X"00006D7C";
    when 16#01B62# => romdata <= X"00006D7C";
    when 16#01B63# => romdata <= X"00006D84";
    when 16#01B64# => romdata <= X"00006D84";
    when 16#01B65# => romdata <= X"00006D8C";
    when 16#01B66# => romdata <= X"00006D8C";
    when 16#01B67# => romdata <= X"00006D94";
    when 16#01B68# => romdata <= X"00006D94";
    when 16#01B69# => romdata <= X"00006D9C";
    when 16#01B6A# => romdata <= X"00006D9C";
    when 16#01B6B# => romdata <= X"00006DA4";
    when 16#01B6C# => romdata <= X"00006DA4";
    when 16#01B6D# => romdata <= X"00006DAC";
    when 16#01B6E# => romdata <= X"00006DAC";
    when 16#01B6F# => romdata <= X"00006DB4";
    when 16#01B70# => romdata <= X"00006DB4";
    when 16#01B71# => romdata <= X"00006DBC";
    when 16#01B72# => romdata <= X"00006DBC";
    when 16#01B73# => romdata <= X"00006DC4";
    when 16#01B74# => romdata <= X"00006DC4";
    when 16#01B75# => romdata <= X"00006DCC";
    when 16#01B76# => romdata <= X"00006DCC";
    when 16#01B77# => romdata <= X"00006DD4";
    when 16#01B78# => romdata <= X"00006DD4";
    when 16#01B79# => romdata <= X"00006DDC";
    when 16#01B7A# => romdata <= X"00006DDC";
    when 16#01B7B# => romdata <= X"00006DE4";
    when 16#01B7C# => romdata <= X"00006DE4";
    when 16#01B7D# => romdata <= X"00006DEC";
    when 16#01B7E# => romdata <= X"00006DEC";
    when 16#01B7F# => romdata <= X"00006DF4";
    when 16#01B80# => romdata <= X"00006DF4";
    when 16#01B81# => romdata <= X"00006DFC";
    when 16#01B82# => romdata <= X"00006DFC";
    when 16#01B83# => romdata <= X"00006E04";
    when 16#01B84# => romdata <= X"00006E04";
    when 16#01B85# => romdata <= X"00006E0C";
    when 16#01B86# => romdata <= X"00006E0C";
    when 16#01B87# => romdata <= X"00006E14";
    when 16#01B88# => romdata <= X"00006E14";
    when 16#01B89# => romdata <= X"00006E1C";
    when 16#01B8A# => romdata <= X"00006E1C";
    when 16#01B8B# => romdata <= X"00006E24";
    when 16#01B8C# => romdata <= X"00006E24";
    when 16#01B8D# => romdata <= X"00006E2C";
    when 16#01B8E# => romdata <= X"00006E2C";
    when 16#01B8F# => romdata <= X"00006E34";
    when 16#01B90# => romdata <= X"00006E34";
    when 16#01B91# => romdata <= X"00006E3C";
    when 16#01B92# => romdata <= X"00006E3C";
    when 16#01B93# => romdata <= X"00006E44";
    when 16#01B94# => romdata <= X"00006E44";
    when 16#01B95# => romdata <= X"00006E44";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
