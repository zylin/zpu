-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80d1d00c",
     3 => x"3a0b0b80",
     4 => x"c9ac0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80c9f72d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80d1",
   162 => x"bc738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8b",
   171 => x"8c2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8c",
   179 => x"be2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80d1cc0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82c73f80",
   257 => x"c8bf3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"fe3d0d0b",
   281 => x"0b80e1b8",
   282 => x"08538413",
   283 => x"0870882a",
   284 => x"70810651",
   285 => x"52527080",
   286 => x"2ef03871",
   287 => x"81ff0680",
   288 => x"0c843d0d",
   289 => x"04ff3d0d",
   290 => x"0b0b80e1",
   291 => x"b8085271",
   292 => x"0870882a",
   293 => x"81327081",
   294 => x"06515151",
   295 => x"70f13873",
   296 => x"720c833d",
   297 => x"0d0480d1",
   298 => x"cc08802e",
   299 => x"a43880d1",
   300 => x"d008822e",
   301 => x"bd388380",
   302 => x"800b0b0b",
   303 => x"80e1b80c",
   304 => x"82a0800b",
   305 => x"80e1bc0c",
   306 => x"8290800b",
   307 => x"80e1c00c",
   308 => x"04f88080",
   309 => x"80a40b0b",
   310 => x"0b80e1b8",
   311 => x"0cf88080",
   312 => x"82800b80",
   313 => x"e1bc0cf8",
   314 => x"80808480",
   315 => x"0b80e1c0",
   316 => x"0c0480c0",
   317 => x"a8808c0b",
   318 => x"0b0b80e1",
   319 => x"b80c80c0",
   320 => x"a880940b",
   321 => x"80e1bc0c",
   322 => x"0b0b80d0",
   323 => x"f40b80e1",
   324 => x"c00c04ff",
   325 => x"3d0d80e1",
   326 => x"c4335170",
   327 => x"a73880d1",
   328 => x"d8087008",
   329 => x"52527080",
   330 => x"2e943884",
   331 => x"1280d1d8",
   332 => x"0c702d80",
   333 => x"d1d80870",
   334 => x"08525270",
   335 => x"ee38810b",
   336 => x"80e1c434",
   337 => x"833d0d04",
   338 => x"04803d0d",
   339 => x"0b0b80e1",
   340 => x"b408802e",
   341 => x"8e380b0b",
   342 => x"0b0b800b",
   343 => x"802e0981",
   344 => x"06853882",
   345 => x"3d0d040b",
   346 => x"0b80e1b4",
   347 => x"510b0b0b",
   348 => x"f58e3f82",
   349 => x"3d0d0404",
   350 => x"803d0d80",
   351 => x"d0f85185",
   352 => x"ed3f80d1",
   353 => x"945185e6",
   354 => x"3f83fd3f",
   355 => x"8c08028c",
   356 => x"0cf93d0d",
   357 => x"800b8c08",
   358 => x"fc050c8c",
   359 => x"08880508",
   360 => x"8025ab38",
   361 => x"8c088805",
   362 => x"08308c08",
   363 => x"88050c80",
   364 => x"0b8c08f4",
   365 => x"050c8c08",
   366 => x"fc050888",
   367 => x"38810b8c",
   368 => x"08f4050c",
   369 => x"8c08f405",
   370 => x"088c08fc",
   371 => x"050c8c08",
   372 => x"8c050880",
   373 => x"25ab388c",
   374 => x"088c0508",
   375 => x"308c088c",
   376 => x"050c800b",
   377 => x"8c08f005",
   378 => x"0c8c08fc",
   379 => x"05088838",
   380 => x"810b8c08",
   381 => x"f0050c8c",
   382 => x"08f00508",
   383 => x"8c08fc05",
   384 => x"0c80538c",
   385 => x"088c0508",
   386 => x"528c0888",
   387 => x"05085181",
   388 => x"a73f8008",
   389 => x"708c08f8",
   390 => x"050c548c",
   391 => x"08fc0508",
   392 => x"802e8c38",
   393 => x"8c08f805",
   394 => x"08308c08",
   395 => x"f8050c8c",
   396 => x"08f80508",
   397 => x"70800c54",
   398 => x"893d0d8c",
   399 => x"0c048c08",
   400 => x"028c0cfb",
   401 => x"3d0d800b",
   402 => x"8c08fc05",
   403 => x"0c8c0888",
   404 => x"05088025",
   405 => x"93388c08",
   406 => x"88050830",
   407 => x"8c088805",
   408 => x"0c810b8c",
   409 => x"08fc050c",
   410 => x"8c088c05",
   411 => x"0880258c",
   412 => x"388c088c",
   413 => x"0508308c",
   414 => x"088c050c",
   415 => x"81538c08",
   416 => x"8c050852",
   417 => x"8c088805",
   418 => x"0851ad3f",
   419 => x"8008708c",
   420 => x"08f8050c",
   421 => x"548c08fc",
   422 => x"0508802e",
   423 => x"8c388c08",
   424 => x"f8050830",
   425 => x"8c08f805",
   426 => x"0c8c08f8",
   427 => x"05087080",
   428 => x"0c54873d",
   429 => x"0d8c0c04",
   430 => x"8c08028c",
   431 => x"0cfd3d0d",
   432 => x"810b8c08",
   433 => x"fc050c80",
   434 => x"0b8c08f8",
   435 => x"050c8c08",
   436 => x"8c05088c",
   437 => x"08880508",
   438 => x"27ac388c",
   439 => x"08fc0508",
   440 => x"802ea338",
   441 => x"800b8c08",
   442 => x"8c050824",
   443 => x"99388c08",
   444 => x"8c050810",
   445 => x"8c088c05",
   446 => x"0c8c08fc",
   447 => x"0508108c",
   448 => x"08fc050c",
   449 => x"c9398c08",
   450 => x"fc050880",
   451 => x"2e80c938",
   452 => x"8c088c05",
   453 => x"088c0888",
   454 => x"050826a1",
   455 => x"388c0888",
   456 => x"05088c08",
   457 => x"8c050831",
   458 => x"8c088805",
   459 => x"0c8c08f8",
   460 => x"05088c08",
   461 => x"fc050807",
   462 => x"8c08f805",
   463 => x"0c8c08fc",
   464 => x"0508812a",
   465 => x"8c08fc05",
   466 => x"0c8c088c",
   467 => x"0508812a",
   468 => x"8c088c05",
   469 => x"0cffaf39",
   470 => x"8c089005",
   471 => x"08802e8f",
   472 => x"388c0888",
   473 => x"0508708c",
   474 => x"08f4050c",
   475 => x"518d398c",
   476 => x"08f80508",
   477 => x"708c08f4",
   478 => x"050c518c",
   479 => x"08f40508",
   480 => x"800c853d",
   481 => x"0d8c0c04",
   482 => x"803d0d86",
   483 => x"5184e73f",
   484 => x"8151bae0",
   485 => x"3ffc3d0d",
   486 => x"7670797b",
   487 => x"55555555",
   488 => x"8f72278c",
   489 => x"38727507",
   490 => x"83065170",
   491 => x"802ea738",
   492 => x"ff125271",
   493 => x"ff2e9838",
   494 => x"72708105",
   495 => x"54337470",
   496 => x"81055634",
   497 => x"ff125271",
   498 => x"ff2e0981",
   499 => x"06ea3874",
   500 => x"800c863d",
   501 => x"0d047451",
   502 => x"72708405",
   503 => x"54087170",
   504 => x"8405530c",
   505 => x"72708405",
   506 => x"54087170",
   507 => x"8405530c",
   508 => x"72708405",
   509 => x"54087170",
   510 => x"8405530c",
   511 => x"72708405",
   512 => x"54087170",
   513 => x"8405530c",
   514 => x"f0125271",
   515 => x"8f26c938",
   516 => x"83722795",
   517 => x"38727084",
   518 => x"05540871",
   519 => x"70840553",
   520 => x"0cfc1252",
   521 => x"718326ed",
   522 => x"387054ff",
   523 => x"8339f73d",
   524 => x"0d7c7052",
   525 => x"5384bd3f",
   526 => x"72548008",
   527 => x"5580d1a8",
   528 => x"56815780",
   529 => x"0881055a",
   530 => x"8b3de411",
   531 => x"59538259",
   532 => x"f413527b",
   533 => x"88110852",
   534 => x"5384f83f",
   535 => x"80083070",
   536 => x"8008079f",
   537 => x"2c8a0780",
   538 => x"0c538b3d",
   539 => x"0d04ff3d",
   540 => x"0d735280",
   541 => x"d1dc0851",
   542 => x"ffb43f83",
   543 => x"3d0d04fd",
   544 => x"3d0d7553",
   545 => x"84d81308",
   546 => x"802e8a38",
   547 => x"80537280",
   548 => x"0c853d0d",
   549 => x"04818052",
   550 => x"72518a9e",
   551 => x"3f800884",
   552 => x"d8140cff",
   553 => x"53800880",
   554 => x"2ee43880",
   555 => x"08549f53",
   556 => x"80747084",
   557 => x"05560cff",
   558 => x"13538073",
   559 => x"24ce3880",
   560 => x"74708405",
   561 => x"560cff13",
   562 => x"53728025",
   563 => x"e338ffbc",
   564 => x"39fd3d0d",
   565 => x"75775553",
   566 => x"9f74278d",
   567 => x"3896730c",
   568 => x"ff527180",
   569 => x"0c853d0d",
   570 => x"0484d813",
   571 => x"08527180",
   572 => x"2e933873",
   573 => x"10101270",
   574 => x"0879720c",
   575 => x"51527180",
   576 => x"0c853d0d",
   577 => x"047251fe",
   578 => x"f63fff52",
   579 => x"8008d338",
   580 => x"84d81308",
   581 => x"74101011",
   582 => x"70087a72",
   583 => x"0c515152",
   584 => x"dd39f93d",
   585 => x"0d797b58",
   586 => x"56769f26",
   587 => x"80e83884",
   588 => x"d8160854",
   589 => x"73802eaa",
   590 => x"38761010",
   591 => x"14700855",
   592 => x"5573802e",
   593 => x"ba388058",
   594 => x"73812e8f",
   595 => x"3873ff2e",
   596 => x"a3388075",
   597 => x"0c765173",
   598 => x"2d805877",
   599 => x"800c893d",
   600 => x"0d047551",
   601 => x"fe993fff",
   602 => x"588008ef",
   603 => x"3884d816",
   604 => x"0854c639",
   605 => x"96760c81",
   606 => x"0b800c89",
   607 => x"3d0d0475",
   608 => x"5181ed3f",
   609 => x"76538008",
   610 => x"52755181",
   611 => x"ad3f8008",
   612 => x"800c893d",
   613 => x"0d049676",
   614 => x"0cff0b80",
   615 => x"0c893d0d",
   616 => x"04fc3d0d",
   617 => x"76785653",
   618 => x"ff54749f",
   619 => x"26b13884",
   620 => x"d8130852",
   621 => x"71802eae",
   622 => x"38741010",
   623 => x"12700853",
   624 => x"53815471",
   625 => x"802e9838",
   626 => x"825471ff",
   627 => x"2e913883",
   628 => x"5471812e",
   629 => x"8a388073",
   630 => x"0c745171",
   631 => x"2d805473",
   632 => x"800c863d",
   633 => x"0d047251",
   634 => x"fd953f80",
   635 => x"08f13884",
   636 => x"d8130852",
   637 => x"c439ff3d",
   638 => x"0d735280",
   639 => x"d1dc0851",
   640 => x"fea03f83",
   641 => x"3d0d04fe",
   642 => x"3d0d7553",
   643 => x"745280d1",
   644 => x"dc0851fd",
   645 => x"bc3f843d",
   646 => x"0d04803d",
   647 => x"0d80d1dc",
   648 => x"0851fcdb",
   649 => x"3f823d0d",
   650 => x"04ff3d0d",
   651 => x"735280d1",
   652 => x"dc0851fe",
   653 => x"ec3f833d",
   654 => x"0d04fc3d",
   655 => x"0d800b80",
   656 => x"e1d00c78",
   657 => x"527751b4",
   658 => x"9d3f8008",
   659 => x"548008ff",
   660 => x"2e883873",
   661 => x"800c863d",
   662 => x"0d0480e1",
   663 => x"d0085574",
   664 => x"802ef038",
   665 => x"7675710c",
   666 => x"5373800c",
   667 => x"863d0d04",
   668 => x"b3ef3f04",
   669 => x"fd3d0d75",
   670 => x"70718306",
   671 => x"53555270",
   672 => x"b8387170",
   673 => x"087009f7",
   674 => x"fbfdff12",
   675 => x"0670f884",
   676 => x"82818006",
   677 => x"51515253",
   678 => x"709d3884",
   679 => x"13700870",
   680 => x"09f7fbfd",
   681 => x"ff120670",
   682 => x"f8848281",
   683 => x"80065151",
   684 => x"52537080",
   685 => x"2ee53872",
   686 => x"52713351",
   687 => x"70802e8a",
   688 => x"38811270",
   689 => x"33525270",
   690 => x"f8387174",
   691 => x"31800c85",
   692 => x"3d0d04f2",
   693 => x"3d0d6062",
   694 => x"88110870",
   695 => x"57575f5a",
   696 => x"74802e81",
   697 => x"90388c1a",
   698 => x"2270832a",
   699 => x"81327081",
   700 => x"06515558",
   701 => x"73863890",
   702 => x"1a089138",
   703 => x"79519ccd",
   704 => x"3fff5480",
   705 => x"0880ee38",
   706 => x"8c1a2258",
   707 => x"7d085780",
   708 => x"7883ffff",
   709 => x"06700a10",
   710 => x"0a708106",
   711 => x"51565755",
   712 => x"73752e80",
   713 => x"d7387490",
   714 => x"38760884",
   715 => x"18088819",
   716 => x"59565974",
   717 => x"802ef238",
   718 => x"74548880",
   719 => x"75278438",
   720 => x"88805473",
   721 => x"5378529c",
   722 => x"1a0851a4",
   723 => x"1a085473",
   724 => x"2d800b80",
   725 => x"082582e6",
   726 => x"38800819",
   727 => x"75800831",
   728 => x"7f880508",
   729 => x"80083170",
   730 => x"6188050c",
   731 => x"56565973",
   732 => x"ffb43880",
   733 => x"5473800c",
   734 => x"903d0d04",
   735 => x"75813270",
   736 => x"81067641",
   737 => x"51547380",
   738 => x"2e81c138",
   739 => x"74903876",
   740 => x"08841808",
   741 => x"88195956",
   742 => x"5974802e",
   743 => x"f238881a",
   744 => x"087883ff",
   745 => x"ff067089",
   746 => x"2a708106",
   747 => x"51565956",
   748 => x"73802e82",
   749 => x"fa387575",
   750 => x"278d3877",
   751 => x"872a7081",
   752 => x"06515473",
   753 => x"82b53874",
   754 => x"76278338",
   755 => x"74567553",
   756 => x"78527908",
   757 => x"5190f83f",
   758 => x"881a0876",
   759 => x"31881b0c",
   760 => x"7908167a",
   761 => x"0c745675",
   762 => x"19757731",
   763 => x"7f880508",
   764 => x"78317061",
   765 => x"88050c56",
   766 => x"56597380",
   767 => x"2efef438",
   768 => x"8c1a2258",
   769 => x"ff863977",
   770 => x"78547953",
   771 => x"7b525690",
   772 => x"be3f881a",
   773 => x"08783188",
   774 => x"1b0c7908",
   775 => x"187a0c7c",
   776 => x"76315d7c",
   777 => x"8e387951",
   778 => x"9c873f80",
   779 => x"08818f38",
   780 => x"80085f75",
   781 => x"19757731",
   782 => x"7f880508",
   783 => x"78317061",
   784 => x"88050c56",
   785 => x"56597380",
   786 => x"2efea838",
   787 => x"74818338",
   788 => x"76088418",
   789 => x"08881959",
   790 => x"56597480",
   791 => x"2ef23874",
   792 => x"538a5278",
   793 => x"518ec93f",
   794 => x"80087931",
   795 => x"81055d80",
   796 => x"08843881",
   797 => x"155d815f",
   798 => x"7c58747d",
   799 => x"27833874",
   800 => x"58941a08",
   801 => x"881b0811",
   802 => x"575c807a",
   803 => x"085c5490",
   804 => x"1a087b27",
   805 => x"83388154",
   806 => x"75782584",
   807 => x"3873ba38",
   808 => x"7b7824fe",
   809 => x"e2387b53",
   810 => x"78529c1a",
   811 => x"0851a41a",
   812 => x"0854732d",
   813 => x"80085680",
   814 => x"088024fe",
   815 => x"e2388c1a",
   816 => x"2280c007",
   817 => x"54738c1b",
   818 => x"23ff5473",
   819 => x"800c903d",
   820 => x"0d047eff",
   821 => x"a338ff87",
   822 => x"39755378",
   823 => x"527a518e",
   824 => x"ee3f7908",
   825 => x"167a0c79",
   826 => x"519ac63f",
   827 => x"8008cf38",
   828 => x"7c76315d",
   829 => x"7cfebc38",
   830 => x"feac3990",
   831 => x"1a087a08",
   832 => x"71317611",
   833 => x"70565a57",
   834 => x"5280d1dc",
   835 => x"08519084",
   836 => x"3f800880",
   837 => x"2effa738",
   838 => x"8008901b",
   839 => x"0c800816",
   840 => x"7a0c7794",
   841 => x"1b0c7488",
   842 => x"1b0c7456",
   843 => x"fd993979",
   844 => x"0858901a",
   845 => x"08782783",
   846 => x"38815475",
   847 => x"75278438",
   848 => x"73b33894",
   849 => x"1a085675",
   850 => x"752680d3",
   851 => x"38755378",
   852 => x"529c1a08",
   853 => x"51a41a08",
   854 => x"54732d80",
   855 => x"08568008",
   856 => x"8024fd83",
   857 => x"388c1a22",
   858 => x"80c00754",
   859 => x"738c1b23",
   860 => x"ff54fed7",
   861 => x"39755378",
   862 => x"5277518d",
   863 => x"d23f7908",
   864 => x"167a0c79",
   865 => x"5199aa3f",
   866 => x"8008802e",
   867 => x"fcd9388c",
   868 => x"1a2280c0",
   869 => x"0754738c",
   870 => x"1b23ff54",
   871 => x"fead3974",
   872 => x"75547953",
   873 => x"7852568d",
   874 => x"a63f881a",
   875 => x"08753188",
   876 => x"1b0c7908",
   877 => x"157a0cfc",
   878 => x"ae39f33d",
   879 => x"0d7f618b",
   880 => x"1170f806",
   881 => x"5c55555e",
   882 => x"72962683",
   883 => x"38905980",
   884 => x"7924747a",
   885 => x"26075380",
   886 => x"5472742e",
   887 => x"09810680",
   888 => x"cb387d51",
   889 => x"8eac3f78",
   890 => x"83f72680",
   891 => x"c6387883",
   892 => x"2a701010",
   893 => x"1080d998",
   894 => x"058c1108",
   895 => x"59595a76",
   896 => x"782e83b0",
   897 => x"38841708",
   898 => x"fc06568c",
   899 => x"17088818",
   900 => x"08718c12",
   901 => x"0c88120c",
   902 => x"58751784",
   903 => x"11088107",
   904 => x"84120c53",
   905 => x"7d518deb",
   906 => x"3f881754",
   907 => x"73800c8f",
   908 => x"3d0d0478",
   909 => x"892a7983",
   910 => x"2a5b5372",
   911 => x"802ebf38",
   912 => x"78862ab8",
   913 => x"055a8473",
   914 => x"27b43880",
   915 => x"db135a94",
   916 => x"7327ab38",
   917 => x"788c2a80",
   918 => x"ee055a80",
   919 => x"d473279e",
   920 => x"38788f2a",
   921 => x"80f7055a",
   922 => x"82d47327",
   923 => x"91387892",
   924 => x"2a80fc05",
   925 => x"5a8ad473",
   926 => x"27843880",
   927 => x"fe5a7910",
   928 => x"101080d9",
   929 => x"98058c11",
   930 => x"08585576",
   931 => x"752ea338",
   932 => x"841708fc",
   933 => x"06707a31",
   934 => x"5556738f",
   935 => x"2488d538",
   936 => x"738025fe",
   937 => x"e6388c17",
   938 => x"08577675",
   939 => x"2e098106",
   940 => x"df38811a",
   941 => x"5a80d9a8",
   942 => x"08577680",
   943 => x"d9a02e82",
   944 => x"c0388417",
   945 => x"08fc0670",
   946 => x"7a315556",
   947 => x"738f2481",
   948 => x"f93880d9",
   949 => x"a00b80d9",
   950 => x"ac0c80d9",
   951 => x"a00b80d9",
   952 => x"a80c7380",
   953 => x"25feb238",
   954 => x"83ff7627",
   955 => x"83df3875",
   956 => x"892a7683",
   957 => x"2a555372",
   958 => x"802ebf38",
   959 => x"75862ab8",
   960 => x"05548473",
   961 => x"27b43880",
   962 => x"db135494",
   963 => x"7327ab38",
   964 => x"758c2a80",
   965 => x"ee055480",
   966 => x"d473279e",
   967 => x"38758f2a",
   968 => x"80f70554",
   969 => x"82d47327",
   970 => x"91387592",
   971 => x"2a80fc05",
   972 => x"548ad473",
   973 => x"27843880",
   974 => x"fe547310",
   975 => x"101080d9",
   976 => x"98058811",
   977 => x"08565874",
   978 => x"782e86cf",
   979 => x"38841508",
   980 => x"fc065375",
   981 => x"73278d38",
   982 => x"88150855",
   983 => x"74782e09",
   984 => x"8106ea38",
   985 => x"8c150880",
   986 => x"d9980b84",
   987 => x"0508718c",
   988 => x"1a0c7688",
   989 => x"1a0c7888",
   990 => x"130c788c",
   991 => x"180c5d58",
   992 => x"7953807a",
   993 => x"2483e638",
   994 => x"72822c81",
   995 => x"712b5c53",
   996 => x"7a7c2681",
   997 => x"98387b7b",
   998 => x"06537282",
   999 => x"f13879fc",
  1000 => x"0684055a",
  1001 => x"7a10707d",
  1002 => x"06545b72",
  1003 => x"82e03884",
  1004 => x"1a5af139",
  1005 => x"88178c11",
  1006 => x"08585876",
  1007 => x"782e0981",
  1008 => x"06fcc238",
  1009 => x"821a5afd",
  1010 => x"ec397817",
  1011 => x"79810784",
  1012 => x"190c7080",
  1013 => x"d9ac0c70",
  1014 => x"80d9a80c",
  1015 => x"80d9a00b",
  1016 => x"8c120c8c",
  1017 => x"11088812",
  1018 => x"0c748107",
  1019 => x"84120c74",
  1020 => x"1175710c",
  1021 => x"51537d51",
  1022 => x"8a993f88",
  1023 => x"1754fcac",
  1024 => x"3980d998",
  1025 => x"0b840508",
  1026 => x"7a545c79",
  1027 => x"8025fef8",
  1028 => x"3882da39",
  1029 => x"7a097c06",
  1030 => x"7080d998",
  1031 => x"0b84050c",
  1032 => x"5c7a105b",
  1033 => x"7a7c2685",
  1034 => x"387a85b8",
  1035 => x"3880d998",
  1036 => x"0b880508",
  1037 => x"70841208",
  1038 => x"fc06707c",
  1039 => x"317c7226",
  1040 => x"8f722507",
  1041 => x"57575c5d",
  1042 => x"5572802e",
  1043 => x"80db3879",
  1044 => x"7a1680d9",
  1045 => x"90081b90",
  1046 => x"115a5557",
  1047 => x"5b80d98c",
  1048 => x"08ff2e88",
  1049 => x"38a08f13",
  1050 => x"e0800657",
  1051 => x"76527d51",
  1052 => x"91a73f80",
  1053 => x"08548008",
  1054 => x"ff2e9038",
  1055 => x"80087627",
  1056 => x"82993874",
  1057 => x"80d9982e",
  1058 => x"82913880",
  1059 => x"d9980b88",
  1060 => x"05085584",
  1061 => x"1508fc06",
  1062 => x"707a317a",
  1063 => x"72268f72",
  1064 => x"25075255",
  1065 => x"537283e6",
  1066 => x"38747981",
  1067 => x"0784170c",
  1068 => x"79167080",
  1069 => x"d9980b88",
  1070 => x"050c7581",
  1071 => x"0784120c",
  1072 => x"547e5257",
  1073 => x"88cd3f88",
  1074 => x"1754fae0",
  1075 => x"3975832a",
  1076 => x"70545480",
  1077 => x"7424819b",
  1078 => x"3872822c",
  1079 => x"81712b80",
  1080 => x"d99c0807",
  1081 => x"7080d998",
  1082 => x"0b84050c",
  1083 => x"75101010",
  1084 => x"80d99805",
  1085 => x"88110858",
  1086 => x"5a5d5377",
  1087 => x"8c180c74",
  1088 => x"88180c76",
  1089 => x"88190c76",
  1090 => x"8c160cfc",
  1091 => x"f339797a",
  1092 => x"10101080",
  1093 => x"d9980570",
  1094 => x"57595d8c",
  1095 => x"15085776",
  1096 => x"752ea338",
  1097 => x"841708fc",
  1098 => x"06707a31",
  1099 => x"5556738f",
  1100 => x"2483ca38",
  1101 => x"73802584",
  1102 => x"81388c17",
  1103 => x"08577675",
  1104 => x"2e098106",
  1105 => x"df388815",
  1106 => x"811b7083",
  1107 => x"06555b55",
  1108 => x"72c9387c",
  1109 => x"83065372",
  1110 => x"802efdb8",
  1111 => x"38ff1df8",
  1112 => x"19595d88",
  1113 => x"1808782e",
  1114 => x"ea38fdb5",
  1115 => x"39831a53",
  1116 => x"fc963983",
  1117 => x"1470822c",
  1118 => x"81712b80",
  1119 => x"d99c0807",
  1120 => x"7080d998",
  1121 => x"0b84050c",
  1122 => x"76101010",
  1123 => x"80d99805",
  1124 => x"88110859",
  1125 => x"5b5e5153",
  1126 => x"fee13980",
  1127 => x"d8dc0817",
  1128 => x"58800876",
  1129 => x"2e818d38",
  1130 => x"80d98c08",
  1131 => x"ff2e83ec",
  1132 => x"38737631",
  1133 => x"1880d8dc",
  1134 => x"0c738706",
  1135 => x"70575372",
  1136 => x"802e8838",
  1137 => x"88733170",
  1138 => x"15555676",
  1139 => x"149fff06",
  1140 => x"a0807131",
  1141 => x"1770547f",
  1142 => x"5357538e",
  1143 => x"bc3f8008",
  1144 => x"538008ff",
  1145 => x"2e81a038",
  1146 => x"80d8dc08",
  1147 => x"167080d8",
  1148 => x"dc0c7475",
  1149 => x"80d9980b",
  1150 => x"88050c74",
  1151 => x"76311870",
  1152 => x"81075155",
  1153 => x"56587b80",
  1154 => x"d9982e83",
  1155 => x"9c38798f",
  1156 => x"2682cb38",
  1157 => x"810b8415",
  1158 => x"0c841508",
  1159 => x"fc06707a",
  1160 => x"317a7226",
  1161 => x"8f722507",
  1162 => x"52555372",
  1163 => x"802efcf9",
  1164 => x"3880db39",
  1165 => x"80089fff",
  1166 => x"065372fe",
  1167 => x"eb387780",
  1168 => x"d8dc0c80",
  1169 => x"d9980b88",
  1170 => x"05087b18",
  1171 => x"81078412",
  1172 => x"0c5580d9",
  1173 => x"88087827",
  1174 => x"86387780",
  1175 => x"d9880c80",
  1176 => x"d9840878",
  1177 => x"27fcac38",
  1178 => x"7780d984",
  1179 => x"0c841508",
  1180 => x"fc06707a",
  1181 => x"317a7226",
  1182 => x"8f722507",
  1183 => x"52555372",
  1184 => x"802efca5",
  1185 => x"38883980",
  1186 => x"745456fe",
  1187 => x"db397d51",
  1188 => x"85813f80",
  1189 => x"0b800c8f",
  1190 => x"3d0d0473",
  1191 => x"53807424",
  1192 => x"a9387282",
  1193 => x"2c81712b",
  1194 => x"80d99c08",
  1195 => x"077080d9",
  1196 => x"980b8405",
  1197 => x"0c5d5377",
  1198 => x"8c180c74",
  1199 => x"88180c76",
  1200 => x"88190c76",
  1201 => x"8c160cf9",
  1202 => x"b7398314",
  1203 => x"70822c81",
  1204 => x"712b80d9",
  1205 => x"9c080770",
  1206 => x"80d9980b",
  1207 => x"84050c5e",
  1208 => x"5153d439",
  1209 => x"7b7b0653",
  1210 => x"72fca338",
  1211 => x"841a7b10",
  1212 => x"5c5af139",
  1213 => x"ff1a8111",
  1214 => x"515af7b9",
  1215 => x"39781779",
  1216 => x"81078419",
  1217 => x"0c8c1808",
  1218 => x"88190871",
  1219 => x"8c120c88",
  1220 => x"120c5970",
  1221 => x"80d9ac0c",
  1222 => x"7080d9a8",
  1223 => x"0c80d9a0",
  1224 => x"0b8c120c",
  1225 => x"8c110888",
  1226 => x"120c7481",
  1227 => x"0784120c",
  1228 => x"74117571",
  1229 => x"0c5153f9",
  1230 => x"bd397517",
  1231 => x"84110881",
  1232 => x"0784120c",
  1233 => x"538c1708",
  1234 => x"88180871",
  1235 => x"8c120c88",
  1236 => x"120c587d",
  1237 => x"5183bc3f",
  1238 => x"881754f5",
  1239 => x"cf397284",
  1240 => x"150cf41a",
  1241 => x"f8067084",
  1242 => x"1e088106",
  1243 => x"07841e0c",
  1244 => x"701d545b",
  1245 => x"850b8414",
  1246 => x"0c850b88",
  1247 => x"140c8f7b",
  1248 => x"27fdcf38",
  1249 => x"881c527d",
  1250 => x"5193ee3f",
  1251 => x"80d9980b",
  1252 => x"88050880",
  1253 => x"d8dc0859",
  1254 => x"55fdb739",
  1255 => x"7780d8dc",
  1256 => x"0c7380d9",
  1257 => x"8c0cfc91",
  1258 => x"39728415",
  1259 => x"0cfda339",
  1260 => x"fa3d0d7a",
  1261 => x"79028805",
  1262 => x"a7053356",
  1263 => x"52538373",
  1264 => x"278a3870",
  1265 => x"83065271",
  1266 => x"802ea838",
  1267 => x"ff135372",
  1268 => x"ff2e9738",
  1269 => x"70335273",
  1270 => x"722e9138",
  1271 => x"8111ff14",
  1272 => x"545172ff",
  1273 => x"2e098106",
  1274 => x"eb388051",
  1275 => x"70800c88",
  1276 => x"3d0d0470",
  1277 => x"72575583",
  1278 => x"51758280",
  1279 => x"2914ff12",
  1280 => x"52567080",
  1281 => x"25f33883",
  1282 => x"7327bf38",
  1283 => x"74087632",
  1284 => x"7009f7fb",
  1285 => x"fdff1206",
  1286 => x"70f88482",
  1287 => x"81800651",
  1288 => x"51517080",
  1289 => x"2e993874",
  1290 => x"51805270",
  1291 => x"33577377",
  1292 => x"2effb938",
  1293 => x"81118113",
  1294 => x"53518372",
  1295 => x"27ed38fc",
  1296 => x"13841656",
  1297 => x"53728326",
  1298 => x"c3387451",
  1299 => x"fefe39fa",
  1300 => x"3d0d787a",
  1301 => x"7c727272",
  1302 => x"57575759",
  1303 => x"56567476",
  1304 => x"27b23876",
  1305 => x"15517571",
  1306 => x"27aa3870",
  1307 => x"7717ff14",
  1308 => x"54555371",
  1309 => x"ff2e9638",
  1310 => x"ff14ff14",
  1311 => x"54547233",
  1312 => x"7434ff12",
  1313 => x"5271ff2e",
  1314 => x"098106ec",
  1315 => x"3875800c",
  1316 => x"883d0d04",
  1317 => x"768f2697",
  1318 => x"38ff1252",
  1319 => x"71ff2eed",
  1320 => x"38727081",
  1321 => x"05543374",
  1322 => x"70810556",
  1323 => x"34eb3974",
  1324 => x"76078306",
  1325 => x"5170e238",
  1326 => x"75755451",
  1327 => x"72708405",
  1328 => x"54087170",
  1329 => x"8405530c",
  1330 => x"72708405",
  1331 => x"54087170",
  1332 => x"8405530c",
  1333 => x"72708405",
  1334 => x"54087170",
  1335 => x"8405530c",
  1336 => x"72708405",
  1337 => x"54087170",
  1338 => x"8405530c",
  1339 => x"f0125271",
  1340 => x"8f26c938",
  1341 => x"83722795",
  1342 => x"38727084",
  1343 => x"05540871",
  1344 => x"70840553",
  1345 => x"0cfc1252",
  1346 => x"718326ed",
  1347 => x"387054ff",
  1348 => x"88390404",
  1349 => x"ef3d0d63",
  1350 => x"6567405d",
  1351 => x"427b802e",
  1352 => x"84f93861",
  1353 => x"51ec3ff8",
  1354 => x"1c708412",
  1355 => x"0870fc06",
  1356 => x"70628b05",
  1357 => x"70f80641",
  1358 => x"59455b5c",
  1359 => x"41579674",
  1360 => x"2782c338",
  1361 => x"807b247e",
  1362 => x"7c260759",
  1363 => x"80547874",
  1364 => x"2e098106",
  1365 => x"82a93877",
  1366 => x"7b2581fc",
  1367 => x"38771780",
  1368 => x"d9980b88",
  1369 => x"05085e56",
  1370 => x"7c762e84",
  1371 => x"bd388416",
  1372 => x"0870fe06",
  1373 => x"17841108",
  1374 => x"81065155",
  1375 => x"5573828b",
  1376 => x"3874fc06",
  1377 => x"597c762e",
  1378 => x"84dd3877",
  1379 => x"195f7e7b",
  1380 => x"2581fd38",
  1381 => x"79810654",
  1382 => x"7382bf38",
  1383 => x"76770831",
  1384 => x"841108fc",
  1385 => x"06565a75",
  1386 => x"802e9138",
  1387 => x"7c762e84",
  1388 => x"ea387419",
  1389 => x"1859787b",
  1390 => x"25848938",
  1391 => x"79802e82",
  1392 => x"99387715",
  1393 => x"567a7624",
  1394 => x"8290388c",
  1395 => x"1a08881b",
  1396 => x"08718c12",
  1397 => x"0c88120c",
  1398 => x"55797659",
  1399 => x"57881761",
  1400 => x"fc055759",
  1401 => x"75a42685",
  1402 => x"ef387b79",
  1403 => x"55559376",
  1404 => x"2780c938",
  1405 => x"7b708405",
  1406 => x"5d087c56",
  1407 => x"790c7470",
  1408 => x"84055608",
  1409 => x"8c180c90",
  1410 => x"17549b76",
  1411 => x"27ae3874",
  1412 => x"70840556",
  1413 => x"08740c74",
  1414 => x"70840556",
  1415 => x"0894180c",
  1416 => x"981754a3",
  1417 => x"76279538",
  1418 => x"74708405",
  1419 => x"5608740c",
  1420 => x"74708405",
  1421 => x"56089c18",
  1422 => x"0ca01754",
  1423 => x"74708405",
  1424 => x"56087470",
  1425 => x"8405560c",
  1426 => x"74708405",
  1427 => x"56087470",
  1428 => x"8405560c",
  1429 => x"7408740c",
  1430 => x"777b3156",
  1431 => x"758f2680",
  1432 => x"c9388417",
  1433 => x"08810678",
  1434 => x"0784180c",
  1435 => x"77178411",
  1436 => x"08810784",
  1437 => x"120c5461",
  1438 => x"51fd983f",
  1439 => x"88175473",
  1440 => x"800c933d",
  1441 => x"0d04905b",
  1442 => x"fdba3978",
  1443 => x"56fe8539",
  1444 => x"8c160888",
  1445 => x"1708718c",
  1446 => x"120c8812",
  1447 => x"0c557e70",
  1448 => x"7c315758",
  1449 => x"8f7627ff",
  1450 => x"b9387a17",
  1451 => x"84180881",
  1452 => x"067c0784",
  1453 => x"190c7681",
  1454 => x"0784120c",
  1455 => x"76118411",
  1456 => x"08810784",
  1457 => x"120c5588",
  1458 => x"05526151",
  1459 => x"8dab3f61",
  1460 => x"51fcc03f",
  1461 => x"881754ff",
  1462 => x"a6397d52",
  1463 => x"6151edda",
  1464 => x"3f800859",
  1465 => x"8008802e",
  1466 => x"81a33880",
  1467 => x"08f80560",
  1468 => x"840508fe",
  1469 => x"06610555",
  1470 => x"5776742e",
  1471 => x"83e638fc",
  1472 => x"185675a4",
  1473 => x"2681aa38",
  1474 => x"7b800855",
  1475 => x"55937627",
  1476 => x"80d83874",
  1477 => x"70840556",
  1478 => x"08800870",
  1479 => x"8405800c",
  1480 => x"0c800875",
  1481 => x"70840557",
  1482 => x"08717084",
  1483 => x"05530c54",
  1484 => x"9b7627b6",
  1485 => x"38747084",
  1486 => x"05560874",
  1487 => x"70840556",
  1488 => x"0c747084",
  1489 => x"05560874",
  1490 => x"70840556",
  1491 => x"0ca37627",
  1492 => x"99387470",
  1493 => x"84055608",
  1494 => x"74708405",
  1495 => x"560c7470",
  1496 => x"84055608",
  1497 => x"74708405",
  1498 => x"560c7470",
  1499 => x"84055608",
  1500 => x"74708405",
  1501 => x"560c7470",
  1502 => x"84055608",
  1503 => x"74708405",
  1504 => x"560c7408",
  1505 => x"740c7b52",
  1506 => x"61518bed",
  1507 => x"3f6151fb",
  1508 => x"823f7854",
  1509 => x"73800c93",
  1510 => x"3d0d047d",
  1511 => x"526151ec",
  1512 => x"993f8008",
  1513 => x"800c933d",
  1514 => x"0d048416",
  1515 => x"0855fbd1",
  1516 => x"3975537b",
  1517 => x"52800851",
  1518 => x"dfdb3f7b",
  1519 => x"5261518b",
  1520 => x"b83fca39",
  1521 => x"8c160888",
  1522 => x"1708718c",
  1523 => x"120c8812",
  1524 => x"0c558c1a",
  1525 => x"08881b08",
  1526 => x"718c120c",
  1527 => x"88120c55",
  1528 => x"79795957",
  1529 => x"fbf73977",
  1530 => x"19901c55",
  1531 => x"55737524",
  1532 => x"fba2387a",
  1533 => x"177080d9",
  1534 => x"980b8805",
  1535 => x"0c757c31",
  1536 => x"81078412",
  1537 => x"0c5d8417",
  1538 => x"0881067b",
  1539 => x"0784180c",
  1540 => x"6151f9ff",
  1541 => x"3f881754",
  1542 => x"fce53974",
  1543 => x"1918901c",
  1544 => x"555d737d",
  1545 => x"24fb9538",
  1546 => x"8c1a0888",
  1547 => x"1b08718c",
  1548 => x"120c8812",
  1549 => x"0c55881a",
  1550 => x"61fc0557",
  1551 => x"5975a426",
  1552 => x"81ae387b",
  1553 => x"79555593",
  1554 => x"762780c9",
  1555 => x"387b7084",
  1556 => x"055d087c",
  1557 => x"56790c74",
  1558 => x"70840556",
  1559 => x"088c1b0c",
  1560 => x"901a549b",
  1561 => x"7627ae38",
  1562 => x"74708405",
  1563 => x"5608740c",
  1564 => x"74708405",
  1565 => x"5608941b",
  1566 => x"0c981a54",
  1567 => x"a3762795",
  1568 => x"38747084",
  1569 => x"05560874",
  1570 => x"0c747084",
  1571 => x"0556089c",
  1572 => x"1b0ca01a",
  1573 => x"54747084",
  1574 => x"05560874",
  1575 => x"70840556",
  1576 => x"0c747084",
  1577 => x"05560874",
  1578 => x"70840556",
  1579 => x"0c740874",
  1580 => x"0c7a1a70",
  1581 => x"80d9980b",
  1582 => x"88050c7d",
  1583 => x"7c318107",
  1584 => x"84120c54",
  1585 => x"841a0881",
  1586 => x"067b0784",
  1587 => x"1b0c6151",
  1588 => x"f8c13f78",
  1589 => x"54fdbd39",
  1590 => x"75537b52",
  1591 => x"7851ddb5",
  1592 => x"3ffaf539",
  1593 => x"841708fc",
  1594 => x"06186058",
  1595 => x"58fae939",
  1596 => x"75537b52",
  1597 => x"7851dd9d",
  1598 => x"3f7a1a70",
  1599 => x"80d9980b",
  1600 => x"88050c7d",
  1601 => x"7c318107",
  1602 => x"84120c54",
  1603 => x"841a0881",
  1604 => x"067b0784",
  1605 => x"1b0cffb6",
  1606 => x"39fd3d0d",
  1607 => x"800b80e1",
  1608 => x"d00c7651",
  1609 => x"96d53f80",
  1610 => x"08538008",
  1611 => x"ff2e8838",
  1612 => x"72800c85",
  1613 => x"3d0d0480",
  1614 => x"e1d00854",
  1615 => x"73802ef0",
  1616 => x"38757471",
  1617 => x"0c527280",
  1618 => x"0c853d0d",
  1619 => x"04fa3d0d",
  1620 => x"7880d1dc",
  1621 => x"085455b8",
  1622 => x"1308802e",
  1623 => x"81b6388c",
  1624 => x"15227083",
  1625 => x"ffff0670",
  1626 => x"832a8132",
  1627 => x"70810651",
  1628 => x"55555672",
  1629 => x"802e80dc",
  1630 => x"3873842a",
  1631 => x"81328106",
  1632 => x"57ff5376",
  1633 => x"80f73873",
  1634 => x"822a7081",
  1635 => x"06515372",
  1636 => x"802eb938",
  1637 => x"b0150854",
  1638 => x"73802e9c",
  1639 => x"3880c015",
  1640 => x"5373732e",
  1641 => x"8f387352",
  1642 => x"80d1dc08",
  1643 => x"5187ca3f",
  1644 => x"8c152256",
  1645 => x"76b0160c",
  1646 => x"75db0653",
  1647 => x"728c1623",
  1648 => x"800b8416",
  1649 => x"0c901508",
  1650 => x"750c7256",
  1651 => x"75880753",
  1652 => x"728c1623",
  1653 => x"90150880",
  1654 => x"2e80c138",
  1655 => x"8c152270",
  1656 => x"81065553",
  1657 => x"739e3872",
  1658 => x"0a100a70",
  1659 => x"81065153",
  1660 => x"72853894",
  1661 => x"15085473",
  1662 => x"88160c80",
  1663 => x"5372800c",
  1664 => x"883d0d04",
  1665 => x"800b8816",
  1666 => x"0c941508",
  1667 => x"3098160c",
  1668 => x"8053ea39",
  1669 => x"725182fb",
  1670 => x"3ffec439",
  1671 => x"74518ce8",
  1672 => x"3f8c1522",
  1673 => x"70810655",
  1674 => x"5373802e",
  1675 => x"ffb938d4",
  1676 => x"39f83d0d",
  1677 => x"7a587780",
  1678 => x"2e819938",
  1679 => x"80d1dc08",
  1680 => x"54b81408",
  1681 => x"802e80ed",
  1682 => x"388c1822",
  1683 => x"70902b70",
  1684 => x"902c7083",
  1685 => x"2a813281",
  1686 => x"065c5157",
  1687 => x"547880cd",
  1688 => x"38901808",
  1689 => x"5776802e",
  1690 => x"80c33877",
  1691 => x"08773177",
  1692 => x"790c7683",
  1693 => x"067a5855",
  1694 => x"55738538",
  1695 => x"94180856",
  1696 => x"7588190c",
  1697 => x"807525a5",
  1698 => x"38745376",
  1699 => x"529c1808",
  1700 => x"51a41808",
  1701 => x"54732d80",
  1702 => x"0b800825",
  1703 => x"80c93880",
  1704 => x"08177580",
  1705 => x"08315657",
  1706 => x"748024dd",
  1707 => x"38800b80",
  1708 => x"0c8a3d0d",
  1709 => x"04735181",
  1710 => x"da3f8c18",
  1711 => x"2270902b",
  1712 => x"70902c70",
  1713 => x"832a8132",
  1714 => x"81065c51",
  1715 => x"575478dd",
  1716 => x"38ff8e39",
  1717 => x"b4b15280",
  1718 => x"d1dc0851",
  1719 => x"89f13f80",
  1720 => x"08800c8a",
  1721 => x"3d0d048c",
  1722 => x"182280c0",
  1723 => x"0754738c",
  1724 => x"1923ff0b",
  1725 => x"800c8a3d",
  1726 => x"0d04803d",
  1727 => x"0d725180",
  1728 => x"710c800b",
  1729 => x"84120c80",
  1730 => x"0b88120c",
  1731 => x"028e0522",
  1732 => x"8c122302",
  1733 => x"9205228e",
  1734 => x"1223800b",
  1735 => x"90120c80",
  1736 => x"0b94120c",
  1737 => x"800b9812",
  1738 => x"0c709c12",
  1739 => x"0c80c49a",
  1740 => x"0ba0120c",
  1741 => x"80c4e60b",
  1742 => x"a4120c80",
  1743 => x"c5e20ba8",
  1744 => x"120c80c6",
  1745 => x"b30bac12",
  1746 => x"0c823d0d",
  1747 => x"04fa3d0d",
  1748 => x"797080dc",
  1749 => x"298c1154",
  1750 => x"7a535657",
  1751 => x"e4dc3f80",
  1752 => x"08800855",
  1753 => x"56800880",
  1754 => x"2ea23880",
  1755 => x"088c0554",
  1756 => x"800b8008",
  1757 => x"0c768008",
  1758 => x"84050c73",
  1759 => x"80088805",
  1760 => x"0c745380",
  1761 => x"5273518c",
  1762 => x"823f7554",
  1763 => x"73800c88",
  1764 => x"3d0d04fc",
  1765 => x"3d0d76b9",
  1766 => x"a60bbc12",
  1767 => x"0c55810b",
  1768 => x"b8160c80",
  1769 => x"0b84dc16",
  1770 => x"0c830b84",
  1771 => x"e0160c84",
  1772 => x"e81584e4",
  1773 => x"160c7454",
  1774 => x"80538452",
  1775 => x"84150851",
  1776 => x"feb83f74",
  1777 => x"54815389",
  1778 => x"52881508",
  1779 => x"51feab3f",
  1780 => x"74548253",
  1781 => x"8a528c15",
  1782 => x"0851fe9e",
  1783 => x"3f863d0d",
  1784 => x"04f93d0d",
  1785 => x"7980d1dc",
  1786 => x"085457b8",
  1787 => x"1308802e",
  1788 => x"80c83884",
  1789 => x"dc135688",
  1790 => x"16088417",
  1791 => x"08ff0555",
  1792 => x"55807424",
  1793 => x"9f388c15",
  1794 => x"2270902b",
  1795 => x"70902c51",
  1796 => x"54587280",
  1797 => x"2e80ca38",
  1798 => x"80dc15ff",
  1799 => x"15555573",
  1800 => x"8025e338",
  1801 => x"75085372",
  1802 => x"802e9f38",
  1803 => x"72568816",
  1804 => x"08841708",
  1805 => x"ff055555",
  1806 => x"c8397251",
  1807 => x"fed53f80",
  1808 => x"d1dc0884",
  1809 => x"dc0556ff",
  1810 => x"ae398452",
  1811 => x"7651fdfd",
  1812 => x"3f800876",
  1813 => x"0c800880",
  1814 => x"2e80c038",
  1815 => x"800856ce",
  1816 => x"39810b8c",
  1817 => x"16237275",
  1818 => x"0c728816",
  1819 => x"0c728416",
  1820 => x"0c729016",
  1821 => x"0c729416",
  1822 => x"0c729816",
  1823 => x"0cff0b8e",
  1824 => x"162372b0",
  1825 => x"160c72b4",
  1826 => x"160c7280",
  1827 => x"c4160c72",
  1828 => x"80c8160c",
  1829 => x"74800c89",
  1830 => x"3d0d048c",
  1831 => x"770c800b",
  1832 => x"800c893d",
  1833 => x"0d04ff3d",
  1834 => x"0db4b152",
  1835 => x"7351869f",
  1836 => x"3f833d0d",
  1837 => x"04803d0d",
  1838 => x"80d1dc08",
  1839 => x"51e83f82",
  1840 => x"3d0d04fb",
  1841 => x"3d0d7770",
  1842 => x"5256f0c6",
  1843 => x"3f80d998",
  1844 => x"0b880508",
  1845 => x"841108fc",
  1846 => x"06707b31",
  1847 => x"9fef05e0",
  1848 => x"8006e080",
  1849 => x"05565653",
  1850 => x"a0807424",
  1851 => x"94388052",
  1852 => x"7551f8a5",
  1853 => x"3f80d9a0",
  1854 => x"08155372",
  1855 => x"80082e8f",
  1856 => x"387551f0",
  1857 => x"8e3f8053",
  1858 => x"72800c87",
  1859 => x"3d0d0473",
  1860 => x"30527551",
  1861 => x"f8833f80",
  1862 => x"08ff2ea8",
  1863 => x"3880d998",
  1864 => x"0b880508",
  1865 => x"75753181",
  1866 => x"0784120c",
  1867 => x"5380d8dc",
  1868 => x"08743180",
  1869 => x"d8dc0c75",
  1870 => x"51efd83f",
  1871 => x"810b800c",
  1872 => x"873d0d04",
  1873 => x"80527551",
  1874 => x"f7cf3f80",
  1875 => x"d9980b88",
  1876 => x"05088008",
  1877 => x"71315653",
  1878 => x"8f7525ff",
  1879 => x"a4388008",
  1880 => x"80d98c08",
  1881 => x"3180d8dc",
  1882 => x"0c748107",
  1883 => x"84140c75",
  1884 => x"51efa03f",
  1885 => x"8053ff90",
  1886 => x"39f63d0d",
  1887 => x"7c7e545b",
  1888 => x"72802e82",
  1889 => x"83387a51",
  1890 => x"ef883ff8",
  1891 => x"13841108",
  1892 => x"70fe0670",
  1893 => x"13841108",
  1894 => x"fc065d58",
  1895 => x"59545880",
  1896 => x"d9a00875",
  1897 => x"2e82de38",
  1898 => x"7884160c",
  1899 => x"80738106",
  1900 => x"545a727a",
  1901 => x"2e81d538",
  1902 => x"78158411",
  1903 => x"08810651",
  1904 => x"5372a038",
  1905 => x"78175779",
  1906 => x"81e63888",
  1907 => x"15085372",
  1908 => x"80d9a02e",
  1909 => x"82f9388c",
  1910 => x"1508708c",
  1911 => x"150c7388",
  1912 => x"120c5676",
  1913 => x"81078419",
  1914 => x"0c761877",
  1915 => x"710c5379",
  1916 => x"81913883",
  1917 => x"ff772781",
  1918 => x"c8387689",
  1919 => x"2a77832a",
  1920 => x"56537280",
  1921 => x"2ebf3876",
  1922 => x"862ab805",
  1923 => x"55847327",
  1924 => x"b43880db",
  1925 => x"13559473",
  1926 => x"27ab3876",
  1927 => x"8c2a80ee",
  1928 => x"055580d4",
  1929 => x"73279e38",
  1930 => x"768f2a80",
  1931 => x"f7055582",
  1932 => x"d4732791",
  1933 => x"3876922a",
  1934 => x"80fc0555",
  1935 => x"8ad47327",
  1936 => x"843880fe",
  1937 => x"55741010",
  1938 => x"1080d998",
  1939 => x"05881108",
  1940 => x"55567376",
  1941 => x"2e82b338",
  1942 => x"841408fc",
  1943 => x"06537673",
  1944 => x"278d3888",
  1945 => x"14085473",
  1946 => x"762e0981",
  1947 => x"06ea388c",
  1948 => x"1408708c",
  1949 => x"1a0c7488",
  1950 => x"1a0c7888",
  1951 => x"120c5677",
  1952 => x"8c150c7a",
  1953 => x"51ed8c3f",
  1954 => x"8c3d0d04",
  1955 => x"77087871",
  1956 => x"31597705",
  1957 => x"88190854",
  1958 => x"577280d9",
  1959 => x"a02e80e0",
  1960 => x"388c1808",
  1961 => x"708c150c",
  1962 => x"7388120c",
  1963 => x"56fe8939",
  1964 => x"8815088c",
  1965 => x"1608708c",
  1966 => x"130c5788",
  1967 => x"170cfea3",
  1968 => x"3976832a",
  1969 => x"70545580",
  1970 => x"75248198",
  1971 => x"3872822c",
  1972 => x"81712b80",
  1973 => x"d99c0807",
  1974 => x"80d9980b",
  1975 => x"84050c53",
  1976 => x"74101010",
  1977 => x"80d99805",
  1978 => x"88110855",
  1979 => x"56758c19",
  1980 => x"0c738819",
  1981 => x"0c778817",
  1982 => x"0c778c15",
  1983 => x"0cff8439",
  1984 => x"815afdb4",
  1985 => x"39781773",
  1986 => x"81065457",
  1987 => x"72983877",
  1988 => x"08787131",
  1989 => x"5977058c",
  1990 => x"1908881a",
  1991 => x"08718c12",
  1992 => x"0c88120c",
  1993 => x"57577681",
  1994 => x"0784190c",
  1995 => x"7780d998",
  1996 => x"0b88050c",
  1997 => x"80d99408",
  1998 => x"7726fec7",
  1999 => x"3880d990",
  2000 => x"08527a51",
  2001 => x"fafd3f7a",
  2002 => x"51ebc83f",
  2003 => x"feba3981",
  2004 => x"788c150c",
  2005 => x"7888150c",
  2006 => x"738c1a0c",
  2007 => x"73881a0c",
  2008 => x"5afd8039",
  2009 => x"83157082",
  2010 => x"2c81712b",
  2011 => x"80d99c08",
  2012 => x"0780d998",
  2013 => x"0b84050c",
  2014 => x"51537410",
  2015 => x"101080d9",
  2016 => x"98058811",
  2017 => x"085556fe",
  2018 => x"e4397453",
  2019 => x"807524a7",
  2020 => x"3872822c",
  2021 => x"81712b80",
  2022 => x"d99c0807",
  2023 => x"80d9980b",
  2024 => x"84050c53",
  2025 => x"758c190c",
  2026 => x"7388190c",
  2027 => x"7788170c",
  2028 => x"778c150c",
  2029 => x"fdcd3983",
  2030 => x"1570822c",
  2031 => x"81712b80",
  2032 => x"d99c0807",
  2033 => x"80d9980b",
  2034 => x"84050c51",
  2035 => x"53d639f9",
  2036 => x"3d0d797b",
  2037 => x"5853800b",
  2038 => x"80d1dc08",
  2039 => x"53567272",
  2040 => x"2e80c038",
  2041 => x"84dc1355",
  2042 => x"74762eb7",
  2043 => x"38881508",
  2044 => x"841608ff",
  2045 => x"05545480",
  2046 => x"73249d38",
  2047 => x"8c142270",
  2048 => x"902b7090",
  2049 => x"2c515358",
  2050 => x"7180d838",
  2051 => x"80dc14ff",
  2052 => x"14545472",
  2053 => x"8025e538",
  2054 => x"74085574",
  2055 => x"d03880d1",
  2056 => x"dc085284",
  2057 => x"dc125574",
  2058 => x"802eb138",
  2059 => x"88150884",
  2060 => x"1608ff05",
  2061 => x"54548073",
  2062 => x"249c388c",
  2063 => x"14227090",
  2064 => x"2b70902c",
  2065 => x"51535871",
  2066 => x"ad3880dc",
  2067 => x"14ff1454",
  2068 => x"54728025",
  2069 => x"e6387408",
  2070 => x"5574d138",
  2071 => x"75800c89",
  2072 => x"3d0d0473",
  2073 => x"51762d75",
  2074 => x"80080780",
  2075 => x"dc15ff15",
  2076 => x"555556ff",
  2077 => x"9e397351",
  2078 => x"762d7580",
  2079 => x"080780dc",
  2080 => x"15ff1555",
  2081 => x"5556ca39",
  2082 => x"ea3d0d68",
  2083 => x"8c112270",
  2084 => x"0a100a81",
  2085 => x"06575856",
  2086 => x"7480e438",
  2087 => x"8e162270",
  2088 => x"902b7090",
  2089 => x"2c515558",
  2090 => x"807424b1",
  2091 => x"38983dc4",
  2092 => x"05537352",
  2093 => x"80d1dc08",
  2094 => x"5186803f",
  2095 => x"800b8008",
  2096 => x"24973879",
  2097 => x"83e08006",
  2098 => x"547380c0",
  2099 => x"802e818f",
  2100 => x"38738280",
  2101 => x"802e8191",
  2102 => x"388c1622",
  2103 => x"57769080",
  2104 => x"0754738c",
  2105 => x"17238880",
  2106 => x"5280d1dc",
  2107 => x"0851d9ca",
  2108 => x"3f80089d",
  2109 => x"388c1622",
  2110 => x"82075473",
  2111 => x"8c172380",
  2112 => x"c3167077",
  2113 => x"0c90170c",
  2114 => x"810b9417",
  2115 => x"0c983d0d",
  2116 => x"0480d1dc",
  2117 => x"08b9a60b",
  2118 => x"bc120c54",
  2119 => x"8c162281",
  2120 => x"80075473",
  2121 => x"8c172380",
  2122 => x"08760c80",
  2123 => x"0890170c",
  2124 => x"88800b94",
  2125 => x"170c7480",
  2126 => x"2ed3388e",
  2127 => x"16227090",
  2128 => x"2b70902c",
  2129 => x"5355588c",
  2130 => x"a13f8008",
  2131 => x"802effbd",
  2132 => x"388c1622",
  2133 => x"81075473",
  2134 => x"8c172398",
  2135 => x"3d0d0481",
  2136 => x"0b8c1722",
  2137 => x"5855fef5",
  2138 => x"39a81608",
  2139 => x"80c5e22e",
  2140 => x"098106fe",
  2141 => x"e4388c16",
  2142 => x"22888007",
  2143 => x"54738c17",
  2144 => x"2388800b",
  2145 => x"80cc170c",
  2146 => x"fedc39fc",
  2147 => x"3d0d7679",
  2148 => x"71028c05",
  2149 => x"9f053357",
  2150 => x"55535583",
  2151 => x"72278a38",
  2152 => x"74830651",
  2153 => x"70802ea2",
  2154 => x"38ff1252",
  2155 => x"71ff2e93",
  2156 => x"38737370",
  2157 => x"81055534",
  2158 => x"ff125271",
  2159 => x"ff2e0981",
  2160 => x"06ef3874",
  2161 => x"800c863d",
  2162 => x"0d047474",
  2163 => x"882b7507",
  2164 => x"7071902b",
  2165 => x"07515451",
  2166 => x"8f7227a5",
  2167 => x"38727170",
  2168 => x"8405530c",
  2169 => x"72717084",
  2170 => x"05530c72",
  2171 => x"71708405",
  2172 => x"530c7271",
  2173 => x"70840553",
  2174 => x"0cf01252",
  2175 => x"718f26dd",
  2176 => x"38837227",
  2177 => x"90387271",
  2178 => x"70840553",
  2179 => x"0cfc1252",
  2180 => x"718326f2",
  2181 => x"387053ff",
  2182 => x"9039f93d",
  2183 => x"0d797c55",
  2184 => x"7b548e11",
  2185 => x"2270902b",
  2186 => x"70902c55",
  2187 => x"5780d1dc",
  2188 => x"08535856",
  2189 => x"83f33f80",
  2190 => x"0857800b",
  2191 => x"80082493",
  2192 => x"3880d016",
  2193 => x"08800805",
  2194 => x"80d0170c",
  2195 => x"76800c89",
  2196 => x"3d0d048c",
  2197 => x"162283df",
  2198 => x"ff065574",
  2199 => x"8c172376",
  2200 => x"800c893d",
  2201 => x"0d04fa3d",
  2202 => x"0d788c11",
  2203 => x"2270882a",
  2204 => x"70810651",
  2205 => x"57585674",
  2206 => x"a9388c16",
  2207 => x"2283dfff",
  2208 => x"0655748c",
  2209 => x"17237a54",
  2210 => x"79538e16",
  2211 => x"2270902b",
  2212 => x"70902c54",
  2213 => x"5680d1dc",
  2214 => x"08525681",
  2215 => x"b23f883d",
  2216 => x"0d048254",
  2217 => x"80538e16",
  2218 => x"2270902b",
  2219 => x"70902c54",
  2220 => x"5680d1dc",
  2221 => x"08525782",
  2222 => x"b83f8c16",
  2223 => x"2283dfff",
  2224 => x"0655748c",
  2225 => x"17237a54",
  2226 => x"79538e16",
  2227 => x"2270902b",
  2228 => x"70902c54",
  2229 => x"5680d1dc",
  2230 => x"08525680",
  2231 => x"f23f883d",
  2232 => x"0d04f93d",
  2233 => x"0d797c55",
  2234 => x"7b548e11",
  2235 => x"2270902b",
  2236 => x"70902c55",
  2237 => x"5780d1dc",
  2238 => x"08535856",
  2239 => x"81f33f80",
  2240 => x"08578008",
  2241 => x"ff2e9938",
  2242 => x"8c1622a0",
  2243 => x"80075574",
  2244 => x"8c172380",
  2245 => x"0880d017",
  2246 => x"0c76800c",
  2247 => x"893d0d04",
  2248 => x"8c162283",
  2249 => x"dfff0655",
  2250 => x"748c1723",
  2251 => x"76800c89",
  2252 => x"3d0d04fe",
  2253 => x"3d0d748e",
  2254 => x"11227090",
  2255 => x"2b70902c",
  2256 => x"55515153",
  2257 => x"80d1dc08",
  2258 => x"51bd3f84",
  2259 => x"3d0d04fb",
  2260 => x"3d0d800b",
  2261 => x"80e1d00c",
  2262 => x"7a537952",
  2263 => x"7851839a",
  2264 => x"3f800855",
  2265 => x"8008ff2e",
  2266 => x"88387480",
  2267 => x"0c873d0d",
  2268 => x"0480e1d0",
  2269 => x"08567580",
  2270 => x"2ef03877",
  2271 => x"76710c54",
  2272 => x"74800c87",
  2273 => x"3d0d04fd",
  2274 => x"3d0d800b",
  2275 => x"80e1d00c",
  2276 => x"765184ef",
  2277 => x"3f800853",
  2278 => x"8008ff2e",
  2279 => x"88387280",
  2280 => x"0c853d0d",
  2281 => x"0480e1d0",
  2282 => x"08547380",
  2283 => x"2ef03875",
  2284 => x"74710c52",
  2285 => x"72800c85",
  2286 => x"3d0d04fc",
  2287 => x"3d0d800b",
  2288 => x"80e1d00c",
  2289 => x"78527751",
  2290 => x"86d73f80",
  2291 => x"08548008",
  2292 => x"ff2e8838",
  2293 => x"73800c86",
  2294 => x"3d0d0480",
  2295 => x"e1d00855",
  2296 => x"74802ef0",
  2297 => x"38767571",
  2298 => x"0c537380",
  2299 => x"0c863d0d",
  2300 => x"04fb3d0d",
  2301 => x"800b80e1",
  2302 => x"d00c7a53",
  2303 => x"79527851",
  2304 => x"84b33f80",
  2305 => x"08558008",
  2306 => x"ff2e8838",
  2307 => x"74800c87",
  2308 => x"3d0d0480",
  2309 => x"e1d00856",
  2310 => x"75802ef0",
  2311 => x"38777671",
  2312 => x"0c547480",
  2313 => x"0c873d0d",
  2314 => x"04fb3d0d",
  2315 => x"800b80e1",
  2316 => x"d00c7a53",
  2317 => x"79527851",
  2318 => x"82b83f80",
  2319 => x"08558008",
  2320 => x"ff2e8838",
  2321 => x"74800c87",
  2322 => x"3d0d0480",
  2323 => x"e1d00856",
  2324 => x"75802ef0",
  2325 => x"38777671",
  2326 => x"0c547480",
  2327 => x"0c873d0d",
  2328 => x"04810b80",
  2329 => x"0c04803d",
  2330 => x"0d72812e",
  2331 => x"8938800b",
  2332 => x"800c823d",
  2333 => x"0d047351",
  2334 => x"80fa3ffe",
  2335 => x"3d0d80e1",
  2336 => x"c8085170",
  2337 => x"8a3880e1",
  2338 => x"d47080e1",
  2339 => x"c80c5170",
  2340 => x"75125252",
  2341 => x"ff537087",
  2342 => x"fb808026",
  2343 => x"88387080",
  2344 => x"e1c80c71",
  2345 => x"5372800c",
  2346 => x"843d0d04",
  2347 => x"fd3d0d80",
  2348 => x"0b80d1d0",
  2349 => x"08545472",
  2350 => x"812e9d38",
  2351 => x"7380e1cc",
  2352 => x"0cffbfe2",
  2353 => x"3fffbeb8",
  2354 => x"3f80e1a0",
  2355 => x"528151c1",
  2356 => x"a73f8008",
  2357 => x"5185ca3f",
  2358 => x"7280e1cc",
  2359 => x"0cffbfc6",
  2360 => x"3fffbe9c",
  2361 => x"3f80e1a0",
  2362 => x"528151c1",
  2363 => x"8b3f8008",
  2364 => x"5185ae3f",
  2365 => x"00ff3900",
  2366 => x"ff39f53d",
  2367 => x"0d7e6080",
  2368 => x"e1cc0870",
  2369 => x"5b585b5b",
  2370 => x"7580c538",
  2371 => x"777a25a2",
  2372 => x"38771b70",
  2373 => x"337081ff",
  2374 => x"06585859",
  2375 => x"758a2e99",
  2376 => x"387681ff",
  2377 => x"0651ffbe",
  2378 => x"dc3f8118",
  2379 => x"58797824",
  2380 => x"e0387980",
  2381 => x"0c8d3d0d",
  2382 => x"048d51ff",
  2383 => x"bec73f78",
  2384 => x"337081ff",
  2385 => x"065257ff",
  2386 => x"bebb3f81",
  2387 => x"1858de39",
  2388 => x"79557a54",
  2389 => x"7d538552",
  2390 => x"8d3dfc05",
  2391 => x"51ffbde2",
  2392 => x"3f800856",
  2393 => x"84b43f7b",
  2394 => x"80080c75",
  2395 => x"800c8d3d",
  2396 => x"0d04f63d",
  2397 => x"0d7d7f80",
  2398 => x"e1cc0870",
  2399 => x"5b585a5a",
  2400 => x"7580c438",
  2401 => x"777925b6",
  2402 => x"38ffbdd4",
  2403 => x"3f800881",
  2404 => x"ff06708d",
  2405 => x"32703070",
  2406 => x"9f2a5151",
  2407 => x"5757768a",
  2408 => x"2e80c638",
  2409 => x"75802e80",
  2410 => x"c038771a",
  2411 => x"56767634",
  2412 => x"7651ffbd",
  2413 => x"d03f8118",
  2414 => x"58787824",
  2415 => x"cc387756",
  2416 => x"75800c8c",
  2417 => x"3d0d0478",
  2418 => x"5579547c",
  2419 => x"5384528c",
  2420 => x"3dfc0551",
  2421 => x"ffbceb3f",
  2422 => x"80085683",
  2423 => x"bd3f7a80",
  2424 => x"080c7580",
  2425 => x"0c8c3d0d",
  2426 => x"04771a56",
  2427 => x"8a763481",
  2428 => x"18588d51",
  2429 => x"ffbd8e3f",
  2430 => x"8a51ffbd",
  2431 => x"883f7756",
  2432 => x"ffbe39fb",
  2433 => x"3d0d80e1",
  2434 => x"cc087056",
  2435 => x"54738838",
  2436 => x"74800c87",
  2437 => x"3d0d0477",
  2438 => x"53835287",
  2439 => x"3dfc0551",
  2440 => x"ffbc9f3f",
  2441 => x"80085482",
  2442 => x"f13f7580",
  2443 => x"080c7380",
  2444 => x"0c873d0d",
  2445 => x"04fa3d0d",
  2446 => x"80e1cc08",
  2447 => x"802ea338",
  2448 => x"7a557954",
  2449 => x"78538652",
  2450 => x"883dfc05",
  2451 => x"51ffbbf2",
  2452 => x"3f800856",
  2453 => x"82c43f76",
  2454 => x"80080c75",
  2455 => x"800c883d",
  2456 => x"0d0482b6",
  2457 => x"3f9d0b80",
  2458 => x"080cff0b",
  2459 => x"800c883d",
  2460 => x"0d04fb3d",
  2461 => x"0d777956",
  2462 => x"56807054",
  2463 => x"54737525",
  2464 => x"9f387410",
  2465 => x"1010f805",
  2466 => x"52721670",
  2467 => x"3370742b",
  2468 => x"76078116",
  2469 => x"f8165656",
  2470 => x"56515174",
  2471 => x"7324ea38",
  2472 => x"73800c87",
  2473 => x"3d0d04fc",
  2474 => x"3d0d7678",
  2475 => x"5555bc53",
  2476 => x"80527351",
  2477 => x"f5d53f84",
  2478 => x"527451ff",
  2479 => x"b53f8008",
  2480 => x"74238452",
  2481 => x"841551ff",
  2482 => x"a93f8008",
  2483 => x"82152384",
  2484 => x"52881551",
  2485 => x"ff9c3f80",
  2486 => x"0884150c",
  2487 => x"84528c15",
  2488 => x"51ff8f3f",
  2489 => x"80088815",
  2490 => x"23845290",
  2491 => x"1551ff82",
  2492 => x"3f80088a",
  2493 => x"15238452",
  2494 => x"941551fe",
  2495 => x"f53f8008",
  2496 => x"8c152384",
  2497 => x"52981551",
  2498 => x"fee83f80",
  2499 => x"088e1523",
  2500 => x"88529c15",
  2501 => x"51fedb3f",
  2502 => x"80089015",
  2503 => x"0c863d0d",
  2504 => x"04e93d0d",
  2505 => x"6a80e1cc",
  2506 => x"08575775",
  2507 => x"933880c0",
  2508 => x"800b8418",
  2509 => x"0c75ac18",
  2510 => x"0c75800c",
  2511 => x"993d0d04",
  2512 => x"893d7055",
  2513 => x"6a54558a",
  2514 => x"52993dff",
  2515 => x"bc0551ff",
  2516 => x"b9f03f80",
  2517 => x"08775375",
  2518 => x"5256fecb",
  2519 => x"3fbc3f77",
  2520 => x"80080c75",
  2521 => x"800c993d",
  2522 => x"0d04fc3d",
  2523 => x"0d815480",
  2524 => x"e1cc0888",
  2525 => x"3873800c",
  2526 => x"863d0d04",
  2527 => x"765397b9",
  2528 => x"52863dfc",
  2529 => x"0551ffb9",
  2530 => x"b93f8008",
  2531 => x"548c3f74",
  2532 => x"80080c73",
  2533 => x"800c863d",
  2534 => x"0d0480d1",
  2535 => x"dc08800c",
  2536 => x"04f73d0d",
  2537 => x"7b80d1dc",
  2538 => x"0882c811",
  2539 => x"085a545a",
  2540 => x"77802e80",
  2541 => x"da388188",
  2542 => x"18841908",
  2543 => x"ff058171",
  2544 => x"2b595559",
  2545 => x"80742480",
  2546 => x"ea388074",
  2547 => x"24b53873",
  2548 => x"822b7811",
  2549 => x"88055656",
  2550 => x"81801908",
  2551 => x"77065372",
  2552 => x"802eb638",
  2553 => x"78167008",
  2554 => x"53537951",
  2555 => x"74085372",
  2556 => x"2dff14fc",
  2557 => x"17fc1779",
  2558 => x"812c5a57",
  2559 => x"57547380",
  2560 => x"25d63877",
  2561 => x"085877ff",
  2562 => x"ad3880d1",
  2563 => x"dc0853bc",
  2564 => x"1308a538",
  2565 => x"7951f9dc",
  2566 => x"3f740853",
  2567 => x"722dff14",
  2568 => x"fc17fc17",
  2569 => x"79812c5a",
  2570 => x"57575473",
  2571 => x"8025ffa8",
  2572 => x"38d13980",
  2573 => x"57ff9339",
  2574 => x"7251bc13",
  2575 => x"0853722d",
  2576 => x"7951f9b0",
  2577 => x"3fff3d0d",
  2578 => x"80e1a80b",
  2579 => x"fc057008",
  2580 => x"525270ff",
  2581 => x"2e913870",
  2582 => x"2dfc1270",
  2583 => x"08525270",
  2584 => x"ff2e0981",
  2585 => x"06f13883",
  2586 => x"3d0d0404",
  2587 => x"ffb9a43f",
  2588 => x"04000000",
  2589 => x"00000040",
  2590 => x"72656164",
  2591 => x"2066726f",
  2592 => x"6d206164",
  2593 => x"72657373",
  2594 => x"20307831",
  2595 => x"3233340a",
  2596 => x"00000000",
  2597 => x"656e6420",
  2598 => x"73696d75",
  2599 => x"6c617469",
  2600 => x"6f6e2e0a",
  2601 => x"00000000",
  2602 => x"0a000000",
  2603 => x"43000000",
  2604 => x"64756d6d",
  2605 => x"792e6578",
  2606 => x"65000000",
  2607 => x"00ffffff",
  2608 => x"ff00ffff",
  2609 => x"ffff00ff",
  2610 => x"ffffff00",
  2611 => x"00000000",
  2612 => x"00000000",
  2613 => x"00000000",
  2614 => x"000030b0",
  2615 => x"000028e0",
  2616 => x"00000000",
  2617 => x"00002b48",
  2618 => x"00002ba4",
  2619 => x"00002c00",
  2620 => x"00000000",
  2621 => x"00000000",
  2622 => x"00000000",
  2623 => x"00000000",
  2624 => x"00000000",
  2625 => x"00000000",
  2626 => x"00000000",
  2627 => x"00000000",
  2628 => x"00000000",
  2629 => x"000028ac",
  2630 => x"00000000",
  2631 => x"00000000",
  2632 => x"00000000",
  2633 => x"00000000",
  2634 => x"00000000",
  2635 => x"00000000",
  2636 => x"00000000",
  2637 => x"00000000",
  2638 => x"00000000",
  2639 => x"00000000",
  2640 => x"00000000",
  2641 => x"00000000",
  2642 => x"00000000",
  2643 => x"00000000",
  2644 => x"00000000",
  2645 => x"00000000",
  2646 => x"00000000",
  2647 => x"00000000",
  2648 => x"00000000",
  2649 => x"00000000",
  2650 => x"00000000",
  2651 => x"00000000",
  2652 => x"00000000",
  2653 => x"00000000",
  2654 => x"00000000",
  2655 => x"00000000",
  2656 => x"00000000",
  2657 => x"00000000",
  2658 => x"00000001",
  2659 => x"330eabcd",
  2660 => x"1234e66d",
  2661 => x"deec0005",
  2662 => x"000b0000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000000",
  2675 => x"00000000",
  2676 => x"00000000",
  2677 => x"00000000",
  2678 => x"00000000",
  2679 => x"00000000",
  2680 => x"00000000",
  2681 => x"00000000",
  2682 => x"00000000",
  2683 => x"00000000",
  2684 => x"00000000",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000000",
  2688 => x"00000000",
  2689 => x"00000000",
  2690 => x"00000000",
  2691 => x"00000000",
  2692 => x"00000000",
  2693 => x"00000000",
  2694 => x"00000000",
  2695 => x"00000000",
  2696 => x"00000000",
  2697 => x"00000000",
  2698 => x"00000000",
  2699 => x"00000000",
  2700 => x"00000000",
  2701 => x"00000000",
  2702 => x"00000000",
  2703 => x"00000000",
  2704 => x"00000000",
  2705 => x"00000000",
  2706 => x"00000000",
  2707 => x"00000000",
  2708 => x"00000000",
  2709 => x"00000000",
  2710 => x"00000000",
  2711 => x"00000000",
  2712 => x"00000000",
  2713 => x"00000000",
  2714 => x"00000000",
  2715 => x"00000000",
  2716 => x"00000000",
  2717 => x"00000000",
  2718 => x"00000000",
  2719 => x"00000000",
  2720 => x"00000000",
  2721 => x"00000000",
  2722 => x"00000000",
  2723 => x"00000000",
  2724 => x"00000000",
  2725 => x"00000000",
  2726 => x"00000000",
  2727 => x"00000000",
  2728 => x"00000000",
  2729 => x"00000000",
  2730 => x"00000000",
  2731 => x"00000000",
  2732 => x"00000000",
  2733 => x"00000000",
  2734 => x"00000000",
  2735 => x"00000000",
  2736 => x"00000000",
  2737 => x"00000000",
  2738 => x"00000000",
  2739 => x"00000000",
  2740 => x"00000000",
  2741 => x"00000000",
  2742 => x"00000000",
  2743 => x"00000000",
  2744 => x"00000000",
  2745 => x"00000000",
  2746 => x"00000000",
  2747 => x"00000000",
  2748 => x"00000000",
  2749 => x"00000000",
  2750 => x"00000000",
  2751 => x"00000000",
  2752 => x"00000000",
  2753 => x"00000000",
  2754 => x"00000000",
  2755 => x"00000000",
  2756 => x"00000000",
  2757 => x"00000000",
  2758 => x"00000000",
  2759 => x"00000000",
  2760 => x"00000000",
  2761 => x"00000000",
  2762 => x"00000000",
  2763 => x"00000000",
  2764 => x"00000000",
  2765 => x"00000000",
  2766 => x"00000000",
  2767 => x"00000000",
  2768 => x"00000000",
  2769 => x"00000000",
  2770 => x"00000000",
  2771 => x"00000000",
  2772 => x"00000000",
  2773 => x"00000000",
  2774 => x"00000000",
  2775 => x"00000000",
  2776 => x"00000000",
  2777 => x"00000000",
  2778 => x"00000000",
  2779 => x"00000000",
  2780 => x"00000000",
  2781 => x"00000000",
  2782 => x"00000000",
  2783 => x"00000000",
  2784 => x"00000000",
  2785 => x"00000000",
  2786 => x"00000000",
  2787 => x"00000000",
  2788 => x"00000000",
  2789 => x"00000000",
  2790 => x"00000000",
  2791 => x"00000000",
  2792 => x"00000000",
  2793 => x"00000000",
  2794 => x"00000000",
  2795 => x"00000000",
  2796 => x"00000000",
  2797 => x"00000000",
  2798 => x"00000000",
  2799 => x"00000000",
  2800 => x"00000000",
  2801 => x"00000000",
  2802 => x"00000000",
  2803 => x"00000000",
  2804 => x"00000000",
  2805 => x"00000000",
  2806 => x"00000000",
  2807 => x"00000000",
  2808 => x"00000000",
  2809 => x"00000000",
  2810 => x"00000000",
  2811 => x"00000000",
  2812 => x"00000000",
  2813 => x"00000000",
  2814 => x"00000000",
  2815 => x"00000000",
  2816 => x"00000000",
  2817 => x"00000000",
  2818 => x"00000000",
  2819 => x"00000000",
  2820 => x"00000000",
  2821 => x"00000000",
  2822 => x"00000000",
  2823 => x"00000000",
  2824 => x"00000000",
  2825 => x"00000000",
  2826 => x"00000000",
  2827 => x"00000000",
  2828 => x"00000000",
  2829 => x"00000000",
  2830 => x"00000000",
  2831 => x"00000000",
  2832 => x"00000000",
  2833 => x"00000000",
  2834 => x"00000000",
  2835 => x"00000000",
  2836 => x"00000000",
  2837 => x"00000000",
  2838 => x"00000000",
  2839 => x"00000000",
  2840 => x"00000000",
  2841 => x"00000000",
  2842 => x"00000000",
  2843 => x"00000000",
  2844 => x"00000000",
  2845 => x"00000000",
  2846 => x"00000000",
  2847 => x"00000000",
  2848 => x"00000000",
  2849 => x"00000000",
  2850 => x"00000000",
  2851 => x"ffffffff",
  2852 => x"00000000",
  2853 => x"00020000",
  2854 => x"00000000",
  2855 => x"00000000",
  2856 => x"00002c98",
  2857 => x"00002c98",
  2858 => x"00002ca0",
  2859 => x"00002ca0",
  2860 => x"00002ca8",
  2861 => x"00002ca8",
  2862 => x"00002cb0",
  2863 => x"00002cb0",
  2864 => x"00002cb8",
  2865 => x"00002cb8",
  2866 => x"00002cc0",
  2867 => x"00002cc0",
  2868 => x"00002cc8",
  2869 => x"00002cc8",
  2870 => x"00002cd0",
  2871 => x"00002cd0",
  2872 => x"00002cd8",
  2873 => x"00002cd8",
  2874 => x"00002ce0",
  2875 => x"00002ce0",
  2876 => x"00002ce8",
  2877 => x"00002ce8",
  2878 => x"00002cf0",
  2879 => x"00002cf0",
  2880 => x"00002cf8",
  2881 => x"00002cf8",
  2882 => x"00002d00",
  2883 => x"00002d00",
  2884 => x"00002d08",
  2885 => x"00002d08",
  2886 => x"00002d10",
  2887 => x"00002d10",
  2888 => x"00002d18",
  2889 => x"00002d18",
  2890 => x"00002d20",
  2891 => x"00002d20",
  2892 => x"00002d28",
  2893 => x"00002d28",
  2894 => x"00002d30",
  2895 => x"00002d30",
  2896 => x"00002d38",
  2897 => x"00002d38",
  2898 => x"00002d40",
  2899 => x"00002d40",
  2900 => x"00002d48",
  2901 => x"00002d48",
  2902 => x"00002d50",
  2903 => x"00002d50",
  2904 => x"00002d58",
  2905 => x"00002d58",
  2906 => x"00002d60",
  2907 => x"00002d60",
  2908 => x"00002d68",
  2909 => x"00002d68",
  2910 => x"00002d70",
  2911 => x"00002d70",
  2912 => x"00002d78",
  2913 => x"00002d78",
  2914 => x"00002d80",
  2915 => x"00002d80",
  2916 => x"00002d88",
  2917 => x"00002d88",
  2918 => x"00002d90",
  2919 => x"00002d90",
  2920 => x"00002d98",
  2921 => x"00002d98",
  2922 => x"00002da0",
  2923 => x"00002da0",
  2924 => x"00002da8",
  2925 => x"00002da8",
  2926 => x"00002db0",
  2927 => x"00002db0",
  2928 => x"00002db8",
  2929 => x"00002db8",
  2930 => x"00002dc0",
  2931 => x"00002dc0",
  2932 => x"00002dc8",
  2933 => x"00002dc8",
  2934 => x"00002dd0",
  2935 => x"00002dd0",
  2936 => x"00002dd8",
  2937 => x"00002dd8",
  2938 => x"00002de0",
  2939 => x"00002de0",
  2940 => x"00002de8",
  2941 => x"00002de8",
  2942 => x"00002df0",
  2943 => x"00002df0",
  2944 => x"00002df8",
  2945 => x"00002df8",
  2946 => x"00002e00",
  2947 => x"00002e00",
  2948 => x"00002e08",
  2949 => x"00002e08",
  2950 => x"00002e10",
  2951 => x"00002e10",
  2952 => x"00002e18",
  2953 => x"00002e18",
  2954 => x"00002e20",
  2955 => x"00002e20",
  2956 => x"00002e28",
  2957 => x"00002e28",
  2958 => x"00002e30",
  2959 => x"00002e30",
  2960 => x"00002e38",
  2961 => x"00002e38",
  2962 => x"00002e40",
  2963 => x"00002e40",
  2964 => x"00002e48",
  2965 => x"00002e48",
  2966 => x"00002e50",
  2967 => x"00002e50",
  2968 => x"00002e58",
  2969 => x"00002e58",
  2970 => x"00002e60",
  2971 => x"00002e60",
  2972 => x"00002e68",
  2973 => x"00002e68",
  2974 => x"00002e70",
  2975 => x"00002e70",
  2976 => x"00002e78",
  2977 => x"00002e78",
  2978 => x"00002e80",
  2979 => x"00002e80",
  2980 => x"00002e88",
  2981 => x"00002e88",
  2982 => x"00002e90",
  2983 => x"00002e90",
  2984 => x"00002e98",
  2985 => x"00002e98",
  2986 => x"00002ea0",
  2987 => x"00002ea0",
  2988 => x"00002ea8",
  2989 => x"00002ea8",
  2990 => x"00002eb0",
  2991 => x"00002eb0",
  2992 => x"00002eb8",
  2993 => x"00002eb8",
  2994 => x"00002ec0",
  2995 => x"00002ec0",
  2996 => x"00002ec8",
  2997 => x"00002ec8",
  2998 => x"00002ed0",
  2999 => x"00002ed0",
  3000 => x"00002ed8",
  3001 => x"00002ed8",
  3002 => x"00002ee0",
  3003 => x"00002ee0",
  3004 => x"00002ee8",
  3005 => x"00002ee8",
  3006 => x"00002ef0",
  3007 => x"00002ef0",
  3008 => x"00002ef8",
  3009 => x"00002ef8",
  3010 => x"00002f00",
  3011 => x"00002f00",
  3012 => x"00002f08",
  3013 => x"00002f08",
  3014 => x"00002f10",
  3015 => x"00002f10",
  3016 => x"00002f18",
  3017 => x"00002f18",
  3018 => x"00002f20",
  3019 => x"00002f20",
  3020 => x"00002f28",
  3021 => x"00002f28",
  3022 => x"00002f30",
  3023 => x"00002f30",
  3024 => x"00002f38",
  3025 => x"00002f38",
  3026 => x"00002f40",
  3027 => x"00002f40",
  3028 => x"00002f48",
  3029 => x"00002f48",
  3030 => x"00002f50",
  3031 => x"00002f50",
  3032 => x"00002f58",
  3033 => x"00002f58",
  3034 => x"00002f60",
  3035 => x"00002f60",
  3036 => x"00002f68",
  3037 => x"00002f68",
  3038 => x"00002f70",
  3039 => x"00002f70",
  3040 => x"00002f78",
  3041 => x"00002f78",
  3042 => x"00002f80",
  3043 => x"00002f80",
  3044 => x"00002f88",
  3045 => x"00002f88",
  3046 => x"00002f90",
  3047 => x"00002f90",
  3048 => x"00002f98",
  3049 => x"00002f98",
  3050 => x"00002fa0",
  3051 => x"00002fa0",
  3052 => x"00002fa8",
  3053 => x"00002fa8",
  3054 => x"00002fb0",
  3055 => x"00002fb0",
  3056 => x"00002fb8",
  3057 => x"00002fb8",
  3058 => x"00002fc0",
  3059 => x"00002fc0",
  3060 => x"00002fc8",
  3061 => x"00002fc8",
  3062 => x"00002fd0",
  3063 => x"00002fd0",
  3064 => x"00002fd8",
  3065 => x"00002fd8",
  3066 => x"00002fe0",
  3067 => x"00002fe0",
  3068 => x"00002fe8",
  3069 => x"00002fe8",
  3070 => x"00002ff0",
  3071 => x"00002ff0",
  3072 => x"00002ff8",
  3073 => x"00002ff8",
  3074 => x"00003000",
  3075 => x"00003000",
  3076 => x"00003008",
  3077 => x"00003008",
  3078 => x"00003010",
  3079 => x"00003010",
  3080 => x"00003018",
  3081 => x"00003018",
  3082 => x"00003020",
  3083 => x"00003020",
  3084 => x"00003028",
  3085 => x"00003028",
  3086 => x"00003030",
  3087 => x"00003030",
  3088 => x"00003038",
  3089 => x"00003038",
  3090 => x"00003040",
  3091 => x"00003040",
  3092 => x"00003048",
  3093 => x"00003048",
  3094 => x"00003050",
  3095 => x"00003050",
  3096 => x"00003058",
  3097 => x"00003058",
  3098 => x"00003060",
  3099 => x"00003060",
  3100 => x"00003068",
  3101 => x"00003068",
  3102 => x"00003070",
  3103 => x"00003070",
  3104 => x"00003078",
  3105 => x"00003078",
  3106 => x"00003080",
  3107 => x"00003080",
  3108 => x"00003088",
  3109 => x"00003088",
  3110 => x"00003090",
  3111 => x"00003090",
  3112 => x"000028b0",
  3113 => x"ffffffff",
  3114 => x"00000000",
  3115 => x"ffffffff",
  3116 => x"00000000",
  3117 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
