-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
    port (
        clk             : in  std_logic;
        --
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memAWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memARead        : out std_logic_vector(wordSize-1 downto 0);
        --
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto minAddrBit);
        memBWrite       : in  std_logic_vector(wordSize-1 downto 0);
        memBRead        : out std_logic_vector(wordSize-1 downto 0)
    );
end entity dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0bb6",
     1 => x"df040000",
     2 => x"00000000",
     3 => x"00000000",
     4 => x"00000000",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"0b0b0bb9",
     9 => x"c4040000",
    10 => x"00000000",
    11 => x"00000000",
    12 => x"00000000",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0bb8",
    73 => x"f8040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0bb8db",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80f4",
   162 => x"b8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"b8de0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"0b0b0bb9",
   169 => x"ac040000",
   170 => x"00000000",
   171 => x"00000000",
   172 => x"00000000",
   173 => x"00000000",
   174 => x"00000000",
   175 => x"00000000",
   176 => x"0b0b0bb9",
   177 => x"94040000",
   178 => x"00000000",
   179 => x"00000000",
   180 => x"00000000",
   181 => x"00000000",
   182 => x"00000000",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80f4c80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"ff3d0d02",
   257 => x"8f053351",
   258 => x"b6d23f71",
   259 => x"b00c833d",
   260 => x"0d04ff3d",
   261 => x"0d80f4d4",
   262 => x"08841108",
   263 => x"70810a07",
   264 => x"84130c53",
   265 => x"84110870",
   266 => x"fe0a0684",
   267 => x"130c5351",
   268 => x"800bb00c",
   269 => x"833d0d04",
   270 => x"fc3d0d8a",
   271 => x"51b1ab3f",
   272 => x"93953fb6",
   273 => x"af530b0b",
   274 => x"80e1e052",
   275 => x"0b0b80e1",
   276 => x"f0519396",
   277 => x"3f8ee153",
   278 => x"0b0b80e1",
   279 => x"f8520b0b",
   280 => x"80e2a851",
   281 => x"93843f8e",
   282 => x"e1530b0b",
   283 => x"80e2ac52",
   284 => x"0b0b80e2",
   285 => x"bc5192f2",
   286 => x"3f8ff753",
   287 => x"0b0b80e2",
   288 => x"c0520b0b",
   289 => x"80e2e051",
   290 => x"92e03f90",
   291 => x"a4530b0b",
   292 => x"80e2e852",
   293 => x"0b0b80e2",
   294 => x"f85192ce",
   295 => x"3f90e153",
   296 => x"0b0b80e2",
   297 => x"fc520b0b",
   298 => x"80e39851",
   299 => x"92bc3f88",
   300 => x"92530b0b",
   301 => x"80e3a052",
   302 => x"0b0b80e3",
   303 => x"c05192aa",
   304 => x"3f90ff53",
   305 => x"0b0b80e3",
   306 => x"c8520b0b",
   307 => x"80e3e851",
   308 => x"92983fb6",
   309 => x"c6530b0b",
   310 => x"80e3f052",
   311 => x"0b0b80e4",
   312 => x"8c519286",
   313 => x"3f92f553",
   314 => x"0b0b80e4",
   315 => x"94520b0b",
   316 => x"80e4b451",
   317 => x"91f43f96",
   318 => x"ef530b0b",
   319 => x"80e4b852",
   320 => x"0b0b80e8",
   321 => x"f45191e2",
   322 => x"3f95ad53",
   323 => x"0b0b80e4",
   324 => x"c4520b0b",
   325 => x"80e4d451",
   326 => x"91d03fb0",
   327 => x"e8530b0b",
   328 => x"80e4d852",
   329 => x"0b0b80e4",
   330 => x"ec5191be",
   331 => x"3fb3f053",
   332 => x"0b0b80e4",
   333 => x"f0520b0b",
   334 => x"80e59851",
   335 => x"91ac3fb4",
   336 => x"aa530b0b",
   337 => x"80e5a052",
   338 => x"0b0b80e5",
   339 => x"ac51919a",
   340 => x"3fb5d953",
   341 => x"0b0b80e5",
   342 => x"b0520b0b",
   343 => x"80e5d851",
   344 => x"91883fb4",
   345 => x"aa530b0b",
   346 => x"80e5e052",
   347 => x"0b0b80e6",
   348 => x"805190f6",
   349 => x"3fb69f53",
   350 => x"0b0b80e6",
   351 => x"84520b0b",
   352 => x"80e69451",
   353 => x"90e43f98",
   354 => x"a9530b0b",
   355 => x"80efd852",
   356 => x"0b0b80e1",
   357 => x"d85190d2",
   358 => x"3f98df3f",
   359 => x"91a93f81",
   360 => x"0b819ca0",
   361 => x"348184b0",
   362 => x"337081ff",
   363 => x"06555573",
   364 => x"80d238b2",
   365 => x"f23fb008",
   366 => x"bc389199",
   367 => x"3f80f4d4",
   368 => x"08700870",
   369 => x"842a7081",
   370 => x"06515155",
   371 => x"5573802e",
   372 => x"97388415",
   373 => x"0870810a",
   374 => x"0784170c",
   375 => x"54841508",
   376 => x"70fe0a06",
   377 => x"84170c54",
   378 => x"819ca033",
   379 => x"5574ffb5",
   380 => x"38863d0d",
   381 => x"04b2c33f",
   382 => x"b00881ff",
   383 => x"065191c3",
   384 => x"3fffb739",
   385 => x"800b8184",
   386 => x"b034998e",
   387 => x"3fb2983f",
   388 => x"b008802e",
   389 => x"ffa438dd",
   390 => x"39fc3d0d",
   391 => x"029b0533",
   392 => x"705254af",
   393 => x"a93f0b0b",
   394 => x"80e6ac51",
   395 => x"add63f73",
   396 => x"10101470",
   397 => x"101080f2",
   398 => x"e8057053",
   399 => x"5455adc4",
   400 => x"3f7251b9",
   401 => x"b93f9052",
   402 => x"b00881ff",
   403 => x"0651b0c7",
   404 => x"3f0b0b80",
   405 => x"e69c51ad",
   406 => x"ab3f7384",
   407 => x"2b80f4b0",
   408 => x"08118411",
   409 => x"08535654",
   410 => x"aee43f88",
   411 => x"52b00881",
   412 => x"ff0651b0",
   413 => x"a23f0b0b",
   414 => x"80e6a851",
   415 => x"ad863f80",
   416 => x"f4b00814",
   417 => x"88110852",
   418 => x"53aec33f",
   419 => x"8852b008",
   420 => x"81ff0651",
   421 => x"b0813f0b",
   422 => x"0b80e6b0",
   423 => x"51ace53f",
   424 => x"80f4b008",
   425 => x"148c1108",
   426 => x"5255aea2",
   427 => x"3f8852b0",
   428 => x"0881ff06",
   429 => x"51afe03f",
   430 => x"0b0b80e6",
   431 => x"b851acc4",
   432 => x"3f800b80",
   433 => x"f4b00815",
   434 => x"70085154",
   435 => x"5572752e",
   436 => x"83388155",
   437 => x"7451adf6",
   438 => x"3f8652b0",
   439 => x"0881ff06",
   440 => x"51afb43f",
   441 => x"80f4b008",
   442 => x"14700870",
   443 => x"9e2a8106",
   444 => x"51545572",
   445 => x"802eaf38",
   446 => x"0b0b80e6",
   447 => x"c451ac84",
   448 => x"3f0b0b80",
   449 => x"e6d051ab",
   450 => x"fb3f80f4",
   451 => x"b0081470",
   452 => x"08515372",
   453 => x"802ead38",
   454 => x"72812eba",
   455 => x"388a51ab",
   456 => x"c93f863d",
   457 => x"0d040b0b",
   458 => x"80e6dc51",
   459 => x"abd63f0b",
   460 => x"0b80e6d0",
   461 => x"51abcd3f",
   462 => x"80f4b008",
   463 => x"14700851",
   464 => x"5372d538",
   465 => x"0b0b80e6",
   466 => x"e851abb8",
   467 => x"3f8a51ab",
   468 => x"993f863d",
   469 => x"0d040b0b",
   470 => x"80e6f051",
   471 => x"aba63fed",
   472 => x"39f93d0d",
   473 => x"815192ae",
   474 => x"3fb00881",
   475 => x"ff065482",
   476 => x"5192a33f",
   477 => x"b0085883",
   478 => x"51929b3f",
   479 => x"b0085784",
   480 => x"5192933f",
   481 => x"b0085685",
   482 => x"51928b3f",
   483 => x"b0085586",
   484 => x"5192833f",
   485 => x"b00881ff",
   486 => x"06527389",
   487 => x"26bb3873",
   488 => x"902980f4",
   489 => x"b0080578",
   490 => x"84120c77",
   491 => x"88120c76",
   492 => x"8c120c53",
   493 => x"80729e2b",
   494 => x"53567176",
   495 => x"2e833881",
   496 => x"56743070",
   497 => x"76079f2a",
   498 => x"7707740c",
   499 => x"745258fc",
   500 => x"c83f73b0",
   501 => x"0c893d0d",
   502 => x"040b0b80",
   503 => x"e6f851aa",
   504 => x"a33f7351",
   505 => x"abe83f0b",
   506 => x"0b80e9ac",
   507 => x"51aa953f",
   508 => x"73b00c89",
   509 => x"3d0d04fd",
   510 => x"3d0d8151",
   511 => x"91983fb0",
   512 => x"0881ff06",
   513 => x"5482518f",
   514 => x"e43fb008",
   515 => x"52731010",
   516 => x"14701010",
   517 => x"80f2e805",
   518 => x"5253b4f5",
   519 => x"3f73b00c",
   520 => x"853d0d04",
   521 => x"ff3d0d81",
   522 => x"5190eb3f",
   523 => x"b00881ff",
   524 => x"06527189",
   525 => x"268d3871",
   526 => x"51fbde3f",
   527 => x"71b00c83",
   528 => x"3d0d040b",
   529 => x"0b80e798",
   530 => x"51a9b93f",
   531 => x"7151aafe",
   532 => x"3f0b0b80",
   533 => x"e9ac51a9",
   534 => x"ab3f71b0",
   535 => x"0c833d0d",
   536 => x"04ff3d0d",
   537 => x"80527151",
   538 => x"fbaf3f81",
   539 => x"127081ff",
   540 => x"06515289",
   541 => x"7227ef38",
   542 => x"71b00c83",
   543 => x"3d0d0480",
   544 => x"3d0d80f4",
   545 => x"b0085180",
   546 => x"c60b8412",
   547 => x"0c940b88",
   548 => x"120c810b",
   549 => x"8c120c81",
   550 => x"710cb40b",
   551 => x"94120c82",
   552 => x"0b98120c",
   553 => x"810b9c12",
   554 => x"0c800b90",
   555 => x"120cb20b",
   556 => x"a4120c81",
   557 => x"0ba8120c",
   558 => x"810bac12",
   559 => x"0c800ba0",
   560 => x"120cb20b",
   561 => x"b4120c81",
   562 => x"0bb8120c",
   563 => x"810bbc12",
   564 => x"0c810bb0",
   565 => x"120cb20b",
   566 => x"80c4120c",
   567 => x"810b80c8",
   568 => x"120c810b",
   569 => x"80cc120c",
   570 => x"800b80c0",
   571 => x"120cb30b",
   572 => x"80d4120c",
   573 => x"820b80d8",
   574 => x"120c820b",
   575 => x"80dc120c",
   576 => x"800b80d0",
   577 => x"120cb40b",
   578 => x"80e4120c",
   579 => x"820b80e8",
   580 => x"120c820b",
   581 => x"80ec120c",
   582 => x"810b80e0",
   583 => x"120c800b",
   584 => x"80f4120c",
   585 => x"810b80f8",
   586 => x"120c810b",
   587 => x"80fc120c",
   588 => x"810b80f0",
   589 => x"120cad0b",
   590 => x"8184120c",
   591 => x"810b8188",
   592 => x"120c810b",
   593 => x"818c120c",
   594 => x"810b8180",
   595 => x"120cb20b",
   596 => x"8194120c",
   597 => x"810b8198",
   598 => x"120c810b",
   599 => x"819c120c",
   600 => x"810b8190",
   601 => x"120c800b",
   602 => x"b00c823d",
   603 => x"0d04810b",
   604 => x"80f2e034",
   605 => x"04fe3d0d",
   606 => x"81518e9a",
   607 => x"3fb00881",
   608 => x"ff065271",
   609 => x"812e8295",
   610 => x"3880f2e4",
   611 => x"08700870",
   612 => x"fdff0651",
   613 => x"53537173",
   614 => x"0c72080b",
   615 => x"0b80e7b8",
   616 => x"5253a6e0",
   617 => x"3f0b0b80",
   618 => x"e7c851a6",
   619 => x"d73f7281",
   620 => x"06527180",
   621 => x"2e81ba38",
   622 => x"0b0b80e7",
   623 => x"d051a6c4",
   624 => x"3f0b0b80",
   625 => x"e7d851a6",
   626 => x"bb3f7281",
   627 => x"2a708106",
   628 => x"51527181",
   629 => x"bc380b0b",
   630 => x"80e7e451",
   631 => x"a6a63f0b",
   632 => x"0b80e7ec",
   633 => x"51a69d3f",
   634 => x"72822a70",
   635 => x"81065152",
   636 => x"71802e80",
   637 => x"f3380b0b",
   638 => x"80e7f051",
   639 => x"a6863f0b",
   640 => x"0b80e888",
   641 => x"51a5fd3f",
   642 => x"72882a70",
   643 => x"81065152",
   644 => x"71802e80",
   645 => x"ca380b0b",
   646 => x"80e89451",
   647 => x"a5e63f0b",
   648 => x"0b80e89c",
   649 => x"51a5dd3f",
   650 => x"72892a70",
   651 => x"81065152",
   652 => x"71802e96",
   653 => x"380b0b80",
   654 => x"e8ac51a5",
   655 => x"c73f8a51",
   656 => x"a5a83f72",
   657 => x"b00c843d",
   658 => x"0d040b0b",
   659 => x"80e8b451",
   660 => x"a5b23f8a",
   661 => x"51a5933f",
   662 => x"72b00c84",
   663 => x"3d0d040b",
   664 => x"0b80e8bc",
   665 => x"51ffb539",
   666 => x"0b0b80e8",
   667 => x"c851ff8c",
   668 => x"390b0b80",
   669 => x"e8dc51a5",
   670 => x"8b3f0b0b",
   671 => x"80e7d851",
   672 => x"a5823f72",
   673 => x"812a7081",
   674 => x"06515271",
   675 => x"802efec6",
   676 => x"380b0b80",
   677 => x"e8e451a4",
   678 => x"eb3ffeba",
   679 => x"3980f2e4",
   680 => x"08700870",
   681 => x"82800751",
   682 => x"5353fdea",
   683 => x"39fd3d0d",
   684 => x"8184ac08",
   685 => x"52f881c0",
   686 => x"8e800b80",
   687 => x"f4d40855",
   688 => x"5371802e",
   689 => x"80f73872",
   690 => x"81ff0684",
   691 => x"150c80f4",
   692 => x"b4337081",
   693 => x"ff065152",
   694 => x"71802e80",
   695 => x"c238729f",
   696 => x"2a731007",
   697 => x"538184b0",
   698 => x"337081ff",
   699 => x"06515271",
   700 => x"802ed438",
   701 => x"800b8184",
   702 => x"b0348f9e",
   703 => x"3f80f2e0",
   704 => x"33547380",
   705 => x"e23880f4",
   706 => x"d4087381",
   707 => x"ff068412",
   708 => x"0c80f4b4",
   709 => x"337081ff",
   710 => x"06515354",
   711 => x"71c03872",
   712 => x"812a739f",
   713 => x"2b0753ff",
   714 => x"bc397281",
   715 => x"2a739f2b",
   716 => x"075380fd",
   717 => x"51a78e3f",
   718 => x"80f4d408",
   719 => x"547281ff",
   720 => x"0684150c",
   721 => x"80f4b433",
   722 => x"7081ff06",
   723 => x"53547180",
   724 => x"2ed83872",
   725 => x"9f2a7310",
   726 => x"075380fd",
   727 => x"51a6e63f",
   728 => x"80f4d408",
   729 => x"54d73980",
   730 => x"0bb00c85",
   731 => x"3d0d04fd",
   732 => x"3d0d0b0b",
   733 => x"80e8ec51",
   734 => x"a38a3f80",
   735 => x"f2e40870",
   736 => x"08828007",
   737 => x"710c7008",
   738 => x"84808007",
   739 => x"710c5372",
   740 => x"0870902a",
   741 => x"81065154",
   742 => x"73f53872",
   743 => x"0870fdff",
   744 => x"06740c52",
   745 => x"0b0b80e8",
   746 => x"fc51a2d8",
   747 => x"3f73b00c",
   748 => x"853d0d04",
   749 => x"803d0d0b",
   750 => x"0b80e984",
   751 => x"51a2c53f",
   752 => x"8c51a2a6",
   753 => x"3f0b0b80",
   754 => x"e98851a2",
   755 => x"b73f8184",
   756 => x"ac08802e",
   757 => x"8e380b0b",
   758 => x"80e9a451",
   759 => x"a2a63f82",
   760 => x"3d0d040b",
   761 => x"0b80e9b0",
   762 => x"51a2993f",
   763 => x"810a51a2",
   764 => x"933f0b0b",
   765 => x"80e9c451",
   766 => x"a28a3f0b",
   767 => x"0b80e9ec",
   768 => x"51a2813f",
   769 => x"80c251a3",
   770 => x"c53f0b0b",
   771 => x"80ea8051",
   772 => x"a1f23f0b",
   773 => x"0b80ea88",
   774 => x"51a1e93f",
   775 => x"0b0b80ea",
   776 => x"9451a1e0",
   777 => x"3f823d0d",
   778 => x"04ff893f",
   779 => x"8bcc3f80",
   780 => x"0bb00c04",
   781 => x"fe3d0d80",
   782 => x"f4d80898",
   783 => x"11087084",
   784 => x"2a708106",
   785 => x"51535353",
   786 => x"70802e8d",
   787 => x"3871ef06",
   788 => x"98140c81",
   789 => x"0b8184b0",
   790 => x"34843d0d",
   791 => x"04fc3d0d",
   792 => x"80f4d408",
   793 => x"7008810a",
   794 => x"068184ac",
   795 => x"0c53a4f9",
   796 => x"3fa59d3f",
   797 => x"8ec13f97",
   798 => x"a83f80f4",
   799 => x"d8089811",
   800 => x"08880798",
   801 => x"120c5481",
   802 => x"84ac0881",
   803 => x"cd388880",
   804 => x"0b819cfc",
   805 => x"0cfe9d3f",
   806 => x"8184ac08",
   807 => x"802e828a",
   808 => x"380b0b80",
   809 => x"e8ec51a0",
   810 => x"db3f80f2",
   811 => x"e4087008",
   812 => x"82800771",
   813 => x"0c700884",
   814 => x"80800771",
   815 => x"0c547308",
   816 => x"70902a81",
   817 => x"06515574",
   818 => x"f5387308",
   819 => x"fdff0674",
   820 => x"0c0b0b80",
   821 => x"e8fc51a0",
   822 => x"ab3f8152",
   823 => x"92ee518c",
   824 => x"993ff881",
   825 => x"c08e800b",
   826 => x"80f4d408",
   827 => x"56548184",
   828 => x"ac08802e",
   829 => x"818a3873",
   830 => x"81ff0684",
   831 => x"160c80f4",
   832 => x"b4337081",
   833 => x"ff065153",
   834 => x"72802e80",
   835 => x"c238739f",
   836 => x"2a741007",
   837 => x"548184b0",
   838 => x"337081ff",
   839 => x"06515372",
   840 => x"802ed438",
   841 => x"800b8184",
   842 => x"b0348aee",
   843 => x"3f80f2e0",
   844 => x"33557481",
   845 => x"9f3880f4",
   846 => x"d4087481",
   847 => x"ff068412",
   848 => x"0c80f4b4",
   849 => x"337081ff",
   850 => x"06515455",
   851 => x"72c03873",
   852 => x"812a749f",
   853 => x"2b0754ff",
   854 => x"bc39b9d4",
   855 => x"0b819cfc",
   856 => x"0cfcd13f",
   857 => x"8184ac08",
   858 => x"feb738be",
   859 => x"3973812a",
   860 => x"749f2b07",
   861 => x"5480fd51",
   862 => x"a2cb3f80",
   863 => x"f4d40855",
   864 => x"7381ff06",
   865 => x"84160c80",
   866 => x"f4b43370",
   867 => x"81ff0654",
   868 => x"5572802e",
   869 => x"d838739f",
   870 => x"2a741007",
   871 => x"5480fd51",
   872 => x"a2a33f80",
   873 => x"f4d40855",
   874 => x"d739bedc",
   875 => x"0b819cfc",
   876 => x"0ced853f",
   877 => x"0b0b80e8",
   878 => x"ec519ec8",
   879 => x"3f80f2e4",
   880 => x"08700882",
   881 => x"8007710c",
   882 => x"70088480",
   883 => x"8007710c",
   884 => x"54fdeb39",
   885 => x"a4a03f80",
   886 => x"0b819c98",
   887 => x"34800b81",
   888 => x"9c943480",
   889 => x"0b819c9c",
   890 => x"0c04fc3d",
   891 => x"0d819c94",
   892 => x"335372a7",
   893 => x"2680c538",
   894 => x"76527210",
   895 => x"10107310",
   896 => x"058184b4",
   897 => x"0551a989",
   898 => x"3f775281",
   899 => x"9c943370",
   900 => x"90297131",
   901 => x"70101081",
   902 => x"87c40553",
   903 => x"5654a8f1",
   904 => x"3f819c94",
   905 => x"33701010",
   906 => x"819aa405",
   907 => x"7a710c54",
   908 => x"81055372",
   909 => x"819c9434",
   910 => x"863d0d04",
   911 => x"80ea9c51",
   912 => x"9dc23f86",
   913 => x"3d0d0480",
   914 => x"3d0d80ea",
   915 => x"b8519db4",
   916 => x"3f823d0d",
   917 => x"04fe3d0d",
   918 => x"819c9c08",
   919 => x"53728538",
   920 => x"843d0d04",
   921 => x"722db008",
   922 => x"53800b81",
   923 => x"9c9c0cb0",
   924 => x"088c3880",
   925 => x"eab8519d",
   926 => x"8b3f843d",
   927 => x"0d0480ee",
   928 => x"f8519d80",
   929 => x"3f7283ff",
   930 => x"ff26aa38",
   931 => x"81ff7327",
   932 => x"96387252",
   933 => x"90519d8f",
   934 => x"3f8a519c",
   935 => x"cd3f80ea",
   936 => x"b8519ce0",
   937 => x"3fd43972",
   938 => x"5288519c",
   939 => x"fa3f8a51",
   940 => x"9cb83fea",
   941 => x"397252a0",
   942 => x"519cec3f",
   943 => x"8a519caa",
   944 => x"3fdc39fa",
   945 => x"3d0d02a3",
   946 => x"05335675",
   947 => x"8d2e80f4",
   948 => x"38758832",
   949 => x"70307780",
   950 => x"ff327030",
   951 => x"72802571",
   952 => x"80250754",
   953 => x"51565855",
   954 => x"7495389f",
   955 => x"76278c38",
   956 => x"819c9833",
   957 => x"5580ce75",
   958 => x"27ae3888",
   959 => x"3d0d0481",
   960 => x"9c983356",
   961 => x"75802ef3",
   962 => x"3888519b",
   963 => x"dd3fa051",
   964 => x"9bd83f88",
   965 => x"519bd33f",
   966 => x"819c9833",
   967 => x"ff055776",
   968 => x"819c9834",
   969 => x"883d0d04",
   970 => x"75519bbe",
   971 => x"3f819c98",
   972 => x"33811155",
   973 => x"5773819c",
   974 => x"98347581",
   975 => x"9bc41834",
   976 => x"883d0d04",
   977 => x"8a519ba2",
   978 => x"3f819c98",
   979 => x"33811156",
   980 => x"5474819c",
   981 => x"9834800b",
   982 => x"819bc415",
   983 => x"34805680",
   984 => x"0b819bc4",
   985 => x"17335654",
   986 => x"74a02e83",
   987 => x"38815474",
   988 => x"802e9038",
   989 => x"73802e8b",
   990 => x"38811670",
   991 => x"81ff0657",
   992 => x"57dd3975",
   993 => x"802ebf38",
   994 => x"800b819c",
   995 => x"94335555",
   996 => x"747427ab",
   997 => x"38735774",
   998 => x"10101075",
   999 => x"10057654",
  1000 => x"819bc453",
  1001 => x"8184b405",
  1002 => x"51a7b23f",
  1003 => x"b008802e",
  1004 => x"a6388115",
  1005 => x"7081ff06",
  1006 => x"56547675",
  1007 => x"26d93880",
  1008 => x"eabc519a",
  1009 => x"bf3f80ea",
  1010 => x"b8519ab8",
  1011 => x"3f800b81",
  1012 => x"9c983488",
  1013 => x"3d0d0474",
  1014 => x"1010819a",
  1015 => x"a4057008",
  1016 => x"819c9c0c",
  1017 => x"56800b81",
  1018 => x"9c9834e7",
  1019 => x"39fb3d0d",
  1020 => x"029f0533",
  1021 => x"56800b81",
  1022 => x"9bc43381",
  1023 => x"9bc45652",
  1024 => x"5370a02e",
  1025 => x"09810696",
  1026 => x"38811370",
  1027 => x"81ff0681",
  1028 => x"9bc41170",
  1029 => x"33535654",
  1030 => x"5170a02e",
  1031 => x"ec388055",
  1032 => x"74762780",
  1033 => x"ea388074",
  1034 => x"33535171",
  1035 => x"712e8338",
  1036 => x"815171a0",
  1037 => x"2e9a3870",
  1038 => x"80c53871",
  1039 => x"a02e9138",
  1040 => x"81157081",
  1041 => x"ff065652",
  1042 => x"757526da",
  1043 => x"3880c039",
  1044 => x"81137081",
  1045 => x"ff06819b",
  1046 => x"c4117033",
  1047 => x"54525454",
  1048 => x"70a02e09",
  1049 => x"8106d938",
  1050 => x"81137081",
  1051 => x"ff06819b",
  1052 => x"c4117033",
  1053 => x"54525454",
  1054 => x"70a02ed4",
  1055 => x"38c23981",
  1056 => x"137081ff",
  1057 => x"06819bc4",
  1058 => x"11565452",
  1059 => x"ff983973",
  1060 => x"b00c873d",
  1061 => x"0d04f73d",
  1062 => x"0d02af05",
  1063 => x"3359800b",
  1064 => x"819bc433",
  1065 => x"819bc459",
  1066 => x"555673a0",
  1067 => x"2e098106",
  1068 => x"96388116",
  1069 => x"7081ff06",
  1070 => x"819bc411",
  1071 => x"70335359",
  1072 => x"575473a0",
  1073 => x"2eec3880",
  1074 => x"58777927",
  1075 => x"80ea3880",
  1076 => x"77335654",
  1077 => x"74742e83",
  1078 => x"38815474",
  1079 => x"a02e9a38",
  1080 => x"7380c538",
  1081 => x"74a02e91",
  1082 => x"38811870",
  1083 => x"81ff0659",
  1084 => x"55787826",
  1085 => x"da3880c0",
  1086 => x"39811670",
  1087 => x"81ff0681",
  1088 => x"9bc41170",
  1089 => x"33575257",
  1090 => x"5773a02e",
  1091 => x"098106d9",
  1092 => x"38811670",
  1093 => x"81ff0681",
  1094 => x"9bc41170",
  1095 => x"33575257",
  1096 => x"5773a02e",
  1097 => x"d438c239",
  1098 => x"81167081",
  1099 => x"ff06819b",
  1100 => x"c4115957",
  1101 => x"55ff9839",
  1102 => x"80538b3d",
  1103 => x"fc055276",
  1104 => x"51a8df3f",
  1105 => x"8b3d0d04",
  1106 => x"f73d0d02",
  1107 => x"af053359",
  1108 => x"800b819b",
  1109 => x"c433819b",
  1110 => x"c4595556",
  1111 => x"73a02e09",
  1112 => x"81069638",
  1113 => x"81167081",
  1114 => x"ff06819b",
  1115 => x"c4117033",
  1116 => x"53595754",
  1117 => x"73a02eec",
  1118 => x"38805877",
  1119 => x"792780ea",
  1120 => x"38807733",
  1121 => x"56547474",
  1122 => x"2e833881",
  1123 => x"5474a02e",
  1124 => x"9a387380",
  1125 => x"c53874a0",
  1126 => x"2e913881",
  1127 => x"187081ff",
  1128 => x"06595578",
  1129 => x"7826da38",
  1130 => x"80c03981",
  1131 => x"167081ff",
  1132 => x"06819bc4",
  1133 => x"11703357",
  1134 => x"52575773",
  1135 => x"a02e0981",
  1136 => x"06d93881",
  1137 => x"167081ff",
  1138 => x"06819bc4",
  1139 => x"11703357",
  1140 => x"52575773",
  1141 => x"a02ed438",
  1142 => x"c2398116",
  1143 => x"7081ff06",
  1144 => x"819bc411",
  1145 => x"595755ff",
  1146 => x"98399053",
  1147 => x"8b3dfc05",
  1148 => x"527651aa",
  1149 => x"ca3f8b3d",
  1150 => x"0d04fc3d",
  1151 => x"0d8a5195",
  1152 => x"e93f80ea",
  1153 => x"d05195fc",
  1154 => x"3f800b81",
  1155 => x"9c943353",
  1156 => x"53727227",
  1157 => x"80f53872",
  1158 => x"10101073",
  1159 => x"10058184",
  1160 => x"b4057052",
  1161 => x"5495dd3f",
  1162 => x"72842b70",
  1163 => x"7431822b",
  1164 => x"8187c411",
  1165 => x"33515355",
  1166 => x"71802eb7",
  1167 => x"387351a1",
  1168 => x"bd3fb008",
  1169 => x"81ff0652",
  1170 => x"71892693",
  1171 => x"38a05195",
  1172 => x"993f8112",
  1173 => x"7081ff06",
  1174 => x"53548972",
  1175 => x"27ef3880",
  1176 => x"eae85195",
  1177 => x"9f3f7473",
  1178 => x"31822b81",
  1179 => x"87c40551",
  1180 => x"95923f8a",
  1181 => x"5194f33f",
  1182 => x"81137081",
  1183 => x"ff06819c",
  1184 => x"94335454",
  1185 => x"55717326",
  1186 => x"ff8d388a",
  1187 => x"5194db3f",
  1188 => x"819c9433",
  1189 => x"b00c863d",
  1190 => x"0d04fe3d",
  1191 => x"0d819cf4",
  1192 => x"22ff0551",
  1193 => x"70819cf4",
  1194 => x"237083ff",
  1195 => x"ff065170",
  1196 => x"80c43881",
  1197 => x"9cf83351",
  1198 => x"7081ff2e",
  1199 => x"b9387010",
  1200 => x"1010819c",
  1201 => x"a4055271",
  1202 => x"33819cf8",
  1203 => x"34fe7234",
  1204 => x"819cf833",
  1205 => x"70101010",
  1206 => x"819ca405",
  1207 => x"52538211",
  1208 => x"22819cf4",
  1209 => x"23841208",
  1210 => x"53722d81",
  1211 => x"9cf42251",
  1212 => x"70802eff",
  1213 => x"be38843d",
  1214 => x"0d04f93d",
  1215 => x"0d02aa05",
  1216 => x"22568055",
  1217 => x"74101010",
  1218 => x"819ca405",
  1219 => x"70335252",
  1220 => x"7081fe2e",
  1221 => x"99388115",
  1222 => x"7081ff06",
  1223 => x"5652748a",
  1224 => x"2e098106",
  1225 => x"df38810b",
  1226 => x"b00c893d",
  1227 => x"0d04819c",
  1228 => x"f8337081",
  1229 => x"ff06819c",
  1230 => x"f4225354",
  1231 => x"587281ff",
  1232 => x"2eb03872",
  1233 => x"832b5470",
  1234 => x"762780de",
  1235 => x"38757131",
  1236 => x"7083ffff",
  1237 => x"0674819c",
  1238 => x"a4173370",
  1239 => x"832b819c",
  1240 => x"a6112256",
  1241 => x"58565257",
  1242 => x"577281ff",
  1243 => x"2e098106",
  1244 => x"d6387272",
  1245 => x"34758213",
  1246 => x"23798413",
  1247 => x"0c7781ff",
  1248 => x"06547373",
  1249 => x"2e963876",
  1250 => x"10101081",
  1251 => x"9ca40553",
  1252 => x"74733480",
  1253 => x"5170b00c",
  1254 => x"893d0d04",
  1255 => x"74819cf8",
  1256 => x"3475819c",
  1257 => x"f4238051",
  1258 => x"ec397076",
  1259 => x"31517081",
  1260 => x"9ca61523",
  1261 => x"ffbc39ff",
  1262 => x"3d0d8a52",
  1263 => x"71101010",
  1264 => x"819c9c05",
  1265 => x"51fe7134",
  1266 => x"ff127081",
  1267 => x"ff065351",
  1268 => x"71ea38ff",
  1269 => x"0b819cf8",
  1270 => x"34833d0d",
  1271 => x"04fe3d0d",
  1272 => x"02930533",
  1273 => x"02840597",
  1274 => x"05335452",
  1275 => x"71842e80",
  1276 => x"e9387184",
  1277 => x"24913871",
  1278 => x"812ead38",
  1279 => x"80eaec51",
  1280 => x"92823f84",
  1281 => x"3d0d0471",
  1282 => x"80d52e09",
  1283 => x"8106ed38",
  1284 => x"80eaf851",
  1285 => x"91ee3f72",
  1286 => x"8a2680ca",
  1287 => x"38721010",
  1288 => x"80efa405",
  1289 => x"52710804",
  1290 => x"80eb8451",
  1291 => x"91d63f72",
  1292 => x"9a2e828b",
  1293 => x"38729a24",
  1294 => x"80c23872",
  1295 => x"8c2e828a",
  1296 => x"38728c24",
  1297 => x"81df3872",
  1298 => x"862e0981",
  1299 => x"06983880",
  1300 => x"eb905191",
  1301 => x"af3f843d",
  1302 => x"0d0480eb",
  1303 => x"a05191a4",
  1304 => x"3f728f2e",
  1305 => x"8c3880eb",
  1306 => x"ac519198",
  1307 => x"3f843d0d",
  1308 => x"0480ebbc",
  1309 => x"51918d3f",
  1310 => x"843d0d04",
  1311 => x"72a82e81",
  1312 => x"d43872a8",
  1313 => x"24818238",
  1314 => x"729d2e09",
  1315 => x"8106d738",
  1316 => x"80ebd451",
  1317 => x"90ee3f84",
  1318 => x"3d0d0480",
  1319 => x"ebf05190",
  1320 => x"e33f843d",
  1321 => x"0d0480ec",
  1322 => x"905190d8",
  1323 => x"3f843d0d",
  1324 => x"0480eca4",
  1325 => x"5190cd3f",
  1326 => x"843d0d04",
  1327 => x"80ecc051",
  1328 => x"90c23f84",
  1329 => x"3d0d0480",
  1330 => x"ecd85190",
  1331 => x"b73f843d",
  1332 => x"0d0480e9",
  1333 => x"905190ac",
  1334 => x"3f843d0d",
  1335 => x"0480ecf0",
  1336 => x"5190a13f",
  1337 => x"843d0d04",
  1338 => x"80ed8051",
  1339 => x"90963f84",
  1340 => x"3d0d0480",
  1341 => x"ed985190",
  1342 => x"8b3f843d",
  1343 => x"0d0480ed",
  1344 => x"ac519080",
  1345 => x"3f843d0d",
  1346 => x"047280c5",
  1347 => x"2e80d138",
  1348 => x"7280e12e",
  1349 => x"098106fe",
  1350 => x"cd3880ed",
  1351 => x"bc518fe4",
  1352 => x"3f843d0d",
  1353 => x"04728f2e",
  1354 => x"80c13872",
  1355 => x"912e0981",
  1356 => x"06feb338",
  1357 => x"80edcc51",
  1358 => x"8fca3f84",
  1359 => x"3d0d0480",
  1360 => x"ede0518f",
  1361 => x"bf3f843d",
  1362 => x"0d0480ed",
  1363 => x"fc518fb4",
  1364 => x"3f843d0d",
  1365 => x"0480ee8c",
  1366 => x"518fa93f",
  1367 => x"843d0d04",
  1368 => x"80eeac51",
  1369 => x"8f9e3f84",
  1370 => x"3d0d0480",
  1371 => x"eec4518f",
  1372 => x"933f843d",
  1373 => x"0d04f73d",
  1374 => x"0d02b305",
  1375 => x"337c7008",
  1376 => x"c0808006",
  1377 => x"59545a80",
  1378 => x"5675832b",
  1379 => x"7707bfe0",
  1380 => x"80077070",
  1381 => x"84055208",
  1382 => x"71088c2a",
  1383 => x"bffe8006",
  1384 => x"79077198",
  1385 => x"2a728c2a",
  1386 => x"9fff0673",
  1387 => x"852a708f",
  1388 => x"06759f06",
  1389 => x"5651585d",
  1390 => x"58525558",
  1391 => x"748d3881",
  1392 => x"16568f76",
  1393 => x"27c3388b",
  1394 => x"3d0d0480",
  1395 => x"eee0518e",
  1396 => x"b33f7551",
  1397 => x"8ff83f84",
  1398 => x"52b00851",
  1399 => x"91b93f80",
  1400 => x"eeec518e",
  1401 => x"9f3f7452",
  1402 => x"88518ebb",
  1403 => x"3f8452b0",
  1404 => x"085191a3",
  1405 => x"3f80eef4",
  1406 => x"518e893f",
  1407 => x"78529051",
  1408 => x"8ea53f86",
  1409 => x"52b00851",
  1410 => x"918d3f80",
  1411 => x"eefc518d",
  1412 => x"f33f7251",
  1413 => x"8fb83f84",
  1414 => x"52b00851",
  1415 => x"90f93f80",
  1416 => x"ef84518d",
  1417 => x"df3f7351",
  1418 => x"8fa43f84",
  1419 => x"52b00851",
  1420 => x"90e53f80",
  1421 => x"ef8c518d",
  1422 => x"cb3f7752",
  1423 => x"a0518de7",
  1424 => x"3f8a52b0",
  1425 => x"085190cf",
  1426 => x"3f799238",
  1427 => x"8a518d9a",
  1428 => x"3f811656",
  1429 => x"8f7627fe",
  1430 => x"b038feeb",
  1431 => x"397881ff",
  1432 => x"06527451",
  1433 => x"faf73f8a",
  1434 => x"518cff3f",
  1435 => x"e439f83d",
  1436 => x"0d02ab05",
  1437 => x"33598056",
  1438 => x"75852be0",
  1439 => x"9011e080",
  1440 => x"12087098",
  1441 => x"2a718c2a",
  1442 => x"9fff0672",
  1443 => x"852a708f",
  1444 => x"06749f06",
  1445 => x"5551585b",
  1446 => x"53565955",
  1447 => x"74802e81",
  1448 => x"a13875bf",
  1449 => x"2681a938",
  1450 => x"80ef9451",
  1451 => x"8cd63f75",
  1452 => x"518e9b3f",
  1453 => x"8652b008",
  1454 => x"518fdc3f",
  1455 => x"80eeec51",
  1456 => x"8cc23f74",
  1457 => x"5288518c",
  1458 => x"de3f8452",
  1459 => x"b008518f",
  1460 => x"c63f80ee",
  1461 => x"f4518cac",
  1462 => x"3f765290",
  1463 => x"518cc83f",
  1464 => x"8652b008",
  1465 => x"518fb03f",
  1466 => x"80eefc51",
  1467 => x"8c963f72",
  1468 => x"518ddb3f",
  1469 => x"8452b008",
  1470 => x"518f9c3f",
  1471 => x"80ef8451",
  1472 => x"8c823f73",
  1473 => x"518dc73f",
  1474 => x"8452b008",
  1475 => x"518f883f",
  1476 => x"80ef8c51",
  1477 => x"8bee3f77",
  1478 => x"08c08080",
  1479 => x"0652a051",
  1480 => x"8c853f8a",
  1481 => x"52b00851",
  1482 => x"8eed3f78",
  1483 => x"81ac388a",
  1484 => x"518bb73f",
  1485 => x"80537481",
  1486 => x"2e81d938",
  1487 => x"76862e81",
  1488 => x"b5388116",
  1489 => x"5680ff76",
  1490 => x"27fead38",
  1491 => x"8a3d0d04",
  1492 => x"80ef9c51",
  1493 => x"8bae3fc0",
  1494 => x"16518cf2",
  1495 => x"3f8652b0",
  1496 => x"08518eb3",
  1497 => x"3f80eeec",
  1498 => x"518b993f",
  1499 => x"74528851",
  1500 => x"8bb53f84",
  1501 => x"52b00851",
  1502 => x"8e9d3f80",
  1503 => x"eef4518b",
  1504 => x"833f7652",
  1505 => x"90518b9f",
  1506 => x"3f8652b0",
  1507 => x"08518e87",
  1508 => x"3f80eefc",
  1509 => x"518aed3f",
  1510 => x"72518cb2",
  1511 => x"3f8452b0",
  1512 => x"08518df3",
  1513 => x"3f80ef84",
  1514 => x"518ad93f",
  1515 => x"73518c9e",
  1516 => x"3f8452b0",
  1517 => x"08518ddf",
  1518 => x"3f80ef8c",
  1519 => x"518ac53f",
  1520 => x"7708c080",
  1521 => x"800652a0",
  1522 => x"518adc3f",
  1523 => x"8a52b008",
  1524 => x"518dc43f",
  1525 => x"78802efe",
  1526 => x"d6387681",
  1527 => x"ff065274",
  1528 => x"51f7fa3f",
  1529 => x"8a518a82",
  1530 => x"3f805374",
  1531 => x"812e0981",
  1532 => x"06fec938",
  1533 => x"9f397281",
  1534 => x"06577680",
  1535 => x"2efec338",
  1536 => x"78527751",
  1537 => x"faf03f81",
  1538 => x"165680ff",
  1539 => x"7627fce8",
  1540 => x"38feb939",
  1541 => x"74537686",
  1542 => x"2e098106",
  1543 => x"fea438d6",
  1544 => x"39803d0d",
  1545 => x"80f4d008",
  1546 => x"51a0710c",
  1547 => x"81800b84",
  1548 => x"120c823d",
  1549 => x"0d04fe3d",
  1550 => x"0d740284",
  1551 => x"05970533",
  1552 => x"0288059b",
  1553 => x"05338813",
  1554 => x"0c8c120c",
  1555 => x"538c1308",
  1556 => x"70812a81",
  1557 => x"06515271",
  1558 => x"f4388c13",
  1559 => x"087081ff",
  1560 => x"06b00c51",
  1561 => x"843d0d04",
  1562 => x"fb3d0d80",
  1563 => x"0b80efd0",
  1564 => x"52568990",
  1565 => x"3f755574",
  1566 => x"105381d0",
  1567 => x"5280f4d0",
  1568 => x"0851ffb2",
  1569 => x"3fb00887",
  1570 => x"2a708106",
  1571 => x"51547380",
  1572 => x"2e993881",
  1573 => x"157081ff",
  1574 => x"0670982b",
  1575 => x"52565473",
  1576 => x"8025d438",
  1577 => x"75b00c87",
  1578 => x"3d0d0480",
  1579 => x"efdc5188",
  1580 => x"d33f7452",
  1581 => x"885188ef",
  1582 => x"3f80efe8",
  1583 => x"5188c53f",
  1584 => x"81167083",
  1585 => x"ffff0681",
  1586 => x"177081ff",
  1587 => x"0670982b",
  1588 => x"52585257",
  1589 => x"54738025",
  1590 => x"ff9d38c8",
  1591 => x"39f33d0d",
  1592 => x"7f028405",
  1593 => x"80c30533",
  1594 => x"02880580",
  1595 => x"c6052280",
  1596 => x"eff8545b",
  1597 => x"5558888c",
  1598 => x"3f785189",
  1599 => x"d13f80f0",
  1600 => x"84518880",
  1601 => x"3f735288",
  1602 => x"51889c3f",
  1603 => x"80e98451",
  1604 => x"87f23f80",
  1605 => x"57767927",
  1606 => x"81913873",
  1607 => x"108e3d5c",
  1608 => x"5a795381",
  1609 => x"90527751",
  1610 => x"fe8c3f76",
  1611 => x"882a5390",
  1612 => x"527751fe",
  1613 => x"813f7681",
  1614 => x"ff065390",
  1615 => x"527751fd",
  1616 => x"f53f811a",
  1617 => x"53819052",
  1618 => x"7751fdea",
  1619 => x"3f805380",
  1620 => x"e0527751",
  1621 => x"fde03fb0",
  1622 => x"08872a81",
  1623 => x"0654738a",
  1624 => x"38881808",
  1625 => x"7081ff06",
  1626 => x"5d567b81",
  1627 => x"ff0680ee",
  1628 => x"f8525687",
  1629 => x"8f3f7552",
  1630 => x"885187ab",
  1631 => x"3f80eba8",
  1632 => x"5187813f",
  1633 => x"e0165480",
  1634 => x"df7427b6",
  1635 => x"38768706",
  1636 => x"701c5755",
  1637 => x"a0763474",
  1638 => x"872eb938",
  1639 => x"81177083",
  1640 => x"ffff0658",
  1641 => x"55787726",
  1642 => x"fef73880",
  1643 => x"e00b8c19",
  1644 => x"0c8c1808",
  1645 => x"70812a81",
  1646 => x"06585a76",
  1647 => x"f4388f3d",
  1648 => x"0d047687",
  1649 => x"06701c55",
  1650 => x"55757434",
  1651 => x"74872e09",
  1652 => x"8106c938",
  1653 => x"7a5186ac",
  1654 => x"3f8a5186",
  1655 => x"8d3f8117",
  1656 => x"7083ffff",
  1657 => x"06585578",
  1658 => x"7726feb5",
  1659 => x"38ffbc39",
  1660 => x"fb3d0d81",
  1661 => x"51ed9f3f",
  1662 => x"8251eecc",
  1663 => x"3fb00881",
  1664 => x"ff065683",
  1665 => x"51ed8f3f",
  1666 => x"b00883ff",
  1667 => x"ff0680f4",
  1668 => x"d0085654",
  1669 => x"73843881",
  1670 => x"80547353",
  1671 => x"75527451",
  1672 => x"fdbb3f73",
  1673 => x"b00c873d",
  1674 => x"0d04fb3d",
  1675 => x"0d8151ee",
  1676 => x"973fb008",
  1677 => x"538251ee",
  1678 => x"8f3fb008",
  1679 => x"56b00883",
  1680 => x"38905672",
  1681 => x"fc065575",
  1682 => x"812e80f1",
  1683 => x"38805473",
  1684 => x"7627aa38",
  1685 => x"73830653",
  1686 => x"72802eae",
  1687 => x"3880eef8",
  1688 => x"5185a13f",
  1689 => x"74708405",
  1690 => x"560852a0",
  1691 => x"5185b83f",
  1692 => x"a05184f6",
  1693 => x"3f811454",
  1694 => x"757426d8",
  1695 => x"388a5184",
  1696 => x"e93f800b",
  1697 => x"b00c873d",
  1698 => x"0d0480f0",
  1699 => x"a05184f4",
  1700 => x"3f7452a0",
  1701 => x"5185903f",
  1702 => x"80f0a451",
  1703 => x"84e63f80",
  1704 => x"eef85184",
  1705 => x"df3f7470",
  1706 => x"84055608",
  1707 => x"52a05184",
  1708 => x"f63fa051",
  1709 => x"84b43f81",
  1710 => x"1454ffbc",
  1711 => x"3980eef8",
  1712 => x"5184c13f",
  1713 => x"740852a0",
  1714 => x"5184dc3f",
  1715 => x"8a51849a",
  1716 => x"3f800bb0",
  1717 => x"0c873d0d",
  1718 => x"04fc3d0d",
  1719 => x"8151ece8",
  1720 => x"3fb00852",
  1721 => x"8251ebae",
  1722 => x"3fb00881",
  1723 => x"ff067256",
  1724 => x"53835472",
  1725 => x"802ea138",
  1726 => x"7351eccc",
  1727 => x"3f811470",
  1728 => x"81ff06ff",
  1729 => x"157081ff",
  1730 => x"06b00879",
  1731 => x"7084055b",
  1732 => x"0c565255",
  1733 => x"5272e138",
  1734 => x"72b00c86",
  1735 => x"3d0d0480",
  1736 => x"3d0d8c51",
  1737 => x"83c43f80",
  1738 => x"0bb00c82",
  1739 => x"3d0d0480",
  1740 => x"3d0d80f4",
  1741 => x"e00851f8",
  1742 => x"bb9586a1",
  1743 => x"710c810b",
  1744 => x"b00c823d",
  1745 => x"0d04803d",
  1746 => x"0d8151ea",
  1747 => x"c93fb008",
  1748 => x"81ff0651",
  1749 => x"f6983f80",
  1750 => x"0bb00c82",
  1751 => x"3d0d04e1",
  1752 => x"fc3f04fb",
  1753 => x"3d0d7779",
  1754 => x"55558056",
  1755 => x"757524ab",
  1756 => x"38807424",
  1757 => x"9d388053",
  1758 => x"73527451",
  1759 => x"80e13fb0",
  1760 => x"08547580",
  1761 => x"2e8538b0",
  1762 => x"08305473",
  1763 => x"b00c873d",
  1764 => x"0d047330",
  1765 => x"76813257",
  1766 => x"54dc3974",
  1767 => x"30558156",
  1768 => x"738025d2",
  1769 => x"38ec39fa",
  1770 => x"3d0d787a",
  1771 => x"57558057",
  1772 => x"767524a4",
  1773 => x"38759f2c",
  1774 => x"54815375",
  1775 => x"74327431",
  1776 => x"5274519b",
  1777 => x"3fb00854",
  1778 => x"76802e85",
  1779 => x"38b00830",
  1780 => x"5473b00c",
  1781 => x"883d0d04",
  1782 => x"74305581",
  1783 => x"57d739fc",
  1784 => x"3d0d7678",
  1785 => x"53548153",
  1786 => x"80747326",
  1787 => x"52557280",
  1788 => x"2e983870",
  1789 => x"802ea938",
  1790 => x"807224a4",
  1791 => x"38711073",
  1792 => x"10757226",
  1793 => x"53545272",
  1794 => x"ea387351",
  1795 => x"78833874",
  1796 => x"5170b00c",
  1797 => x"863d0d04",
  1798 => x"72812a72",
  1799 => x"812a5353",
  1800 => x"72802ee6",
  1801 => x"38717426",
  1802 => x"ef387372",
  1803 => x"31757407",
  1804 => x"74812a74",
  1805 => x"812a5555",
  1806 => x"5654e539",
  1807 => x"10101010",
  1808 => x"10101010",
  1809 => x"10101010",
  1810 => x"10101010",
  1811 => x"10101010",
  1812 => x"10101010",
  1813 => x"10101010",
  1814 => x"10101053",
  1815 => x"51047381",
  1816 => x"ff067383",
  1817 => x"06098105",
  1818 => x"83051010",
  1819 => x"102b0772",
  1820 => x"fc060c51",
  1821 => x"51043c04",
  1822 => x"72728072",
  1823 => x"8106ff05",
  1824 => x"09720605",
  1825 => x"71105272",
  1826 => x"0a100a53",
  1827 => x"72ed3851",
  1828 => x"51535104",
  1829 => x"b008b408",
  1830 => x"b8087575",
  1831 => x"b7a72d50",
  1832 => x"50b00856",
  1833 => x"b80cb40c",
  1834 => x"b00c5104",
  1835 => x"b008b408",
  1836 => x"b8087575",
  1837 => x"b6e32d50",
  1838 => x"50b00856",
  1839 => x"b80cb40c",
  1840 => x"b00c5104",
  1841 => x"b008b408",
  1842 => x"b80898b4",
  1843 => x"2db80cb4",
  1844 => x"0cb00c04",
  1845 => x"ff3d0d02",
  1846 => x"8f053380",
  1847 => x"f4e40852",
  1848 => x"710c800b",
  1849 => x"b00c833d",
  1850 => x"0d04ff3d",
  1851 => x"0d028f05",
  1852 => x"3351819c",
  1853 => x"fc085271",
  1854 => x"2db00881",
  1855 => x"ff06b00c",
  1856 => x"833d0d04",
  1857 => x"fe3d0d74",
  1858 => x"70335353",
  1859 => x"71802e93",
  1860 => x"38811372",
  1861 => x"52819cfc",
  1862 => x"08535371",
  1863 => x"2d723352",
  1864 => x"71ef3884",
  1865 => x"3d0d04f4",
  1866 => x"3d0d7f02",
  1867 => x"8405bb05",
  1868 => x"33555788",
  1869 => x"0b8c3d5b",
  1870 => x"59895380",
  1871 => x"f0cc5279",
  1872 => x"5185c03f",
  1873 => x"73792e80",
  1874 => x"ff387856",
  1875 => x"73902e80",
  1876 => x"ec3802a7",
  1877 => x"0558768f",
  1878 => x"06547389",
  1879 => x"2680c238",
  1880 => x"7518b015",
  1881 => x"55557375",
  1882 => x"3476842a",
  1883 => x"ff177081",
  1884 => x"ff065855",
  1885 => x"5775df38",
  1886 => x"781a5575",
  1887 => x"75347970",
  1888 => x"33555573",
  1889 => x"802e9338",
  1890 => x"81157452",
  1891 => x"819cfc08",
  1892 => x"5755752d",
  1893 => x"74335473",
  1894 => x"ef3878b0",
  1895 => x"0c8e3d0d",
  1896 => x"047518b7",
  1897 => x"15555573",
  1898 => x"75347684",
  1899 => x"2aff1770",
  1900 => x"81ff0658",
  1901 => x"555775ff",
  1902 => x"9d38ffbc",
  1903 => x"39847057",
  1904 => x"5902a705",
  1905 => x"58ff8f39",
  1906 => x"82705759",
  1907 => x"f439f13d",
  1908 => x"0d618d3d",
  1909 => x"705b5c5a",
  1910 => x"807a5657",
  1911 => x"767a2481",
  1912 => x"85387817",
  1913 => x"548a5274",
  1914 => x"5183e63f",
  1915 => x"b008b005",
  1916 => x"53727434",
  1917 => x"8117578a",
  1918 => x"52745183",
  1919 => x"af3fb008",
  1920 => x"55b008de",
  1921 => x"38b00877",
  1922 => x"9f2a1870",
  1923 => x"812c5a56",
  1924 => x"56807825",
  1925 => x"9e387817",
  1926 => x"ff055575",
  1927 => x"19703355",
  1928 => x"53743373",
  1929 => x"34737534",
  1930 => x"8116ff16",
  1931 => x"56567776",
  1932 => x"24e93876",
  1933 => x"19588078",
  1934 => x"34807a24",
  1935 => x"177081ff",
  1936 => x"067c7033",
  1937 => x"56575556",
  1938 => x"72802e93",
  1939 => x"38811573",
  1940 => x"52819cfc",
  1941 => x"08585576",
  1942 => x"2d743353",
  1943 => x"72ef3873",
  1944 => x"b00c913d",
  1945 => x"0d04ad7b",
  1946 => x"3402ad05",
  1947 => x"7a307119",
  1948 => x"5656598a",
  1949 => x"52745182",
  1950 => x"d83fb008",
  1951 => x"b0055372",
  1952 => x"74348117",
  1953 => x"578a5274",
  1954 => x"5182a13f",
  1955 => x"b00855b0",
  1956 => x"08fecf38",
  1957 => x"feef39fd",
  1958 => x"3d0d0297",
  1959 => x"05330284",
  1960 => x"059b0533",
  1961 => x"55537274",
  1962 => x"279738a0",
  1963 => x"51819cfc",
  1964 => x"0852712d",
  1965 => x"81137081",
  1966 => x"ff065452",
  1967 => x"737326eb",
  1968 => x"38853d0d",
  1969 => x"04fd3d0d",
  1970 => x"80f4d808",
  1971 => x"7680c18d",
  1972 => x"2994120c",
  1973 => x"54850b98",
  1974 => x"150c9814",
  1975 => x"08708106",
  1976 => x"515372f6",
  1977 => x"38853d0d",
  1978 => x"04803d0d",
  1979 => x"80f4d808",
  1980 => x"51870b84",
  1981 => x"120cff0b",
  1982 => x"a4120ca7",
  1983 => x"0ba8120c",
  1984 => x"80c18d0b",
  1985 => x"94120c87",
  1986 => x"0b98120c",
  1987 => x"823d0d04",
  1988 => x"803d0d80",
  1989 => x"f4dc0851",
  1990 => x"80c80b8c",
  1991 => x"120c830b",
  1992 => x"88120c82",
  1993 => x"3d0d0480",
  1994 => x"3d0d80f4",
  1995 => x"dc088411",
  1996 => x"088106b0",
  1997 => x"0c51823d",
  1998 => x"0d04ff3d",
  1999 => x"0d80f4dc",
  2000 => x"08528412",
  2001 => x"08708106",
  2002 => x"51517080",
  2003 => x"2ef43871",
  2004 => x"087081ff",
  2005 => x"06b00c51",
  2006 => x"833d0d04",
  2007 => x"fe3d0d02",
  2008 => x"93053353",
  2009 => x"728a2e9c",
  2010 => x"3880f4dc",
  2011 => x"08528412",
  2012 => x"0870892a",
  2013 => x"70810651",
  2014 => x"515170f2",
  2015 => x"3872720c",
  2016 => x"843d0d04",
  2017 => x"80f4dc08",
  2018 => x"52841208",
  2019 => x"70892a70",
  2020 => x"81065151",
  2021 => x"5170f238",
  2022 => x"8d720c84",
  2023 => x"12087089",
  2024 => x"2a708106",
  2025 => x"51515170",
  2026 => x"c538d239",
  2027 => x"bc0802bc",
  2028 => x"0cfd3d0d",
  2029 => x"8053bc08",
  2030 => x"8c050852",
  2031 => x"bc088805",
  2032 => x"0851f89b",
  2033 => x"3fb00870",
  2034 => x"b00c5485",
  2035 => x"3d0dbc0c",
  2036 => x"04bc0802",
  2037 => x"bc0cfd3d",
  2038 => x"0d8153bc",
  2039 => x"088c0508",
  2040 => x"52bc0888",
  2041 => x"050851f7",
  2042 => x"f63fb008",
  2043 => x"70b00c54",
  2044 => x"853d0dbc",
  2045 => x"0c04803d",
  2046 => x"0d865184",
  2047 => x"963f8151",
  2048 => x"a1d33ffc",
  2049 => x"3d0d7670",
  2050 => x"797b5555",
  2051 => x"55558f72",
  2052 => x"278c3872",
  2053 => x"75078306",
  2054 => x"5170802e",
  2055 => x"a738ff12",
  2056 => x"5271ff2e",
  2057 => x"98387270",
  2058 => x"81055433",
  2059 => x"74708105",
  2060 => x"5634ff12",
  2061 => x"5271ff2e",
  2062 => x"098106ea",
  2063 => x"3874b00c",
  2064 => x"863d0d04",
  2065 => x"74517270",
  2066 => x"84055408",
  2067 => x"71708405",
  2068 => x"530c7270",
  2069 => x"84055408",
  2070 => x"71708405",
  2071 => x"530c7270",
  2072 => x"84055408",
  2073 => x"71708405",
  2074 => x"530c7270",
  2075 => x"84055408",
  2076 => x"71708405",
  2077 => x"530cf012",
  2078 => x"52718f26",
  2079 => x"c9388372",
  2080 => x"27953872",
  2081 => x"70840554",
  2082 => x"08717084",
  2083 => x"05530cfc",
  2084 => x"12527183",
  2085 => x"26ed3870",
  2086 => x"54ff8339",
  2087 => x"fd3d0d75",
  2088 => x"5384d813",
  2089 => x"08802e8a",
  2090 => x"38805372",
  2091 => x"b00c853d",
  2092 => x"0d048180",
  2093 => x"5272518d",
  2094 => x"9b3fb008",
  2095 => x"84d8140c",
  2096 => x"ff53b008",
  2097 => x"802ee438",
  2098 => x"b008549f",
  2099 => x"53807470",
  2100 => x"8405560c",
  2101 => x"ff135380",
  2102 => x"7324ce38",
  2103 => x"80747084",
  2104 => x"05560cff",
  2105 => x"13537280",
  2106 => x"25e338ff",
  2107 => x"bc39fd3d",
  2108 => x"0d757755",
  2109 => x"539f7427",
  2110 => x"8d389673",
  2111 => x"0cff5271",
  2112 => x"b00c853d",
  2113 => x"0d0484d8",
  2114 => x"13085271",
  2115 => x"802e9338",
  2116 => x"73101012",
  2117 => x"70087972",
  2118 => x"0c515271",
  2119 => x"b00c853d",
  2120 => x"0d047251",
  2121 => x"fef63fff",
  2122 => x"52b008d3",
  2123 => x"3884d813",
  2124 => x"08741010",
  2125 => x"1170087a",
  2126 => x"720c5151",
  2127 => x"52dd39f9",
  2128 => x"3d0d797b",
  2129 => x"5856769f",
  2130 => x"2680e838",
  2131 => x"84d81608",
  2132 => x"5473802e",
  2133 => x"aa387610",
  2134 => x"10147008",
  2135 => x"55557380",
  2136 => x"2eba3880",
  2137 => x"5873812e",
  2138 => x"8f3873ff",
  2139 => x"2ea33880",
  2140 => x"750c7651",
  2141 => x"732d8058",
  2142 => x"77b00c89",
  2143 => x"3d0d0475",
  2144 => x"51fe993f",
  2145 => x"ff58b008",
  2146 => x"ef3884d8",
  2147 => x"160854c6",
  2148 => x"3996760c",
  2149 => x"810bb00c",
  2150 => x"893d0d04",
  2151 => x"755181ed",
  2152 => x"3f7653b0",
  2153 => x"08527551",
  2154 => x"81ad3fb0",
  2155 => x"08b00c89",
  2156 => x"3d0d0496",
  2157 => x"760cff0b",
  2158 => x"b00c893d",
  2159 => x"0d04fc3d",
  2160 => x"0d767856",
  2161 => x"53ff5474",
  2162 => x"9f26b138",
  2163 => x"84d81308",
  2164 => x"5271802e",
  2165 => x"ae387410",
  2166 => x"10127008",
  2167 => x"53538154",
  2168 => x"71802e98",
  2169 => x"38825471",
  2170 => x"ff2e9138",
  2171 => x"83547181",
  2172 => x"2e8a3880",
  2173 => x"730c7451",
  2174 => x"712d8054",
  2175 => x"73b00c86",
  2176 => x"3d0d0472",
  2177 => x"51fd953f",
  2178 => x"b008f138",
  2179 => x"84d81308",
  2180 => x"52c439ff",
  2181 => x"3d0d7352",
  2182 => x"80f4e808",
  2183 => x"51fea03f",
  2184 => x"833d0d04",
  2185 => x"fe3d0d75",
  2186 => x"53745280",
  2187 => x"f4e80851",
  2188 => x"fdbc3f84",
  2189 => x"3d0d0480",
  2190 => x"3d0d80f4",
  2191 => x"e80851fc",
  2192 => x"db3f823d",
  2193 => x"0d04ff3d",
  2194 => x"0d735280",
  2195 => x"f4e80851",
  2196 => x"feec3f83",
  2197 => x"3d0d04fc",
  2198 => x"3d0d800b",
  2199 => x"819d840c",
  2200 => x"78527751",
  2201 => x"9caa3fb0",
  2202 => x"0854b008",
  2203 => x"ff2e8838",
  2204 => x"73b00c86",
  2205 => x"3d0d0481",
  2206 => x"9d840855",
  2207 => x"74802ef0",
  2208 => x"38767571",
  2209 => x"0c5373b0",
  2210 => x"0c863d0d",
  2211 => x"049bfc3f",
  2212 => x"04fc3d0d",
  2213 => x"76707970",
  2214 => x"73078306",
  2215 => x"54545455",
  2216 => x"7080c338",
  2217 => x"71700870",
  2218 => x"0970f7fb",
  2219 => x"fdff1306",
  2220 => x"70f88482",
  2221 => x"81800651",
  2222 => x"51535354",
  2223 => x"70a63884",
  2224 => x"14727470",
  2225 => x"8405560c",
  2226 => x"70087009",
  2227 => x"70f7fbfd",
  2228 => x"ff130670",
  2229 => x"f8848281",
  2230 => x"80065151",
  2231 => x"53535470",
  2232 => x"802edc38",
  2233 => x"73527170",
  2234 => x"81055333",
  2235 => x"51707370",
  2236 => x"81055534",
  2237 => x"70f03874",
  2238 => x"b00c863d",
  2239 => x"0d04fd3d",
  2240 => x"0d757071",
  2241 => x"83065355",
  2242 => x"5270b838",
  2243 => x"71700870",
  2244 => x"09f7fbfd",
  2245 => x"ff120670",
  2246 => x"f8848281",
  2247 => x"80065151",
  2248 => x"5253709d",
  2249 => x"38841370",
  2250 => x"087009f7",
  2251 => x"fbfdff12",
  2252 => x"0670f884",
  2253 => x"82818006",
  2254 => x"51515253",
  2255 => x"70802ee5",
  2256 => x"38725271",
  2257 => x"33517080",
  2258 => x"2e8a3881",
  2259 => x"12703352",
  2260 => x"5270f838",
  2261 => x"717431b0",
  2262 => x"0c853d0d",
  2263 => x"04fa3d0d",
  2264 => x"787a7c70",
  2265 => x"54555552",
  2266 => x"72802e80",
  2267 => x"d9387174",
  2268 => x"07830651",
  2269 => x"70802e80",
  2270 => x"d438ff13",
  2271 => x"5372ff2e",
  2272 => x"b1387133",
  2273 => x"74335651",
  2274 => x"74712e09",
  2275 => x"8106a938",
  2276 => x"72802e81",
  2277 => x"87387081",
  2278 => x"ff065170",
  2279 => x"802e80fc",
  2280 => x"38811281",
  2281 => x"15ff1555",
  2282 => x"555272ff",
  2283 => x"2e098106",
  2284 => x"d1387133",
  2285 => x"74335651",
  2286 => x"7081ff06",
  2287 => x"7581ff06",
  2288 => x"71713151",
  2289 => x"525270b0",
  2290 => x"0c883d0d",
  2291 => x"04717457",
  2292 => x"55837327",
  2293 => x"88387108",
  2294 => x"74082e88",
  2295 => x"38747655",
  2296 => x"52ff9739",
  2297 => x"fc135372",
  2298 => x"802eb138",
  2299 => x"74087009",
  2300 => x"f7fbfdff",
  2301 => x"120670f8",
  2302 => x"84828180",
  2303 => x"06515151",
  2304 => x"709a3884",
  2305 => x"15841757",
  2306 => x"55837327",
  2307 => x"d0387408",
  2308 => x"76082ed0",
  2309 => x"38747655",
  2310 => x"52fedf39",
  2311 => x"800bb00c",
  2312 => x"883d0d04",
  2313 => x"f33d0d60",
  2314 => x"6264725a",
  2315 => x"5a5e5e80",
  2316 => x"5c767081",
  2317 => x"05583380",
  2318 => x"f0d91133",
  2319 => x"70832a70",
  2320 => x"81065155",
  2321 => x"555672e9",
  2322 => x"3875ad2e",
  2323 => x"82883875",
  2324 => x"ab2e8284",
  2325 => x"38773070",
  2326 => x"79078025",
  2327 => x"79903270",
  2328 => x"30707207",
  2329 => x"80257307",
  2330 => x"53575751",
  2331 => x"5372802e",
  2332 => x"873875b0",
  2333 => x"2e81eb38",
  2334 => x"778a3888",
  2335 => x"5875b02e",
  2336 => x"83388a58",
  2337 => x"810a5a7b",
  2338 => x"8438fe0a",
  2339 => x"5a775279",
  2340 => x"51f6be3f",
  2341 => x"b0087853",
  2342 => x"7a525bf6",
  2343 => x"8f3fb008",
  2344 => x"5a807080",
  2345 => x"f0d91833",
  2346 => x"70822a70",
  2347 => x"81065156",
  2348 => x"565a5572",
  2349 => x"802e80c1",
  2350 => x"38d01656",
  2351 => x"75782580",
  2352 => x"d7388079",
  2353 => x"24757b26",
  2354 => x"07537293",
  2355 => x"38747a2e",
  2356 => x"80eb387a",
  2357 => x"762580ed",
  2358 => x"3872802e",
  2359 => x"80e738ff",
  2360 => x"77708105",
  2361 => x"59335759",
  2362 => x"80f0d916",
  2363 => x"3370822a",
  2364 => x"70810651",
  2365 => x"545472c1",
  2366 => x"38738306",
  2367 => x"5372802e",
  2368 => x"97387381",
  2369 => x"06c91755",
  2370 => x"53728538",
  2371 => x"ffa91654",
  2372 => x"73567776",
  2373 => x"24ffab38",
  2374 => x"80792480",
  2375 => x"f0387b80",
  2376 => x"2e843874",
  2377 => x"30557c80",
  2378 => x"2e8c38ff",
  2379 => x"17537883",
  2380 => x"387d5372",
  2381 => x"7d0c74b0",
  2382 => x"0c8f3d0d",
  2383 => x"04815375",
  2384 => x"7b24ff95",
  2385 => x"38817579",
  2386 => x"29177870",
  2387 => x"81055a33",
  2388 => x"585659ff",
  2389 => x"9339815c",
  2390 => x"76708105",
  2391 => x"583356fd",
  2392 => x"f4398077",
  2393 => x"33545472",
  2394 => x"80f82eb2",
  2395 => x"387280d8",
  2396 => x"32703070",
  2397 => x"80257607",
  2398 => x"51515372",
  2399 => x"802efdf8",
  2400 => x"38811733",
  2401 => x"82185856",
  2402 => x"9058fdf8",
  2403 => x"39810a55",
  2404 => x"7b8438fe",
  2405 => x"0a557f53",
  2406 => x"a2730cff",
  2407 => x"89398154",
  2408 => x"cc39fd3d",
  2409 => x"0d775476",
  2410 => x"53755280",
  2411 => x"f4e80851",
  2412 => x"fcf23f85",
  2413 => x"3d0d04f3",
  2414 => x"3d0d6062",
  2415 => x"64725a5a",
  2416 => x"5d5d805e",
  2417 => x"76708105",
  2418 => x"583380f0",
  2419 => x"d9113370",
  2420 => x"832a7081",
  2421 => x"06515555",
  2422 => x"5672e938",
  2423 => x"75ad2e81",
  2424 => x"ff3875ab",
  2425 => x"2e81fb38",
  2426 => x"77307079",
  2427 => x"07802579",
  2428 => x"90327030",
  2429 => x"70720780",
  2430 => x"25730753",
  2431 => x"57575153",
  2432 => x"72802e87",
  2433 => x"3875b02e",
  2434 => x"81e23877",
  2435 => x"8a388858",
  2436 => x"75b02e83",
  2437 => x"388a5877",
  2438 => x"52ff51f3",
  2439 => x"8f3fb008",
  2440 => x"78535aff",
  2441 => x"51f3aa3f",
  2442 => x"b0085b80",
  2443 => x"705a5580",
  2444 => x"f0d91633",
  2445 => x"70822a70",
  2446 => x"81065154",
  2447 => x"5472802e",
  2448 => x"80c138d0",
  2449 => x"16567578",
  2450 => x"2580d738",
  2451 => x"80792475",
  2452 => x"7b260753",
  2453 => x"72933874",
  2454 => x"7a2e80eb",
  2455 => x"387a7625",
  2456 => x"80ed3872",
  2457 => x"802e80e7",
  2458 => x"38ff7770",
  2459 => x"81055933",
  2460 => x"575980f0",
  2461 => x"d9163370",
  2462 => x"822a7081",
  2463 => x"06515454",
  2464 => x"72c13873",
  2465 => x"83065372",
  2466 => x"802e9738",
  2467 => x"738106c9",
  2468 => x"17555372",
  2469 => x"8538ffa9",
  2470 => x"16547356",
  2471 => x"777624ff",
  2472 => x"ab388079",
  2473 => x"24818938",
  2474 => x"7d802e84",
  2475 => x"38743055",
  2476 => x"7b802e8c",
  2477 => x"38ff1753",
  2478 => x"7883387c",
  2479 => x"53727c0c",
  2480 => x"74b00c8f",
  2481 => x"3d0d0481",
  2482 => x"53757b24",
  2483 => x"ff953881",
  2484 => x"75792917",
  2485 => x"78708105",
  2486 => x"5a335856",
  2487 => x"59ff9339",
  2488 => x"815e7670",
  2489 => x"81055833",
  2490 => x"56fdfd39",
  2491 => x"80773354",
  2492 => x"547280f8",
  2493 => x"2e80c338",
  2494 => x"7280d832",
  2495 => x"70307080",
  2496 => x"25760751",
  2497 => x"51537280",
  2498 => x"2efe8038",
  2499 => x"81173382",
  2500 => x"18585690",
  2501 => x"705358ff",
  2502 => x"51f1913f",
  2503 => x"b0087853",
  2504 => x"5aff51f1",
  2505 => x"ac3fb008",
  2506 => x"5b80705a",
  2507 => x"55fe8039",
  2508 => x"ff605455",
  2509 => x"a2730cfe",
  2510 => x"f7398154",
  2511 => x"ffba39fd",
  2512 => x"3d0d7754",
  2513 => x"76537552",
  2514 => x"80f4e808",
  2515 => x"51fce83f",
  2516 => x"853d0d04",
  2517 => x"f33d0d7f",
  2518 => x"618b1170",
  2519 => x"f8065c55",
  2520 => x"555e7296",
  2521 => x"26833890",
  2522 => x"59807924",
  2523 => x"747a2607",
  2524 => x"53805472",
  2525 => x"742e0981",
  2526 => x"0680cb38",
  2527 => x"7d518bca",
  2528 => x"3f7883f7",
  2529 => x"2680c638",
  2530 => x"78832a70",
  2531 => x"10101080",
  2532 => x"fca4058c",
  2533 => x"11085959",
  2534 => x"5a76782e",
  2535 => x"83b03884",
  2536 => x"1708fc06",
  2537 => x"568c1708",
  2538 => x"88180871",
  2539 => x"8c120c88",
  2540 => x"120c5875",
  2541 => x"17841108",
  2542 => x"81078412",
  2543 => x"0c537d51",
  2544 => x"8b893f88",
  2545 => x"175473b0",
  2546 => x"0c8f3d0d",
  2547 => x"0478892a",
  2548 => x"79832a5b",
  2549 => x"5372802e",
  2550 => x"bf387886",
  2551 => x"2ab8055a",
  2552 => x"847327b4",
  2553 => x"3880db13",
  2554 => x"5a947327",
  2555 => x"ab38788c",
  2556 => x"2a80ee05",
  2557 => x"5a80d473",
  2558 => x"279e3878",
  2559 => x"8f2a80f7",
  2560 => x"055a82d4",
  2561 => x"73279138",
  2562 => x"78922a80",
  2563 => x"fc055a8a",
  2564 => x"d4732784",
  2565 => x"3880fe5a",
  2566 => x"79101010",
  2567 => x"80fca405",
  2568 => x"8c110858",
  2569 => x"5576752e",
  2570 => x"a3388417",
  2571 => x"08fc0670",
  2572 => x"7a315556",
  2573 => x"738f2488",
  2574 => x"d5387380",
  2575 => x"25fee638",
  2576 => x"8c170857",
  2577 => x"76752e09",
  2578 => x"8106df38",
  2579 => x"811a5a80",
  2580 => x"fcb40857",
  2581 => x"7680fcac",
  2582 => x"2e82c038",
  2583 => x"841708fc",
  2584 => x"06707a31",
  2585 => x"5556738f",
  2586 => x"2481f938",
  2587 => x"80fcac0b",
  2588 => x"80fcb80c",
  2589 => x"80fcac0b",
  2590 => x"80fcb40c",
  2591 => x"738025fe",
  2592 => x"b23883ff",
  2593 => x"762783df",
  2594 => x"3875892a",
  2595 => x"76832a55",
  2596 => x"5372802e",
  2597 => x"bf387586",
  2598 => x"2ab80554",
  2599 => x"847327b4",
  2600 => x"3880db13",
  2601 => x"54947327",
  2602 => x"ab38758c",
  2603 => x"2a80ee05",
  2604 => x"5480d473",
  2605 => x"279e3875",
  2606 => x"8f2a80f7",
  2607 => x"055482d4",
  2608 => x"73279138",
  2609 => x"75922a80",
  2610 => x"fc05548a",
  2611 => x"d4732784",
  2612 => x"3880fe54",
  2613 => x"73101010",
  2614 => x"80fca405",
  2615 => x"88110856",
  2616 => x"5874782e",
  2617 => x"86cf3884",
  2618 => x"1508fc06",
  2619 => x"53757327",
  2620 => x"8d388815",
  2621 => x"08557478",
  2622 => x"2e098106",
  2623 => x"ea388c15",
  2624 => x"0880fca4",
  2625 => x"0b840508",
  2626 => x"718c1a0c",
  2627 => x"76881a0c",
  2628 => x"7888130c",
  2629 => x"788c180c",
  2630 => x"5d587953",
  2631 => x"807a2483",
  2632 => x"e6387282",
  2633 => x"2c81712b",
  2634 => x"5c537a7c",
  2635 => x"26819838",
  2636 => x"7b7b0653",
  2637 => x"7282f138",
  2638 => x"79fc0684",
  2639 => x"055a7a10",
  2640 => x"707d0654",
  2641 => x"5b7282e0",
  2642 => x"38841a5a",
  2643 => x"f1398817",
  2644 => x"8c110858",
  2645 => x"5876782e",
  2646 => x"098106fc",
  2647 => x"c238821a",
  2648 => x"5afdec39",
  2649 => x"78177981",
  2650 => x"0784190c",
  2651 => x"7080fcb8",
  2652 => x"0c7080fc",
  2653 => x"b40c80fc",
  2654 => x"ac0b8c12",
  2655 => x"0c8c1108",
  2656 => x"88120c74",
  2657 => x"81078412",
  2658 => x"0c741175",
  2659 => x"710c5153",
  2660 => x"7d5187b7",
  2661 => x"3f881754",
  2662 => x"fcac3980",
  2663 => x"fca40b84",
  2664 => x"05087a54",
  2665 => x"5c798025",
  2666 => x"fef83882",
  2667 => x"da397a09",
  2668 => x"7c067080",
  2669 => x"fca40b84",
  2670 => x"050c5c7a",
  2671 => x"105b7a7c",
  2672 => x"2685387a",
  2673 => x"85b83880",
  2674 => x"fca40b88",
  2675 => x"05087084",
  2676 => x"1208fc06",
  2677 => x"707c317c",
  2678 => x"72268f72",
  2679 => x"25075757",
  2680 => x"5c5d5572",
  2681 => x"802e80db",
  2682 => x"38797a16",
  2683 => x"80fc9c08",
  2684 => x"1b90115a",
  2685 => x"55575b80",
  2686 => x"fc9808ff",
  2687 => x"2e8838a0",
  2688 => x"8f13e080",
  2689 => x"06577652",
  2690 => x"7d5186c0",
  2691 => x"3fb00854",
  2692 => x"b008ff2e",
  2693 => x"9038b008",
  2694 => x"76278299",
  2695 => x"387480fc",
  2696 => x"a42e8291",
  2697 => x"3880fca4",
  2698 => x"0b880508",
  2699 => x"55841508",
  2700 => x"fc06707a",
  2701 => x"317a7226",
  2702 => x"8f722507",
  2703 => x"52555372",
  2704 => x"83e63874",
  2705 => x"79810784",
  2706 => x"170c7916",
  2707 => x"7080fca4",
  2708 => x"0b88050c",
  2709 => x"75810784",
  2710 => x"120c547e",
  2711 => x"525785eb",
  2712 => x"3f881754",
  2713 => x"fae03975",
  2714 => x"832a7054",
  2715 => x"54807424",
  2716 => x"819b3872",
  2717 => x"822c8171",
  2718 => x"2b80fca8",
  2719 => x"08077080",
  2720 => x"fca40b84",
  2721 => x"050c7510",
  2722 => x"101080fc",
  2723 => x"a4058811",
  2724 => x"08585a5d",
  2725 => x"53778c18",
  2726 => x"0c748818",
  2727 => x"0c768819",
  2728 => x"0c768c16",
  2729 => x"0cfcf339",
  2730 => x"797a1010",
  2731 => x"1080fca4",
  2732 => x"05705759",
  2733 => x"5d8c1508",
  2734 => x"5776752e",
  2735 => x"a3388417",
  2736 => x"08fc0670",
  2737 => x"7a315556",
  2738 => x"738f2483",
  2739 => x"ca387380",
  2740 => x"25848138",
  2741 => x"8c170857",
  2742 => x"76752e09",
  2743 => x"8106df38",
  2744 => x"8815811b",
  2745 => x"70830655",
  2746 => x"5b5572c9",
  2747 => x"387c8306",
  2748 => x"5372802e",
  2749 => x"fdb838ff",
  2750 => x"1df81959",
  2751 => x"5d881808",
  2752 => x"782eea38",
  2753 => x"fdb53983",
  2754 => x"1a53fc96",
  2755 => x"39831470",
  2756 => x"822c8171",
  2757 => x"2b80fca8",
  2758 => x"08077080",
  2759 => x"fca40b84",
  2760 => x"050c7610",
  2761 => x"101080fc",
  2762 => x"a4058811",
  2763 => x"08595b5e",
  2764 => x"5153fee1",
  2765 => x"3980fbe8",
  2766 => x"081758b0",
  2767 => x"08762e81",
  2768 => x"8d3880fc",
  2769 => x"9808ff2e",
  2770 => x"83ec3873",
  2771 => x"76311880",
  2772 => x"fbe80c73",
  2773 => x"87067057",
  2774 => x"5372802e",
  2775 => x"88388873",
  2776 => x"31701555",
  2777 => x"5676149f",
  2778 => x"ff06a080",
  2779 => x"71311770",
  2780 => x"547f5357",
  2781 => x"5383d53f",
  2782 => x"b00853b0",
  2783 => x"08ff2e81",
  2784 => x"a03880fb",
  2785 => x"e8081670",
  2786 => x"80fbe80c",
  2787 => x"747580fc",
  2788 => x"a40b8805",
  2789 => x"0c747631",
  2790 => x"18708107",
  2791 => x"51555658",
  2792 => x"7b80fca4",
  2793 => x"2e839c38",
  2794 => x"798f2682",
  2795 => x"cb38810b",
  2796 => x"84150c84",
  2797 => x"1508fc06",
  2798 => x"707a317a",
  2799 => x"72268f72",
  2800 => x"25075255",
  2801 => x"5372802e",
  2802 => x"fcf93880",
  2803 => x"db39b008",
  2804 => x"9fff0653",
  2805 => x"72feeb38",
  2806 => x"7780fbe8",
  2807 => x"0c80fca4",
  2808 => x"0b880508",
  2809 => x"7b188107",
  2810 => x"84120c55",
  2811 => x"80fc9408",
  2812 => x"78278638",
  2813 => x"7780fc94",
  2814 => x"0c80fc90",
  2815 => x"087827fc",
  2816 => x"ac387780",
  2817 => x"fc900c84",
  2818 => x"1508fc06",
  2819 => x"707a317a",
  2820 => x"72268f72",
  2821 => x"25075255",
  2822 => x"5372802e",
  2823 => x"fca53888",
  2824 => x"39807454",
  2825 => x"56fedb39",
  2826 => x"7d51829f",
  2827 => x"3f800bb0",
  2828 => x"0c8f3d0d",
  2829 => x"04735380",
  2830 => x"7424a938",
  2831 => x"72822c81",
  2832 => x"712b80fc",
  2833 => x"a8080770",
  2834 => x"80fca40b",
  2835 => x"84050c5d",
  2836 => x"53778c18",
  2837 => x"0c748818",
  2838 => x"0c768819",
  2839 => x"0c768c16",
  2840 => x"0cf9b739",
  2841 => x"83147082",
  2842 => x"2c81712b",
  2843 => x"80fca808",
  2844 => x"077080fc",
  2845 => x"a40b8405",
  2846 => x"0c5e5153",
  2847 => x"d4397b7b",
  2848 => x"065372fc",
  2849 => x"a338841a",
  2850 => x"7b105c5a",
  2851 => x"f139ff1a",
  2852 => x"8111515a",
  2853 => x"f7b93978",
  2854 => x"17798107",
  2855 => x"84190c8c",
  2856 => x"18088819",
  2857 => x"08718c12",
  2858 => x"0c88120c",
  2859 => x"597080fc",
  2860 => x"b80c7080",
  2861 => x"fcb40c80",
  2862 => x"fcac0b8c",
  2863 => x"120c8c11",
  2864 => x"0888120c",
  2865 => x"74810784",
  2866 => x"120c7411",
  2867 => x"75710c51",
  2868 => x"53f9bd39",
  2869 => x"75178411",
  2870 => x"08810784",
  2871 => x"120c538c",
  2872 => x"17088818",
  2873 => x"08718c12",
  2874 => x"0c88120c",
  2875 => x"587d5180",
  2876 => x"da3f8817",
  2877 => x"54f5cf39",
  2878 => x"7284150c",
  2879 => x"f41af806",
  2880 => x"70841e08",
  2881 => x"81060784",
  2882 => x"1e0c701d",
  2883 => x"545b850b",
  2884 => x"84140c85",
  2885 => x"0b88140c",
  2886 => x"8f7b27fd",
  2887 => x"cf38881c",
  2888 => x"527d5182",
  2889 => x"903f80fc",
  2890 => x"a40b8805",
  2891 => x"0880fbe8",
  2892 => x"085955fd",
  2893 => x"b7397780",
  2894 => x"fbe80c73",
  2895 => x"80fc980c",
  2896 => x"fc913972",
  2897 => x"84150cfd",
  2898 => x"a3390404",
  2899 => x"fd3d0d80",
  2900 => x"0b819d84",
  2901 => x"0c765186",
  2902 => x"cb3fb008",
  2903 => x"53b008ff",
  2904 => x"2e883872",
  2905 => x"b00c853d",
  2906 => x"0d04819d",
  2907 => x"84085473",
  2908 => x"802ef038",
  2909 => x"7574710c",
  2910 => x"5272b00c",
  2911 => x"853d0d04",
  2912 => x"fb3d0d77",
  2913 => x"705256c2",
  2914 => x"3f80fca4",
  2915 => x"0b880508",
  2916 => x"841108fc",
  2917 => x"06707b31",
  2918 => x"9fef05e0",
  2919 => x"8006e080",
  2920 => x"05565653",
  2921 => x"a0807424",
  2922 => x"94388052",
  2923 => x"7551ff9c",
  2924 => x"3f80fcac",
  2925 => x"08155372",
  2926 => x"b0082e8f",
  2927 => x"387551ff",
  2928 => x"8a3f8053",
  2929 => x"72b00c87",
  2930 => x"3d0d0473",
  2931 => x"30527551",
  2932 => x"fefa3fb0",
  2933 => x"08ff2ea8",
  2934 => x"3880fca4",
  2935 => x"0b880508",
  2936 => x"75753181",
  2937 => x"0784120c",
  2938 => x"5380fbe8",
  2939 => x"08743180",
  2940 => x"fbe80c75",
  2941 => x"51fed43f",
  2942 => x"810bb00c",
  2943 => x"873d0d04",
  2944 => x"80527551",
  2945 => x"fec63f80",
  2946 => x"fca40b88",
  2947 => x"0508b008",
  2948 => x"71315653",
  2949 => x"8f7525ff",
  2950 => x"a438b008",
  2951 => x"80fc9808",
  2952 => x"3180fbe8",
  2953 => x"0c748107",
  2954 => x"84140c75",
  2955 => x"51fe9c3f",
  2956 => x"8053ff90",
  2957 => x"39f63d0d",
  2958 => x"7c7e545b",
  2959 => x"72802e82",
  2960 => x"83387a51",
  2961 => x"fe843ff8",
  2962 => x"13841108",
  2963 => x"70fe0670",
  2964 => x"13841108",
  2965 => x"fc065d58",
  2966 => x"59545880",
  2967 => x"fcac0875",
  2968 => x"2e82de38",
  2969 => x"7884160c",
  2970 => x"80738106",
  2971 => x"545a727a",
  2972 => x"2e81d538",
  2973 => x"78158411",
  2974 => x"08810651",
  2975 => x"5372a038",
  2976 => x"78175779",
  2977 => x"81e63888",
  2978 => x"15085372",
  2979 => x"80fcac2e",
  2980 => x"82f9388c",
  2981 => x"1508708c",
  2982 => x"150c7388",
  2983 => x"120c5676",
  2984 => x"81078419",
  2985 => x"0c761877",
  2986 => x"710c5379",
  2987 => x"81913883",
  2988 => x"ff772781",
  2989 => x"c8387689",
  2990 => x"2a77832a",
  2991 => x"56537280",
  2992 => x"2ebf3876",
  2993 => x"862ab805",
  2994 => x"55847327",
  2995 => x"b43880db",
  2996 => x"13559473",
  2997 => x"27ab3876",
  2998 => x"8c2a80ee",
  2999 => x"055580d4",
  3000 => x"73279e38",
  3001 => x"768f2a80",
  3002 => x"f7055582",
  3003 => x"d4732791",
  3004 => x"3876922a",
  3005 => x"80fc0555",
  3006 => x"8ad47327",
  3007 => x"843880fe",
  3008 => x"55741010",
  3009 => x"1080fca4",
  3010 => x"05881108",
  3011 => x"55567376",
  3012 => x"2e82b338",
  3013 => x"841408fc",
  3014 => x"06537673",
  3015 => x"278d3888",
  3016 => x"14085473",
  3017 => x"762e0981",
  3018 => x"06ea388c",
  3019 => x"1408708c",
  3020 => x"1a0c7488",
  3021 => x"1a0c7888",
  3022 => x"120c5677",
  3023 => x"8c150c7a",
  3024 => x"51fc883f",
  3025 => x"8c3d0d04",
  3026 => x"77087871",
  3027 => x"31597705",
  3028 => x"88190854",
  3029 => x"577280fc",
  3030 => x"ac2e80e0",
  3031 => x"388c1808",
  3032 => x"708c150c",
  3033 => x"7388120c",
  3034 => x"56fe8939",
  3035 => x"8815088c",
  3036 => x"1608708c",
  3037 => x"130c5788",
  3038 => x"170cfea3",
  3039 => x"3976832a",
  3040 => x"70545580",
  3041 => x"75248198",
  3042 => x"3872822c",
  3043 => x"81712b80",
  3044 => x"fca80807",
  3045 => x"80fca40b",
  3046 => x"84050c53",
  3047 => x"74101010",
  3048 => x"80fca405",
  3049 => x"88110855",
  3050 => x"56758c19",
  3051 => x"0c738819",
  3052 => x"0c778817",
  3053 => x"0c778c15",
  3054 => x"0cff8439",
  3055 => x"815afdb4",
  3056 => x"39781773",
  3057 => x"81065457",
  3058 => x"72983877",
  3059 => x"08787131",
  3060 => x"5977058c",
  3061 => x"1908881a",
  3062 => x"08718c12",
  3063 => x"0c88120c",
  3064 => x"57577681",
  3065 => x"0784190c",
  3066 => x"7780fca4",
  3067 => x"0b88050c",
  3068 => x"80fca008",
  3069 => x"7726fec7",
  3070 => x"3880fc9c",
  3071 => x"08527a51",
  3072 => x"fafe3f7a",
  3073 => x"51fac43f",
  3074 => x"feba3981",
  3075 => x"788c150c",
  3076 => x"7888150c",
  3077 => x"738c1a0c",
  3078 => x"73881a0c",
  3079 => x"5afd8039",
  3080 => x"83157082",
  3081 => x"2c81712b",
  3082 => x"80fca808",
  3083 => x"0780fca4",
  3084 => x"0b84050c",
  3085 => x"51537410",
  3086 => x"101080fc",
  3087 => x"a4058811",
  3088 => x"085556fe",
  3089 => x"e4397453",
  3090 => x"807524a7",
  3091 => x"3872822c",
  3092 => x"81712b80",
  3093 => x"fca80807",
  3094 => x"80fca40b",
  3095 => x"84050c53",
  3096 => x"758c190c",
  3097 => x"7388190c",
  3098 => x"7788170c",
  3099 => x"778c150c",
  3100 => x"fdcd3983",
  3101 => x"1570822c",
  3102 => x"81712b80",
  3103 => x"fca80807",
  3104 => x"80fca40b",
  3105 => x"84050c51",
  3106 => x"53d63981",
  3107 => x"0bb00c04",
  3108 => x"803d0d72",
  3109 => x"812e8938",
  3110 => x"800bb00c",
  3111 => x"823d0d04",
  3112 => x"7351b23f",
  3113 => x"fe3d0d81",
  3114 => x"9d800851",
  3115 => x"708a3881",
  3116 => x"9d887081",
  3117 => x"9d800c51",
  3118 => x"70751252",
  3119 => x"52ff5370",
  3120 => x"87fb8080",
  3121 => x"26883870",
  3122 => x"819d800c",
  3123 => x"715372b0",
  3124 => x"0c843d0d",
  3125 => x"0400ff39",
  3126 => x"68656c70",
  3127 => x"00000000",
  3128 => x"73797374",
  3129 => x"656d2072",
  3130 => x"65736574",
  3131 => x"00000000",
  3132 => x"72657365",
  3133 => x"74000000",
  3134 => x"73657420",
  3135 => x"3c636861",
  3136 => x"6e6e656c",
  3137 => x"3e203c77",
  3138 => x"6169743e",
  3139 => x"203c6f6e",
  3140 => x"3e203c6f",
  3141 => x"66663e20",
  3142 => x"3c636f75",
  3143 => x"6e743e20",
  3144 => x"3c676174",
  3145 => x"653e0000",
  3146 => x"73657400",
  3147 => x"616c6961",
  3148 => x"7320666f",
  3149 => x"72207365",
  3150 => x"74000000",
  3151 => x"63680000",
  3152 => x"6e616d65",
  3153 => x"203c6368",
  3154 => x"616e6e65",
  3155 => x"6c3e203c",
  3156 => x"6368616e",
  3157 => x"6e656c5f",
  3158 => x"6e616d65",
  3159 => x"3e000000",
  3160 => x"6e616d65",
  3161 => x"00000000",
  3162 => x"67657420",
  3163 => x"3c636861",
  3164 => x"6e6e656c",
  3165 => x"3e000000",
  3166 => x"67657400",
  3167 => x"67657420",
  3168 => x"616c6c20",
  3169 => x"6368616e",
  3170 => x"6e656c20",
  3171 => x"73657474",
  3172 => x"696e6773",
  3173 => x"00000000",
  3174 => x"73746174",
  3175 => x"75730000",
  3176 => x"75706461",
  3177 => x"74652073",
  3178 => x"69676e61",
  3179 => x"6c73206f",
  3180 => x"6e20616c",
  3181 => x"6c206368",
  3182 => x"616e6e65",
  3183 => x"6c730000",
  3184 => x"75706461",
  3185 => x"74650000",
  3186 => x"73657420",
  3187 => x"64656d6f",
  3188 => x"6e737472",
  3189 => x"6174696f",
  3190 => x"6e20636f",
  3191 => x"6e666967",
  3192 => x"75726174",
  3193 => x"696f6e00",
  3194 => x"64656d6f",
  3195 => x"00000000",
  3196 => x"73686f77",
  3197 => x"20737973",
  3198 => x"74656d20",
  3199 => x"696e666f",
  3200 => x"203c7665",
  3201 => x"72626f73",
  3202 => x"653e0000",
  3203 => x"73797369",
  3204 => x"6e666f00",
  3205 => x"72656164",
  3206 => x"2f736574",
  3207 => x"20736670",
  3208 => x"20737461",
  3209 => x"74757320",
  3210 => x"3c6f6e2f",
  3211 => x"6f66663e",
  3212 => x"00000000",
  3213 => x"73667000",
  3214 => x"53465020",
  3215 => x"54582074",
  3216 => x"65737400",
  3217 => x"72756e6e",
  3218 => x"696e6720",
  3219 => x"6c696768",
  3220 => x"74000000",
  3221 => x"72756e00",
  3222 => x"63686563",
  3223 => x"6b204932",
  3224 => x"43206164",
  3225 => x"64726573",
  3226 => x"73000000",
  3227 => x"69326300",
  3228 => x"72656164",
  3229 => x"20454550",
  3230 => x"524f4d20",
  3231 => x"3c627573",
  3232 => x"3e203c69",
  3233 => x"32635f61",
  3234 => x"6464723e",
  3235 => x"203c6c65",
  3236 => x"6e677468",
  3237 => x"3e000000",
  3238 => x"65657072",
  3239 => x"6f6d0000",
  3240 => x"616c6961",
  3241 => x"7320666f",
  3242 => x"72207800",
  3243 => x"6d656d00",
  3244 => x"77726974",
  3245 => x"6520776f",
  3246 => x"7264203c",
  3247 => x"61646472",
  3248 => x"3e203c6c",
  3249 => x"656e6774",
  3250 => x"683e203c",
  3251 => x"76616c75",
  3252 => x"65287329",
  3253 => x"3e000000",
  3254 => x"776d656d",
  3255 => x"00000000",
  3256 => x"6558616d",
  3257 => x"696e6520",
  3258 => x"6d656d6f",
  3259 => x"7279203c",
  3260 => x"61646472",
  3261 => x"3e203c6c",
  3262 => x"656e6774",
  3263 => x"683e0000",
  3264 => x"78000000",
  3265 => x"636c6561",
  3266 => x"72207363",
  3267 => x"7265656e",
  3268 => x"00000000",
  3269 => x"636c6561",
  3270 => x"72000000",
  3271 => x"20207761",
  3272 => x"69743a20",
  3273 => x"00000000",
  3274 => x"20206f6e",
  3275 => x"3a200000",
  3276 => x"20206f66",
  3277 => x"663a2000",
  3278 => x"2020636f",
  3279 => x"756e743a",
  3280 => x"20000000",
  3281 => x"20206761",
  3282 => x"74656420",
  3283 => x"00000000",
  3284 => x"20207374",
  3285 => x"61747573",
  3286 => x"3a200000",
  3287 => x"20206469",
  3288 => x"72656374",
  3289 => x"00000000",
  3290 => x"69646c65",
  3291 => x"00000000",
  3292 => x"61637469",
  3293 => x"76650000",
  3294 => x"4572726f",
  3295 => x"723a2069",
  3296 => x"6e76616c",
  3297 => x"69642063",
  3298 => x"68616e6e",
  3299 => x"656c206e",
  3300 => x"756d6265",
  3301 => x"72202800",
  3302 => x"4572726f",
  3303 => x"723a2077",
  3304 => x"726f6e67",
  3305 => x"20636861",
  3306 => x"6e6e656c",
  3307 => x"206e756d",
  3308 => x"62657220",
  3309 => x"28000000",
  3310 => x"53465020",
  3311 => x"73746174",
  3312 => x"75733a20",
  3313 => x"00000000",
  3314 => x"0a202054",
  3315 => x"58200000",
  3316 => x"6661756c",
  3317 => x"74000000",
  3318 => x"0a20206d",
  3319 => x"6f64756c",
  3320 => x"65200000",
  3321 => x"70726573",
  3322 => x"656e7400",
  3323 => x"0a202000",
  3324 => x"6c6f7373",
  3325 => x"206f6620",
  3326 => x"72656365",
  3327 => x"69766572",
  3328 => x"20536967",
  3329 => x"6e616c00",
  3330 => x"0a202053",
  3331 => x"46502074",
  3332 => x"78200000",
  3333 => x"656e6162",
  3334 => x"6c656400",
  3335 => x"0a202062",
  3336 => x"616e6477",
  3337 => x"69746820",
  3338 => x"00000000",
  3339 => x"66756c6c",
  3340 => x"00000000",
  3341 => x"72656475",
  3342 => x"63656400",
  3343 => x"64697361",
  3344 => x"626c6564",
  3345 => x"00000000",
  3346 => x"6e6f726d",
  3347 => x"616c206f",
  3348 => x"70657261",
  3349 => x"74696f6e",
  3350 => x"00000000",
  3351 => x"6e6f726d",
  3352 => x"616c0000",
  3353 => x"6e6f7420",
  3354 => x"00000000",
  3355 => x"0a534654",
  3356 => x"20545820",
  3357 => x"74657374",
  3358 => x"00000000",
  3359 => x"0a646f6e",
  3360 => x"652e0000",
  3361 => x"0a0a0000",
  3362 => x"63656e74",
  3363 => x"72616c20",
  3364 => x"74726967",
  3365 => x"67657220",
  3366 => x"67656e65",
  3367 => x"7261746f",
  3368 => x"72000000",
  3369 => x"20286f6e",
  3370 => x"2073696d",
  3371 => x"290a0000",
  3372 => x"0a485720",
  3373 => x"73796e74",
  3374 => x"68657369",
  3375 => x"7a65643a",
  3376 => x"20000000",
  3377 => x"0a535720",
  3378 => x"636f6d70",
  3379 => x"696c6564",
  3380 => x"2020203a",
  3381 => x"204e6f76",
  3382 => x"20203420",
  3383 => x"32303131",
  3384 => x"20203135",
  3385 => x"3a35363a",
  3386 => x"31320000",
  3387 => x"0a737973",
  3388 => x"74656d20",
  3389 => x"636c6f63",
  3390 => x"6b20203a",
  3391 => x"20000000",
  3392 => x"204d487a",
  3393 => x"0a000000",
  3394 => x"44454255",
  3395 => x"47204d4f",
  3396 => x"44450000",
  3397 => x"204f4e0a",
  3398 => x"00000000",
  3399 => x"4552524f",
  3400 => x"523a2074",
  3401 => x"6f6f206d",
  3402 => x"75636820",
  3403 => x"636f6d6d",
  3404 => x"616e6473",
  3405 => x"2e0a0000",
  3406 => x"3e200000",
  3407 => x"636f6d6d",
  3408 => x"616e6420",
  3409 => x"6e6f7420",
  3410 => x"666f756e",
  3411 => x"642e0a00",
  3412 => x"73757070",
  3413 => x"6f727465",
  3414 => x"6420636f",
  3415 => x"6d6d616e",
  3416 => x"64733a0a",
  3417 => x"0a000000",
  3418 => x"202d2000",
  3419 => x"76656e64",
  3420 => x"6f723f20",
  3421 => x"20000000",
  3422 => x"485a4452",
  3423 => x"20202020",
  3424 => x"20000000",
  3425 => x"67616973",
  3426 => x"6c657220",
  3427 => x"20000000",
  3428 => x"4148422f",
  3429 => x"41504220",
  3430 => x"42726964",
  3431 => x"67650000",
  3432 => x"45534120",
  3433 => x"20202020",
  3434 => x"20000000",
  3435 => x"756e6b6e",
  3436 => x"6f776e20",
  3437 => x"64657669",
  3438 => x"63650000",
  3439 => x"4c656f6e",
  3440 => x"32204d65",
  3441 => x"6d6f7279",
  3442 => x"20436f6e",
  3443 => x"74726f6c",
  3444 => x"6c657200",
  3445 => x"47522031",
  3446 => x"302f3130",
  3447 => x"30204d62",
  3448 => x"69742045",
  3449 => x"74686572",
  3450 => x"6e657420",
  3451 => x"4d414300",
  3452 => x"64696666",
  3453 => x"6572656e",
  3454 => x"7469616c",
  3455 => x"20637572",
  3456 => x"72656e74",
  3457 => x"206d6f6e",
  3458 => x"69746f72",
  3459 => x"00000000",
  3460 => x"64656275",
  3461 => x"67207472",
  3462 => x"61636572",
  3463 => x"206d656d",
  3464 => x"6f727900",
  3465 => x"4541444f",
  3466 => x"47533130",
  3467 => x"32206469",
  3468 => x"73706c61",
  3469 => x"79206472",
  3470 => x"69766572",
  3471 => x"00000000",
  3472 => x"64656275",
  3473 => x"67206275",
  3474 => x"66666572",
  3475 => x"20636f6e",
  3476 => x"74726f6c",
  3477 => x"00000000",
  3478 => x"6265616d",
  3479 => x"20706f73",
  3480 => x"6974696f",
  3481 => x"6e206d6f",
  3482 => x"6e69746f",
  3483 => x"72000000",
  3484 => x"64656275",
  3485 => x"6720636f",
  3486 => x"6e736f6c",
  3487 => x"65000000",
  3488 => x"44434d20",
  3489 => x"70686173",
  3490 => x"65207368",
  3491 => x"69667420",
  3492 => x"636f6e74",
  3493 => x"726f6c00",
  3494 => x"5a505520",
  3495 => x"4d656d6f",
  3496 => x"72792077",
  3497 => x"72617070",
  3498 => x"65720000",
  3499 => x"5a505520",
  3500 => x"41484220",
  3501 => x"57726170",
  3502 => x"70657200",
  3503 => x"56474120",
  3504 => x"636f6e74",
  3505 => x"726f6c6c",
  3506 => x"65720000",
  3507 => x"4d6f6475",
  3508 => x"6c617220",
  3509 => x"54696d65",
  3510 => x"7220556e",
  3511 => x"69740000",
  3512 => x"47656e65",
  3513 => x"72616c20",
  3514 => x"50757270",
  3515 => x"6f736520",
  3516 => x"492f4f20",
  3517 => x"706f7274",
  3518 => x"00000000",
  3519 => x"47656e65",
  3520 => x"72696320",
  3521 => x"55415254",
  3522 => x"00000000",
  3523 => x"414d4241",
  3524 => x"20577261",
  3525 => x"70706572",
  3526 => x"20666f72",
  3527 => x"204f4320",
  3528 => x"4932432d",
  3529 => x"6d617374",
  3530 => x"65720000",
  3531 => x"53504920",
  3532 => x"4d656d6f",
  3533 => x"72792043",
  3534 => x"6f6e7472",
  3535 => x"6f6c6c65",
  3536 => x"72000000",
  3537 => x"4475616c",
  3538 => x"2d706f72",
  3539 => x"74204148",
  3540 => x"42205352",
  3541 => x"414d206d",
  3542 => x"6f64756c",
  3543 => x"65000000",
  3544 => x"20206170",
  3545 => x"62736c76",
  3546 => x"00000000",
  3547 => x"76656e64",
  3548 => x"20307800",
  3549 => x"64657620",
  3550 => x"30780000",
  3551 => x"76657220",
  3552 => x"00000000",
  3553 => x"69727120",
  3554 => x"00000000",
  3555 => x"61646472",
  3556 => x"20307800",
  3557 => x"6168626d",
  3558 => x"73740000",
  3559 => x"61686273",
  3560 => x"6c760000",
  3561 => x"00001466",
  3562 => x"000014fe",
  3563 => x"000014f3",
  3564 => x"000014e8",
  3565 => x"000014dd",
  3566 => x"000014d2",
  3567 => x"000014c7",
  3568 => x"000014bc",
  3569 => x"000014b1",
  3570 => x"000014a6",
  3571 => x"0000149b",
  3572 => x"69326320",
  3573 => x"464d430a",
  3574 => x"00000000",
  3575 => x"61646472",
  3576 => x"6573733a",
  3577 => x"20307800",
  3578 => x"2020202d",
  3579 => x"2d3e2020",
  3580 => x"2041434b",
  3581 => x"0a000000",
  3582 => x"72656164",
  3583 => x"20646174",
  3584 => x"61202800",
  3585 => x"20627974",
  3586 => x"65732920",
  3587 => x"66726f6d",
  3588 => x"20493243",
  3589 => x"2d616464",
  3590 => x"72657373",
  3591 => x"20307800",
  3592 => x"0a307800",
  3593 => x"203a2000",
  3594 => x"30622020",
  3595 => x"20202020",
  3596 => x"20202020",
  3597 => x"20202020",
  3598 => x"20202020",
  3599 => x"20202020",
  3600 => x"20202020",
  3601 => x"20202020",
  3602 => x"20200000",
  3603 => x"20202020",
  3604 => x"20202020",
  3605 => x"00000000",
  3606 => x"00202020",
  3607 => x"20202020",
  3608 => x"20202828",
  3609 => x"28282820",
  3610 => x"20202020",
  3611 => x"20202020",
  3612 => x"20202020",
  3613 => x"20202020",
  3614 => x"20881010",
  3615 => x"10101010",
  3616 => x"10101010",
  3617 => x"10101010",
  3618 => x"10040404",
  3619 => x"04040404",
  3620 => x"04040410",
  3621 => x"10101010",
  3622 => x"10104141",
  3623 => x"41414141",
  3624 => x"01010101",
  3625 => x"01010101",
  3626 => x"01010101",
  3627 => x"01010101",
  3628 => x"01010101",
  3629 => x"10101010",
  3630 => x"10104242",
  3631 => x"42424242",
  3632 => x"02020202",
  3633 => x"02020202",
  3634 => x"02020202",
  3635 => x"02020202",
  3636 => x"02020202",
  3637 => x"10101010",
  3638 => x"20000000",
  3639 => x"00000000",
  3640 => x"00000000",
  3641 => x"00000000",
  3642 => x"00000000",
  3643 => x"00000000",
  3644 => x"00000000",
  3645 => x"00000000",
  3646 => x"00000000",
  3647 => x"00000000",
  3648 => x"00000000",
  3649 => x"00000000",
  3650 => x"00000000",
  3651 => x"00000000",
  3652 => x"00000000",
  3653 => x"00000000",
  3654 => x"00000000",
  3655 => x"00000000",
  3656 => x"00000000",
  3657 => x"00000000",
  3658 => x"00000000",
  3659 => x"00000000",
  3660 => x"00000000",
  3661 => x"00000000",
  3662 => x"00000000",
  3663 => x"00000000",
  3664 => x"00000000",
  3665 => x"00000000",
  3666 => x"00000000",
  3667 => x"00000000",
  3668 => x"00000000",
  3669 => x"00000000",
  3670 => x"00000000",
  3671 => x"43000000",
  3672 => x"00000000",
  3673 => x"80000900",
  3674 => x"6368616e",
  3675 => x"6e656c20",
  3676 => x"30000000",
  3677 => x"00000000",
  3678 => x"00000000",
  3679 => x"6368616e",
  3680 => x"6e656c20",
  3681 => x"31000000",
  3682 => x"00000000",
  3683 => x"00000000",
  3684 => x"6368616e",
  3685 => x"6e656c20",
  3686 => x"32000000",
  3687 => x"00000000",
  3688 => x"00000000",
  3689 => x"6368616e",
  3690 => x"6e656c20",
  3691 => x"33000000",
  3692 => x"00000000",
  3693 => x"00000000",
  3694 => x"00000000",
  3695 => x"00000000",
  3696 => x"00000000",
  3697 => x"00000000",
  3698 => x"00000000",
  3699 => x"00000000",
  3700 => x"00000000",
  3701 => x"00000000",
  3702 => x"00000000",
  3703 => x"00000000",
  3704 => x"00000000",
  3705 => x"00000000",
  3706 => x"00000000",
  3707 => x"00000000",
  3708 => x"00000000",
  3709 => x"00000000",
  3710 => x"00000000",
  3711 => x"00000000",
  3712 => x"00000000",
  3713 => x"00000000",
  3714 => x"00000000",
  3715 => x"00000000",
  3716 => x"00000000",
  3717 => x"00000000",
  3718 => x"00000000",
  3719 => x"00000000",
  3720 => x"00000000",
  3721 => x"00000000",
  3722 => x"00000000",
  3723 => x"00000000",
  3724 => x"80000800",
  3725 => x"00000000",
  3726 => x"00ffffff",
  3727 => x"ff00ffff",
  3728 => x"ffff00ff",
  3729 => x"ffffff00",
  3730 => x"00000000",
  3731 => x"00000000",
  3732 => x"80000a00",
  3733 => x"80000400",
  3734 => x"80000200",
  3735 => x"80000100",
  3736 => x"80000004",
  3737 => x"80000000",
  3738 => x"00003a6c",
  3739 => x"00000000",
  3740 => x"00003cd4",
  3741 => x"00003d30",
  3742 => x"00003d8c",
  3743 => x"00000000",
  3744 => x"00000000",
  3745 => x"00000000",
  3746 => x"00000000",
  3747 => x"00000000",
  3748 => x"00000000",
  3749 => x"00000000",
  3750 => x"00000000",
  3751 => x"00000000",
  3752 => x"0000395c",
  3753 => x"00000000",
  3754 => x"00000000",
  3755 => x"00000000",
  3756 => x"00000000",
  3757 => x"00000000",
  3758 => x"00000000",
  3759 => x"00000000",
  3760 => x"00000000",
  3761 => x"00000000",
  3762 => x"00000000",
  3763 => x"00000000",
  3764 => x"00000000",
  3765 => x"00000000",
  3766 => x"00000000",
  3767 => x"00000000",
  3768 => x"00000000",
  3769 => x"00000000",
  3770 => x"00000000",
  3771 => x"00000000",
  3772 => x"00000000",
  3773 => x"00000000",
  3774 => x"00000000",
  3775 => x"00000000",
  3776 => x"00000000",
  3777 => x"00000000",
  3778 => x"00000000",
  3779 => x"00000000",
  3780 => x"00000000",
  3781 => x"00000001",
  3782 => x"330eabcd",
  3783 => x"1234e66d",
  3784 => x"deec0005",
  3785 => x"000b0000",
  3786 => x"00000000",
  3787 => x"00000000",
  3788 => x"00000000",
  3789 => x"00000000",
  3790 => x"00000000",
  3791 => x"00000000",
  3792 => x"00000000",
  3793 => x"00000000",
  3794 => x"00000000",
  3795 => x"00000000",
  3796 => x"00000000",
  3797 => x"00000000",
  3798 => x"00000000",
  3799 => x"00000000",
  3800 => x"00000000",
  3801 => x"00000000",
  3802 => x"00000000",
  3803 => x"00000000",
  3804 => x"00000000",
  3805 => x"00000000",
  3806 => x"00000000",
  3807 => x"00000000",
  3808 => x"00000000",
  3809 => x"00000000",
  3810 => x"00000000",
  3811 => x"00000000",
  3812 => x"00000000",
  3813 => x"00000000",
  3814 => x"00000000",
  3815 => x"00000000",
  3816 => x"00000000",
  3817 => x"00000000",
  3818 => x"00000000",
  3819 => x"00000000",
  3820 => x"00000000",
  3821 => x"00000000",
  3822 => x"00000000",
  3823 => x"00000000",
  3824 => x"00000000",
  3825 => x"00000000",
  3826 => x"00000000",
  3827 => x"00000000",
  3828 => x"00000000",
  3829 => x"00000000",
  3830 => x"00000000",
  3831 => x"00000000",
  3832 => x"00000000",
  3833 => x"00000000",
  3834 => x"00000000",
  3835 => x"00000000",
  3836 => x"00000000",
  3837 => x"00000000",
  3838 => x"00000000",
  3839 => x"00000000",
  3840 => x"00000000",
  3841 => x"00000000",
  3842 => x"00000000",
  3843 => x"00000000",
  3844 => x"00000000",
  3845 => x"00000000",
  3846 => x"00000000",
  3847 => x"00000000",
  3848 => x"00000000",
  3849 => x"00000000",
  3850 => x"00000000",
  3851 => x"00000000",
  3852 => x"00000000",
  3853 => x"00000000",
  3854 => x"00000000",
  3855 => x"00000000",
  3856 => x"00000000",
  3857 => x"00000000",
  3858 => x"00000000",
  3859 => x"00000000",
  3860 => x"00000000",
  3861 => x"00000000",
  3862 => x"00000000",
  3863 => x"00000000",
  3864 => x"00000000",
  3865 => x"00000000",
  3866 => x"00000000",
  3867 => x"00000000",
  3868 => x"00000000",
  3869 => x"00000000",
  3870 => x"00000000",
  3871 => x"00000000",
  3872 => x"00000000",
  3873 => x"00000000",
  3874 => x"00000000",
  3875 => x"00000000",
  3876 => x"00000000",
  3877 => x"00000000",
  3878 => x"00000000",
  3879 => x"00000000",
  3880 => x"00000000",
  3881 => x"00000000",
  3882 => x"00000000",
  3883 => x"00000000",
  3884 => x"00000000",
  3885 => x"00000000",
  3886 => x"00000000",
  3887 => x"00000000",
  3888 => x"00000000",
  3889 => x"00000000",
  3890 => x"00000000",
  3891 => x"00000000",
  3892 => x"00000000",
  3893 => x"00000000",
  3894 => x"00000000",
  3895 => x"00000000",
  3896 => x"00000000",
  3897 => x"00000000",
  3898 => x"00000000",
  3899 => x"00000000",
  3900 => x"00000000",
  3901 => x"00000000",
  3902 => x"00000000",
  3903 => x"00000000",
  3904 => x"00000000",
  3905 => x"00000000",
  3906 => x"00000000",
  3907 => x"00000000",
  3908 => x"00000000",
  3909 => x"00000000",
  3910 => x"00000000",
  3911 => x"00000000",
  3912 => x"00000000",
  3913 => x"00000000",
  3914 => x"00000000",
  3915 => x"00000000",
  3916 => x"00000000",
  3917 => x"00000000",
  3918 => x"00000000",
  3919 => x"00000000",
  3920 => x"00000000",
  3921 => x"00000000",
  3922 => x"00000000",
  3923 => x"00000000",
  3924 => x"00000000",
  3925 => x"00000000",
  3926 => x"00000000",
  3927 => x"00000000",
  3928 => x"00000000",
  3929 => x"00000000",
  3930 => x"00000000",
  3931 => x"00000000",
  3932 => x"00000000",
  3933 => x"00000000",
  3934 => x"00000000",
  3935 => x"00000000",
  3936 => x"00000000",
  3937 => x"00000000",
  3938 => x"00000000",
  3939 => x"00000000",
  3940 => x"00000000",
  3941 => x"00000000",
  3942 => x"00000000",
  3943 => x"00000000",
  3944 => x"00000000",
  3945 => x"00000000",
  3946 => x"00000000",
  3947 => x"00000000",
  3948 => x"00000000",
  3949 => x"00000000",
  3950 => x"00000000",
  3951 => x"00000000",
  3952 => x"00000000",
  3953 => x"00000000",
  3954 => x"00000000",
  3955 => x"00000000",
  3956 => x"00000000",
  3957 => x"00000000",
  3958 => x"00000000",
  3959 => x"00000000",
  3960 => x"00000000",
  3961 => x"00000000",
  3962 => x"00000000",
  3963 => x"00000000",
  3964 => x"00000000",
  3965 => x"00000000",
  3966 => x"00000000",
  3967 => x"00000000",
  3968 => x"00000000",
  3969 => x"00000000",
  3970 => x"00000000",
  3971 => x"00000000",
  3972 => x"00000000",
  3973 => x"00000000",
  3974 => x"ffffffff",
  3975 => x"00000000",
  3976 => x"00020000",
  3977 => x"00000000",
  3978 => x"00000000",
  3979 => x"00003e24",
  3980 => x"00003e24",
  3981 => x"00003e2c",
  3982 => x"00003e2c",
  3983 => x"00003e34",
  3984 => x"00003e34",
  3985 => x"00003e3c",
  3986 => x"00003e3c",
  3987 => x"00003e44",
  3988 => x"00003e44",
  3989 => x"00003e4c",
  3990 => x"00003e4c",
  3991 => x"00003e54",
  3992 => x"00003e54",
  3993 => x"00003e5c",
  3994 => x"00003e5c",
  3995 => x"00003e64",
  3996 => x"00003e64",
  3997 => x"00003e6c",
  3998 => x"00003e6c",
  3999 => x"00003e74",
  4000 => x"00003e74",
  4001 => x"00003e7c",
  4002 => x"00003e7c",
  4003 => x"00003e84",
  4004 => x"00003e84",
  4005 => x"00003e8c",
  4006 => x"00003e8c",
  4007 => x"00003e94",
  4008 => x"00003e94",
  4009 => x"00003e9c",
  4010 => x"00003e9c",
  4011 => x"00003ea4",
  4012 => x"00003ea4",
  4013 => x"00003eac",
  4014 => x"00003eac",
  4015 => x"00003eb4",
  4016 => x"00003eb4",
  4017 => x"00003ebc",
  4018 => x"00003ebc",
  4019 => x"00003ec4",
  4020 => x"00003ec4",
  4021 => x"00003ecc",
  4022 => x"00003ecc",
  4023 => x"00003ed4",
  4024 => x"00003ed4",
  4025 => x"00003edc",
  4026 => x"00003edc",
  4027 => x"00003ee4",
  4028 => x"00003ee4",
  4029 => x"00003eec",
  4030 => x"00003eec",
  4031 => x"00003ef4",
  4032 => x"00003ef4",
  4033 => x"00003efc",
  4034 => x"00003efc",
  4035 => x"00003f04",
  4036 => x"00003f04",
  4037 => x"00003f0c",
  4038 => x"00003f0c",
  4039 => x"00003f14",
  4040 => x"00003f14",
  4041 => x"00003f1c",
  4042 => x"00003f1c",
  4043 => x"00003f24",
  4044 => x"00003f24",
  4045 => x"00003f2c",
  4046 => x"00003f2c",
  4047 => x"00003f34",
  4048 => x"00003f34",
  4049 => x"00003f3c",
  4050 => x"00003f3c",
  4051 => x"00003f44",
  4052 => x"00003f44",
  4053 => x"00003f4c",
  4054 => x"00003f4c",
  4055 => x"00003f54",
  4056 => x"00003f54",
  4057 => x"00003f5c",
  4058 => x"00003f5c",
  4059 => x"00003f64",
  4060 => x"00003f64",
  4061 => x"00003f6c",
  4062 => x"00003f6c",
  4063 => x"00003f74",
  4064 => x"00003f74",
  4065 => x"00003f7c",
  4066 => x"00003f7c",
  4067 => x"00003f84",
  4068 => x"00003f84",
  4069 => x"00003f8c",
  4070 => x"00003f8c",
  4071 => x"00003f94",
  4072 => x"00003f94",
  4073 => x"00003f9c",
  4074 => x"00003f9c",
  4075 => x"00003fa4",
  4076 => x"00003fa4",
  4077 => x"00003fac",
  4078 => x"00003fac",
  4079 => x"00003fb4",
  4080 => x"00003fb4",
  4081 => x"00003fbc",
  4082 => x"00003fbc",
  4083 => x"00003fc4",
  4084 => x"00003fc4",
  4085 => x"00003fcc",
  4086 => x"00003fcc",
  4087 => x"00003fd4",
  4088 => x"00003fd4",
  4089 => x"00003fdc",
  4090 => x"00003fdc",
  4091 => x"00003fe4",
  4092 => x"00003fe4",
  4093 => x"00003fec",
  4094 => x"00003fec",
  4095 => x"00003ff4",
  4096 => x"00003ff4",
  4097 => x"00003ffc",
  4098 => x"00003ffc",
  4099 => x"00004004",
  4100 => x"00004004",
  4101 => x"0000400c",
  4102 => x"0000400c",
  4103 => x"00004014",
  4104 => x"00004014",
  4105 => x"0000401c",
  4106 => x"0000401c",
  4107 => x"00004024",
  4108 => x"00004024",
  4109 => x"0000402c",
  4110 => x"0000402c",
  4111 => x"00004034",
  4112 => x"00004034",
  4113 => x"0000403c",
  4114 => x"0000403c",
  4115 => x"00004044",
  4116 => x"00004044",
  4117 => x"0000404c",
  4118 => x"0000404c",
  4119 => x"00004054",
  4120 => x"00004054",
  4121 => x"0000405c",
  4122 => x"0000405c",
  4123 => x"00004064",
  4124 => x"00004064",
  4125 => x"0000406c",
  4126 => x"0000406c",
  4127 => x"00004074",
  4128 => x"00004074",
  4129 => x"0000407c",
  4130 => x"0000407c",
  4131 => x"00004084",
  4132 => x"00004084",
  4133 => x"0000408c",
  4134 => x"0000408c",
  4135 => x"00004094",
  4136 => x"00004094",
  4137 => x"0000409c",
  4138 => x"0000409c",
  4139 => x"000040a4",
  4140 => x"000040a4",
  4141 => x"000040ac",
  4142 => x"000040ac",
  4143 => x"000040b4",
  4144 => x"000040b4",
  4145 => x"000040bc",
  4146 => x"000040bc",
  4147 => x"000040c4",
  4148 => x"000040c4",
  4149 => x"000040cc",
  4150 => x"000040cc",
  4151 => x"000040d4",
  4152 => x"000040d4",
  4153 => x"000040dc",
  4154 => x"000040dc",
  4155 => x"000040e4",
  4156 => x"000040e4",
  4157 => x"000040ec",
  4158 => x"000040ec",
  4159 => x"000040f4",
  4160 => x"000040f4",
  4161 => x"000040fc",
  4162 => x"000040fc",
  4163 => x"00004104",
  4164 => x"00004104",
  4165 => x"0000410c",
  4166 => x"0000410c",
  4167 => x"00004114",
  4168 => x"00004114",
  4169 => x"0000411c",
  4170 => x"0000411c",
  4171 => x"00004124",
  4172 => x"00004124",
  4173 => x"0000412c",
  4174 => x"0000412c",
  4175 => x"00004134",
  4176 => x"00004134",
  4177 => x"0000413c",
  4178 => x"0000413c",
  4179 => x"00004144",
  4180 => x"00004144",
  4181 => x"0000414c",
  4182 => x"0000414c",
  4183 => x"00004154",
  4184 => x"00004154",
  4185 => x"0000415c",
  4186 => x"0000415c",
  4187 => x"00004164",
  4188 => x"00004164",
  4189 => x"0000416c",
  4190 => x"0000416c",
  4191 => x"00004174",
  4192 => x"00004174",
  4193 => x"0000417c",
  4194 => x"0000417c",
  4195 => x"00004184",
  4196 => x"00004184",
  4197 => x"0000418c",
  4198 => x"0000418c",
  4199 => x"00004194",
  4200 => x"00004194",
  4201 => x"0000419c",
  4202 => x"0000419c",
  4203 => x"000041a4",
  4204 => x"000041a4",
  4205 => x"000041ac",
  4206 => x"000041ac",
  4207 => x"000041b4",
  4208 => x"000041b4",
  4209 => x"000041bc",
  4210 => x"000041bc",
  4211 => x"000041c4",
  4212 => x"000041c4",
  4213 => x"000041cc",
  4214 => x"000041cc",
  4215 => x"000041d4",
  4216 => x"000041d4",
  4217 => x"000041dc",
  4218 => x"000041dc",
  4219 => x"000041e4",
  4220 => x"000041e4",
  4221 => x"000041ec",
  4222 => x"000041ec",
  4223 => x"000041f4",
  4224 => x"000041f4",
  4225 => x"000041fc",
  4226 => x"000041fc",
  4227 => x"00004204",
  4228 => x"00004204",
  4229 => x"0000420c",
  4230 => x"0000420c",
  4231 => x"00004214",
  4232 => x"00004214",
  4233 => x"0000421c",
  4234 => x"0000421c",
	others => x"00dead00" -- mask for mem check
	--others => x"00000000"
);

begin

-- port A
process
begin
    wait until rising_edge( clk);

    -- check 
    if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
        report "write collision" severity failure;
    end if;

    if memAWriteEnable = '1' then
        ram( to_integer( unsigned( memAAddr))) := memAWrite;
        memARead <= memAWrite;
    else
        memARead <= ram( to_integer( unsigned( memAAddr)));
    end if;

end process;


-- port B
process
begin
    wait until rising_edge( clk);

    if memBWriteEnable = '1' then
        ram( to_integer( unsigned( memBAddr))) := memBWrite;
        memBRead <= memBWrite;
    else
        memBRead <= ram(to_integer(unsigned(memBAddr)));
    end if;

end process;




end dualport_ram_arch;
