-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0b92e80c",
     3 => x"3a0b0b0b",
     4 => x"90af0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b90ef2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b92",
   162 => x"d4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b8c",
   171 => x"b32d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b8d",
   179 => x"e52d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0b92e40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f8a",
   257 => x"8f3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"53510492",
   280 => x"e408802e",
   281 => x"a13892e8",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"9a980c82",
   286 => x"a0800b9a",
   287 => x"9c0c8290",
   288 => x"800b9aa0",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0b9a",
   292 => x"980cf880",
   293 => x"8082800b",
   294 => x"9a9c0cf8",
   295 => x"80808480",
   296 => x"0b9aa00c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0b9a98",
   300 => x"0c80c0a8",
   301 => x"80940b9a",
   302 => x"9c0c0b0b",
   303 => x"0b92c00b",
   304 => x"9aa00c04",
   305 => x"ff3d0d9a",
   306 => x"a4335170",
   307 => x"a33892f0",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"92f00c70",
   312 => x"2d92f008",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0b9aa434",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0b9a",
   319 => x"9408802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0b9a94",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"fd3d0d92",
   330 => x"f80876b0",
   331 => x"ea299412",
   332 => x"0c54850b",
   333 => x"98150c98",
   334 => x"14087081",
   335 => x"06515372",
   336 => x"f638853d",
   337 => x"0d04ff3d",
   338 => x"0d92f808",
   339 => x"74101075",
   340 => x"10059412",
   341 => x"0c52850b",
   342 => x"98130c98",
   343 => x"12087081",
   344 => x"06515170",
   345 => x"f638833d",
   346 => x"0d04803d",
   347 => x"0d725180",
   348 => x"71278738",
   349 => x"ff115170",
   350 => x"fb38823d",
   351 => x"0d04803d",
   352 => x"0d92f808",
   353 => x"51870b84",
   354 => x"120c823d",
   355 => x"0d04803d",
   356 => x"0d92f408",
   357 => x"5181ff0b",
   358 => x"88120c82",
   359 => x"3d0d04fb",
   360 => x"3d0d8880",
   361 => x"e0870b92",
   362 => x"f40892f8",
   363 => x"08728413",
   364 => x"0c565755",
   365 => x"afd7c20b",
   366 => x"94150c85",
   367 => x"0b98150c",
   368 => x"98140870",
   369 => x"81065153",
   370 => x"72f63874",
   371 => x"9f2a7510",
   372 => x"07708418",
   373 => x"0c55afd7",
   374 => x"c20b9415",
   375 => x"0c850b98",
   376 => x"150cdd39",
   377 => x"fb3d0d92",
   378 => x"f8085487",
   379 => x"0b84150c",
   380 => x"92f40856",
   381 => x"81ff0b88",
   382 => x"170c8880",
   383 => x"e0877084",
   384 => x"180c55af",
   385 => x"d7c20b94",
   386 => x"150c850b",
   387 => x"98150c98",
   388 => x"14087081",
   389 => x"06515372",
   390 => x"f638749f",
   391 => x"2a751007",
   392 => x"7084180c",
   393 => x"55afd7c2",
   394 => x"0b94150c",
   395 => x"850b9815",
   396 => x"0cdd398c",
   397 => x"08028c0c",
   398 => x"f93d0d80",
   399 => x"0b8c08fc",
   400 => x"050c8c08",
   401 => x"88050880",
   402 => x"25ab388c",
   403 => x"08880508",
   404 => x"308c0888",
   405 => x"050c800b",
   406 => x"8c08f405",
   407 => x"0c8c08fc",
   408 => x"05088838",
   409 => x"810b8c08",
   410 => x"f4050c8c",
   411 => x"08f40508",
   412 => x"8c08fc05",
   413 => x"0c8c088c",
   414 => x"05088025",
   415 => x"ab388c08",
   416 => x"8c050830",
   417 => x"8c088c05",
   418 => x"0c800b8c",
   419 => x"08f0050c",
   420 => x"8c08fc05",
   421 => x"08883881",
   422 => x"0b8c08f0",
   423 => x"050c8c08",
   424 => x"f005088c",
   425 => x"08fc050c",
   426 => x"80538c08",
   427 => x"8c050852",
   428 => x"8c088805",
   429 => x"085181a7",
   430 => x"3f800870",
   431 => x"8c08f805",
   432 => x"0c548c08",
   433 => x"fc050880",
   434 => x"2e8c388c",
   435 => x"08f80508",
   436 => x"308c08f8",
   437 => x"050c8c08",
   438 => x"f8050870",
   439 => x"800c5489",
   440 => x"3d0d8c0c",
   441 => x"048c0802",
   442 => x"8c0cfb3d",
   443 => x"0d800b8c",
   444 => x"08fc050c",
   445 => x"8c088805",
   446 => x"08802593",
   447 => x"388c0888",
   448 => x"0508308c",
   449 => x"0888050c",
   450 => x"810b8c08",
   451 => x"fc050c8c",
   452 => x"088c0508",
   453 => x"80258c38",
   454 => x"8c088c05",
   455 => x"08308c08",
   456 => x"8c050c81",
   457 => x"538c088c",
   458 => x"0508528c",
   459 => x"08880508",
   460 => x"51ad3f80",
   461 => x"08708c08",
   462 => x"f8050c54",
   463 => x"8c08fc05",
   464 => x"08802e8c",
   465 => x"388c08f8",
   466 => x"0508308c",
   467 => x"08f8050c",
   468 => x"8c08f805",
   469 => x"0870800c",
   470 => x"54873d0d",
   471 => x"8c0c048c",
   472 => x"08028c0c",
   473 => x"fd3d0d81",
   474 => x"0b8c08fc",
   475 => x"050c800b",
   476 => x"8c08f805",
   477 => x"0c8c088c",
   478 => x"05088c08",
   479 => x"88050827",
   480 => x"ac388c08",
   481 => x"fc050880",
   482 => x"2ea33880",
   483 => x"0b8c088c",
   484 => x"05082499",
   485 => x"388c088c",
   486 => x"0508108c",
   487 => x"088c050c",
   488 => x"8c08fc05",
   489 => x"08108c08",
   490 => x"fc050cc9",
   491 => x"398c08fc",
   492 => x"0508802e",
   493 => x"80c9388c",
   494 => x"088c0508",
   495 => x"8c088805",
   496 => x"0826a138",
   497 => x"8c088805",
   498 => x"088c088c",
   499 => x"0508318c",
   500 => x"0888050c",
   501 => x"8c08f805",
   502 => x"088c08fc",
   503 => x"0508078c",
   504 => x"08f8050c",
   505 => x"8c08fc05",
   506 => x"08812a8c",
   507 => x"08fc050c",
   508 => x"8c088c05",
   509 => x"08812a8c",
   510 => x"088c050c",
   511 => x"ffaf398c",
   512 => x"08900508",
   513 => x"802e8f38",
   514 => x"8c088805",
   515 => x"08708c08",
   516 => x"f4050c51",
   517 => x"8d398c08",
   518 => x"f8050870",
   519 => x"8c08f405",
   520 => x"0c518c08",
   521 => x"f4050880",
   522 => x"0c853d0d",
   523 => x"8c0c04fd",
   524 => x"3d0d800b",
   525 => x"92e80854",
   526 => x"5472812e",
   527 => x"9838739a",
   528 => x"a80cf89b",
   529 => x"3ff7b93f",
   530 => x"93805281",
   531 => x"51fb953f",
   532 => x"8008519e",
   533 => x"3f729aa8",
   534 => x"0cf8843f",
   535 => x"f7a23f93",
   536 => x"80528151",
   537 => x"fafe3f80",
   538 => x"0851873f",
   539 => x"00ff3900",
   540 => x"ff39f73d",
   541 => x"0d7b9384",
   542 => x"0882c811",
   543 => x"085a545a",
   544 => x"77802e80",
   545 => x"d9388188",
   546 => x"18841908",
   547 => x"ff058171",
   548 => x"2b595559",
   549 => x"80742480",
   550 => x"e9388074",
   551 => x"24b53873",
   552 => x"822b7811",
   553 => x"88055656",
   554 => x"81801908",
   555 => x"77065372",
   556 => x"802eb538",
   557 => x"78167008",
   558 => x"53537951",
   559 => x"74085372",
   560 => x"2dff14fc",
   561 => x"17fc1779",
   562 => x"812c5a57",
   563 => x"57547380",
   564 => x"25d63877",
   565 => x"085877ff",
   566 => x"ad389384",
   567 => x"0853bc13",
   568 => x"08a53879",
   569 => x"51ff853f",
   570 => x"74085372",
   571 => x"2dff14fc",
   572 => x"17fc1779",
   573 => x"812c5a57",
   574 => x"57547380",
   575 => x"25ffa938",
   576 => x"d2398057",
   577 => x"ff943972",
   578 => x"51bc1308",
   579 => x"53722d79",
   580 => x"51fed93f",
   581 => x"ff3d0d9a",
   582 => x"880bfc05",
   583 => x"70085252",
   584 => x"70ff2e91",
   585 => x"38702dfc",
   586 => x"12700852",
   587 => x"5270ff2e",
   588 => x"098106f1",
   589 => x"38833d0d",
   590 => x"0404f788",
   591 => x"3f040000",
   592 => x"00000040",
   593 => x"64756d6d",
   594 => x"792e6578",
   595 => x"65000000",
   596 => x"43000000",
   597 => x"00ffffff",
   598 => x"ff00ffff",
   599 => x"ffff00ff",
   600 => x"ffffff00",
   601 => x"00000000",
   602 => x"00000000",
   603 => x"00000000",
   604 => x"00000d10",
   605 => x"80000800",
   606 => x"80000200",
   607 => x"80000100",
   608 => x"00000944",
   609 => x"00000988",
   610 => x"00000000",
   611 => x"00000bf0",
   612 => x"00000c4c",
   613 => x"00000ca8",
   614 => x"00000000",
   615 => x"00000000",
   616 => x"00000000",
   617 => x"00000000",
   618 => x"00000000",
   619 => x"00000000",
   620 => x"00000000",
   621 => x"00000000",
   622 => x"00000000",
   623 => x"00000950",
   624 => x"00000000",
   625 => x"00000000",
   626 => x"00000000",
   627 => x"00000000",
   628 => x"00000000",
   629 => x"00000000",
   630 => x"00000000",
   631 => x"00000000",
   632 => x"00000000",
   633 => x"00000000",
   634 => x"00000000",
   635 => x"00000000",
   636 => x"00000000",
   637 => x"00000000",
   638 => x"00000000",
   639 => x"00000000",
   640 => x"00000000",
   641 => x"00000000",
   642 => x"00000000",
   643 => x"00000000",
   644 => x"00000000",
   645 => x"00000000",
   646 => x"00000000",
   647 => x"00000000",
   648 => x"00000000",
   649 => x"00000000",
   650 => x"00000000",
   651 => x"00000000",
   652 => x"00000001",
   653 => x"330eabcd",
   654 => x"1234e66d",
   655 => x"deec0005",
   656 => x"000b0000",
   657 => x"00000000",
   658 => x"00000000",
   659 => x"00000000",
   660 => x"00000000",
   661 => x"00000000",
   662 => x"00000000",
   663 => x"00000000",
   664 => x"00000000",
   665 => x"00000000",
   666 => x"00000000",
   667 => x"00000000",
   668 => x"00000000",
   669 => x"00000000",
   670 => x"00000000",
   671 => x"00000000",
   672 => x"00000000",
   673 => x"00000000",
   674 => x"00000000",
   675 => x"00000000",
   676 => x"00000000",
   677 => x"00000000",
   678 => x"00000000",
   679 => x"00000000",
   680 => x"00000000",
   681 => x"00000000",
   682 => x"00000000",
   683 => x"00000000",
   684 => x"00000000",
   685 => x"00000000",
   686 => x"00000000",
   687 => x"00000000",
   688 => x"00000000",
   689 => x"00000000",
   690 => x"00000000",
   691 => x"00000000",
   692 => x"00000000",
   693 => x"00000000",
   694 => x"00000000",
   695 => x"00000000",
   696 => x"00000000",
   697 => x"00000000",
   698 => x"00000000",
   699 => x"00000000",
   700 => x"00000000",
   701 => x"00000000",
   702 => x"00000000",
   703 => x"00000000",
   704 => x"00000000",
   705 => x"00000000",
   706 => x"00000000",
   707 => x"00000000",
   708 => x"00000000",
   709 => x"00000000",
   710 => x"00000000",
   711 => x"00000000",
   712 => x"00000000",
   713 => x"00000000",
   714 => x"00000000",
   715 => x"00000000",
   716 => x"00000000",
   717 => x"00000000",
   718 => x"00000000",
   719 => x"00000000",
   720 => x"00000000",
   721 => x"00000000",
   722 => x"00000000",
   723 => x"00000000",
   724 => x"00000000",
   725 => x"00000000",
   726 => x"00000000",
   727 => x"00000000",
   728 => x"00000000",
   729 => x"00000000",
   730 => x"00000000",
   731 => x"00000000",
   732 => x"00000000",
   733 => x"00000000",
   734 => x"00000000",
   735 => x"00000000",
   736 => x"00000000",
   737 => x"00000000",
   738 => x"00000000",
   739 => x"00000000",
   740 => x"00000000",
   741 => x"00000000",
   742 => x"00000000",
   743 => x"00000000",
   744 => x"00000000",
   745 => x"00000000",
   746 => x"00000000",
   747 => x"00000000",
   748 => x"00000000",
   749 => x"00000000",
   750 => x"00000000",
   751 => x"00000000",
   752 => x"00000000",
   753 => x"00000000",
   754 => x"00000000",
   755 => x"00000000",
   756 => x"00000000",
   757 => x"00000000",
   758 => x"00000000",
   759 => x"00000000",
   760 => x"00000000",
   761 => x"00000000",
   762 => x"00000000",
   763 => x"00000000",
   764 => x"00000000",
   765 => x"00000000",
   766 => x"00000000",
   767 => x"00000000",
   768 => x"00000000",
   769 => x"00000000",
   770 => x"00000000",
   771 => x"00000000",
   772 => x"00000000",
   773 => x"00000000",
   774 => x"00000000",
   775 => x"00000000",
   776 => x"00000000",
   777 => x"00000000",
   778 => x"00000000",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000000",
   783 => x"00000000",
   784 => x"00000000",
   785 => x"00000000",
   786 => x"00000000",
   787 => x"00000000",
   788 => x"00000000",
   789 => x"00000000",
   790 => x"00000000",
   791 => x"00000000",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
   799 => x"00000000",
   800 => x"00000000",
   801 => x"00000000",
   802 => x"00000000",
   803 => x"00000000",
   804 => x"00000000",
   805 => x"00000000",
   806 => x"00000000",
   807 => x"00000000",
   808 => x"00000000",
   809 => x"00000000",
   810 => x"00000000",
   811 => x"00000000",
   812 => x"00000000",
   813 => x"00000000",
   814 => x"00000000",
   815 => x"00000000",
   816 => x"00000000",
   817 => x"00000000",
   818 => x"00000000",
   819 => x"00000000",
   820 => x"00000000",
   821 => x"00000000",
   822 => x"00000000",
   823 => x"00000000",
   824 => x"00000000",
   825 => x"00000000",
   826 => x"00000000",
   827 => x"00000000",
   828 => x"00000000",
   829 => x"00000000",
   830 => x"00000000",
   831 => x"00000000",
   832 => x"00000000",
   833 => x"ffffffff",
   834 => x"00000000",
   835 => x"ffffffff",
   836 => x"00000000",
   837 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
