-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80e0f40c",
     3 => x"3a0b0b80",
     4 => x"d9f40400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80dabd2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80e0",
   162 => x"e0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0bbd",
   171 => x"db2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bbf",
   179 => x"8d2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80e0f00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"d3de3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80e0f008",
   281 => x"802ea438",
   282 => x"80e0f408",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80f0",
   286 => x"ec0c82a0",
   287 => x"800b80f0",
   288 => x"f00c8290",
   289 => x"800b80f0",
   290 => x"f40c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"f0ec0cf8",
   294 => x"80808280",
   295 => x"0b80f0f0",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"f0f40c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80f0ec0c",
   302 => x"80c0a880",
   303 => x"940b80f0",
   304 => x"f00c0b0b",
   305 => x"80dc900b",
   306 => x"80f0f40c",
   307 => x"04ff3d0d",
   308 => x"80f0f833",
   309 => x"5170a738",
   310 => x"80e0fc08",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"e0fc0c70",
   315 => x"2d80e0fc",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80f0",
   319 => x"f834833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80f0e808",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"f0e8510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404fd3d",
   333 => x"0d80e188",
   334 => x"0876b0ea",
   335 => x"2994120c",
   336 => x"54850b98",
   337 => x"150c9814",
   338 => x"08708106",
   339 => x"515372f6",
   340 => x"38853d0d",
   341 => x"04ff3d0d",
   342 => x"80e18808",
   343 => x"74101075",
   344 => x"10059412",
   345 => x"0c52850b",
   346 => x"98130c98",
   347 => x"12087081",
   348 => x"06515170",
   349 => x"f638833d",
   350 => x"0d04803d",
   351 => x"0d725180",
   352 => x"71278738",
   353 => x"ff115170",
   354 => x"fb38823d",
   355 => x"0d04803d",
   356 => x"0d80e188",
   357 => x"0851870b",
   358 => x"84120c82",
   359 => x"3d0d0480",
   360 => x"3d0d80e1",
   361 => x"8c0851b6",
   362 => x"0b8c120c",
   363 => x"830b8812",
   364 => x"0c823d0d",
   365 => x"04ff3d0d",
   366 => x"80e18c08",
   367 => x"52841208",
   368 => x"70810651",
   369 => x"5170802e",
   370 => x"f4387108",
   371 => x"7081ff06",
   372 => x"800c5183",
   373 => x"3d0d04fe",
   374 => x"3d0d0293",
   375 => x"053380e1",
   376 => x"8c085353",
   377 => x"84120870",
   378 => x"892a7081",
   379 => x"06515151",
   380 => x"70f23872",
   381 => x"720c843d",
   382 => x"0d04fe3d",
   383 => x"0d029305",
   384 => x"3353728a",
   385 => x"2e9c3880",
   386 => x"e18c0852",
   387 => x"84120870",
   388 => x"892a7081",
   389 => x"06515151",
   390 => x"70f23872",
   391 => x"720c843d",
   392 => x"0d0480e1",
   393 => x"8c085284",
   394 => x"12087089",
   395 => x"2a708106",
   396 => x"51515170",
   397 => x"f2388d72",
   398 => x"0c841208",
   399 => x"70892a70",
   400 => x"81065151",
   401 => x"5170c538",
   402 => x"d239fd3d",
   403 => x"0d757033",
   404 => x"52547080",
   405 => x"2ea83870",
   406 => x"80e18c08",
   407 => x"53538114",
   408 => x"54728a2e",
   409 => x"9d388412",
   410 => x"0870892a",
   411 => x"70810651",
   412 => x"515170f2",
   413 => x"3872720c",
   414 => x"73335372",
   415 => x"e138853d",
   416 => x"0d048412",
   417 => x"0870892a",
   418 => x"70810651",
   419 => x"515170f2",
   420 => x"388d720c",
   421 => x"84120870",
   422 => x"892a7081",
   423 => x"06515151",
   424 => x"70c438d1",
   425 => x"39f53d0d",
   426 => x"7e028405",
   427 => x"b705338c",
   428 => x"3d5b5557",
   429 => x"8b5380dc",
   430 => x"94527851",
   431 => x"b4a63f82",
   432 => x"5673882e",
   433 => x"96388456",
   434 => x"73902e8f",
   435 => x"38885673",
   436 => x"a02e8838",
   437 => x"74567480",
   438 => x"2ea73802",
   439 => x"a5055876",
   440 => x"8f065473",
   441 => x"892680cc",
   442 => x"387518b0",
   443 => x"15555573",
   444 => x"75347684",
   445 => x"2aff1770",
   446 => x"81ff0658",
   447 => x"555775df",
   448 => x"38787933",
   449 => x"55577380",
   450 => x"2ea63873",
   451 => x"80e18c08",
   452 => x"56568117",
   453 => x"57758a2e",
   454 => x"b7388415",
   455 => x"0870892a",
   456 => x"81065954",
   457 => x"77f43875",
   458 => x"750c7633",
   459 => x"5675e338",
   460 => x"8d3d0d04",
   461 => x"7518b715",
   462 => x"55557375",
   463 => x"3476842a",
   464 => x"ff177081",
   465 => x"ff065855",
   466 => x"5775ff93",
   467 => x"38ffb239",
   468 => x"84150870",
   469 => x"892a8106",
   470 => x"595477f4",
   471 => x"388d750c",
   472 => x"84150870",
   473 => x"892a8106",
   474 => x"595477ff",
   475 => x"ad38ffb7",
   476 => x"39f83d0d",
   477 => x"7a7c5953",
   478 => x"80735657",
   479 => x"76732480",
   480 => x"dc387717",
   481 => x"548a5274",
   482 => x"51aeab3f",
   483 => x"8008b005",
   484 => x"53727434",
   485 => x"8117578a",
   486 => x"527451ad",
   487 => x"f43f8008",
   488 => x"558008de",
   489 => x"38800877",
   490 => x"9f2a1870",
   491 => x"812c5b56",
   492 => x"56807925",
   493 => x"9e387717",
   494 => x"ff055575",
   495 => x"18703355",
   496 => x"53743373",
   497 => x"34737534",
   498 => x"8116ff16",
   499 => x"56567876",
   500 => x"24e93876",
   501 => x"18568076",
   502 => x"348a3d0d",
   503 => x"04ad7870",
   504 => x"81055a34",
   505 => x"72307818",
   506 => x"55558a52",
   507 => x"7451adc6",
   508 => x"3f8008b0",
   509 => x"05537274",
   510 => x"34811757",
   511 => x"8a527451",
   512 => x"ad8f3f80",
   513 => x"08558008",
   514 => x"fef838ff",
   515 => x"9839803d",
   516 => x"0d80e184",
   517 => x"085181ff",
   518 => x"0b88120c",
   519 => x"823d0d04",
   520 => x"f83d0d7a",
   521 => x"59f881c0",
   522 => x"8e8055a0",
   523 => x"0b80e184",
   524 => x"0880e188",
   525 => x"085a5856",
   526 => x"7484180c",
   527 => x"749f2a75",
   528 => x"10075578",
   529 => x"802e9738",
   530 => x"75802ebb",
   531 => x"38ff1675",
   532 => x"84190c75",
   533 => x"9f2a7610",
   534 => x"07565678",
   535 => x"eb387754",
   536 => x"afd7c20b",
   537 => x"94190c85",
   538 => x"0b98190c",
   539 => x"98140870",
   540 => x"81065153",
   541 => x"72802ec0",
   542 => x"38981408",
   543 => x"70810651",
   544 => x"5372e938",
   545 => x"ffb2398a",
   546 => x"3d0d04fd",
   547 => x"3d0d80e1",
   548 => x"84085480",
   549 => x"d50b8415",
   550 => x"0c80e18c",
   551 => x"08528412",
   552 => x"08810651",
   553 => x"70802ef6",
   554 => x"38710870",
   555 => x"81ff06f6",
   556 => x"11525451",
   557 => x"70ae268c",
   558 => x"38701010",
   559 => x"80df9405",
   560 => x"51700804",
   561 => x"84120870",
   562 => x"892a7081",
   563 => x"06515151",
   564 => x"70f238ab",
   565 => x"720c728a",
   566 => x"2ea63884",
   567 => x"12087089",
   568 => x"2a708106",
   569 => x"51515170",
   570 => x"f2387272",
   571 => x"0c841208",
   572 => x"70892a81",
   573 => x"06515372",
   574 => x"f438ad72",
   575 => x"0cff9f39",
   576 => x"84120870",
   577 => x"892a7081",
   578 => x"06515151",
   579 => x"70f2388d",
   580 => x"720c8412",
   581 => x"0870892a",
   582 => x"70810651",
   583 => x"515170ff",
   584 => x"ba38c739",
   585 => x"81ff0b84",
   586 => x"150cfef2",
   587 => x"3980ff0b",
   588 => x"84150cfe",
   589 => x"e939bf0b",
   590 => x"84150cfe",
   591 => x"e1399f0b",
   592 => x"84150cfe",
   593 => x"d9398f0b",
   594 => x"84150cfe",
   595 => x"d139870b",
   596 => x"84150cfe",
   597 => x"c939830b",
   598 => x"84150cfe",
   599 => x"c139810b",
   600 => x"84150cfe",
   601 => x"b939800b",
   602 => x"84150cfe",
   603 => x"b139ff3d",
   604 => x"0d80e184",
   605 => x"08527108",
   606 => x"708f0670",
   607 => x"71842b07",
   608 => x"84150c51",
   609 => x"51710870",
   610 => x"8f067071",
   611 => x"842b0784",
   612 => x"150c5151",
   613 => x"e139fc3d",
   614 => x"0d029a05",
   615 => x"22028405",
   616 => x"9e052202",
   617 => x"8805a205",
   618 => x"2280e180",
   619 => x"08555654",
   620 => x"55901208",
   621 => x"70832a70",
   622 => x"81065151",
   623 => x"5170f238",
   624 => x"74902b73",
   625 => x"8b2b0774",
   626 => x"862b0781",
   627 => x"0790130c",
   628 => x"863d0d04",
   629 => x"fd3d0d02",
   630 => x"96052202",
   631 => x"84059a05",
   632 => x"2280e180",
   633 => x"08545454",
   634 => x"90120870",
   635 => x"832a7081",
   636 => x"06515151",
   637 => x"70f23873",
   638 => x"8b2b7386",
   639 => x"2b078207",
   640 => x"90130c90",
   641 => x"12087083",
   642 => x"2a810655",
   643 => x"5173f438",
   644 => x"90120870",
   645 => x"902a800c",
   646 => x"54853d0d",
   647 => x"04ff3d0d",
   648 => x"80e18008",
   649 => x"52ff0b84",
   650 => x"130cfc94",
   651 => x"800b8813",
   652 => x"0c82d0af",
   653 => x"fdfb0b8c",
   654 => x"130c80c0",
   655 => x"720c7108",
   656 => x"70862a70",
   657 => x"81065151",
   658 => x"5170f338",
   659 => x"90120870",
   660 => x"832a7081",
   661 => x"06515151",
   662 => x"70f23881",
   663 => x"fc80810b",
   664 => x"90130c90",
   665 => x"12087083",
   666 => x"2a708106",
   667 => x"51515170",
   668 => x"f23880fd",
   669 => x"c0810b90",
   670 => x"130c833d",
   671 => x"0d04d53d",
   672 => x"0d80e180",
   673 => x"0858ff0b",
   674 => x"84190cfc",
   675 => x"809b0b88",
   676 => x"190c828b",
   677 => x"a1968a0b",
   678 => x"8c190ca4",
   679 => x"b40b9419",
   680 => x"0c8186a1",
   681 => x"0b98190c",
   682 => x"80dca00b",
   683 => x"80dca033",
   684 => x"55577380",
   685 => x"2ea73873",
   686 => x"80e18c08",
   687 => x"56568117",
   688 => x"57758a2e",
   689 => x"8db93884",
   690 => x"15087089",
   691 => x"2a810651",
   692 => x"5978f438",
   693 => x"75750c76",
   694 => x"335675e2",
   695 => x"3880dcb4",
   696 => x"0b80dcb4",
   697 => x"33555773",
   698 => x"802ea738",
   699 => x"80e18c08",
   700 => x"74575581",
   701 => x"1757758a",
   702 => x"2e8da538",
   703 => x"84150870",
   704 => x"892a8106",
   705 => x"515978f4",
   706 => x"3875750c",
   707 => x"76335675",
   708 => x"e2387708",
   709 => x"a63d5a56",
   710 => x"8b5380dc",
   711 => x"94527851",
   712 => x"abc23f88",
   713 => x"02840581",
   714 => x"91055957",
   715 => x"758f0654",
   716 => x"7389268d",
   717 => x"8c387618",
   718 => x"b0155555",
   719 => x"73753475",
   720 => x"842aff18",
   721 => x"7081ff06",
   722 => x"59565676",
   723 => x"df387879",
   724 => x"33555773",
   725 => x"802ea738",
   726 => x"80e18c08",
   727 => x"74575581",
   728 => x"1757758a",
   729 => x"2e8cf638",
   730 => x"84150870",
   731 => x"892a8106",
   732 => x"595977f4",
   733 => x"3875750c",
   734 => x"76335675",
   735 => x"e23880dc",
   736 => x"c40b80dc",
   737 => x"c4335557",
   738 => x"73802ea7",
   739 => x"3880e18c",
   740 => x"08745755",
   741 => x"81175775",
   742 => x"8a2e8ce2",
   743 => x"38841508",
   744 => x"70892a81",
   745 => x"06595977",
   746 => x"f4387575",
   747 => x"0c763356",
   748 => x"75e23880",
   749 => x"e1800884",
   750 => x"1108a43d",
   751 => x"5b57578b",
   752 => x"5380dc94",
   753 => x"527851aa",
   754 => x"9b3f8802",
   755 => x"84058185",
   756 => x"05595775",
   757 => x"8f065473",
   758 => x"892691bc",
   759 => x"387618b0",
   760 => x"15555573",
   761 => x"75347584",
   762 => x"2aff1870",
   763 => x"81ff0659",
   764 => x"565676df",
   765 => x"38787933",
   766 => x"55577380",
   767 => x"2ea73880",
   768 => x"e18c0874",
   769 => x"57558117",
   770 => x"57758a2e",
   771 => x"8c913884",
   772 => x"15087089",
   773 => x"2a810659",
   774 => x"5977f438",
   775 => x"75750c76",
   776 => x"335675e2",
   777 => x"3880dcd4",
   778 => x"0b80dcd4",
   779 => x"33555773",
   780 => x"802ea738",
   781 => x"80e18c08",
   782 => x"74575581",
   783 => x"1757758a",
   784 => x"2e8bfd38",
   785 => x"84150870",
   786 => x"892a8106",
   787 => x"595977f4",
   788 => x"3875750c",
   789 => x"76335675",
   790 => x"e23880e1",
   791 => x"80088811",
   792 => x"08a13d5b",
   793 => x"57578b53",
   794 => x"80dc9452",
   795 => x"7851a8f4",
   796 => x"3f880284",
   797 => x"0580f905",
   798 => x"5957758f",
   799 => x"06547389",
   800 => x"26908c38",
   801 => x"7618b015",
   802 => x"55557375",
   803 => x"3475842a",
   804 => x"ff187081",
   805 => x"ff065956",
   806 => x"5676df38",
   807 => x"78793355",
   808 => x"5773802e",
   809 => x"a73880e1",
   810 => x"8c087457",
   811 => x"55811757",
   812 => x"758a2e8b",
   813 => x"ac388415",
   814 => x"0870892a",
   815 => x"81065959",
   816 => x"77f43875",
   817 => x"750c7633",
   818 => x"5675e238",
   819 => x"80dce40b",
   820 => x"80dce433",
   821 => x"55577380",
   822 => x"2ea73880",
   823 => x"e18c0874",
   824 => x"57558117",
   825 => x"57758a2e",
   826 => x"8b983884",
   827 => x"15087089",
   828 => x"2a810659",
   829 => x"5977f438",
   830 => x"75750c76",
   831 => x"335675e2",
   832 => x"3880e180",
   833 => x"088c1108",
   834 => x"9e3d5b57",
   835 => x"578b5380",
   836 => x"dc945278",
   837 => x"51a7cd3f",
   838 => x"88028405",
   839 => x"80ed0559",
   840 => x"57758f06",
   841 => x"54738926",
   842 => x"8edc3876",
   843 => x"18b01555",
   844 => x"55737534",
   845 => x"75842aff",
   846 => x"187081ff",
   847 => x"06595656",
   848 => x"76df3878",
   849 => x"79335557",
   850 => x"73802ea7",
   851 => x"3880e18c",
   852 => x"08745755",
   853 => x"81175775",
   854 => x"8a2e8ac7",
   855 => x"38841508",
   856 => x"70892a81",
   857 => x"06595977",
   858 => x"f4387575",
   859 => x"0c763356",
   860 => x"75e23880",
   861 => x"dcf40b80",
   862 => x"dcf43355",
   863 => x"5773802e",
   864 => x"a73880e1",
   865 => x"8c087457",
   866 => x"55811757",
   867 => x"758a2e8a",
   868 => x"b3388415",
   869 => x"0870892a",
   870 => x"81065959",
   871 => x"77f43875",
   872 => x"750c7633",
   873 => x"5675e238",
   874 => x"80e18008",
   875 => x"9011089b",
   876 => x"3d5b5757",
   877 => x"8b5380dc",
   878 => x"94527851",
   879 => x"a6a63f88",
   880 => x"02840580",
   881 => x"e1055957",
   882 => x"758f0654",
   883 => x"7389268d",
   884 => x"ac387618",
   885 => x"b0155555",
   886 => x"73753475",
   887 => x"842aff18",
   888 => x"7081ff06",
   889 => x"59565676",
   890 => x"df387879",
   891 => x"33555773",
   892 => x"802ea738",
   893 => x"80e18c08",
   894 => x"74575581",
   895 => x"1757758a",
   896 => x"2e89e238",
   897 => x"84150870",
   898 => x"892a8106",
   899 => x"595977f4",
   900 => x"3875750c",
   901 => x"76335675",
   902 => x"e23880dd",
   903 => x"840b80dd",
   904 => x"84335557",
   905 => x"73802ea7",
   906 => x"3880e18c",
   907 => x"08745755",
   908 => x"81175775",
   909 => x"8a2e89ce",
   910 => x"38841508",
   911 => x"70892a81",
   912 => x"06595977",
   913 => x"f4387575",
   914 => x"0c763356",
   915 => x"75e23880",
   916 => x"e1800894",
   917 => x"1108983d",
   918 => x"5b57578b",
   919 => x"5380dc94",
   920 => x"527851a4",
   921 => x"ff3f8802",
   922 => x"840580d5",
   923 => x"05595775",
   924 => x"8f065473",
   925 => x"89268bfc",
   926 => x"387618b0",
   927 => x"15555573",
   928 => x"75347584",
   929 => x"2aff1870",
   930 => x"81ff0659",
   931 => x"565676df",
   932 => x"38787933",
   933 => x"55577380",
   934 => x"2ea73880",
   935 => x"e18c0874",
   936 => x"57558117",
   937 => x"57758a2e",
   938 => x"88fd3884",
   939 => x"15087089",
   940 => x"2a810659",
   941 => x"5977f438",
   942 => x"75750c76",
   943 => x"335675e2",
   944 => x"3880dd94",
   945 => x"0b80dd94",
   946 => x"33555773",
   947 => x"802ea738",
   948 => x"80e18c08",
   949 => x"74575581",
   950 => x"1757758a",
   951 => x"2e88e938",
   952 => x"84150870",
   953 => x"892a8106",
   954 => x"595977f4",
   955 => x"3875750c",
   956 => x"76335675",
   957 => x"e23880e1",
   958 => x"80089811",
   959 => x"08953d5b",
   960 => x"57578b53",
   961 => x"80dc9452",
   962 => x"7851a3d8",
   963 => x"3f880284",
   964 => x"0580c905",
   965 => x"5957758f",
   966 => x"06547389",
   967 => x"268acc38",
   968 => x"7618b015",
   969 => x"55557375",
   970 => x"3475842a",
   971 => x"ff187081",
   972 => x"ff065956",
   973 => x"5676df38",
   974 => x"78793355",
   975 => x"5773802e",
   976 => x"a73880e1",
   977 => x"8c087457",
   978 => x"55811757",
   979 => x"758a2e88",
   980 => x"98388415",
   981 => x"0870892a",
   982 => x"81065959",
   983 => x"77f43875",
   984 => x"750c7633",
   985 => x"5675e238",
   986 => x"80dda40b",
   987 => x"80dda433",
   988 => x"55577380",
   989 => x"2ea73880",
   990 => x"e18c0874",
   991 => x"57558117",
   992 => x"57758a2e",
   993 => x"88843884",
   994 => x"15087089",
   995 => x"2a810659",
   996 => x"5977f438",
   997 => x"75750c76",
   998 => x"335675e2",
   999 => x"3880e180",
  1000 => x"089c1108",
  1001 => x"923d5b57",
  1002 => x"578b5380",
  1003 => x"dc945278",
  1004 => x"51a2b13f",
  1005 => x"88028405",
  1006 => x"bd055957",
  1007 => x"758f0654",
  1008 => x"73892689",
  1009 => x"9d387618",
  1010 => x"b0155555",
  1011 => x"73753475",
  1012 => x"842aff18",
  1013 => x"7081ff06",
  1014 => x"59565676",
  1015 => x"df387879",
  1016 => x"33555773",
  1017 => x"802ea738",
  1018 => x"80e18c08",
  1019 => x"74575581",
  1020 => x"1757758a",
  1021 => x"2e87b438",
  1022 => x"84150870",
  1023 => x"892a8106",
  1024 => x"595977f4",
  1025 => x"3875750c",
  1026 => x"76335675",
  1027 => x"e23880dd",
  1028 => x"b40b80dd",
  1029 => x"b4335557",
  1030 => x"73802ea7",
  1031 => x"3880e18c",
  1032 => x"08745755",
  1033 => x"81175775",
  1034 => x"8a2e87a0",
  1035 => x"38841508",
  1036 => x"70892a81",
  1037 => x"06595977",
  1038 => x"f4387575",
  1039 => x"0c763356",
  1040 => x"75e23880",
  1041 => x"e18008a0",
  1042 => x"11088f3d",
  1043 => x"5b57578b",
  1044 => x"5380dc94",
  1045 => x"527851a1",
  1046 => x"8b3f8802",
  1047 => x"8405b105",
  1048 => x"5957758f",
  1049 => x"06547389",
  1050 => x"2687ee38",
  1051 => x"7618b015",
  1052 => x"55557375",
  1053 => x"3475842a",
  1054 => x"ff187081",
  1055 => x"ff065956",
  1056 => x"5676df38",
  1057 => x"78793355",
  1058 => x"5773802e",
  1059 => x"a73880e1",
  1060 => x"8c087457",
  1061 => x"55811757",
  1062 => x"758a2e86",
  1063 => x"d0388415",
  1064 => x"0870892a",
  1065 => x"81065959",
  1066 => x"77f43875",
  1067 => x"750c7633",
  1068 => x"5675e238",
  1069 => x"80ddc40b",
  1070 => x"80ddc433",
  1071 => x"55577380",
  1072 => x"2ea73880",
  1073 => x"e18c0874",
  1074 => x"57558117",
  1075 => x"57758a2e",
  1076 => x"86bc3884",
  1077 => x"15087089",
  1078 => x"2a810659",
  1079 => x"5977f438",
  1080 => x"75750c76",
  1081 => x"335675e2",
  1082 => x"3880e180",
  1083 => x"08a41108",
  1084 => x"8c3d5b57",
  1085 => x"578b5380",
  1086 => x"dc945278",
  1087 => x"519fe53f",
  1088 => x"88028405",
  1089 => x"a5055957",
  1090 => x"758f0654",
  1091 => x"73892686",
  1092 => x"bf387618",
  1093 => x"b0155555",
  1094 => x"73753475",
  1095 => x"842aff18",
  1096 => x"7081ff06",
  1097 => x"59565676",
  1098 => x"df387879",
  1099 => x"33555773",
  1100 => x"802e86ed",
  1101 => x"3880e18c",
  1102 => x"08745755",
  1103 => x"81175775",
  1104 => x"8a2e85eb",
  1105 => x"38841508",
  1106 => x"70892a81",
  1107 => x"06595977",
  1108 => x"f4387575",
  1109 => x"0c763356",
  1110 => x"75e23884",
  1111 => x"15087089",
  1112 => x"2a810657",
  1113 => x"5875f438",
  1114 => x"8d750c84",
  1115 => x"15087089",
  1116 => x"2a810655",
  1117 => x"5673f438",
  1118 => x"8a750cad",
  1119 => x"3d0d0484",
  1120 => x"15087089",
  1121 => x"2a810651",
  1122 => x"5473f438",
  1123 => x"8d750c84",
  1124 => x"15087089",
  1125 => x"2a810651",
  1126 => x"5978f2ab",
  1127 => x"38f2b539",
  1128 => x"84150870",
  1129 => x"892a8106",
  1130 => x"515473f4",
  1131 => x"388d750c",
  1132 => x"84150870",
  1133 => x"892a8106",
  1134 => x"515978f2",
  1135 => x"bf38f2c9",
  1136 => x"397618b7",
  1137 => x"15555573",
  1138 => x"75347584",
  1139 => x"2aff1870",
  1140 => x"81ff0659",
  1141 => x"565676f2",
  1142 => x"d338f2f2",
  1143 => x"39841508",
  1144 => x"70892a81",
  1145 => x"06595977",
  1146 => x"f4388d75",
  1147 => x"0c841508",
  1148 => x"70892a81",
  1149 => x"06595977",
  1150 => x"f2ee38f2",
  1151 => x"f8398415",
  1152 => x"0870892a",
  1153 => x"81065959",
  1154 => x"77f4388d",
  1155 => x"750c8415",
  1156 => x"0870892a",
  1157 => x"81065959",
  1158 => x"77f38238",
  1159 => x"f38c3984",
  1160 => x"15087089",
  1161 => x"2a810659",
  1162 => x"5977f438",
  1163 => x"8d750c84",
  1164 => x"15087089",
  1165 => x"2a810659",
  1166 => x"5977f3d3",
  1167 => x"38f3dd39",
  1168 => x"84150870",
  1169 => x"892a8106",
  1170 => x"595977f4",
  1171 => x"388d750c",
  1172 => x"84150870",
  1173 => x"892a8106",
  1174 => x"595977f3",
  1175 => x"e738f3f1",
  1176 => x"39841508",
  1177 => x"70892a81",
  1178 => x"06595977",
  1179 => x"f4388d75",
  1180 => x"0c841508",
  1181 => x"70892a81",
  1182 => x"06595977",
  1183 => x"f4b838f4",
  1184 => x"c2398415",
  1185 => x"0870892a",
  1186 => x"81065959",
  1187 => x"77f4388d",
  1188 => x"750c8415",
  1189 => x"0870892a",
  1190 => x"81065959",
  1191 => x"77f4cc38",
  1192 => x"f4d63984",
  1193 => x"15087089",
  1194 => x"2a810659",
  1195 => x"5977f438",
  1196 => x"8d750c84",
  1197 => x"15087089",
  1198 => x"2a810659",
  1199 => x"5977f59d",
  1200 => x"38f5a739",
  1201 => x"84150870",
  1202 => x"892a8106",
  1203 => x"595977f4",
  1204 => x"388d750c",
  1205 => x"84150870",
  1206 => x"892a8106",
  1207 => x"595977f5",
  1208 => x"b138f5bb",
  1209 => x"39841508",
  1210 => x"70892a81",
  1211 => x"06595977",
  1212 => x"f4388d75",
  1213 => x"0c841508",
  1214 => x"70892a81",
  1215 => x"06595977",
  1216 => x"f68238f6",
  1217 => x"8c398415",
  1218 => x"0870892a",
  1219 => x"81065959",
  1220 => x"77f4388d",
  1221 => x"750c8415",
  1222 => x"0870892a",
  1223 => x"81065959",
  1224 => x"77f69638",
  1225 => x"f6a03984",
  1226 => x"15087089",
  1227 => x"2a810659",
  1228 => x"5977f438",
  1229 => x"8d750c84",
  1230 => x"15087089",
  1231 => x"2a810659",
  1232 => x"5977f6e7",
  1233 => x"38f6f139",
  1234 => x"84150870",
  1235 => x"892a8106",
  1236 => x"595977f4",
  1237 => x"388d750c",
  1238 => x"84150870",
  1239 => x"892a8106",
  1240 => x"595977f6",
  1241 => x"fb38f785",
  1242 => x"39841508",
  1243 => x"70892a81",
  1244 => x"06595977",
  1245 => x"f4388d75",
  1246 => x"0c841508",
  1247 => x"70892a81",
  1248 => x"06595977",
  1249 => x"f7cc38f7",
  1250 => x"d6398415",
  1251 => x"0870892a",
  1252 => x"81065959",
  1253 => x"77f4388d",
  1254 => x"750c8415",
  1255 => x"0870892a",
  1256 => x"81065959",
  1257 => x"77f7e038",
  1258 => x"f7ea3984",
  1259 => x"15087089",
  1260 => x"2a810659",
  1261 => x"5977f438",
  1262 => x"8d750c84",
  1263 => x"15087089",
  1264 => x"2a810659",
  1265 => x"5977f8b0",
  1266 => x"38f8ba39",
  1267 => x"84150870",
  1268 => x"892a8106",
  1269 => x"595977f4",
  1270 => x"388d750c",
  1271 => x"84150870",
  1272 => x"892a8106",
  1273 => x"595977f8",
  1274 => x"c438f8ce",
  1275 => x"39841508",
  1276 => x"70892a81",
  1277 => x"06595977",
  1278 => x"f4388d75",
  1279 => x"0c841508",
  1280 => x"70892a81",
  1281 => x"06595977",
  1282 => x"f99438f9",
  1283 => x"9e398415",
  1284 => x"0870892a",
  1285 => x"81065959",
  1286 => x"77f4388d",
  1287 => x"750c8415",
  1288 => x"0870892a",
  1289 => x"81065959",
  1290 => x"77f9a838",
  1291 => x"f9b23984",
  1292 => x"15087089",
  1293 => x"2a810659",
  1294 => x"5977f438",
  1295 => x"8d750c84",
  1296 => x"15087089",
  1297 => x"2a810659",
  1298 => x"5977f9f9",
  1299 => x"38fa8339",
  1300 => x"7618b715",
  1301 => x"5555f9c0",
  1302 => x"397618b7",
  1303 => x"155555f8",
  1304 => x"91397618",
  1305 => x"b7155555",
  1306 => x"f6e23976",
  1307 => x"18b71555",
  1308 => x"55f5b339",
  1309 => x"7618b715",
  1310 => x"5555f483",
  1311 => x"397618b7",
  1312 => x"155555f2",
  1313 => x"d3397618",
  1314 => x"b7155555",
  1315 => x"f1a33976",
  1316 => x"18b71555",
  1317 => x"55eff339",
  1318 => x"7618b715",
  1319 => x"5555eec3",
  1320 => x"3980e18c",
  1321 => x"08841108",
  1322 => x"70892a81",
  1323 => x"06585955",
  1324 => x"75f9a838",
  1325 => x"f9b239e4",
  1326 => x"3d0d80dd",
  1327 => x"d40b80dd",
  1328 => x"d4335557",
  1329 => x"73802ea7",
  1330 => x"387380e1",
  1331 => x"8c085656",
  1332 => x"81175775",
  1333 => x"8a2e85b1",
  1334 => x"38841508",
  1335 => x"70892a81",
  1336 => x"065b5c79",
  1337 => x"f4387575",
  1338 => x"0c763356",
  1339 => x"75e2389f",
  1340 => x"0b973d02",
  1341 => x"880580d5",
  1342 => x"059c3d97",
  1343 => x"3d029405",
  1344 => x"80c90541",
  1345 => x"44404442",
  1346 => x"5f80dde8",
  1347 => x"0b80dde8",
  1348 => x"33555773",
  1349 => x"802ea738",
  1350 => x"80e18c08",
  1351 => x"74575581",
  1352 => x"1757758a",
  1353 => x"2e858338",
  1354 => x"84150870",
  1355 => x"892a8106",
  1356 => x"5a5b78f4",
  1357 => x"3875750c",
  1358 => x"76335675",
  1359 => x"e2387e56",
  1360 => x"8b5380dc",
  1361 => x"94526051",
  1362 => x"979a3f82",
  1363 => x"57758f06",
  1364 => x"54738926",
  1365 => x"84f53861",
  1366 => x"17b01555",
  1367 => x"55737534",
  1368 => x"75842aff",
  1369 => x"187081ff",
  1370 => x"06595656",
  1371 => x"76df3860",
  1372 => x"61335557",
  1373 => x"73802ea7",
  1374 => x"3880e18c",
  1375 => x"08745755",
  1376 => x"81175775",
  1377 => x"8a2e84df",
  1378 => x"38841508",
  1379 => x"70892a81",
  1380 => x"065a5b78",
  1381 => x"f4387575",
  1382 => x"0c763356",
  1383 => x"75e23880",
  1384 => x"7f83ffff",
  1385 => x"065f5b7a",
  1386 => x"872e86a0",
  1387 => x"387a932e",
  1388 => x"869f387a",
  1389 => x"982e8686",
  1390 => x"3880ddf8",
  1391 => x"0b80ddf8",
  1392 => x"33555773",
  1393 => x"802ea738",
  1394 => x"80e18c08",
  1395 => x"74575581",
  1396 => x"1757758a",
  1397 => x"2e84b138",
  1398 => x"84150870",
  1399 => x"892a8106",
  1400 => x"5b5879f4",
  1401 => x"3875750c",
  1402 => x"76335675",
  1403 => x"e2387c5a",
  1404 => x"807b5758",
  1405 => x"777b2485",
  1406 => x"93387918",
  1407 => x"578a5275",
  1408 => x"5191b33f",
  1409 => x"8008b005",
  1410 => x"55747734",
  1411 => x"8118588a",
  1412 => x"52755190",
  1413 => x"fc3f8008",
  1414 => x"568008de",
  1415 => x"38800878",
  1416 => x"9f2a1970",
  1417 => x"812c5b57",
  1418 => x"57807925",
  1419 => x"9e387918",
  1420 => x"ff055676",
  1421 => x"1a703356",
  1422 => x"54753374",
  1423 => x"34747634",
  1424 => x"8117ff17",
  1425 => x"57577877",
  1426 => x"24e93877",
  1427 => x"1a598079",
  1428 => x"347c7d33",
  1429 => x"55577380",
  1430 => x"2ea73880",
  1431 => x"e18c0874",
  1432 => x"57558117",
  1433 => x"57758a2e",
  1434 => x"83bf3884",
  1435 => x"15087089",
  1436 => x"2a81065a",
  1437 => x"5878f438",
  1438 => x"75750c76",
  1439 => x"335675e2",
  1440 => x"3880de84",
  1441 => x"0b80de84",
  1442 => x"33555773",
  1443 => x"802ea738",
  1444 => x"80e18c08",
  1445 => x"74575581",
  1446 => x"1757758a",
  1447 => x"2e83ab38",
  1448 => x"84150870",
  1449 => x"892a8106",
  1450 => x"595977f4",
  1451 => x"3875750c",
  1452 => x"76335675",
  1453 => x"e2387a83",
  1454 => x"ffff0680",
  1455 => x"e1800856",
  1456 => x"56901508",
  1457 => x"70832a81",
  1458 => x"06585876",
  1459 => x"f4387d8b",
  1460 => x"2b76862b",
  1461 => x"07820790",
  1462 => x"160c9015",
  1463 => x"0870832a",
  1464 => x"81065a5a",
  1465 => x"78f43890",
  1466 => x"15087090",
  1467 => x"2a57588b",
  1468 => x"5380dc94",
  1469 => x"527f5193",
  1470 => x"eb3f8457",
  1471 => x"758f0654",
  1472 => x"73892683",
  1473 => x"be38761c",
  1474 => x"b0155555",
  1475 => x"73753475",
  1476 => x"842aff18",
  1477 => x"7081ff06",
  1478 => x"59565676",
  1479 => x"df387f60",
  1480 => x"33555773",
  1481 => x"802ea738",
  1482 => x"80e18c08",
  1483 => x"74575581",
  1484 => x"1757758a",
  1485 => x"2e82b438",
  1486 => x"84150870",
  1487 => x"892a8106",
  1488 => x"595977f4",
  1489 => x"3875750c",
  1490 => x"76335675",
  1491 => x"e238811b",
  1492 => x"5b9f7b27",
  1493 => x"fcd13881",
  1494 => x"1f5f9f7f",
  1495 => x"27fbaa38",
  1496 => x"80e18c08",
  1497 => x"55841508",
  1498 => x"70892a81",
  1499 => x"065e407c",
  1500 => x"f4388d75",
  1501 => x"0c841508",
  1502 => x"70892a81",
  1503 => x"06425c60",
  1504 => x"f4388a75",
  1505 => x"0c9e3d0d",
  1506 => x"04841508",
  1507 => x"70892a81",
  1508 => x"06555973",
  1509 => x"f4388d75",
  1510 => x"0c841508",
  1511 => x"70892a81",
  1512 => x"065b5c79",
  1513 => x"fab338fa",
  1514 => x"bd398415",
  1515 => x"0870892a",
  1516 => x"81065f58",
  1517 => x"7df4388d",
  1518 => x"750c8415",
  1519 => x"0870892a",
  1520 => x"81065a5b",
  1521 => x"78fae138",
  1522 => x"faeb3961",
  1523 => x"17b71555",
  1524 => x"55737534",
  1525 => x"75842aff",
  1526 => x"187081ff",
  1527 => x"06595656",
  1528 => x"76faea38",
  1529 => x"fb893984",
  1530 => x"15087089",
  1531 => x"2a81065f",
  1532 => x"587df438",
  1533 => x"8d750c84",
  1534 => x"15087089",
  1535 => x"2a81065a",
  1536 => x"5b78fb85",
  1537 => x"38fb8f39",
  1538 => x"84150870",
  1539 => x"892a8106",
  1540 => x"555973f4",
  1541 => x"388d750c",
  1542 => x"84150870",
  1543 => x"892a8106",
  1544 => x"5b5879fb",
  1545 => x"b338fbbd",
  1546 => x"39841508",
  1547 => x"70892a81",
  1548 => x"065b5479",
  1549 => x"f4388d75",
  1550 => x"0c841508",
  1551 => x"70892a81",
  1552 => x"065a5878",
  1553 => x"fca538fc",
  1554 => x"af398415",
  1555 => x"0870892a",
  1556 => x"8106555a",
  1557 => x"73f4388d",
  1558 => x"750c8415",
  1559 => x"0870892a",
  1560 => x"81065959",
  1561 => x"77fcb938",
  1562 => x"fcc33984",
  1563 => x"15087089",
  1564 => x"2a810655",
  1565 => x"5a73f438",
  1566 => x"8d750c84",
  1567 => x"15087089",
  1568 => x"2a810659",
  1569 => x"5977fdb0",
  1570 => x"38fdba39",
  1571 => x"ad7d3402",
  1572 => x"80e1057b",
  1573 => x"30711a59",
  1574 => x"575a8a52",
  1575 => x"75518c96",
  1576 => x"3f8008b0",
  1577 => x"05557477",
  1578 => x"34811858",
  1579 => x"8a527551",
  1580 => x"8bdf3f80",
  1581 => x"08568008",
  1582 => x"fac038fa",
  1583 => x"e0399b5b",
  1584 => x"f9f73976",
  1585 => x"1cb71555",
  1586 => x"55fcc139",
  1587 => x"905bf9e9",
  1588 => x"39945bf9",
  1589 => x"e439ef3d",
  1590 => x"0d80e184",
  1591 => x"0857810b",
  1592 => x"84180c80",
  1593 => x"55fa8080",
  1594 => x"82805680",
  1595 => x"e4753176",
  1596 => x"70840558",
  1597 => x"0c811555",
  1598 => x"80c07526",
  1599 => x"ee38830b",
  1600 => x"84180cfa",
  1601 => x"80808280",
  1602 => x"0bfa8080",
  1603 => x"80840cb0",
  1604 => x"c00b850a",
  1605 => x"0c80e180",
  1606 => x"0858850a",
  1607 => x"0b94190c",
  1608 => x"91780c80",
  1609 => x"f59754ff",
  1610 => x"b5145473",
  1611 => x"8025f838",
  1612 => x"80de880b",
  1613 => x"80de8833",
  1614 => x"55577380",
  1615 => x"2ea73873",
  1616 => x"80e18c08",
  1617 => x"56568117",
  1618 => x"57758a2e",
  1619 => x"83d03884",
  1620 => x"15087089",
  1621 => x"2a810651",
  1622 => x"5473f438",
  1623 => x"75750c76",
  1624 => x"335675e2",
  1625 => x"38770891",
  1626 => x"3d5a568b",
  1627 => x"5380dc94",
  1628 => x"5278518e",
  1629 => x"ef3f8802",
  1630 => x"8405bd05",
  1631 => x"5957758f",
  1632 => x"06547389",
  1633 => x"2684ef38",
  1634 => x"7618b015",
  1635 => x"55557375",
  1636 => x"3475842a",
  1637 => x"ff187081",
  1638 => x"ff065956",
  1639 => x"5676df38",
  1640 => x"78793355",
  1641 => x"5773802e",
  1642 => x"a73880e1",
  1643 => x"8c087457",
  1644 => x"55811757",
  1645 => x"758a2e83",
  1646 => x"86388415",
  1647 => x"0870892a",
  1648 => x"81065954",
  1649 => x"77f43875",
  1650 => x"750c7633",
  1651 => x"5675e238",
  1652 => x"80de9c0b",
  1653 => x"80de9c33",
  1654 => x"55577380",
  1655 => x"2ea73880",
  1656 => x"e18c0874",
  1657 => x"57558117",
  1658 => x"57758a2e",
  1659 => x"82f23884",
  1660 => x"15087089",
  1661 => x"2a810659",
  1662 => x"5477f438",
  1663 => x"75750c76",
  1664 => x"335675e2",
  1665 => x"3880e180",
  1666 => x"08841108",
  1667 => x"8f3d5b57",
  1668 => x"578b5380",
  1669 => x"dc945278",
  1670 => x"518dc93f",
  1671 => x"88028405",
  1672 => x"b1055957",
  1673 => x"758f0654",
  1674 => x"73892683",
  1675 => x"c0387618",
  1676 => x"b0155555",
  1677 => x"73753475",
  1678 => x"842aff18",
  1679 => x"7081ff06",
  1680 => x"59565676",
  1681 => x"df387879",
  1682 => x"33555773",
  1683 => x"802ea738",
  1684 => x"80e18c08",
  1685 => x"74575581",
  1686 => x"1757758a",
  1687 => x"2e82a238",
  1688 => x"84150870",
  1689 => x"892a8106",
  1690 => x"595477f4",
  1691 => x"3875750c",
  1692 => x"76335675",
  1693 => x"e23880de",
  1694 => x"b00b80de",
  1695 => x"b0335557",
  1696 => x"73802ea7",
  1697 => x"3880e18c",
  1698 => x"08745755",
  1699 => x"81175775",
  1700 => x"8a2e828e",
  1701 => x"38841508",
  1702 => x"70892a81",
  1703 => x"06595477",
  1704 => x"f4387575",
  1705 => x"0c763356",
  1706 => x"75e23885",
  1707 => x"0a088b3d",
  1708 => x"5a568b53",
  1709 => x"80dc9452",
  1710 => x"78518ca8",
  1711 => x"3f880284",
  1712 => x"05a50559",
  1713 => x"57758f06",
  1714 => x"54738926",
  1715 => x"82963876",
  1716 => x"18b01555",
  1717 => x"55737534",
  1718 => x"75842aff",
  1719 => x"187081ff",
  1720 => x"06595656",
  1721 => x"76df3878",
  1722 => x"79335557",
  1723 => x"73802ea7",
  1724 => x"3880e18c",
  1725 => x"08745755",
  1726 => x"81175775",
  1727 => x"8a2e81c3",
  1728 => x"38841508",
  1729 => x"70892a81",
  1730 => x"06595477",
  1731 => x"f4387575",
  1732 => x"0c763356",
  1733 => x"75e238f3",
  1734 => x"9e3f933d",
  1735 => x"0d048415",
  1736 => x"0870892a",
  1737 => x"81065159",
  1738 => x"78f4388d",
  1739 => x"750c8415",
  1740 => x"0870892a",
  1741 => x"81065154",
  1742 => x"73fc9438",
  1743 => x"fc9e3984",
  1744 => x"15087089",
  1745 => x"2a810659",
  1746 => x"5477f438",
  1747 => x"8d750c84",
  1748 => x"15087089",
  1749 => x"2a810659",
  1750 => x"5477fcde",
  1751 => x"38fce839",
  1752 => x"84150870",
  1753 => x"892a8106",
  1754 => x"595477f4",
  1755 => x"388d750c",
  1756 => x"84150870",
  1757 => x"892a8106",
  1758 => x"595477fc",
  1759 => x"f238fcfc",
  1760 => x"39841508",
  1761 => x"70892a81",
  1762 => x"06595477",
  1763 => x"f4388d75",
  1764 => x"0c841508",
  1765 => x"70892a81",
  1766 => x"06595477",
  1767 => x"fdc238fd",
  1768 => x"cc398415",
  1769 => x"0870892a",
  1770 => x"81065954",
  1771 => x"77f4388d",
  1772 => x"750c8415",
  1773 => x"0870892a",
  1774 => x"81065954",
  1775 => x"77fdd638",
  1776 => x"fde03984",
  1777 => x"15087089",
  1778 => x"2a810659",
  1779 => x"5477f438",
  1780 => x"8d750c84",
  1781 => x"15087089",
  1782 => x"2a810659",
  1783 => x"5477fea1",
  1784 => x"38feab39",
  1785 => x"7618b715",
  1786 => x"5555fde9",
  1787 => x"397618b7",
  1788 => x"155555fc",
  1789 => x"bf397618",
  1790 => x"b7155555",
  1791 => x"fb9039f8",
  1792 => x"3d0d80e1",
  1793 => x"84087008",
  1794 => x"810a0680",
  1795 => x"e1880856",
  1796 => x"5a53870b",
  1797 => x"84150c80",
  1798 => x"e18c0854",
  1799 => x"b60b8c15",
  1800 => x"0c830b88",
  1801 => x"150c81ff",
  1802 => x"0b88140c",
  1803 => x"80e18008",
  1804 => x"55ff0b84",
  1805 => x"160cfc94",
  1806 => x"800b8816",
  1807 => x"0c82d0af",
  1808 => x"fdfb0b8c",
  1809 => x"160c80c0",
  1810 => x"750c7408",
  1811 => x"70862a81",
  1812 => x"06575875",
  1813 => x"f5389015",
  1814 => x"0870832a",
  1815 => x"81065457",
  1816 => x"72f43881",
  1817 => x"fc80810b",
  1818 => x"90160c90",
  1819 => x"15087083",
  1820 => x"2a810659",
  1821 => x"5677f438",
  1822 => x"80fdc081",
  1823 => x"0b90160c",
  1824 => x"80dec40b",
  1825 => x"80dec433",
  1826 => x"54567280",
  1827 => x"2ea23872",
  1828 => x"55811656",
  1829 => x"748a2e82",
  1830 => x"94388414",
  1831 => x"0870892a",
  1832 => x"81065853",
  1833 => x"76f43874",
  1834 => x"740c7533",
  1835 => x"5574e238",
  1836 => x"80dec80b",
  1837 => x"80dec833",
  1838 => x"54567280",
  1839 => x"2ea23872",
  1840 => x"55811656",
  1841 => x"748a2e82",
  1842 => x"85388414",
  1843 => x"0870892a",
  1844 => x"81065853",
  1845 => x"76f43874",
  1846 => x"740c7533",
  1847 => x"5574e238",
  1848 => x"78802e82",
  1849 => x"cf3880de",
  1850 => x"d00b80de",
  1851 => x"d0335456",
  1852 => x"72802ea2",
  1853 => x"38725581",
  1854 => x"1656748a",
  1855 => x"2e81f038",
  1856 => x"84140870",
  1857 => x"892a8106",
  1858 => x"585376f4",
  1859 => x"3874740c",
  1860 => x"75335574",
  1861 => x"e23880de",
  1862 => x"e00b80de",
  1863 => x"e0335456",
  1864 => x"72802ea2",
  1865 => x"38725581",
  1866 => x"1656748a",
  1867 => x"2e81e138",
  1868 => x"84140870",
  1869 => x"892a8106",
  1870 => x"585376f4",
  1871 => x"3874740c",
  1872 => x"75335574",
  1873 => x"e238f78e",
  1874 => x"3ff881c0",
  1875 => x"8e8055a0",
  1876 => x"0b80e184",
  1877 => x"0880e188",
  1878 => x"085a5856",
  1879 => x"7484180c",
  1880 => x"749f2a75",
  1881 => x"10075578",
  1882 => x"802e9838",
  1883 => x"75802e81",
  1884 => x"c038ff16",
  1885 => x"7584190c",
  1886 => x"759f2a76",
  1887 => x"10075656",
  1888 => x"78ea3877",
  1889 => x"54afd7c2",
  1890 => x"0b94190c",
  1891 => x"850b9819",
  1892 => x"0c981408",
  1893 => x"70810651",
  1894 => x"5372802e",
  1895 => x"ffbe3898",
  1896 => x"14087081",
  1897 => x"06515372",
  1898 => x"e838ffb0",
  1899 => x"39841408",
  1900 => x"70892a81",
  1901 => x"06585376",
  1902 => x"f4388d74",
  1903 => x"0c841408",
  1904 => x"70892a81",
  1905 => x"06585376",
  1906 => x"fdd038fd",
  1907 => x"da398414",
  1908 => x"0870892a",
  1909 => x"81065853",
  1910 => x"76f4388d",
  1911 => x"740c8414",
  1912 => x"0870892a",
  1913 => x"81065853",
  1914 => x"76fddf38",
  1915 => x"fde93984",
  1916 => x"14087089",
  1917 => x"2a810658",
  1918 => x"5376f438",
  1919 => x"8d740c84",
  1920 => x"14087089",
  1921 => x"2a810658",
  1922 => x"5376fdf4",
  1923 => x"38fdfe39",
  1924 => x"84140870",
  1925 => x"892a8106",
  1926 => x"585376f4",
  1927 => x"388d740c",
  1928 => x"84140870",
  1929 => x"892a8106",
  1930 => x"585376fe",
  1931 => x"8338fe8d",
  1932 => x"3985a43f",
  1933 => x"80df840b",
  1934 => x"80df8433",
  1935 => x"54567280",
  1936 => x"2efdd338",
  1937 => x"72811757",
  1938 => x"55748a2e",
  1939 => x"a5388414",
  1940 => x"0870892a",
  1941 => x"81065853",
  1942 => x"76f43874",
  1943 => x"740c7533",
  1944 => x"5574802e",
  1945 => x"fdb03881",
  1946 => x"1656748a",
  1947 => x"2e098106",
  1948 => x"dd388414",
  1949 => x"0870892a",
  1950 => x"81065853",
  1951 => x"76f4388d",
  1952 => x"740c8414",
  1953 => x"0870892a",
  1954 => x"81065853",
  1955 => x"76c038cb",
  1956 => x"398c0802",
  1957 => x"8c0cfd3d",
  1958 => x"0d80538c",
  1959 => x"088c0508",
  1960 => x"528c0888",
  1961 => x"05085182",
  1962 => x"de3f8008",
  1963 => x"70800c54",
  1964 => x"853d0d8c",
  1965 => x"0c048c08",
  1966 => x"028c0cfd",
  1967 => x"3d0d8153",
  1968 => x"8c088c05",
  1969 => x"08528c08",
  1970 => x"88050851",
  1971 => x"82b93f80",
  1972 => x"0870800c",
  1973 => x"54853d0d",
  1974 => x"8c0c048c",
  1975 => x"08028c0c",
  1976 => x"f93d0d80",
  1977 => x"0b8c08fc",
  1978 => x"050c8c08",
  1979 => x"88050880",
  1980 => x"25ab388c",
  1981 => x"08880508",
  1982 => x"308c0888",
  1983 => x"050c800b",
  1984 => x"8c08f405",
  1985 => x"0c8c08fc",
  1986 => x"05088838",
  1987 => x"810b8c08",
  1988 => x"f4050c8c",
  1989 => x"08f40508",
  1990 => x"8c08fc05",
  1991 => x"0c8c088c",
  1992 => x"05088025",
  1993 => x"ab388c08",
  1994 => x"8c050830",
  1995 => x"8c088c05",
  1996 => x"0c800b8c",
  1997 => x"08f0050c",
  1998 => x"8c08fc05",
  1999 => x"08883881",
  2000 => x"0b8c08f0",
  2001 => x"050c8c08",
  2002 => x"f005088c",
  2003 => x"08fc050c",
  2004 => x"80538c08",
  2005 => x"8c050852",
  2006 => x"8c088805",
  2007 => x"085181a7",
  2008 => x"3f800870",
  2009 => x"8c08f805",
  2010 => x"0c548c08",
  2011 => x"fc050880",
  2012 => x"2e8c388c",
  2013 => x"08f80508",
  2014 => x"308c08f8",
  2015 => x"050c8c08",
  2016 => x"f8050870",
  2017 => x"800c5489",
  2018 => x"3d0d8c0c",
  2019 => x"048c0802",
  2020 => x"8c0cfb3d",
  2021 => x"0d800b8c",
  2022 => x"08fc050c",
  2023 => x"8c088805",
  2024 => x"08802593",
  2025 => x"388c0888",
  2026 => x"0508308c",
  2027 => x"0888050c",
  2028 => x"810b8c08",
  2029 => x"fc050c8c",
  2030 => x"088c0508",
  2031 => x"80258c38",
  2032 => x"8c088c05",
  2033 => x"08308c08",
  2034 => x"8c050c81",
  2035 => x"538c088c",
  2036 => x"0508528c",
  2037 => x"08880508",
  2038 => x"51ad3f80",
  2039 => x"08708c08",
  2040 => x"f8050c54",
  2041 => x"8c08fc05",
  2042 => x"08802e8c",
  2043 => x"388c08f8",
  2044 => x"0508308c",
  2045 => x"08f8050c",
  2046 => x"8c08f805",
  2047 => x"0870800c",
  2048 => x"54873d0d",
  2049 => x"8c0c048c",
  2050 => x"08028c0c",
  2051 => x"fd3d0d81",
  2052 => x"0b8c08fc",
  2053 => x"050c800b",
  2054 => x"8c08f805",
  2055 => x"0c8c088c",
  2056 => x"05088c08",
  2057 => x"88050827",
  2058 => x"ac388c08",
  2059 => x"fc050880",
  2060 => x"2ea33880",
  2061 => x"0b8c088c",
  2062 => x"05082499",
  2063 => x"388c088c",
  2064 => x"0508108c",
  2065 => x"088c050c",
  2066 => x"8c08fc05",
  2067 => x"08108c08",
  2068 => x"fc050cc9",
  2069 => x"398c08fc",
  2070 => x"0508802e",
  2071 => x"80c9388c",
  2072 => x"088c0508",
  2073 => x"8c088805",
  2074 => x"0826a138",
  2075 => x"8c088805",
  2076 => x"088c088c",
  2077 => x"0508318c",
  2078 => x"0888050c",
  2079 => x"8c08f805",
  2080 => x"088c08fc",
  2081 => x"0508078c",
  2082 => x"08f8050c",
  2083 => x"8c08fc05",
  2084 => x"08812a8c",
  2085 => x"08fc050c",
  2086 => x"8c088c05",
  2087 => x"08812a8c",
  2088 => x"088c050c",
  2089 => x"ffaf398c",
  2090 => x"08900508",
  2091 => x"802e8f38",
  2092 => x"8c088805",
  2093 => x"08708c08",
  2094 => x"f4050c51",
  2095 => x"8d398c08",
  2096 => x"f8050870",
  2097 => x"8c08f405",
  2098 => x"0c518c08",
  2099 => x"f4050880",
  2100 => x"0c853d0d",
  2101 => x"8c0c0480",
  2102 => x"3d0d8651",
  2103 => x"84963f81",
  2104 => x"5198d73f",
  2105 => x"fc3d0d76",
  2106 => x"70797b55",
  2107 => x"5555558f",
  2108 => x"72278c38",
  2109 => x"72750783",
  2110 => x"06517080",
  2111 => x"2ea738ff",
  2112 => x"125271ff",
  2113 => x"2e983872",
  2114 => x"70810554",
  2115 => x"33747081",
  2116 => x"055634ff",
  2117 => x"125271ff",
  2118 => x"2e098106",
  2119 => x"ea387480",
  2120 => x"0c863d0d",
  2121 => x"04745172",
  2122 => x"70840554",
  2123 => x"08717084",
  2124 => x"05530c72",
  2125 => x"70840554",
  2126 => x"08717084",
  2127 => x"05530c72",
  2128 => x"70840554",
  2129 => x"08717084",
  2130 => x"05530c72",
  2131 => x"70840554",
  2132 => x"08717084",
  2133 => x"05530cf0",
  2134 => x"1252718f",
  2135 => x"26c93883",
  2136 => x"72279538",
  2137 => x"72708405",
  2138 => x"54087170",
  2139 => x"8405530c",
  2140 => x"fc125271",
  2141 => x"8326ed38",
  2142 => x"7054ff83",
  2143 => x"39fd3d0d",
  2144 => x"755384d8",
  2145 => x"1308802e",
  2146 => x"8a388053",
  2147 => x"72800c85",
  2148 => x"3d0d0481",
  2149 => x"80527251",
  2150 => x"83d83f80",
  2151 => x"0884d814",
  2152 => x"0cff5380",
  2153 => x"08802ee4",
  2154 => x"38800854",
  2155 => x"9f538074",
  2156 => x"70840556",
  2157 => x"0cff1353",
  2158 => x"807324ce",
  2159 => x"38807470",
  2160 => x"8405560c",
  2161 => x"ff135372",
  2162 => x"8025e338",
  2163 => x"ffbc39fd",
  2164 => x"3d0d7577",
  2165 => x"55539f74",
  2166 => x"278d3896",
  2167 => x"730cff52",
  2168 => x"71800c85",
  2169 => x"3d0d0484",
  2170 => x"d8130852",
  2171 => x"71802e93",
  2172 => x"38731010",
  2173 => x"12700879",
  2174 => x"720c5152",
  2175 => x"71800c85",
  2176 => x"3d0d0472",
  2177 => x"51fef63f",
  2178 => x"ff528008",
  2179 => x"d33884d8",
  2180 => x"13087410",
  2181 => x"10117008",
  2182 => x"7a720c51",
  2183 => x"5152dd39",
  2184 => x"f93d0d79",
  2185 => x"7b585676",
  2186 => x"9f2680e8",
  2187 => x"3884d816",
  2188 => x"08547380",
  2189 => x"2eaa3876",
  2190 => x"10101470",
  2191 => x"08555573",
  2192 => x"802eba38",
  2193 => x"80587381",
  2194 => x"2e8f3873",
  2195 => x"ff2ea338",
  2196 => x"80750c76",
  2197 => x"51732d80",
  2198 => x"5877800c",
  2199 => x"893d0d04",
  2200 => x"7551fe99",
  2201 => x"3fff5880",
  2202 => x"08ef3884",
  2203 => x"d8160854",
  2204 => x"c6399676",
  2205 => x"0c810b80",
  2206 => x"0c893d0d",
  2207 => x"04755181",
  2208 => x"ed3f7653",
  2209 => x"80085275",
  2210 => x"5181ad3f",
  2211 => x"8008800c",
  2212 => x"893d0d04",
  2213 => x"96760cff",
  2214 => x"0b800c89",
  2215 => x"3d0d04fc",
  2216 => x"3d0d7678",
  2217 => x"5653ff54",
  2218 => x"749f26b1",
  2219 => x"3884d813",
  2220 => x"08527180",
  2221 => x"2eae3874",
  2222 => x"10101270",
  2223 => x"08535381",
  2224 => x"5471802e",
  2225 => x"98388254",
  2226 => x"71ff2e91",
  2227 => x"38835471",
  2228 => x"812e8a38",
  2229 => x"80730c74",
  2230 => x"51712d80",
  2231 => x"5473800c",
  2232 => x"863d0d04",
  2233 => x"7251fd95",
  2234 => x"3f8008f1",
  2235 => x"3884d813",
  2236 => x"0852c439",
  2237 => x"ff3d0d73",
  2238 => x"5280e190",
  2239 => x"0851fea0",
  2240 => x"3f833d0d",
  2241 => x"04fe3d0d",
  2242 => x"75537452",
  2243 => x"80e19008",
  2244 => x"51fdbc3f",
  2245 => x"843d0d04",
  2246 => x"803d0d80",
  2247 => x"e1900851",
  2248 => x"fcdb3f82",
  2249 => x"3d0d04ff",
  2250 => x"3d0d7352",
  2251 => x"80e19008",
  2252 => x"51feec3f",
  2253 => x"833d0d04",
  2254 => x"fc3d0d80",
  2255 => x"0b80f184",
  2256 => x"0c785277",
  2257 => x"5192e73f",
  2258 => x"80085480",
  2259 => x"08ff2e88",
  2260 => x"3873800c",
  2261 => x"863d0d04",
  2262 => x"80f18408",
  2263 => x"5574802e",
  2264 => x"f0387675",
  2265 => x"710c5373",
  2266 => x"800c863d",
  2267 => x"0d0492b9",
  2268 => x"3f04f33d",
  2269 => x"0d7f618b",
  2270 => x"1170f806",
  2271 => x"5c55555e",
  2272 => x"72962683",
  2273 => x"38905980",
  2274 => x"7924747a",
  2275 => x"26075380",
  2276 => x"5472742e",
  2277 => x"09810680",
  2278 => x"cb387d51",
  2279 => x"8bca3f78",
  2280 => x"83f72680",
  2281 => x"c6387883",
  2282 => x"2a701010",
  2283 => x"1080e8cc",
  2284 => x"058c1108",
  2285 => x"59595a76",
  2286 => x"782e83b0",
  2287 => x"38841708",
  2288 => x"fc06568c",
  2289 => x"17088818",
  2290 => x"08718c12",
  2291 => x"0c88120c",
  2292 => x"58751784",
  2293 => x"11088107",
  2294 => x"84120c53",
  2295 => x"7d518b89",
  2296 => x"3f881754",
  2297 => x"73800c8f",
  2298 => x"3d0d0478",
  2299 => x"892a7983",
  2300 => x"2a5b5372",
  2301 => x"802ebf38",
  2302 => x"78862ab8",
  2303 => x"055a8473",
  2304 => x"27b43880",
  2305 => x"db135a94",
  2306 => x"7327ab38",
  2307 => x"788c2a80",
  2308 => x"ee055a80",
  2309 => x"d473279e",
  2310 => x"38788f2a",
  2311 => x"80f7055a",
  2312 => x"82d47327",
  2313 => x"91387892",
  2314 => x"2a80fc05",
  2315 => x"5a8ad473",
  2316 => x"27843880",
  2317 => x"fe5a7910",
  2318 => x"101080e8",
  2319 => x"cc058c11",
  2320 => x"08585576",
  2321 => x"752ea338",
  2322 => x"841708fc",
  2323 => x"06707a31",
  2324 => x"5556738f",
  2325 => x"2488d538",
  2326 => x"738025fe",
  2327 => x"e6388c17",
  2328 => x"08577675",
  2329 => x"2e098106",
  2330 => x"df38811a",
  2331 => x"5a80e8dc",
  2332 => x"08577680",
  2333 => x"e8d42e82",
  2334 => x"c0388417",
  2335 => x"08fc0670",
  2336 => x"7a315556",
  2337 => x"738f2481",
  2338 => x"f93880e8",
  2339 => x"d40b80e8",
  2340 => x"e00c80e8",
  2341 => x"d40b80e8",
  2342 => x"dc0c7380",
  2343 => x"25feb238",
  2344 => x"83ff7627",
  2345 => x"83df3875",
  2346 => x"892a7683",
  2347 => x"2a555372",
  2348 => x"802ebf38",
  2349 => x"75862ab8",
  2350 => x"05548473",
  2351 => x"27b43880",
  2352 => x"db135494",
  2353 => x"7327ab38",
  2354 => x"758c2a80",
  2355 => x"ee055480",
  2356 => x"d473279e",
  2357 => x"38758f2a",
  2358 => x"80f70554",
  2359 => x"82d47327",
  2360 => x"91387592",
  2361 => x"2a80fc05",
  2362 => x"548ad473",
  2363 => x"27843880",
  2364 => x"fe547310",
  2365 => x"101080e8",
  2366 => x"cc058811",
  2367 => x"08565874",
  2368 => x"782e86cf",
  2369 => x"38841508",
  2370 => x"fc065375",
  2371 => x"73278d38",
  2372 => x"88150855",
  2373 => x"74782e09",
  2374 => x"8106ea38",
  2375 => x"8c150880",
  2376 => x"e8cc0b84",
  2377 => x"0508718c",
  2378 => x"1a0c7688",
  2379 => x"1a0c7888",
  2380 => x"130c788c",
  2381 => x"180c5d58",
  2382 => x"7953807a",
  2383 => x"2483e638",
  2384 => x"72822c81",
  2385 => x"712b5c53",
  2386 => x"7a7c2681",
  2387 => x"98387b7b",
  2388 => x"06537282",
  2389 => x"f13879fc",
  2390 => x"0684055a",
  2391 => x"7a10707d",
  2392 => x"06545b72",
  2393 => x"82e03884",
  2394 => x"1a5af139",
  2395 => x"88178c11",
  2396 => x"08585876",
  2397 => x"782e0981",
  2398 => x"06fcc238",
  2399 => x"821a5afd",
  2400 => x"ec397817",
  2401 => x"79810784",
  2402 => x"190c7080",
  2403 => x"e8e00c70",
  2404 => x"80e8dc0c",
  2405 => x"80e8d40b",
  2406 => x"8c120c8c",
  2407 => x"11088812",
  2408 => x"0c748107",
  2409 => x"84120c74",
  2410 => x"1175710c",
  2411 => x"51537d51",
  2412 => x"87b73f88",
  2413 => x"1754fcac",
  2414 => x"3980e8cc",
  2415 => x"0b840508",
  2416 => x"7a545c79",
  2417 => x"8025fef8",
  2418 => x"3882da39",
  2419 => x"7a097c06",
  2420 => x"7080e8cc",
  2421 => x"0b84050c",
  2422 => x"5c7a105b",
  2423 => x"7a7c2685",
  2424 => x"387a85b8",
  2425 => x"3880e8cc",
  2426 => x"0b880508",
  2427 => x"70841208",
  2428 => x"fc06707c",
  2429 => x"317c7226",
  2430 => x"8f722507",
  2431 => x"57575c5d",
  2432 => x"5572802e",
  2433 => x"80db3879",
  2434 => x"7a1680e8",
  2435 => x"c4081b90",
  2436 => x"115a5557",
  2437 => x"5b80e8c0",
  2438 => x"08ff2e88",
  2439 => x"38a08f13",
  2440 => x"e0800657",
  2441 => x"76527d51",
  2442 => x"86c03f80",
  2443 => x"08548008",
  2444 => x"ff2e9038",
  2445 => x"80087627",
  2446 => x"82993874",
  2447 => x"80e8cc2e",
  2448 => x"82913880",
  2449 => x"e8cc0b88",
  2450 => x"05085584",
  2451 => x"1508fc06",
  2452 => x"707a317a",
  2453 => x"72268f72",
  2454 => x"25075255",
  2455 => x"537283e6",
  2456 => x"38747981",
  2457 => x"0784170c",
  2458 => x"79167080",
  2459 => x"e8cc0b88",
  2460 => x"050c7581",
  2461 => x"0784120c",
  2462 => x"547e5257",
  2463 => x"85eb3f88",
  2464 => x"1754fae0",
  2465 => x"3975832a",
  2466 => x"70545480",
  2467 => x"7424819b",
  2468 => x"3872822c",
  2469 => x"81712b80",
  2470 => x"e8d00807",
  2471 => x"7080e8cc",
  2472 => x"0b84050c",
  2473 => x"75101010",
  2474 => x"80e8cc05",
  2475 => x"88110858",
  2476 => x"5a5d5377",
  2477 => x"8c180c74",
  2478 => x"88180c76",
  2479 => x"88190c76",
  2480 => x"8c160cfc",
  2481 => x"f339797a",
  2482 => x"10101080",
  2483 => x"e8cc0570",
  2484 => x"57595d8c",
  2485 => x"15085776",
  2486 => x"752ea338",
  2487 => x"841708fc",
  2488 => x"06707a31",
  2489 => x"5556738f",
  2490 => x"2483ca38",
  2491 => x"73802584",
  2492 => x"81388c17",
  2493 => x"08577675",
  2494 => x"2e098106",
  2495 => x"df388815",
  2496 => x"811b7083",
  2497 => x"06555b55",
  2498 => x"72c9387c",
  2499 => x"83065372",
  2500 => x"802efdb8",
  2501 => x"38ff1df8",
  2502 => x"19595d88",
  2503 => x"1808782e",
  2504 => x"ea38fdb5",
  2505 => x"39831a53",
  2506 => x"fc963983",
  2507 => x"1470822c",
  2508 => x"81712b80",
  2509 => x"e8d00807",
  2510 => x"7080e8cc",
  2511 => x"0b84050c",
  2512 => x"76101010",
  2513 => x"80e8cc05",
  2514 => x"88110859",
  2515 => x"5b5e5153",
  2516 => x"fee13980",
  2517 => x"e8900817",
  2518 => x"58800876",
  2519 => x"2e818d38",
  2520 => x"80e8c008",
  2521 => x"ff2e83ec",
  2522 => x"38737631",
  2523 => x"1880e890",
  2524 => x"0c738706",
  2525 => x"70575372",
  2526 => x"802e8838",
  2527 => x"88733170",
  2528 => x"15555676",
  2529 => x"149fff06",
  2530 => x"a0807131",
  2531 => x"1770547f",
  2532 => x"53575383",
  2533 => x"d53f8008",
  2534 => x"538008ff",
  2535 => x"2e81a038",
  2536 => x"80e89008",
  2537 => x"167080e8",
  2538 => x"900c7475",
  2539 => x"80e8cc0b",
  2540 => x"88050c74",
  2541 => x"76311870",
  2542 => x"81075155",
  2543 => x"56587b80",
  2544 => x"e8cc2e83",
  2545 => x"9c38798f",
  2546 => x"2682cb38",
  2547 => x"810b8415",
  2548 => x"0c841508",
  2549 => x"fc06707a",
  2550 => x"317a7226",
  2551 => x"8f722507",
  2552 => x"52555372",
  2553 => x"802efcf9",
  2554 => x"3880db39",
  2555 => x"80089fff",
  2556 => x"065372fe",
  2557 => x"eb387780",
  2558 => x"e8900c80",
  2559 => x"e8cc0b88",
  2560 => x"05087b18",
  2561 => x"81078412",
  2562 => x"0c5580e8",
  2563 => x"bc087827",
  2564 => x"86387780",
  2565 => x"e8bc0c80",
  2566 => x"e8b80878",
  2567 => x"27fcac38",
  2568 => x"7780e8b8",
  2569 => x"0c841508",
  2570 => x"fc06707a",
  2571 => x"317a7226",
  2572 => x"8f722507",
  2573 => x"52555372",
  2574 => x"802efca5",
  2575 => x"38883980",
  2576 => x"745456fe",
  2577 => x"db397d51",
  2578 => x"829f3f80",
  2579 => x"0b800c8f",
  2580 => x"3d0d0473",
  2581 => x"53807424",
  2582 => x"a9387282",
  2583 => x"2c81712b",
  2584 => x"80e8d008",
  2585 => x"077080e8",
  2586 => x"cc0b8405",
  2587 => x"0c5d5377",
  2588 => x"8c180c74",
  2589 => x"88180c76",
  2590 => x"88190c76",
  2591 => x"8c160cf9",
  2592 => x"b7398314",
  2593 => x"70822c81",
  2594 => x"712b80e8",
  2595 => x"d0080770",
  2596 => x"80e8cc0b",
  2597 => x"84050c5e",
  2598 => x"5153d439",
  2599 => x"7b7b0653",
  2600 => x"72fca338",
  2601 => x"841a7b10",
  2602 => x"5c5af139",
  2603 => x"ff1a8111",
  2604 => x"515af7b9",
  2605 => x"39781779",
  2606 => x"81078419",
  2607 => x"0c8c1808",
  2608 => x"88190871",
  2609 => x"8c120c88",
  2610 => x"120c5970",
  2611 => x"80e8e00c",
  2612 => x"7080e8dc",
  2613 => x"0c80e8d4",
  2614 => x"0b8c120c",
  2615 => x"8c110888",
  2616 => x"120c7481",
  2617 => x"0784120c",
  2618 => x"74117571",
  2619 => x"0c5153f9",
  2620 => x"bd397517",
  2621 => x"84110881",
  2622 => x"0784120c",
  2623 => x"538c1708",
  2624 => x"88180871",
  2625 => x"8c120c88",
  2626 => x"120c587d",
  2627 => x"5180da3f",
  2628 => x"881754f5",
  2629 => x"cf397284",
  2630 => x"150cf41a",
  2631 => x"f8067084",
  2632 => x"1e088106",
  2633 => x"07841e0c",
  2634 => x"701d545b",
  2635 => x"850b8414",
  2636 => x"0c850b88",
  2637 => x"140c8f7b",
  2638 => x"27fdcf38",
  2639 => x"881c527d",
  2640 => x"5182903f",
  2641 => x"80e8cc0b",
  2642 => x"88050880",
  2643 => x"e8900859",
  2644 => x"55fdb739",
  2645 => x"7780e890",
  2646 => x"0c7380e8",
  2647 => x"c00cfc91",
  2648 => x"39728415",
  2649 => x"0cfda339",
  2650 => x"0404fd3d",
  2651 => x"0d800b80",
  2652 => x"f1840c76",
  2653 => x"5186cc3f",
  2654 => x"80085380",
  2655 => x"08ff2e88",
  2656 => x"3872800c",
  2657 => x"853d0d04",
  2658 => x"80f18408",
  2659 => x"5473802e",
  2660 => x"f0387574",
  2661 => x"710c5272",
  2662 => x"800c853d",
  2663 => x"0d04fb3d",
  2664 => x"0d777052",
  2665 => x"56c23f80",
  2666 => x"e8cc0b88",
  2667 => x"05088411",
  2668 => x"08fc0670",
  2669 => x"7b319fef",
  2670 => x"05e08006",
  2671 => x"e0800556",
  2672 => x"5653a080",
  2673 => x"74249438",
  2674 => x"80527551",
  2675 => x"ff9c3f80",
  2676 => x"e8d40815",
  2677 => x"53728008",
  2678 => x"2e8f3875",
  2679 => x"51ff8a3f",
  2680 => x"80537280",
  2681 => x"0c873d0d",
  2682 => x"04733052",
  2683 => x"7551fefa",
  2684 => x"3f8008ff",
  2685 => x"2ea83880",
  2686 => x"e8cc0b88",
  2687 => x"05087575",
  2688 => x"31810784",
  2689 => x"120c5380",
  2690 => x"e8900874",
  2691 => x"3180e890",
  2692 => x"0c7551fe",
  2693 => x"d43f810b",
  2694 => x"800c873d",
  2695 => x"0d048052",
  2696 => x"7551fec6",
  2697 => x"3f80e8cc",
  2698 => x"0b880508",
  2699 => x"80087131",
  2700 => x"56538f75",
  2701 => x"25ffa438",
  2702 => x"800880e8",
  2703 => x"c0083180",
  2704 => x"e8900c74",
  2705 => x"81078414",
  2706 => x"0c7551fe",
  2707 => x"9c3f8053",
  2708 => x"ff9039f6",
  2709 => x"3d0d7c7e",
  2710 => x"545b7280",
  2711 => x"2e828338",
  2712 => x"7a51fe84",
  2713 => x"3ff81384",
  2714 => x"110870fe",
  2715 => x"06701384",
  2716 => x"1108fc06",
  2717 => x"5d585954",
  2718 => x"5880e8d4",
  2719 => x"08752e82",
  2720 => x"de387884",
  2721 => x"160c8073",
  2722 => x"8106545a",
  2723 => x"727a2e81",
  2724 => x"d5387815",
  2725 => x"84110881",
  2726 => x"06515372",
  2727 => x"a0387817",
  2728 => x"577981e6",
  2729 => x"38881508",
  2730 => x"537280e8",
  2731 => x"d42e82f9",
  2732 => x"388c1508",
  2733 => x"708c150c",
  2734 => x"7388120c",
  2735 => x"56768107",
  2736 => x"84190c76",
  2737 => x"1877710c",
  2738 => x"53798191",
  2739 => x"3883ff77",
  2740 => x"2781c838",
  2741 => x"76892a77",
  2742 => x"832a5653",
  2743 => x"72802ebf",
  2744 => x"3876862a",
  2745 => x"b8055584",
  2746 => x"7327b438",
  2747 => x"80db1355",
  2748 => x"947327ab",
  2749 => x"38768c2a",
  2750 => x"80ee0555",
  2751 => x"80d47327",
  2752 => x"9e38768f",
  2753 => x"2a80f705",
  2754 => x"5582d473",
  2755 => x"27913876",
  2756 => x"922a80fc",
  2757 => x"05558ad4",
  2758 => x"73278438",
  2759 => x"80fe5574",
  2760 => x"10101080",
  2761 => x"e8cc0588",
  2762 => x"11085556",
  2763 => x"73762e82",
  2764 => x"b3388414",
  2765 => x"08fc0653",
  2766 => x"7673278d",
  2767 => x"38881408",
  2768 => x"5473762e",
  2769 => x"098106ea",
  2770 => x"388c1408",
  2771 => x"708c1a0c",
  2772 => x"74881a0c",
  2773 => x"7888120c",
  2774 => x"56778c15",
  2775 => x"0c7a51fc",
  2776 => x"883f8c3d",
  2777 => x"0d047708",
  2778 => x"78713159",
  2779 => x"77058819",
  2780 => x"08545772",
  2781 => x"80e8d42e",
  2782 => x"80e0388c",
  2783 => x"1808708c",
  2784 => x"150c7388",
  2785 => x"120c56fe",
  2786 => x"89398815",
  2787 => x"088c1608",
  2788 => x"708c130c",
  2789 => x"5788170c",
  2790 => x"fea33976",
  2791 => x"832a7054",
  2792 => x"55807524",
  2793 => x"81983872",
  2794 => x"822c8171",
  2795 => x"2b80e8d0",
  2796 => x"080780e8",
  2797 => x"cc0b8405",
  2798 => x"0c537410",
  2799 => x"101080e8",
  2800 => x"cc058811",
  2801 => x"08555675",
  2802 => x"8c190c73",
  2803 => x"88190c77",
  2804 => x"88170c77",
  2805 => x"8c150cff",
  2806 => x"8439815a",
  2807 => x"fdb43978",
  2808 => x"17738106",
  2809 => x"54577298",
  2810 => x"38770878",
  2811 => x"71315977",
  2812 => x"058c1908",
  2813 => x"881a0871",
  2814 => x"8c120c88",
  2815 => x"120c5757",
  2816 => x"76810784",
  2817 => x"190c7780",
  2818 => x"e8cc0b88",
  2819 => x"050c80e8",
  2820 => x"c8087726",
  2821 => x"fec73880",
  2822 => x"e8c40852",
  2823 => x"7a51fafe",
  2824 => x"3f7a51fa",
  2825 => x"c43ffeba",
  2826 => x"3981788c",
  2827 => x"150c7888",
  2828 => x"150c738c",
  2829 => x"1a0c7388",
  2830 => x"1a0c5afd",
  2831 => x"80398315",
  2832 => x"70822c81",
  2833 => x"712b80e8",
  2834 => x"d0080780",
  2835 => x"e8cc0b84",
  2836 => x"050c5153",
  2837 => x"74101010",
  2838 => x"80e8cc05",
  2839 => x"88110855",
  2840 => x"56fee439",
  2841 => x"74538075",
  2842 => x"24a73872",
  2843 => x"822c8171",
  2844 => x"2b80e8d0",
  2845 => x"080780e8",
  2846 => x"cc0b8405",
  2847 => x"0c53758c",
  2848 => x"190c7388",
  2849 => x"190c7788",
  2850 => x"170c778c",
  2851 => x"150cfdcd",
  2852 => x"39831570",
  2853 => x"822c8171",
  2854 => x"2b80e8d0",
  2855 => x"080780e8",
  2856 => x"cc0b8405",
  2857 => x"0c5153d6",
  2858 => x"39810b80",
  2859 => x"0c04803d",
  2860 => x"0d72812e",
  2861 => x"8938800b",
  2862 => x"800c823d",
  2863 => x"0d047351",
  2864 => x"80f83ffe",
  2865 => x"3d0d80f0",
  2866 => x"fc085170",
  2867 => x"8a3880f1",
  2868 => x"887080f0",
  2869 => x"fc0c5170",
  2870 => x"75125252",
  2871 => x"ff537087",
  2872 => x"fb808026",
  2873 => x"88387080",
  2874 => x"f0fc0c71",
  2875 => x"5372800c",
  2876 => x"843d0d04",
  2877 => x"fd3d0d80",
  2878 => x"0b80e0f4",
  2879 => x"08545472",
  2880 => x"812e9c38",
  2881 => x"7380f180",
  2882 => x"0cffaed4",
  2883 => x"3fffadf0",
  2884 => x"3f80f0d4",
  2885 => x"528151dd",
  2886 => x"e63f8008",
  2887 => x"51a23f72",
  2888 => x"80f1800c",
  2889 => x"ffaeb93f",
  2890 => x"ffadd53f",
  2891 => x"80f0d452",
  2892 => x"8151ddcb",
  2893 => x"3f800851",
  2894 => x"873f00ff",
  2895 => x"3900ff39",
  2896 => x"f73d0d7b",
  2897 => x"80e19008",
  2898 => x"82c81108",
  2899 => x"5a545a77",
  2900 => x"802e80da",
  2901 => x"38818818",
  2902 => x"841908ff",
  2903 => x"0581712b",
  2904 => x"59555980",
  2905 => x"742480ea",
  2906 => x"38807424",
  2907 => x"b5387382",
  2908 => x"2b781188",
  2909 => x"05565681",
  2910 => x"80190877",
  2911 => x"06537280",
  2912 => x"2eb63878",
  2913 => x"16700853",
  2914 => x"53795174",
  2915 => x"0853722d",
  2916 => x"ff14fc17",
  2917 => x"fc177981",
  2918 => x"2c5a5757",
  2919 => x"54738025",
  2920 => x"d6387708",
  2921 => x"5877ffad",
  2922 => x"3880e190",
  2923 => x"0853bc13",
  2924 => x"08a53879",
  2925 => x"51ff833f",
  2926 => x"74085372",
  2927 => x"2dff14fc",
  2928 => x"17fc1779",
  2929 => x"812c5a57",
  2930 => x"57547380",
  2931 => x"25ffa838",
  2932 => x"d1398057",
  2933 => x"ff933972",
  2934 => x"51bc1308",
  2935 => x"53722d79",
  2936 => x"51fed73f",
  2937 => x"ff3d0d80",
  2938 => x"f0dc0bfc",
  2939 => x"05700852",
  2940 => x"5270ff2e",
  2941 => x"9138702d",
  2942 => x"fc127008",
  2943 => x"525270ff",
  2944 => x"2e098106",
  2945 => x"f138833d",
  2946 => x"0d0404ff",
  2947 => x"adbf3f04",
  2948 => x"00000040",
  2949 => x"30782020",
  2950 => x"20202020",
  2951 => x"20200000",
  2952 => x"0a677265",
  2953 => x"74682072",
  2954 => x"65676973",
  2955 => x"74657273",
  2956 => x"3a000000",
  2957 => x"0a636f6e",
  2958 => x"74726f6c",
  2959 => x"3a202020",
  2960 => x"20202000",
  2961 => x"0a737461",
  2962 => x"7475733a",
  2963 => x"20202020",
  2964 => x"20202000",
  2965 => x"0a6d6163",
  2966 => x"5f6d7362",
  2967 => x"3a202020",
  2968 => x"20202000",
  2969 => x"0a6d6163",
  2970 => x"5f6c7362",
  2971 => x"3a202020",
  2972 => x"20202000",
  2973 => x"0a6d6469",
  2974 => x"6f5f636f",
  2975 => x"6e74726f",
  2976 => x"6c3a2000",
  2977 => x"0a74785f",
  2978 => x"706f696e",
  2979 => x"7465723a",
  2980 => x"20202000",
  2981 => x"0a72785f",
  2982 => x"706f696e",
  2983 => x"7465723a",
  2984 => x"20202000",
  2985 => x"0a656463",
  2986 => x"6c5f6970",
  2987 => x"3a202020",
  2988 => x"20202000",
  2989 => x"0a686173",
  2990 => x"685f6d73",
  2991 => x"623a2020",
  2992 => x"20202000",
  2993 => x"0a686173",
  2994 => x"685f6c73",
  2995 => x"623a2020",
  2996 => x"20202000",
  2997 => x"0a6d6469",
  2998 => x"6f207068",
  2999 => x"79207265",
  3000 => x"67697374",
  3001 => x"65727300",
  3002 => x"0a206d64",
  3003 => x"696f2070",
  3004 => x"68793a20",
  3005 => x"00000000",
  3006 => x"0a202072",
  3007 => x"65673a20",
  3008 => x"00000000",
  3009 => x"2d3e2000",
  3010 => x"0a677265",
  3011 => x"74682d3e",
  3012 => x"636f6e74",
  3013 => x"726f6c20",
  3014 => x"3a000000",
  3015 => x"0a677265",
  3016 => x"74682d3e",
  3017 => x"73746174",
  3018 => x"75732020",
  3019 => x"3a000000",
  3020 => x"0a646573",
  3021 => x"63722d3e",
  3022 => x"636f6e74",
  3023 => x"726f6c20",
  3024 => x"3a000000",
  3025 => x"0a0a0000",
  3026 => x"74657374",
  3027 => x"2e632000",
  3028 => x"286f6e20",
  3029 => x"73696d75",
  3030 => x"6c61746f",
  3031 => x"72290a00",
  3032 => x"636f6d70",
  3033 => x"696c6564",
  3034 => x"3a204175",
  3035 => x"67203132",
  3036 => x"20323031",
  3037 => x"30202031",
  3038 => x"373a3036",
  3039 => x"3a34330a",
  3040 => x"00000000",
  3041 => x"286f6e20",
  3042 => x"68617264",
  3043 => x"77617265",
  3044 => x"290a0000",
  3045 => x"0000089e",
  3046 => x"000008c4",
  3047 => x"000008c4",
  3048 => x"0000089e",
  3049 => x"000008c4",
  3050 => x"000008c4",
  3051 => x"000008c4",
  3052 => x"000008c4",
  3053 => x"000008c4",
  3054 => x"000008c4",
  3055 => x"000008c4",
  3056 => x"000008c4",
  3057 => x"000008c4",
  3058 => x"000008c4",
  3059 => x"000008c4",
  3060 => x"000008c4",
  3061 => x"000008c4",
  3062 => x"000008c4",
  3063 => x"000008c4",
  3064 => x"000008c4",
  3065 => x"000008c4",
  3066 => x"000008c4",
  3067 => x"000008c4",
  3068 => x"000008c4",
  3069 => x"000008c4",
  3070 => x"000008c4",
  3071 => x"000008c4",
  3072 => x"000008c4",
  3073 => x"000008c4",
  3074 => x"000008c4",
  3075 => x"000008c4",
  3076 => x"000008c4",
  3077 => x"000008c4",
  3078 => x"000008c4",
  3079 => x"000008c4",
  3080 => x"000008c4",
  3081 => x"000008c4",
  3082 => x"000008c4",
  3083 => x"00000966",
  3084 => x"0000095e",
  3085 => x"00000956",
  3086 => x"0000094e",
  3087 => x"00000946",
  3088 => x"0000093e",
  3089 => x"00000936",
  3090 => x"0000092d",
  3091 => x"00000924",
  3092 => x"43000000",
  3093 => x"64756d6d",
  3094 => x"792e6578",
  3095 => x"65000000",
  3096 => x"00ffffff",
  3097 => x"ff00ffff",
  3098 => x"ffff00ff",
  3099 => x"ffffff00",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00000000",
  3103 => x"00003864",
  3104 => x"80000c00",
  3105 => x"80000800",
  3106 => x"80000200",
  3107 => x"80000100",
  3108 => x"00003094",
  3109 => x"00000000",
  3110 => x"000032fc",
  3111 => x"00003358",
  3112 => x"000033b4",
  3113 => x"00000000",
  3114 => x"00000000",
  3115 => x"00000000",
  3116 => x"00000000",
  3117 => x"00000000",
  3118 => x"00000000",
  3119 => x"00000000",
  3120 => x"00000000",
  3121 => x"00000000",
  3122 => x"00003050",
  3123 => x"00000000",
  3124 => x"00000000",
  3125 => x"00000000",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000000",
  3151 => x"00000001",
  3152 => x"330eabcd",
  3153 => x"1234e66d",
  3154 => x"deec0005",
  3155 => x"000b0000",
  3156 => x"00000000",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"00000000",
  3161 => x"00000000",
  3162 => x"00000000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"00000000",
  3166 => x"00000000",
  3167 => x"00000000",
  3168 => x"00000000",
  3169 => x"00000000",
  3170 => x"00000000",
  3171 => x"00000000",
  3172 => x"00000000",
  3173 => x"00000000",
  3174 => x"00000000",
  3175 => x"00000000",
  3176 => x"00000000",
  3177 => x"00000000",
  3178 => x"00000000",
  3179 => x"00000000",
  3180 => x"00000000",
  3181 => x"00000000",
  3182 => x"00000000",
  3183 => x"00000000",
  3184 => x"00000000",
  3185 => x"00000000",
  3186 => x"00000000",
  3187 => x"00000000",
  3188 => x"00000000",
  3189 => x"00000000",
  3190 => x"00000000",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00000000",
  3195 => x"00000000",
  3196 => x"00000000",
  3197 => x"00000000",
  3198 => x"00000000",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"00000000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000000",
  3246 => x"00000000",
  3247 => x"00000000",
  3248 => x"00000000",
  3249 => x"00000000",
  3250 => x"00000000",
  3251 => x"00000000",
  3252 => x"00000000",
  3253 => x"00000000",
  3254 => x"00000000",
  3255 => x"00000000",
  3256 => x"00000000",
  3257 => x"00000000",
  3258 => x"00000000",
  3259 => x"00000000",
  3260 => x"00000000",
  3261 => x"00000000",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00000000",
  3265 => x"00000000",
  3266 => x"00000000",
  3267 => x"00000000",
  3268 => x"00000000",
  3269 => x"00000000",
  3270 => x"00000000",
  3271 => x"00000000",
  3272 => x"00000000",
  3273 => x"00000000",
  3274 => x"00000000",
  3275 => x"00000000",
  3276 => x"00000000",
  3277 => x"00000000",
  3278 => x"00000000",
  3279 => x"00000000",
  3280 => x"00000000",
  3281 => x"00000000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"00000000",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00000000",
  3288 => x"00000000",
  3289 => x"00000000",
  3290 => x"00000000",
  3291 => x"00000000",
  3292 => x"00000000",
  3293 => x"00000000",
  3294 => x"00000000",
  3295 => x"00000000",
  3296 => x"00000000",
  3297 => x"00000000",
  3298 => x"00000000",
  3299 => x"00000000",
  3300 => x"00000000",
  3301 => x"00000000",
  3302 => x"00000000",
  3303 => x"00000000",
  3304 => x"00000000",
  3305 => x"00000000",
  3306 => x"00000000",
  3307 => x"00000000",
  3308 => x"00000000",
  3309 => x"00000000",
  3310 => x"00000000",
  3311 => x"00000000",
  3312 => x"00000000",
  3313 => x"00000000",
  3314 => x"00000000",
  3315 => x"00000000",
  3316 => x"00000000",
  3317 => x"00000000",
  3318 => x"00000000",
  3319 => x"00000000",
  3320 => x"00000000",
  3321 => x"00000000",
  3322 => x"00000000",
  3323 => x"00000000",
  3324 => x"00000000",
  3325 => x"00000000",
  3326 => x"00000000",
  3327 => x"00000000",
  3328 => x"00000000",
  3329 => x"00000000",
  3330 => x"00000000",
  3331 => x"00000000",
  3332 => x"00000000",
  3333 => x"00000000",
  3334 => x"00000000",
  3335 => x"00000000",
  3336 => x"00000000",
  3337 => x"00000000",
  3338 => x"00000000",
  3339 => x"00000000",
  3340 => x"00000000",
  3341 => x"00000000",
  3342 => x"00000000",
  3343 => x"00000000",
  3344 => x"ffffffff",
  3345 => x"00000000",
  3346 => x"00020000",
  3347 => x"00000000",
  3348 => x"00000000",
  3349 => x"0000344c",
  3350 => x"0000344c",
  3351 => x"00003454",
  3352 => x"00003454",
  3353 => x"0000345c",
  3354 => x"0000345c",
  3355 => x"00003464",
  3356 => x"00003464",
  3357 => x"0000346c",
  3358 => x"0000346c",
  3359 => x"00003474",
  3360 => x"00003474",
  3361 => x"0000347c",
  3362 => x"0000347c",
  3363 => x"00003484",
  3364 => x"00003484",
  3365 => x"0000348c",
  3366 => x"0000348c",
  3367 => x"00003494",
  3368 => x"00003494",
  3369 => x"0000349c",
  3370 => x"0000349c",
  3371 => x"000034a4",
  3372 => x"000034a4",
  3373 => x"000034ac",
  3374 => x"000034ac",
  3375 => x"000034b4",
  3376 => x"000034b4",
  3377 => x"000034bc",
  3378 => x"000034bc",
  3379 => x"000034c4",
  3380 => x"000034c4",
  3381 => x"000034cc",
  3382 => x"000034cc",
  3383 => x"000034d4",
  3384 => x"000034d4",
  3385 => x"000034dc",
  3386 => x"000034dc",
  3387 => x"000034e4",
  3388 => x"000034e4",
  3389 => x"000034ec",
  3390 => x"000034ec",
  3391 => x"000034f4",
  3392 => x"000034f4",
  3393 => x"000034fc",
  3394 => x"000034fc",
  3395 => x"00003504",
  3396 => x"00003504",
  3397 => x"0000350c",
  3398 => x"0000350c",
  3399 => x"00003514",
  3400 => x"00003514",
  3401 => x"0000351c",
  3402 => x"0000351c",
  3403 => x"00003524",
  3404 => x"00003524",
  3405 => x"0000352c",
  3406 => x"0000352c",
  3407 => x"00003534",
  3408 => x"00003534",
  3409 => x"0000353c",
  3410 => x"0000353c",
  3411 => x"00003544",
  3412 => x"00003544",
  3413 => x"0000354c",
  3414 => x"0000354c",
  3415 => x"00003554",
  3416 => x"00003554",
  3417 => x"0000355c",
  3418 => x"0000355c",
  3419 => x"00003564",
  3420 => x"00003564",
  3421 => x"0000356c",
  3422 => x"0000356c",
  3423 => x"00003574",
  3424 => x"00003574",
  3425 => x"0000357c",
  3426 => x"0000357c",
  3427 => x"00003584",
  3428 => x"00003584",
  3429 => x"0000358c",
  3430 => x"0000358c",
  3431 => x"00003594",
  3432 => x"00003594",
  3433 => x"0000359c",
  3434 => x"0000359c",
  3435 => x"000035a4",
  3436 => x"000035a4",
  3437 => x"000035ac",
  3438 => x"000035ac",
  3439 => x"000035b4",
  3440 => x"000035b4",
  3441 => x"000035bc",
  3442 => x"000035bc",
  3443 => x"000035c4",
  3444 => x"000035c4",
  3445 => x"000035cc",
  3446 => x"000035cc",
  3447 => x"000035d4",
  3448 => x"000035d4",
  3449 => x"000035dc",
  3450 => x"000035dc",
  3451 => x"000035e4",
  3452 => x"000035e4",
  3453 => x"000035ec",
  3454 => x"000035ec",
  3455 => x"000035f4",
  3456 => x"000035f4",
  3457 => x"000035fc",
  3458 => x"000035fc",
  3459 => x"00003604",
  3460 => x"00003604",
  3461 => x"0000360c",
  3462 => x"0000360c",
  3463 => x"00003614",
  3464 => x"00003614",
  3465 => x"0000361c",
  3466 => x"0000361c",
  3467 => x"00003624",
  3468 => x"00003624",
  3469 => x"0000362c",
  3470 => x"0000362c",
  3471 => x"00003634",
  3472 => x"00003634",
  3473 => x"0000363c",
  3474 => x"0000363c",
  3475 => x"00003644",
  3476 => x"00003644",
  3477 => x"0000364c",
  3478 => x"0000364c",
  3479 => x"00003654",
  3480 => x"00003654",
  3481 => x"0000365c",
  3482 => x"0000365c",
  3483 => x"00003664",
  3484 => x"00003664",
  3485 => x"0000366c",
  3486 => x"0000366c",
  3487 => x"00003674",
  3488 => x"00003674",
  3489 => x"0000367c",
  3490 => x"0000367c",
  3491 => x"00003684",
  3492 => x"00003684",
  3493 => x"0000368c",
  3494 => x"0000368c",
  3495 => x"00003694",
  3496 => x"00003694",
  3497 => x"0000369c",
  3498 => x"0000369c",
  3499 => x"000036a4",
  3500 => x"000036a4",
  3501 => x"000036ac",
  3502 => x"000036ac",
  3503 => x"000036b4",
  3504 => x"000036b4",
  3505 => x"000036bc",
  3506 => x"000036bc",
  3507 => x"000036c4",
  3508 => x"000036c4",
  3509 => x"000036cc",
  3510 => x"000036cc",
  3511 => x"000036d4",
  3512 => x"000036d4",
  3513 => x"000036dc",
  3514 => x"000036dc",
  3515 => x"000036e4",
  3516 => x"000036e4",
  3517 => x"000036ec",
  3518 => x"000036ec",
  3519 => x"000036f4",
  3520 => x"000036f4",
  3521 => x"000036fc",
  3522 => x"000036fc",
  3523 => x"00003704",
  3524 => x"00003704",
  3525 => x"0000370c",
  3526 => x"0000370c",
  3527 => x"00003714",
  3528 => x"00003714",
  3529 => x"0000371c",
  3530 => x"0000371c",
  3531 => x"00003724",
  3532 => x"00003724",
  3533 => x"0000372c",
  3534 => x"0000372c",
  3535 => x"00003734",
  3536 => x"00003734",
  3537 => x"0000373c",
  3538 => x"0000373c",
  3539 => x"00003744",
  3540 => x"00003744",
  3541 => x"0000374c",
  3542 => x"0000374c",
  3543 => x"00003754",
  3544 => x"00003754",
  3545 => x"0000375c",
  3546 => x"0000375c",
  3547 => x"00003764",
  3548 => x"00003764",
  3549 => x"0000376c",
  3550 => x"0000376c",
  3551 => x"00003774",
  3552 => x"00003774",
  3553 => x"0000377c",
  3554 => x"0000377c",
  3555 => x"00003784",
  3556 => x"00003784",
  3557 => x"0000378c",
  3558 => x"0000378c",
  3559 => x"00003794",
  3560 => x"00003794",
  3561 => x"0000379c",
  3562 => x"0000379c",
  3563 => x"000037a4",
  3564 => x"000037a4",
  3565 => x"000037ac",
  3566 => x"000037ac",
  3567 => x"000037b4",
  3568 => x"000037b4",
  3569 => x"000037bc",
  3570 => x"000037bc",
  3571 => x"000037c4",
  3572 => x"000037c4",
  3573 => x"000037cc",
  3574 => x"000037cc",
  3575 => x"000037d4",
  3576 => x"000037d4",
  3577 => x"000037dc",
  3578 => x"000037dc",
  3579 => x"000037e4",
  3580 => x"000037e4",
  3581 => x"000037ec",
  3582 => x"000037ec",
  3583 => x"000037f4",
  3584 => x"000037f4",
  3585 => x"000037fc",
  3586 => x"000037fc",
  3587 => x"00003804",
  3588 => x"00003804",
  3589 => x"0000380c",
  3590 => x"0000380c",
  3591 => x"00003814",
  3592 => x"00003814",
  3593 => x"0000381c",
  3594 => x"0000381c",
  3595 => x"00003824",
  3596 => x"00003824",
  3597 => x"0000382c",
  3598 => x"0000382c",
  3599 => x"00003834",
  3600 => x"00003834",
  3601 => x"0000383c",
  3602 => x"0000383c",
  3603 => x"00003844",
  3604 => x"00003844",
  3605 => x"00003054",
  3606 => x"ffffffff",
  3607 => x"00000000",
  3608 => x"ffffffff",
  3609 => x"00000000",
  3610 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
