-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80e5f80c",
     3 => x"3a0b0b80",
     4 => x"def50400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80dfbe2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80e5",
   162 => x"e4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80c2",
   171 => x"dc2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80c4",
   179 => x"8e2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80e5f40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"d8df3f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80e5f408",
   281 => x"802ea438",
   282 => x"80e5f808",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80f5",
   286 => x"f40c82a0",
   287 => x"800b80f5",
   288 => x"f80c8290",
   289 => x"800b80f5",
   290 => x"fc0c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"f5f40cf8",
   294 => x"80808280",
   295 => x"0b80f5f8",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"f5fc0c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80f5f40c",
   302 => x"80c0a880",
   303 => x"940b80f5",
   304 => x"f80c0b0b",
   305 => x"80e1940b",
   306 => x"80f5fc0c",
   307 => x"04ff3d0d",
   308 => x"80f68033",
   309 => x"5170a738",
   310 => x"80e68008",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"e6800c70",
   315 => x"2d80e680",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80f6",
   319 => x"8034833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80f5f008",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"f5f0510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404fd3d",
   333 => x"0d80e68c",
   334 => x"0876b0ea",
   335 => x"2994120c",
   336 => x"54850b98",
   337 => x"150c9814",
   338 => x"08708106",
   339 => x"515372f6",
   340 => x"38853d0d",
   341 => x"04ff3d0d",
   342 => x"80e68c08",
   343 => x"74101075",
   344 => x"10059412",
   345 => x"0c52850b",
   346 => x"98130c98",
   347 => x"12087081",
   348 => x"06515170",
   349 => x"f638833d",
   350 => x"0d04803d",
   351 => x"0d725180",
   352 => x"71278738",
   353 => x"ff115170",
   354 => x"fb38823d",
   355 => x"0d04803d",
   356 => x"0d80e68c",
   357 => x"0851870b",
   358 => x"84120c82",
   359 => x"3d0d0480",
   360 => x"3d0d80e6",
   361 => x"900851b6",
   362 => x"0b8c120c",
   363 => x"830b8812",
   364 => x"0c823d0d",
   365 => x"04ff3d0d",
   366 => x"80e69008",
   367 => x"52841208",
   368 => x"70810651",
   369 => x"5170802e",
   370 => x"f4387108",
   371 => x"7081ff06",
   372 => x"800c5183",
   373 => x"3d0d04fe",
   374 => x"3d0d0293",
   375 => x"053380e6",
   376 => x"90085353",
   377 => x"84120870",
   378 => x"822a7081",
   379 => x"06515151",
   380 => x"70802ef0",
   381 => x"3872720c",
   382 => x"843d0d04",
   383 => x"fe3d0d02",
   384 => x"93053353",
   385 => x"728a2e9e",
   386 => x"3880e690",
   387 => x"08528412",
   388 => x"0870822a",
   389 => x"70810651",
   390 => x"51517080",
   391 => x"2ef03872",
   392 => x"720c843d",
   393 => x"0d0480e6",
   394 => x"90085284",
   395 => x"12087082",
   396 => x"2a708106",
   397 => x"51515170",
   398 => x"802ef038",
   399 => x"8d720c84",
   400 => x"12087082",
   401 => x"2a708106",
   402 => x"51515170",
   403 => x"802effbe",
   404 => x"38cd39fd",
   405 => x"3d0d7570",
   406 => x"33525470",
   407 => x"802eaa38",
   408 => x"7080e690",
   409 => x"08535381",
   410 => x"1454728a",
   411 => x"2e9f3884",
   412 => x"12087082",
   413 => x"2a708106",
   414 => x"51515170",
   415 => x"802ef038",
   416 => x"72720c73",
   417 => x"335372df",
   418 => x"38853d0d",
   419 => x"04841208",
   420 => x"70822a70",
   421 => x"81065151",
   422 => x"5170802e",
   423 => x"f0388d72",
   424 => x"0c841208",
   425 => x"70822a70",
   426 => x"81065151",
   427 => x"5170802e",
   428 => x"ffbd38cc",
   429 => x"39f53d0d",
   430 => x"7e028405",
   431 => x"b705338c",
   432 => x"3d5b5557",
   433 => x"8b5380e1",
   434 => x"98527851",
   435 => x"b9973f82",
   436 => x"5673882e",
   437 => x"96388456",
   438 => x"73902e8f",
   439 => x"38885673",
   440 => x"a02e8838",
   441 => x"74567480",
   442 => x"2ea73802",
   443 => x"a5055876",
   444 => x"8f065473",
   445 => x"892680ce",
   446 => x"387518b0",
   447 => x"15555573",
   448 => x"75347684",
   449 => x"2aff1770",
   450 => x"81ff0658",
   451 => x"555775df",
   452 => x"38787933",
   453 => x"55577380",
   454 => x"2ea83873",
   455 => x"80e69008",
   456 => x"56568117",
   457 => x"57758a2e",
   458 => x"b9388415",
   459 => x"0870822a",
   460 => x"81065954",
   461 => x"77802ef2",
   462 => x"3875750c",
   463 => x"76335675",
   464 => x"e1388d3d",
   465 => x"0d047518",
   466 => x"b7155555",
   467 => x"73753476",
   468 => x"842aff17",
   469 => x"7081ff06",
   470 => x"58555775",
   471 => x"ff9138ff",
   472 => x"b0398415",
   473 => x"0870822a",
   474 => x"81065954",
   475 => x"77802ef2",
   476 => x"388d750c",
   477 => x"84150870",
   478 => x"822a8106",
   479 => x"59547780",
   480 => x"2effa738",
   481 => x"ffb339f8",
   482 => x"3d0d7a7c",
   483 => x"59538073",
   484 => x"56577673",
   485 => x"2480dc38",
   486 => x"7717548a",
   487 => x"527451b3",
   488 => x"963f8008",
   489 => x"b0055372",
   490 => x"74348117",
   491 => x"578a5274",
   492 => x"51b2df3f",
   493 => x"80085580",
   494 => x"08de3880",
   495 => x"08779f2a",
   496 => x"1870812c",
   497 => x"5b565680",
   498 => x"79259e38",
   499 => x"7717ff05",
   500 => x"55751870",
   501 => x"33555374",
   502 => x"33733473",
   503 => x"75348116",
   504 => x"ff165656",
   505 => x"787624e9",
   506 => x"38761856",
   507 => x"8076348a",
   508 => x"3d0d04ad",
   509 => x"78708105",
   510 => x"5a347230",
   511 => x"78185555",
   512 => x"8a527451",
   513 => x"b2b13f80",
   514 => x"08b00553",
   515 => x"72743481",
   516 => x"17578a52",
   517 => x"7451b1fa",
   518 => x"3f800855",
   519 => x"8008fef8",
   520 => x"38ff9839",
   521 => x"803d0d80",
   522 => x"e6880851",
   523 => x"81ff0b88",
   524 => x"120c823d",
   525 => x"0d04f83d",
   526 => x"0d7a59f8",
   527 => x"81c08e80",
   528 => x"55a00b80",
   529 => x"e6880880",
   530 => x"e68c085a",
   531 => x"58567484",
   532 => x"180c749f",
   533 => x"2a751007",
   534 => x"5578802e",
   535 => x"97387580",
   536 => x"2ebb38ff",
   537 => x"16758419",
   538 => x"0c759f2a",
   539 => x"76100756",
   540 => x"5678eb38",
   541 => x"7754afd7",
   542 => x"c20b9419",
   543 => x"0c850b98",
   544 => x"190c9814",
   545 => x"08708106",
   546 => x"51537280",
   547 => x"2ec03898",
   548 => x"14087081",
   549 => x"06515372",
   550 => x"e938ffb2",
   551 => x"398a3d0d",
   552 => x"04fd3d0d",
   553 => x"80e68808",
   554 => x"5480d50b",
   555 => x"84150c80",
   556 => x"e6900852",
   557 => x"84120881",
   558 => x"06517080",
   559 => x"2ef63871",
   560 => x"087081ff",
   561 => x"06f61152",
   562 => x"545170ae",
   563 => x"268c3870",
   564 => x"101080e4",
   565 => x"98055170",
   566 => x"08048412",
   567 => x"0870822a",
   568 => x"70810651",
   569 => x"51517080",
   570 => x"2ef038ab",
   571 => x"720c728a",
   572 => x"2eaa3884",
   573 => x"12087082",
   574 => x"2a708106",
   575 => x"51515170",
   576 => x"802ef038",
   577 => x"72720c84",
   578 => x"12087082",
   579 => x"2a810651",
   580 => x"5372802e",
   581 => x"f238ad72",
   582 => x"0cff9939",
   583 => x"84120870",
   584 => x"822a7081",
   585 => x"06515151",
   586 => x"70802ef0",
   587 => x"388d720c",
   588 => x"84120870",
   589 => x"822a7081",
   590 => x"06515151",
   591 => x"70802eff",
   592 => x"b238c139",
   593 => x"81ff0b84",
   594 => x"150cfee8",
   595 => x"3980ff0b",
   596 => x"84150cfe",
   597 => x"df39bf0b",
   598 => x"84150cfe",
   599 => x"d7399f0b",
   600 => x"84150cfe",
   601 => x"cf398f0b",
   602 => x"84150cfe",
   603 => x"c739870b",
   604 => x"84150cfe",
   605 => x"bf39830b",
   606 => x"84150cfe",
   607 => x"b739810b",
   608 => x"84150cfe",
   609 => x"af39800b",
   610 => x"84150cfe",
   611 => x"a739ff3d",
   612 => x"0d80e688",
   613 => x"08527108",
   614 => x"708f0670",
   615 => x"71842b07",
   616 => x"84150c51",
   617 => x"51710870",
   618 => x"8f067071",
   619 => x"842b0784",
   620 => x"150c5151",
   621 => x"e139fc3d",
   622 => x"0d029a05",
   623 => x"22028405",
   624 => x"9e052202",
   625 => x"8805a205",
   626 => x"2280e684",
   627 => x"08555654",
   628 => x"55901208",
   629 => x"70832a70",
   630 => x"81065151",
   631 => x"5170f238",
   632 => x"74902b73",
   633 => x"8b2b0774",
   634 => x"862b0781",
   635 => x"0790130c",
   636 => x"863d0d04",
   637 => x"fd3d0d02",
   638 => x"96052202",
   639 => x"84059a05",
   640 => x"2280e684",
   641 => x"08545454",
   642 => x"90120870",
   643 => x"832a7081",
   644 => x"06515151",
   645 => x"70f23873",
   646 => x"8b2b7386",
   647 => x"2b078207",
   648 => x"90130c90",
   649 => x"12087083",
   650 => x"2a810655",
   651 => x"5173f438",
   652 => x"90120870",
   653 => x"902a800c",
   654 => x"54853d0d",
   655 => x"04ff3d0d",
   656 => x"80e68408",
   657 => x"52ff0b84",
   658 => x"130cfc94",
   659 => x"800b8813",
   660 => x"0c82d0af",
   661 => x"fdfb0b8c",
   662 => x"130c80c0",
   663 => x"720c7108",
   664 => x"70862a70",
   665 => x"81065151",
   666 => x"5170f338",
   667 => x"90120870",
   668 => x"832a7081",
   669 => x"06515151",
   670 => x"70f23881",
   671 => x"fc80810b",
   672 => x"90130c90",
   673 => x"12087083",
   674 => x"2a708106",
   675 => x"51515170",
   676 => x"f23880fd",
   677 => x"c0810b90",
   678 => x"130c833d",
   679 => x"0d04d53d",
   680 => x"0d80e684",
   681 => x"0858ff0b",
   682 => x"84190cfc",
   683 => x"809b0b88",
   684 => x"190c828b",
   685 => x"a1968a0b",
   686 => x"8c190ca4",
   687 => x"b40b9419",
   688 => x"0c8186a1",
   689 => x"0b98190c",
   690 => x"80e1a40b",
   691 => x"80e1a433",
   692 => x"55577380",
   693 => x"2ea93873",
   694 => x"80e69008",
   695 => x"56568117",
   696 => x"57758a2e",
   697 => x"8de73884",
   698 => x"15087082",
   699 => x"2a810651",
   700 => x"5978802e",
   701 => x"f2387575",
   702 => x"0c763356",
   703 => x"75e03880",
   704 => x"e1b80b80",
   705 => x"e1b83355",
   706 => x"5773802e",
   707 => x"a93880e6",
   708 => x"90087457",
   709 => x"55811757",
   710 => x"758a2e8d",
   711 => x"d5388415",
   712 => x"0870822a",
   713 => x"81065159",
   714 => x"78802ef2",
   715 => x"3875750c",
   716 => x"76335675",
   717 => x"e0387708",
   718 => x"a63d5a56",
   719 => x"8b5380e1",
   720 => x"98527851",
   721 => x"b09f3f88",
   722 => x"02840581",
   723 => x"91055957",
   724 => x"758f0654",
   725 => x"7389268d",
   726 => x"be387618",
   727 => x"b0155555",
   728 => x"73753475",
   729 => x"842aff18",
   730 => x"7081ff06",
   731 => x"59565676",
   732 => x"df387879",
   733 => x"33555773",
   734 => x"802ea938",
   735 => x"80e69008",
   736 => x"74575581",
   737 => x"1757758a",
   738 => x"2e8da838",
   739 => x"84150870",
   740 => x"822a8106",
   741 => x"59597780",
   742 => x"2ef23875",
   743 => x"750c7633",
   744 => x"5675e038",
   745 => x"80e1c80b",
   746 => x"80e1c833",
   747 => x"55577380",
   748 => x"2ea93880",
   749 => x"e6900874",
   750 => x"57558117",
   751 => x"57758a2e",
   752 => x"8d963884",
   753 => x"15087082",
   754 => x"2a810659",
   755 => x"5977802e",
   756 => x"f2387575",
   757 => x"0c763356",
   758 => x"75e03880",
   759 => x"e6840884",
   760 => x"1108a43d",
   761 => x"5b57578b",
   762 => x"5380e198",
   763 => x"527851ae",
   764 => x"f43f8802",
   765 => x"84058185",
   766 => x"05595775",
   767 => x"8f065473",
   768 => x"892692b6",
   769 => x"387618b0",
   770 => x"15555573",
   771 => x"75347584",
   772 => x"2aff1870",
   773 => x"81ff0659",
   774 => x"565676df",
   775 => x"38787933",
   776 => x"55577380",
   777 => x"2ea93880",
   778 => x"e6900874",
   779 => x"57558117",
   780 => x"57758a2e",
   781 => x"8cc73884",
   782 => x"15087082",
   783 => x"2a810659",
   784 => x"5977802e",
   785 => x"f2387575",
   786 => x"0c763356",
   787 => x"75e03880",
   788 => x"e1d80b80",
   789 => x"e1d83355",
   790 => x"5773802e",
   791 => x"a93880e6",
   792 => x"90087457",
   793 => x"55811757",
   794 => x"758a2e8c",
   795 => x"b5388415",
   796 => x"0870822a",
   797 => x"81065959",
   798 => x"77802ef2",
   799 => x"3875750c",
   800 => x"76335675",
   801 => x"e03880e6",
   802 => x"84088811",
   803 => x"08a13d5b",
   804 => x"57578b53",
   805 => x"80e19852",
   806 => x"7851adc9",
   807 => x"3f880284",
   808 => x"0580f905",
   809 => x"5957758f",
   810 => x"06547389",
   811 => x"26918238",
   812 => x"7618b015",
   813 => x"55557375",
   814 => x"3475842a",
   815 => x"ff187081",
   816 => x"ff065956",
   817 => x"5676df38",
   818 => x"78793355",
   819 => x"5773802e",
   820 => x"a93880e6",
   821 => x"90087457",
   822 => x"55811757",
   823 => x"758a2e8b",
   824 => x"e6388415",
   825 => x"0870822a",
   826 => x"81065959",
   827 => x"77802ef2",
   828 => x"3875750c",
   829 => x"76335675",
   830 => x"e03880e1",
   831 => x"e80b80e1",
   832 => x"e8335557",
   833 => x"73802ea9",
   834 => x"3880e690",
   835 => x"08745755",
   836 => x"81175775",
   837 => x"8a2e8bd4",
   838 => x"38841508",
   839 => x"70822a81",
   840 => x"06595977",
   841 => x"802ef238",
   842 => x"75750c76",
   843 => x"335675e0",
   844 => x"3880e684",
   845 => x"088c1108",
   846 => x"9e3d5b57",
   847 => x"578b5380",
   848 => x"e1985278",
   849 => x"51ac9e3f",
   850 => x"88028405",
   851 => x"80ed0559",
   852 => x"57758f06",
   853 => x"54738926",
   854 => x"8fce3876",
   855 => x"18b01555",
   856 => x"55737534",
   857 => x"75842aff",
   858 => x"187081ff",
   859 => x"06595656",
   860 => x"76df3878",
   861 => x"79335557",
   862 => x"73802ea9",
   863 => x"3880e690",
   864 => x"08745755",
   865 => x"81175775",
   866 => x"8a2e8b85",
   867 => x"38841508",
   868 => x"70822a81",
   869 => x"06595977",
   870 => x"802ef238",
   871 => x"75750c76",
   872 => x"335675e0",
   873 => x"3880e1f8",
   874 => x"0b80e1f8",
   875 => x"33555773",
   876 => x"802ea938",
   877 => x"80e69008",
   878 => x"74575581",
   879 => x"1757758a",
   880 => x"2e8af338",
   881 => x"84150870",
   882 => x"822a8106",
   883 => x"59597780",
   884 => x"2ef23875",
   885 => x"750c7633",
   886 => x"5675e038",
   887 => x"80e68408",
   888 => x"9011089b",
   889 => x"3d5b5757",
   890 => x"8b5380e1",
   891 => x"98527851",
   892 => x"aaf33f88",
   893 => x"02840580",
   894 => x"e1055957",
   895 => x"758f0654",
   896 => x"7389268e",
   897 => x"9a387618",
   898 => x"b0155555",
   899 => x"73753475",
   900 => x"842aff18",
   901 => x"7081ff06",
   902 => x"59565676",
   903 => x"df387879",
   904 => x"33555773",
   905 => x"802ea938",
   906 => x"80e69008",
   907 => x"74575581",
   908 => x"1757758a",
   909 => x"2e8aa438",
   910 => x"84150870",
   911 => x"822a8106",
   912 => x"59597780",
   913 => x"2ef23875",
   914 => x"750c7633",
   915 => x"5675e038",
   916 => x"80e2880b",
   917 => x"80e28833",
   918 => x"55577380",
   919 => x"2ea93880",
   920 => x"e6900874",
   921 => x"57558117",
   922 => x"57758a2e",
   923 => x"8a923884",
   924 => x"15087082",
   925 => x"2a810659",
   926 => x"5977802e",
   927 => x"f2387575",
   928 => x"0c763356",
   929 => x"75e03880",
   930 => x"e6840894",
   931 => x"1108983d",
   932 => x"5b57578b",
   933 => x"5380e198",
   934 => x"527851a9",
   935 => x"c83f8802",
   936 => x"840580d5",
   937 => x"05595775",
   938 => x"8f065473",
   939 => x"89268ce6",
   940 => x"387618b0",
   941 => x"15555573",
   942 => x"75347584",
   943 => x"2aff1870",
   944 => x"81ff0659",
   945 => x"565676df",
   946 => x"38787933",
   947 => x"55577380",
   948 => x"2ea93880",
   949 => x"e6900874",
   950 => x"57558117",
   951 => x"57758a2e",
   952 => x"89c33884",
   953 => x"15087082",
   954 => x"2a810659",
   955 => x"5977802e",
   956 => x"f2387575",
   957 => x"0c763356",
   958 => x"75e03880",
   959 => x"e2980b80",
   960 => x"e2983355",
   961 => x"5773802e",
   962 => x"a93880e6",
   963 => x"90087457",
   964 => x"55811757",
   965 => x"758a2e89",
   966 => x"b1388415",
   967 => x"0870822a",
   968 => x"81065959",
   969 => x"77802ef2",
   970 => x"3875750c",
   971 => x"76335675",
   972 => x"e03880e6",
   973 => x"84089811",
   974 => x"08953d5b",
   975 => x"57578b53",
   976 => x"80e19852",
   977 => x"7851a89d",
   978 => x"3f880284",
   979 => x"0580c905",
   980 => x"5957758f",
   981 => x"06547389",
   982 => x"268bb238",
   983 => x"7618b015",
   984 => x"55557375",
   985 => x"3475842a",
   986 => x"ff187081",
   987 => x"ff065956",
   988 => x"5676df38",
   989 => x"78793355",
   990 => x"5773802e",
   991 => x"a93880e6",
   992 => x"90087457",
   993 => x"55811757",
   994 => x"758a2e88",
   995 => x"e2388415",
   996 => x"0870822a",
   997 => x"81065959",
   998 => x"77802ef2",
   999 => x"3875750c",
  1000 => x"76335675",
  1001 => x"e03880e2",
  1002 => x"a80b80e2",
  1003 => x"a8335557",
  1004 => x"73802ea9",
  1005 => x"3880e690",
  1006 => x"08745755",
  1007 => x"81175775",
  1008 => x"8a2e88d0",
  1009 => x"38841508",
  1010 => x"70822a81",
  1011 => x"06595977",
  1012 => x"802ef238",
  1013 => x"75750c76",
  1014 => x"335675e0",
  1015 => x"3880e684",
  1016 => x"089c1108",
  1017 => x"923d5b57",
  1018 => x"578b5380",
  1019 => x"e1985278",
  1020 => x"51a6f23f",
  1021 => x"88028405",
  1022 => x"bd055957",
  1023 => x"758f0654",
  1024 => x"73892689",
  1025 => x"ff387618",
  1026 => x"b0155555",
  1027 => x"73753475",
  1028 => x"842aff18",
  1029 => x"7081ff06",
  1030 => x"59565676",
  1031 => x"df387879",
  1032 => x"33555773",
  1033 => x"802ea938",
  1034 => x"80e69008",
  1035 => x"74575581",
  1036 => x"1757758a",
  1037 => x"2e888238",
  1038 => x"84150870",
  1039 => x"822a8106",
  1040 => x"59597780",
  1041 => x"2ef23875",
  1042 => x"750c7633",
  1043 => x"5675e038",
  1044 => x"80e2b80b",
  1045 => x"80e2b833",
  1046 => x"55577380",
  1047 => x"2ea93880",
  1048 => x"e6900874",
  1049 => x"57558117",
  1050 => x"57758a2e",
  1051 => x"87f03884",
  1052 => x"15087082",
  1053 => x"2a810659",
  1054 => x"5977802e",
  1055 => x"f2387575",
  1056 => x"0c763356",
  1057 => x"75e03880",
  1058 => x"e68408a0",
  1059 => x"11088f3d",
  1060 => x"5b57578b",
  1061 => x"5380e198",
  1062 => x"527851a5",
  1063 => x"c83f8802",
  1064 => x"8405b105",
  1065 => x"5957758f",
  1066 => x"06547389",
  1067 => x"2688cc38",
  1068 => x"7618b015",
  1069 => x"55557375",
  1070 => x"3475842a",
  1071 => x"ff187081",
  1072 => x"ff065956",
  1073 => x"5676df38",
  1074 => x"78793355",
  1075 => x"5773802e",
  1076 => x"a93880e6",
  1077 => x"90087457",
  1078 => x"55811757",
  1079 => x"758a2e87",
  1080 => x"a2388415",
  1081 => x"0870822a",
  1082 => x"81065959",
  1083 => x"77802ef2",
  1084 => x"3875750c",
  1085 => x"76335675",
  1086 => x"e03880e2",
  1087 => x"c80b80e2",
  1088 => x"c8335557",
  1089 => x"73802ea9",
  1090 => x"3880e690",
  1091 => x"08745755",
  1092 => x"81175775",
  1093 => x"8a2e8790",
  1094 => x"38841508",
  1095 => x"70822a81",
  1096 => x"06595977",
  1097 => x"802ef238",
  1098 => x"75750c76",
  1099 => x"335675e0",
  1100 => x"3880e684",
  1101 => x"08a41108",
  1102 => x"8c3d5b57",
  1103 => x"578b5380",
  1104 => x"e1985278",
  1105 => x"51a49e3f",
  1106 => x"88028405",
  1107 => x"a5055957",
  1108 => x"758f0654",
  1109 => x"73892687",
  1110 => x"99387618",
  1111 => x"b0155555",
  1112 => x"73753475",
  1113 => x"842aff18",
  1114 => x"7081ff06",
  1115 => x"59565676",
  1116 => x"df387879",
  1117 => x"33555773",
  1118 => x"802e87c7",
  1119 => x"3880e690",
  1120 => x"08745755",
  1121 => x"81175775",
  1122 => x"8a2e86c1",
  1123 => x"38841508",
  1124 => x"70822a81",
  1125 => x"06595977",
  1126 => x"802ef238",
  1127 => x"75750c76",
  1128 => x"335675e0",
  1129 => x"38841508",
  1130 => x"70822a81",
  1131 => x"06575875",
  1132 => x"802ef238",
  1133 => x"8d750c84",
  1134 => x"15087082",
  1135 => x"2a810655",
  1136 => x"5673802e",
  1137 => x"f2388a75",
  1138 => x"0cad3d0d",
  1139 => x"04841508",
  1140 => x"70822a81",
  1141 => x"06515473",
  1142 => x"802ef238",
  1143 => x"8d750c84",
  1144 => x"15087082",
  1145 => x"2a810651",
  1146 => x"5978802e",
  1147 => x"f1f938f2",
  1148 => x"85398415",
  1149 => x"0870822a",
  1150 => x"81065154",
  1151 => x"73802ef2",
  1152 => x"388d750c",
  1153 => x"84150870",
  1154 => x"822a8106",
  1155 => x"51597880",
  1156 => x"2ef28b38",
  1157 => x"f2973976",
  1158 => x"18b71555",
  1159 => x"55737534",
  1160 => x"75842aff",
  1161 => x"187081ff",
  1162 => x"06595656",
  1163 => x"76f2a138",
  1164 => x"f2c03984",
  1165 => x"15087082",
  1166 => x"2a810659",
  1167 => x"5977802e",
  1168 => x"f2388d75",
  1169 => x"0c841508",
  1170 => x"70822a81",
  1171 => x"06595977",
  1172 => x"802ef2b8",
  1173 => x"38f2c439",
  1174 => x"84150870",
  1175 => x"822a8106",
  1176 => x"59597780",
  1177 => x"2ef2388d",
  1178 => x"750c8415",
  1179 => x"0870822a",
  1180 => x"81065959",
  1181 => x"77802ef2",
  1182 => x"ca38f2d6",
  1183 => x"39841508",
  1184 => x"70822a81",
  1185 => x"06595977",
  1186 => x"802ef238",
  1187 => x"8d750c84",
  1188 => x"15087082",
  1189 => x"2a810659",
  1190 => x"5977802e",
  1191 => x"f39938f3",
  1192 => x"a5398415",
  1193 => x"0870822a",
  1194 => x"81065959",
  1195 => x"77802ef2",
  1196 => x"388d750c",
  1197 => x"84150870",
  1198 => x"822a8106",
  1199 => x"59597780",
  1200 => x"2ef3ab38",
  1201 => x"f3b73984",
  1202 => x"15087082",
  1203 => x"2a810659",
  1204 => x"5977802e",
  1205 => x"f2388d75",
  1206 => x"0c841508",
  1207 => x"70822a81",
  1208 => x"06595977",
  1209 => x"802ef3fa",
  1210 => x"38f48639",
  1211 => x"84150870",
  1212 => x"822a8106",
  1213 => x"59597780",
  1214 => x"2ef2388d",
  1215 => x"750c8415",
  1216 => x"0870822a",
  1217 => x"81065959",
  1218 => x"77802ef4",
  1219 => x"8c38f498",
  1220 => x"39841508",
  1221 => x"70822a81",
  1222 => x"06595977",
  1223 => x"802ef238",
  1224 => x"8d750c84",
  1225 => x"15087082",
  1226 => x"2a810659",
  1227 => x"5977802e",
  1228 => x"f4db38f4",
  1229 => x"e7398415",
  1230 => x"0870822a",
  1231 => x"81065959",
  1232 => x"77802ef2",
  1233 => x"388d750c",
  1234 => x"84150870",
  1235 => x"822a8106",
  1236 => x"59597780",
  1237 => x"2ef4ed38",
  1238 => x"f4f93984",
  1239 => x"15087082",
  1240 => x"2a810659",
  1241 => x"5977802e",
  1242 => x"f2388d75",
  1243 => x"0c841508",
  1244 => x"70822a81",
  1245 => x"06595977",
  1246 => x"802ef5bc",
  1247 => x"38f5c839",
  1248 => x"84150870",
  1249 => x"822a8106",
  1250 => x"59597780",
  1251 => x"2ef2388d",
  1252 => x"750c8415",
  1253 => x"0870822a",
  1254 => x"81065959",
  1255 => x"77802ef5",
  1256 => x"ce38f5da",
  1257 => x"39841508",
  1258 => x"70822a81",
  1259 => x"06595977",
  1260 => x"802ef238",
  1261 => x"8d750c84",
  1262 => x"15087082",
  1263 => x"2a810659",
  1264 => x"5977802e",
  1265 => x"f69d38f6",
  1266 => x"a9398415",
  1267 => x"0870822a",
  1268 => x"81065959",
  1269 => x"77802ef2",
  1270 => x"388d750c",
  1271 => x"84150870",
  1272 => x"822a8106",
  1273 => x"59597780",
  1274 => x"2ef6af38",
  1275 => x"f6bb3984",
  1276 => x"15087082",
  1277 => x"2a810659",
  1278 => x"5977802e",
  1279 => x"f2388d75",
  1280 => x"0c841508",
  1281 => x"70822a81",
  1282 => x"06595977",
  1283 => x"802ef6fe",
  1284 => x"38f78a39",
  1285 => x"84150870",
  1286 => x"822a8106",
  1287 => x"59597780",
  1288 => x"2ef2388d",
  1289 => x"750c8415",
  1290 => x"0870822a",
  1291 => x"81065959",
  1292 => x"77802ef7",
  1293 => x"9038f79c",
  1294 => x"39841508",
  1295 => x"70822a81",
  1296 => x"06595977",
  1297 => x"802ef238",
  1298 => x"8d750c84",
  1299 => x"15087082",
  1300 => x"2a810659",
  1301 => x"5977802e",
  1302 => x"f7de38f7",
  1303 => x"ea398415",
  1304 => x"0870822a",
  1305 => x"81065959",
  1306 => x"77802ef2",
  1307 => x"388d750c",
  1308 => x"84150870",
  1309 => x"822a8106",
  1310 => x"59597780",
  1311 => x"2ef7f038",
  1312 => x"f7fc3984",
  1313 => x"15087082",
  1314 => x"2a810659",
  1315 => x"5977802e",
  1316 => x"f2388d75",
  1317 => x"0c841508",
  1318 => x"70822a81",
  1319 => x"06595977",
  1320 => x"802ef8be",
  1321 => x"38f8ca39",
  1322 => x"84150870",
  1323 => x"822a8106",
  1324 => x"59597780",
  1325 => x"2ef2388d",
  1326 => x"750c8415",
  1327 => x"0870822a",
  1328 => x"81065959",
  1329 => x"77802ef8",
  1330 => x"d038f8dc",
  1331 => x"39841508",
  1332 => x"70822a81",
  1333 => x"06595977",
  1334 => x"802ef238",
  1335 => x"8d750c84",
  1336 => x"15087082",
  1337 => x"2a810659",
  1338 => x"5977802e",
  1339 => x"f99f38f9",
  1340 => x"ab397618",
  1341 => x"b7155555",
  1342 => x"f8e63976",
  1343 => x"18b71555",
  1344 => x"55f7b339",
  1345 => x"7618b715",
  1346 => x"5555f680",
  1347 => x"397618b7",
  1348 => x"155555f4",
  1349 => x"cd397618",
  1350 => x"b7155555",
  1351 => x"f3993976",
  1352 => x"18b71555",
  1353 => x"55f1e539",
  1354 => x"7618b715",
  1355 => x"5555f0b1",
  1356 => x"397618b7",
  1357 => x"155555ee",
  1358 => x"fd397618",
  1359 => x"b7155555",
  1360 => x"edc93980",
  1361 => x"e6900884",
  1362 => x"11087082",
  1363 => x"2a810658",
  1364 => x"59557580",
  1365 => x"2ef8ce38",
  1366 => x"f8da39e4",
  1367 => x"3d0d80e2",
  1368 => x"d80b80e2",
  1369 => x"d8335557",
  1370 => x"73802ea9",
  1371 => x"387380e6",
  1372 => x"90085656",
  1373 => x"81175775",
  1374 => x"8a2e85c3",
  1375 => x"38841508",
  1376 => x"70822a81",
  1377 => x"065b5c79",
  1378 => x"802ef238",
  1379 => x"75750c76",
  1380 => x"335675e0",
  1381 => x"389f0b97",
  1382 => x"3d028805",
  1383 => x"80d5059c",
  1384 => x"3d973d02",
  1385 => x"940580c9",
  1386 => x"05414440",
  1387 => x"44425f80",
  1388 => x"e2ec0b80",
  1389 => x"e2ec3355",
  1390 => x"5773802e",
  1391 => x"a93880e6",
  1392 => x"90087457",
  1393 => x"55811757",
  1394 => x"758a2e85",
  1395 => x"97388415",
  1396 => x"0870822a",
  1397 => x"81065a5b",
  1398 => x"78802ef2",
  1399 => x"3875750c",
  1400 => x"76335675",
  1401 => x"e0387e56",
  1402 => x"8b5380e1",
  1403 => x"98526051",
  1404 => x"9af33f82",
  1405 => x"57758f06",
  1406 => x"54738926",
  1407 => x"858b3861",
  1408 => x"17b01555",
  1409 => x"55737534",
  1410 => x"75842aff",
  1411 => x"187081ff",
  1412 => x"06595656",
  1413 => x"76df3860",
  1414 => x"61335557",
  1415 => x"73802ea9",
  1416 => x"3880e690",
  1417 => x"08745755",
  1418 => x"81175775",
  1419 => x"8a2e84f5",
  1420 => x"38841508",
  1421 => x"70822a81",
  1422 => x"065a5b78",
  1423 => x"802ef238",
  1424 => x"75750c76",
  1425 => x"335675e0",
  1426 => x"38807f83",
  1427 => x"ffff065f",
  1428 => x"5b7a872e",
  1429 => x"86c8387a",
  1430 => x"932e86c7",
  1431 => x"387a982e",
  1432 => x"86ae3880",
  1433 => x"e2fc0b80",
  1434 => x"e2fc3355",
  1435 => x"5773802e",
  1436 => x"a93880e6",
  1437 => x"90087457",
  1438 => x"55811757",
  1439 => x"758a2e84",
  1440 => x"c9388415",
  1441 => x"0870822a",
  1442 => x"81065b58",
  1443 => x"79802ef2",
  1444 => x"3875750c",
  1445 => x"76335675",
  1446 => x"e0387c5a",
  1447 => x"807b5758",
  1448 => x"777b2485",
  1449 => x"b9387918",
  1450 => x"578a5275",
  1451 => x"5195883f",
  1452 => x"8008b005",
  1453 => x"55747734",
  1454 => x"8118588a",
  1455 => x"52755194",
  1456 => x"d13f8008",
  1457 => x"568008de",
  1458 => x"38800878",
  1459 => x"9f2a1970",
  1460 => x"812c5b57",
  1461 => x"57807925",
  1462 => x"9e387918",
  1463 => x"ff055676",
  1464 => x"1a703356",
  1465 => x"54753374",
  1466 => x"34747634",
  1467 => x"8117ff17",
  1468 => x"57577877",
  1469 => x"24e93877",
  1470 => x"1a598079",
  1471 => x"347c7d33",
  1472 => x"55577380",
  1473 => x"2ea93880",
  1474 => x"e6900874",
  1475 => x"57558117",
  1476 => x"57758a2e",
  1477 => x"83d93884",
  1478 => x"15087082",
  1479 => x"2a81065a",
  1480 => x"5878802e",
  1481 => x"f2387575",
  1482 => x"0c763356",
  1483 => x"75e03880",
  1484 => x"e3880b80",
  1485 => x"e3883355",
  1486 => x"5773802e",
  1487 => x"a93880e6",
  1488 => x"90087457",
  1489 => x"55811757",
  1490 => x"758a2e83",
  1491 => x"c7388415",
  1492 => x"0870822a",
  1493 => x"81065959",
  1494 => x"77802ef2",
  1495 => x"3875750c",
  1496 => x"76335675",
  1497 => x"e0387a83",
  1498 => x"ffff0680",
  1499 => x"e6840856",
  1500 => x"56901508",
  1501 => x"70832a81",
  1502 => x"06585876",
  1503 => x"f4387d8b",
  1504 => x"2b76862b",
  1505 => x"07820790",
  1506 => x"160c9015",
  1507 => x"0870832a",
  1508 => x"81065a5a",
  1509 => x"78f43890",
  1510 => x"15087090",
  1511 => x"2a57588b",
  1512 => x"5380e198",
  1513 => x"527f5197",
  1514 => x"bc3f8457",
  1515 => x"758f0654",
  1516 => x"73892683",
  1517 => x"e038761c",
  1518 => x"b0155555",
  1519 => x"73753475",
  1520 => x"842aff18",
  1521 => x"7081ff06",
  1522 => x"59565676",
  1523 => x"df387f60",
  1524 => x"33555773",
  1525 => x"802ea938",
  1526 => x"80e69008",
  1527 => x"74575581",
  1528 => x"1757758a",
  1529 => x"2e82d238",
  1530 => x"84150870",
  1531 => x"822a8106",
  1532 => x"59597780",
  1533 => x"2ef23875",
  1534 => x"750c7633",
  1535 => x"5675e038",
  1536 => x"811b5b9f",
  1537 => x"7b27fcc9",
  1538 => x"38811f5f",
  1539 => x"9f7f27fb",
  1540 => x"9e3880e6",
  1541 => x"90085584",
  1542 => x"15087082",
  1543 => x"2a81065e",
  1544 => x"407c802e",
  1545 => x"f2388d75",
  1546 => x"0c841508",
  1547 => x"70822a81",
  1548 => x"06425c60",
  1549 => x"802ef238",
  1550 => x"8a750c9e",
  1551 => x"3d0d0484",
  1552 => x"15087082",
  1553 => x"2a810655",
  1554 => x"5973802e",
  1555 => x"f2388d75",
  1556 => x"0c841508",
  1557 => x"70822a81",
  1558 => x"065b5c79",
  1559 => x"802efa9d",
  1560 => x"38faa939",
  1561 => x"84150870",
  1562 => x"822a8106",
  1563 => x"5f587d80",
  1564 => x"2ef2388d",
  1565 => x"750c8415",
  1566 => x"0870822a",
  1567 => x"81065a5b",
  1568 => x"78802efa",
  1569 => x"c938fad5",
  1570 => x"396117b7",
  1571 => x"15555573",
  1572 => x"75347584",
  1573 => x"2aff1870",
  1574 => x"81ff0659",
  1575 => x"565676fa",
  1576 => x"d438faf3",
  1577 => x"39841508",
  1578 => x"70822a81",
  1579 => x"065f587d",
  1580 => x"802ef238",
  1581 => x"8d750c84",
  1582 => x"15087082",
  1583 => x"2a81065a",
  1584 => x"5b78802e",
  1585 => x"faeb38fa",
  1586 => x"f7398415",
  1587 => x"0870822a",
  1588 => x"81065559",
  1589 => x"73802ef2",
  1590 => x"388d750c",
  1591 => x"84150870",
  1592 => x"822a8106",
  1593 => x"5b587980",
  1594 => x"2efb9738",
  1595 => x"fba33984",
  1596 => x"15087082",
  1597 => x"2a81065b",
  1598 => x"5479802e",
  1599 => x"f2388d75",
  1600 => x"0c841508",
  1601 => x"70822a81",
  1602 => x"065a5878",
  1603 => x"802efc87",
  1604 => x"38fc9339",
  1605 => x"84150870",
  1606 => x"822a8106",
  1607 => x"555a7380",
  1608 => x"2ef2388d",
  1609 => x"750c8415",
  1610 => x"0870822a",
  1611 => x"81065959",
  1612 => x"77802efc",
  1613 => x"9938fca5",
  1614 => x"39841508",
  1615 => x"70822a81",
  1616 => x"06555a73",
  1617 => x"802ef238",
  1618 => x"8d750c84",
  1619 => x"15087082",
  1620 => x"2a810659",
  1621 => x"5977802e",
  1622 => x"fd8e38fd",
  1623 => x"9a39ad7d",
  1624 => x"340280e1",
  1625 => x"057b3071",
  1626 => x"1a59575a",
  1627 => x"8a527551",
  1628 => x"8fc53f80",
  1629 => x"08b00555",
  1630 => x"74773481",
  1631 => x"18588a52",
  1632 => x"75518f8e",
  1633 => x"3f800856",
  1634 => x"8008fa9a",
  1635 => x"38faba39",
  1636 => x"9b5bf9cf",
  1637 => x"39761cb7",
  1638 => x"155555fc",
  1639 => x"9f39905b",
  1640 => x"f9c13994",
  1641 => x"5bf9bc39",
  1642 => x"ef3d0d80",
  1643 => x"0b80e694",
  1644 => x"08575574",
  1645 => x"76279a38",
  1646 => x"75753154",
  1647 => x"73fa8080",
  1648 => x"82aa1634",
  1649 => x"811580e6",
  1650 => x"94085755",
  1651 => x"757526e8",
  1652 => x"38800bfa",
  1653 => x"80808280",
  1654 => x"349b0bfa",
  1655 => x"80808281",
  1656 => x"34a10bfa",
  1657 => x"80808282",
  1658 => x"3480e80b",
  1659 => x"fa808082",
  1660 => x"833480cb",
  1661 => x"0bfa8080",
  1662 => x"8284348a",
  1663 => x"0bfa8080",
  1664 => x"828534de",
  1665 => x"0bfa8080",
  1666 => x"828634ff",
  1667 => x"ad0bfa80",
  1668 => x"80828734",
  1669 => x"ffbe0bfa",
  1670 => x"80808288",
  1671 => x"34ef0bfa",
  1672 => x"80808289",
  1673 => x"34800bfa",
  1674 => x"8080828a",
  1675 => x"34a00bfa",
  1676 => x"8080828b",
  1677 => x"34880bfa",
  1678 => x"8080828c",
  1679 => x"34800bfa",
  1680 => x"8080828d",
  1681 => x"3480c50b",
  1682 => x"fa808082",
  1683 => x"8e34800b",
  1684 => x"fa808082",
  1685 => x"8f349d16",
  1686 => x"7083ffff",
  1687 => x"0670882a",
  1688 => x"57555774",
  1689 => x"fa808082",
  1690 => x"903473fa",
  1691 => x"80808291",
  1692 => x"34800bfa",
  1693 => x"80808292",
  1694 => x"34800bfa",
  1695 => x"80808293",
  1696 => x"3480c00b",
  1697 => x"fa808082",
  1698 => x"9434800b",
  1699 => x"fa808082",
  1700 => x"9534ff0b",
  1701 => x"fa808082",
  1702 => x"9634910b",
  1703 => x"fa808082",
  1704 => x"973480e7",
  1705 => x"0bfa8080",
  1706 => x"829834ff",
  1707 => x"8d0bfa80",
  1708 => x"80829934",
  1709 => x"8a0bfa80",
  1710 => x"80829a34",
  1711 => x"800bfa80",
  1712 => x"80829b34",
  1713 => x"800bfa80",
  1714 => x"80829c34",
  1715 => x"820bfa80",
  1716 => x"80829d34",
  1717 => x"8a0bfa80",
  1718 => x"80829e34",
  1719 => x"800bfa80",
  1720 => x"80829f34",
  1721 => x"800bfa80",
  1722 => x"8082a034",
  1723 => x"810bfa80",
  1724 => x"8082a134",
  1725 => x"930bfa80",
  1726 => x"8082a234",
  1727 => x"ffba0bfa",
  1728 => x"808082a3",
  1729 => x"34930bfa",
  1730 => x"808082a4",
  1731 => x"34ffba0b",
  1732 => x"fa808082",
  1733 => x"a5348816",
  1734 => x"7083ffff",
  1735 => x"0670882a",
  1736 => x"5a585977",
  1737 => x"fa808082",
  1738 => x"a63476fa",
  1739 => x"808082a7",
  1740 => x"34ff9f0b",
  1741 => x"fa808082",
  1742 => x"a834e30b",
  1743 => x"fa808082",
  1744 => x"a934fa80",
  1745 => x"8082800b",
  1746 => x"fa808080",
  1747 => x"840caa16",
  1748 => x"b0800785",
  1749 => x"0a0c80e6",
  1750 => x"84085885",
  1751 => x"0a0b9419",
  1752 => x"0c91780c",
  1753 => x"850a0870",
  1754 => x"8b2a8106",
  1755 => x"575475f4",
  1756 => x"3880e38c",
  1757 => x"0b80e38c",
  1758 => x"33555773",
  1759 => x"802ea938",
  1760 => x"7380e690",
  1761 => x"08565681",
  1762 => x"1757758a",
  1763 => x"2e83d938",
  1764 => x"84150870",
  1765 => x"822a8106",
  1766 => x"51547380",
  1767 => x"2ef23875",
  1768 => x"750c7633",
  1769 => x"5675e038",
  1770 => x"7708913d",
  1771 => x"5a568b53",
  1772 => x"80e19852",
  1773 => x"78518fad",
  1774 => x"3f880284",
  1775 => x"05bd0559",
  1776 => x"57758f06",
  1777 => x"54738926",
  1778 => x"858e3876",
  1779 => x"18b01555",
  1780 => x"55737534",
  1781 => x"75842aff",
  1782 => x"187081ff",
  1783 => x"06595656",
  1784 => x"76df3878",
  1785 => x"79335557",
  1786 => x"73802ea9",
  1787 => x"3880e690",
  1788 => x"08745755",
  1789 => x"81175775",
  1790 => x"8a2e8391",
  1791 => x"38841508",
  1792 => x"70822a81",
  1793 => x"06595477",
  1794 => x"802ef238",
  1795 => x"75750c76",
  1796 => x"335675e0",
  1797 => x"3880e3a0",
  1798 => x"0b80e3a0",
  1799 => x"33555773",
  1800 => x"802ea938",
  1801 => x"80e69008",
  1802 => x"74575581",
  1803 => x"1757758a",
  1804 => x"2e82ff38",
  1805 => x"84150870",
  1806 => x"822a8106",
  1807 => x"59547780",
  1808 => x"2ef23875",
  1809 => x"750c7633",
  1810 => x"5675e038",
  1811 => x"80e68408",
  1812 => x"8411088f",
  1813 => x"3d5b5757",
  1814 => x"8b5380e1",
  1815 => x"98527851",
  1816 => x"8e833f88",
  1817 => x"028405b1",
  1818 => x"05595775",
  1819 => x"8f065473",
  1820 => x"892683db",
  1821 => x"387618b0",
  1822 => x"15555573",
  1823 => x"75347584",
  1824 => x"2aff1870",
  1825 => x"81ff0659",
  1826 => x"565676df",
  1827 => x"38787933",
  1828 => x"55577380",
  1829 => x"2ea93880",
  1830 => x"e6900874",
  1831 => x"57558117",
  1832 => x"57758a2e",
  1833 => x"82b13884",
  1834 => x"15087082",
  1835 => x"2a810659",
  1836 => x"5477802e",
  1837 => x"f2387575",
  1838 => x"0c763356",
  1839 => x"75e03880",
  1840 => x"e3b40b80",
  1841 => x"e3b43355",
  1842 => x"5773802e",
  1843 => x"a93880e6",
  1844 => x"90087457",
  1845 => x"55811757",
  1846 => x"758a2e82",
  1847 => x"9f388415",
  1848 => x"0870822a",
  1849 => x"81065954",
  1850 => x"77802ef2",
  1851 => x"3875750c",
  1852 => x"76335675",
  1853 => x"e038850a",
  1854 => x"088b3d5a",
  1855 => x"568b5380",
  1856 => x"e1985278",
  1857 => x"518cde3f",
  1858 => x"88028405",
  1859 => x"a5055957",
  1860 => x"758f0654",
  1861 => x"73892682",
  1862 => x"ad387618",
  1863 => x"b0155555",
  1864 => x"73753475",
  1865 => x"842aff18",
  1866 => x"7081ff06",
  1867 => x"59565676",
  1868 => x"df387879",
  1869 => x"33555773",
  1870 => x"802ea938",
  1871 => x"80e69008",
  1872 => x"74575581",
  1873 => x"1757758a",
  1874 => x"2e81d638",
  1875 => x"84150870",
  1876 => x"822a8106",
  1877 => x"59547780",
  1878 => x"2ef23875",
  1879 => x"750c7633",
  1880 => x"5675e038",
  1881 => x"933d0d04",
  1882 => x"84150870",
  1883 => x"822a8106",
  1884 => x"51597880",
  1885 => x"2ef2388d",
  1886 => x"750c8415",
  1887 => x"0870822a",
  1888 => x"81065154",
  1889 => x"73802efc",
  1890 => x"8738fc93",
  1891 => x"39841508",
  1892 => x"70822a81",
  1893 => x"06595477",
  1894 => x"802ef238",
  1895 => x"8d750c84",
  1896 => x"15087082",
  1897 => x"2a810659",
  1898 => x"5477802e",
  1899 => x"fccf38fc",
  1900 => x"db398415",
  1901 => x"0870822a",
  1902 => x"81065954",
  1903 => x"77802ef2",
  1904 => x"388d750c",
  1905 => x"84150870",
  1906 => x"822a8106",
  1907 => x"59547780",
  1908 => x"2efce138",
  1909 => x"fced3984",
  1910 => x"15087082",
  1911 => x"2a810659",
  1912 => x"5477802e",
  1913 => x"f2388d75",
  1914 => x"0c841508",
  1915 => x"70822a81",
  1916 => x"06595477",
  1917 => x"802efdaf",
  1918 => x"38fdbb39",
  1919 => x"84150870",
  1920 => x"822a8106",
  1921 => x"59547780",
  1922 => x"2ef2388d",
  1923 => x"750c8415",
  1924 => x"0870822a",
  1925 => x"81065954",
  1926 => x"77802efd",
  1927 => x"c138fdcd",
  1928 => x"39841508",
  1929 => x"70822a81",
  1930 => x"06595477",
  1931 => x"802ef238",
  1932 => x"8d750c84",
  1933 => x"15087082",
  1934 => x"2a810659",
  1935 => x"5477802e",
  1936 => x"fe8a38fe",
  1937 => x"96397618",
  1938 => x"b7155555",
  1939 => x"fdd23976",
  1940 => x"18b71555",
  1941 => x"55fca439",
  1942 => x"7618b715",
  1943 => x"5555faf1",
  1944 => x"39f83d0d",
  1945 => x"80e68808",
  1946 => x"7008810a",
  1947 => x"0680e68c",
  1948 => x"08565a53",
  1949 => x"870b8415",
  1950 => x"0c80e690",
  1951 => x"0854b60b",
  1952 => x"8c150c83",
  1953 => x"0b88150c",
  1954 => x"81ff0b88",
  1955 => x"140c80e6",
  1956 => x"840855ff",
  1957 => x"0b84160c",
  1958 => x"fc94800b",
  1959 => x"88160c82",
  1960 => x"d0affdfb",
  1961 => x"0b8c160c",
  1962 => x"80c0750c",
  1963 => x"74087086",
  1964 => x"2a810657",
  1965 => x"5875f538",
  1966 => x"90150870",
  1967 => x"832a8106",
  1968 => x"545772f4",
  1969 => x"3881fc80",
  1970 => x"810b9016",
  1971 => x"0c901508",
  1972 => x"70832a81",
  1973 => x"06595677",
  1974 => x"f43880fd",
  1975 => x"c0810b90",
  1976 => x"160c80e3",
  1977 => x"c80b80e3",
  1978 => x"c8335456",
  1979 => x"72802ea4",
  1980 => x"38725581",
  1981 => x"1656748a",
  1982 => x"2e829c38",
  1983 => x"84140870",
  1984 => x"822a8106",
  1985 => x"58537680",
  1986 => x"2ef23874",
  1987 => x"740c7533",
  1988 => x"5574e038",
  1989 => x"80e3cc0b",
  1990 => x"80e3cc33",
  1991 => x"54567280",
  1992 => x"2ea43872",
  1993 => x"55811656",
  1994 => x"748a2e82",
  1995 => x"8f388414",
  1996 => x"0870822a",
  1997 => x"81065853",
  1998 => x"76802ef2",
  1999 => x"3874740c",
  2000 => x"75335574",
  2001 => x"e0387880",
  2002 => x"2e82e338",
  2003 => x"80e3d40b",
  2004 => x"80e3d433",
  2005 => x"54567280",
  2006 => x"2ea43872",
  2007 => x"55811656",
  2008 => x"748a2e81",
  2009 => x"fc388414",
  2010 => x"0870822a",
  2011 => x"81065853",
  2012 => x"76802ef2",
  2013 => x"3874740c",
  2014 => x"75335574",
  2015 => x"e03880e3",
  2016 => x"e40b80e3",
  2017 => x"e4335456",
  2018 => x"72802ea4",
  2019 => x"38725581",
  2020 => x"1656748a",
  2021 => x"2e81ef38",
  2022 => x"84140870",
  2023 => x"822a8106",
  2024 => x"58537680",
  2025 => x"2ef23874",
  2026 => x"740c7533",
  2027 => x"5574e038",
  2028 => x"f3f63ff8",
  2029 => x"81c08e80",
  2030 => x"55a00b80",
  2031 => x"e6880880",
  2032 => x"e68c085a",
  2033 => x"58567484",
  2034 => x"180c749f",
  2035 => x"2a751007",
  2036 => x"5578802e",
  2037 => x"98387580",
  2038 => x"2e81d038",
  2039 => x"ff167584",
  2040 => x"190c759f",
  2041 => x"2a761007",
  2042 => x"565678ea",
  2043 => x"387754af",
  2044 => x"d7c20b94",
  2045 => x"190c850b",
  2046 => x"98190c98",
  2047 => x"14087081",
  2048 => x"06515372",
  2049 => x"802effbe",
  2050 => x"38981408",
  2051 => x"70810651",
  2052 => x"5372e838",
  2053 => x"ffb03984",
  2054 => x"14087082",
  2055 => x"2a810658",
  2056 => x"5376802e",
  2057 => x"f2388d74",
  2058 => x"0c841408",
  2059 => x"70822a81",
  2060 => x"06585376",
  2061 => x"802efdc4",
  2062 => x"38fdd039",
  2063 => x"84140870",
  2064 => x"822a8106",
  2065 => x"58537680",
  2066 => x"2ef2388d",
  2067 => x"740c8414",
  2068 => x"0870822a",
  2069 => x"81065853",
  2070 => x"76802efd",
  2071 => x"d138fddd",
  2072 => x"39841408",
  2073 => x"70822a81",
  2074 => x"06585376",
  2075 => x"802ef238",
  2076 => x"8d740c84",
  2077 => x"14087082",
  2078 => x"2a810658",
  2079 => x"5376802e",
  2080 => x"fde438fd",
  2081 => x"f0398414",
  2082 => x"0870822a",
  2083 => x"81065853",
  2084 => x"76802ef2",
  2085 => x"388d740c",
  2086 => x"84140870",
  2087 => x"822a8106",
  2088 => x"58537680",
  2089 => x"2efdf138",
  2090 => x"fdfd3985",
  2091 => x"ab3f80e4",
  2092 => x"880b80e4",
  2093 => x"88335456",
  2094 => x"72802efd",
  2095 => x"c1387281",
  2096 => x"17575574",
  2097 => x"8a2ea738",
  2098 => x"84140870",
  2099 => x"822a8106",
  2100 => x"58537680",
  2101 => x"2ef23874",
  2102 => x"740c7533",
  2103 => x"5574802e",
  2104 => x"fd9c3881",
  2105 => x"1656748a",
  2106 => x"2e098106",
  2107 => x"db388414",
  2108 => x"0870822a",
  2109 => x"81065853",
  2110 => x"76802ef2",
  2111 => x"388d740c",
  2112 => x"84140870",
  2113 => x"822a8106",
  2114 => x"58537680",
  2115 => x"2effb938",
  2116 => x"c6398c08",
  2117 => x"028c0cfd",
  2118 => x"3d0d8053",
  2119 => x"8c088c05",
  2120 => x"08528c08",
  2121 => x"88050851",
  2122 => x"82de3f80",
  2123 => x"0870800c",
  2124 => x"54853d0d",
  2125 => x"8c0c048c",
  2126 => x"08028c0c",
  2127 => x"fd3d0d81",
  2128 => x"538c088c",
  2129 => x"0508528c",
  2130 => x"08880508",
  2131 => x"5182b93f",
  2132 => x"80087080",
  2133 => x"0c54853d",
  2134 => x"0d8c0c04",
  2135 => x"8c08028c",
  2136 => x"0cf93d0d",
  2137 => x"800b8c08",
  2138 => x"fc050c8c",
  2139 => x"08880508",
  2140 => x"8025ab38",
  2141 => x"8c088805",
  2142 => x"08308c08",
  2143 => x"88050c80",
  2144 => x"0b8c08f4",
  2145 => x"050c8c08",
  2146 => x"fc050888",
  2147 => x"38810b8c",
  2148 => x"08f4050c",
  2149 => x"8c08f405",
  2150 => x"088c08fc",
  2151 => x"050c8c08",
  2152 => x"8c050880",
  2153 => x"25ab388c",
  2154 => x"088c0508",
  2155 => x"308c088c",
  2156 => x"050c800b",
  2157 => x"8c08f005",
  2158 => x"0c8c08fc",
  2159 => x"05088838",
  2160 => x"810b8c08",
  2161 => x"f0050c8c",
  2162 => x"08f00508",
  2163 => x"8c08fc05",
  2164 => x"0c80538c",
  2165 => x"088c0508",
  2166 => x"528c0888",
  2167 => x"05085181",
  2168 => x"a73f8008",
  2169 => x"708c08f8",
  2170 => x"050c548c",
  2171 => x"08fc0508",
  2172 => x"802e8c38",
  2173 => x"8c08f805",
  2174 => x"08308c08",
  2175 => x"f8050c8c",
  2176 => x"08f80508",
  2177 => x"70800c54",
  2178 => x"893d0d8c",
  2179 => x"0c048c08",
  2180 => x"028c0cfb",
  2181 => x"3d0d800b",
  2182 => x"8c08fc05",
  2183 => x"0c8c0888",
  2184 => x"05088025",
  2185 => x"93388c08",
  2186 => x"88050830",
  2187 => x"8c088805",
  2188 => x"0c810b8c",
  2189 => x"08fc050c",
  2190 => x"8c088c05",
  2191 => x"0880258c",
  2192 => x"388c088c",
  2193 => x"0508308c",
  2194 => x"088c050c",
  2195 => x"81538c08",
  2196 => x"8c050852",
  2197 => x"8c088805",
  2198 => x"0851ad3f",
  2199 => x"8008708c",
  2200 => x"08f8050c",
  2201 => x"548c08fc",
  2202 => x"0508802e",
  2203 => x"8c388c08",
  2204 => x"f8050830",
  2205 => x"8c08f805",
  2206 => x"0c8c08f8",
  2207 => x"05087080",
  2208 => x"0c54873d",
  2209 => x"0d8c0c04",
  2210 => x"8c08028c",
  2211 => x"0cfd3d0d",
  2212 => x"810b8c08",
  2213 => x"fc050c80",
  2214 => x"0b8c08f8",
  2215 => x"050c8c08",
  2216 => x"8c05088c",
  2217 => x"08880508",
  2218 => x"27ac388c",
  2219 => x"08fc0508",
  2220 => x"802ea338",
  2221 => x"800b8c08",
  2222 => x"8c050824",
  2223 => x"99388c08",
  2224 => x"8c050810",
  2225 => x"8c088c05",
  2226 => x"0c8c08fc",
  2227 => x"0508108c",
  2228 => x"08fc050c",
  2229 => x"c9398c08",
  2230 => x"fc050880",
  2231 => x"2e80c938",
  2232 => x"8c088c05",
  2233 => x"088c0888",
  2234 => x"050826a1",
  2235 => x"388c0888",
  2236 => x"05088c08",
  2237 => x"8c050831",
  2238 => x"8c088805",
  2239 => x"0c8c08f8",
  2240 => x"05088c08",
  2241 => x"fc050807",
  2242 => x"8c08f805",
  2243 => x"0c8c08fc",
  2244 => x"0508812a",
  2245 => x"8c08fc05",
  2246 => x"0c8c088c",
  2247 => x"0508812a",
  2248 => x"8c088c05",
  2249 => x"0cffaf39",
  2250 => x"8c089005",
  2251 => x"08802e8f",
  2252 => x"388c0888",
  2253 => x"0508708c",
  2254 => x"08f4050c",
  2255 => x"518d398c",
  2256 => x"08f80508",
  2257 => x"708c08f4",
  2258 => x"050c518c",
  2259 => x"08f40508",
  2260 => x"800c853d",
  2261 => x"0d8c0c04",
  2262 => x"803d0d86",
  2263 => x"5184963f",
  2264 => x"815198d7",
  2265 => x"3ffc3d0d",
  2266 => x"7670797b",
  2267 => x"55555555",
  2268 => x"8f72278c",
  2269 => x"38727507",
  2270 => x"83065170",
  2271 => x"802ea738",
  2272 => x"ff125271",
  2273 => x"ff2e9838",
  2274 => x"72708105",
  2275 => x"54337470",
  2276 => x"81055634",
  2277 => x"ff125271",
  2278 => x"ff2e0981",
  2279 => x"06ea3874",
  2280 => x"800c863d",
  2281 => x"0d047451",
  2282 => x"72708405",
  2283 => x"54087170",
  2284 => x"8405530c",
  2285 => x"72708405",
  2286 => x"54087170",
  2287 => x"8405530c",
  2288 => x"72708405",
  2289 => x"54087170",
  2290 => x"8405530c",
  2291 => x"72708405",
  2292 => x"54087170",
  2293 => x"8405530c",
  2294 => x"f0125271",
  2295 => x"8f26c938",
  2296 => x"83722795",
  2297 => x"38727084",
  2298 => x"05540871",
  2299 => x"70840553",
  2300 => x"0cfc1252",
  2301 => x"718326ed",
  2302 => x"387054ff",
  2303 => x"8339fd3d",
  2304 => x"0d755384",
  2305 => x"d8130880",
  2306 => x"2e8a3880",
  2307 => x"5372800c",
  2308 => x"853d0d04",
  2309 => x"81805272",
  2310 => x"5183d83f",
  2311 => x"800884d8",
  2312 => x"140cff53",
  2313 => x"8008802e",
  2314 => x"e4388008",
  2315 => x"549f5380",
  2316 => x"74708405",
  2317 => x"560cff13",
  2318 => x"53807324",
  2319 => x"ce388074",
  2320 => x"70840556",
  2321 => x"0cff1353",
  2322 => x"728025e3",
  2323 => x"38ffbc39",
  2324 => x"fd3d0d75",
  2325 => x"7755539f",
  2326 => x"74278d38",
  2327 => x"96730cff",
  2328 => x"5271800c",
  2329 => x"853d0d04",
  2330 => x"84d81308",
  2331 => x"5271802e",
  2332 => x"93387310",
  2333 => x"10127008",
  2334 => x"79720c51",
  2335 => x"5271800c",
  2336 => x"853d0d04",
  2337 => x"7251fef6",
  2338 => x"3fff5280",
  2339 => x"08d33884",
  2340 => x"d8130874",
  2341 => x"10101170",
  2342 => x"087a720c",
  2343 => x"515152dd",
  2344 => x"39f93d0d",
  2345 => x"797b5856",
  2346 => x"769f2680",
  2347 => x"e83884d8",
  2348 => x"16085473",
  2349 => x"802eaa38",
  2350 => x"76101014",
  2351 => x"70085555",
  2352 => x"73802eba",
  2353 => x"38805873",
  2354 => x"812e8f38",
  2355 => x"73ff2ea3",
  2356 => x"3880750c",
  2357 => x"7651732d",
  2358 => x"80587780",
  2359 => x"0c893d0d",
  2360 => x"047551fe",
  2361 => x"993fff58",
  2362 => x"8008ef38",
  2363 => x"84d81608",
  2364 => x"54c63996",
  2365 => x"760c810b",
  2366 => x"800c893d",
  2367 => x"0d047551",
  2368 => x"81ed3f76",
  2369 => x"53800852",
  2370 => x"755181ad",
  2371 => x"3f800880",
  2372 => x"0c893d0d",
  2373 => x"0496760c",
  2374 => x"ff0b800c",
  2375 => x"893d0d04",
  2376 => x"fc3d0d76",
  2377 => x"785653ff",
  2378 => x"54749f26",
  2379 => x"b13884d8",
  2380 => x"13085271",
  2381 => x"802eae38",
  2382 => x"74101012",
  2383 => x"70085353",
  2384 => x"81547180",
  2385 => x"2e983882",
  2386 => x"5471ff2e",
  2387 => x"91388354",
  2388 => x"71812e8a",
  2389 => x"3880730c",
  2390 => x"7451712d",
  2391 => x"80547380",
  2392 => x"0c863d0d",
  2393 => x"047251fd",
  2394 => x"953f8008",
  2395 => x"f13884d8",
  2396 => x"130852c4",
  2397 => x"39ff3d0d",
  2398 => x"735280e6",
  2399 => x"980851fe",
  2400 => x"a03f833d",
  2401 => x"0d04fe3d",
  2402 => x"0d755374",
  2403 => x"5280e698",
  2404 => x"0851fdbc",
  2405 => x"3f843d0d",
  2406 => x"04803d0d",
  2407 => x"80e69808",
  2408 => x"51fcdb3f",
  2409 => x"823d0d04",
  2410 => x"ff3d0d73",
  2411 => x"5280e698",
  2412 => x"0851feec",
  2413 => x"3f833d0d",
  2414 => x"04fc3d0d",
  2415 => x"800b80f6",
  2416 => x"8c0c7852",
  2417 => x"775192e7",
  2418 => x"3f800854",
  2419 => x"8008ff2e",
  2420 => x"88387380",
  2421 => x"0c863d0d",
  2422 => x"0480f68c",
  2423 => x"08557480",
  2424 => x"2ef03876",
  2425 => x"75710c53",
  2426 => x"73800c86",
  2427 => x"3d0d0492",
  2428 => x"b93f04f3",
  2429 => x"3d0d7f61",
  2430 => x"8b1170f8",
  2431 => x"065c5555",
  2432 => x"5e729626",
  2433 => x"83389059",
  2434 => x"80792474",
  2435 => x"7a260753",
  2436 => x"80547274",
  2437 => x"2e098106",
  2438 => x"80cb387d",
  2439 => x"518bca3f",
  2440 => x"7883f726",
  2441 => x"80c63878",
  2442 => x"832a7010",
  2443 => x"101080ed",
  2444 => x"d4058c11",
  2445 => x"0859595a",
  2446 => x"76782e83",
  2447 => x"b0388417",
  2448 => x"08fc0656",
  2449 => x"8c170888",
  2450 => x"1808718c",
  2451 => x"120c8812",
  2452 => x"0c587517",
  2453 => x"84110881",
  2454 => x"0784120c",
  2455 => x"537d518b",
  2456 => x"893f8817",
  2457 => x"5473800c",
  2458 => x"8f3d0d04",
  2459 => x"78892a79",
  2460 => x"832a5b53",
  2461 => x"72802ebf",
  2462 => x"3878862a",
  2463 => x"b8055a84",
  2464 => x"7327b438",
  2465 => x"80db135a",
  2466 => x"947327ab",
  2467 => x"38788c2a",
  2468 => x"80ee055a",
  2469 => x"80d47327",
  2470 => x"9e38788f",
  2471 => x"2a80f705",
  2472 => x"5a82d473",
  2473 => x"27913878",
  2474 => x"922a80fc",
  2475 => x"055a8ad4",
  2476 => x"73278438",
  2477 => x"80fe5a79",
  2478 => x"10101080",
  2479 => x"edd4058c",
  2480 => x"11085855",
  2481 => x"76752ea3",
  2482 => x"38841708",
  2483 => x"fc06707a",
  2484 => x"31555673",
  2485 => x"8f2488d5",
  2486 => x"38738025",
  2487 => x"fee6388c",
  2488 => x"17085776",
  2489 => x"752e0981",
  2490 => x"06df3881",
  2491 => x"1a5a80ed",
  2492 => x"e4085776",
  2493 => x"80eddc2e",
  2494 => x"82c03884",
  2495 => x"1708fc06",
  2496 => x"707a3155",
  2497 => x"56738f24",
  2498 => x"81f93880",
  2499 => x"eddc0b80",
  2500 => x"ede80c80",
  2501 => x"eddc0b80",
  2502 => x"ede40c73",
  2503 => x"8025feb2",
  2504 => x"3883ff76",
  2505 => x"2783df38",
  2506 => x"75892a76",
  2507 => x"832a5553",
  2508 => x"72802ebf",
  2509 => x"3875862a",
  2510 => x"b8055484",
  2511 => x"7327b438",
  2512 => x"80db1354",
  2513 => x"947327ab",
  2514 => x"38758c2a",
  2515 => x"80ee0554",
  2516 => x"80d47327",
  2517 => x"9e38758f",
  2518 => x"2a80f705",
  2519 => x"5482d473",
  2520 => x"27913875",
  2521 => x"922a80fc",
  2522 => x"05548ad4",
  2523 => x"73278438",
  2524 => x"80fe5473",
  2525 => x"10101080",
  2526 => x"edd40588",
  2527 => x"11085658",
  2528 => x"74782e86",
  2529 => x"cf388415",
  2530 => x"08fc0653",
  2531 => x"7573278d",
  2532 => x"38881508",
  2533 => x"5574782e",
  2534 => x"098106ea",
  2535 => x"388c1508",
  2536 => x"80edd40b",
  2537 => x"84050871",
  2538 => x"8c1a0c76",
  2539 => x"881a0c78",
  2540 => x"88130c78",
  2541 => x"8c180c5d",
  2542 => x"58795380",
  2543 => x"7a2483e6",
  2544 => x"3872822c",
  2545 => x"81712b5c",
  2546 => x"537a7c26",
  2547 => x"8198387b",
  2548 => x"7b065372",
  2549 => x"82f13879",
  2550 => x"fc068405",
  2551 => x"5a7a1070",
  2552 => x"7d06545b",
  2553 => x"7282e038",
  2554 => x"841a5af1",
  2555 => x"3988178c",
  2556 => x"11085858",
  2557 => x"76782e09",
  2558 => x"8106fcc2",
  2559 => x"38821a5a",
  2560 => x"fdec3978",
  2561 => x"17798107",
  2562 => x"84190c70",
  2563 => x"80ede80c",
  2564 => x"7080ede4",
  2565 => x"0c80eddc",
  2566 => x"0b8c120c",
  2567 => x"8c110888",
  2568 => x"120c7481",
  2569 => x"0784120c",
  2570 => x"74117571",
  2571 => x"0c51537d",
  2572 => x"5187b73f",
  2573 => x"881754fc",
  2574 => x"ac3980ed",
  2575 => x"d40b8405",
  2576 => x"087a545c",
  2577 => x"798025fe",
  2578 => x"f83882da",
  2579 => x"397a097c",
  2580 => x"067080ed",
  2581 => x"d40b8405",
  2582 => x"0c5c7a10",
  2583 => x"5b7a7c26",
  2584 => x"85387a85",
  2585 => x"b83880ed",
  2586 => x"d40b8805",
  2587 => x"08708412",
  2588 => x"08fc0670",
  2589 => x"7c317c72",
  2590 => x"268f7225",
  2591 => x"0757575c",
  2592 => x"5d557280",
  2593 => x"2e80db38",
  2594 => x"797a1680",
  2595 => x"edcc081b",
  2596 => x"90115a55",
  2597 => x"575b80ed",
  2598 => x"c808ff2e",
  2599 => x"8838a08f",
  2600 => x"13e08006",
  2601 => x"5776527d",
  2602 => x"5186c03f",
  2603 => x"80085480",
  2604 => x"08ff2e90",
  2605 => x"38800876",
  2606 => x"27829938",
  2607 => x"7480edd4",
  2608 => x"2e829138",
  2609 => x"80edd40b",
  2610 => x"88050855",
  2611 => x"841508fc",
  2612 => x"06707a31",
  2613 => x"7a72268f",
  2614 => x"72250752",
  2615 => x"55537283",
  2616 => x"e6387479",
  2617 => x"81078417",
  2618 => x"0c791670",
  2619 => x"80edd40b",
  2620 => x"88050c75",
  2621 => x"81078412",
  2622 => x"0c547e52",
  2623 => x"5785eb3f",
  2624 => x"881754fa",
  2625 => x"e0397583",
  2626 => x"2a705454",
  2627 => x"80742481",
  2628 => x"9b387282",
  2629 => x"2c81712b",
  2630 => x"80edd808",
  2631 => x"077080ed",
  2632 => x"d40b8405",
  2633 => x"0c751010",
  2634 => x"1080edd4",
  2635 => x"05881108",
  2636 => x"585a5d53",
  2637 => x"778c180c",
  2638 => x"7488180c",
  2639 => x"7688190c",
  2640 => x"768c160c",
  2641 => x"fcf33979",
  2642 => x"7a101010",
  2643 => x"80edd405",
  2644 => x"7057595d",
  2645 => x"8c150857",
  2646 => x"76752ea3",
  2647 => x"38841708",
  2648 => x"fc06707a",
  2649 => x"31555673",
  2650 => x"8f2483ca",
  2651 => x"38738025",
  2652 => x"8481388c",
  2653 => x"17085776",
  2654 => x"752e0981",
  2655 => x"06df3888",
  2656 => x"15811b70",
  2657 => x"8306555b",
  2658 => x"5572c938",
  2659 => x"7c830653",
  2660 => x"72802efd",
  2661 => x"b838ff1d",
  2662 => x"f819595d",
  2663 => x"88180878",
  2664 => x"2eea38fd",
  2665 => x"b539831a",
  2666 => x"53fc9639",
  2667 => x"83147082",
  2668 => x"2c81712b",
  2669 => x"80edd808",
  2670 => x"077080ed",
  2671 => x"d40b8405",
  2672 => x"0c761010",
  2673 => x"1080edd4",
  2674 => x"05881108",
  2675 => x"595b5e51",
  2676 => x"53fee139",
  2677 => x"80ed9808",
  2678 => x"17588008",
  2679 => x"762e818d",
  2680 => x"3880edc8",
  2681 => x"08ff2e83",
  2682 => x"ec387376",
  2683 => x"311880ed",
  2684 => x"980c7387",
  2685 => x"06705753",
  2686 => x"72802e88",
  2687 => x"38887331",
  2688 => x"70155556",
  2689 => x"76149fff",
  2690 => x"06a08071",
  2691 => x"31177054",
  2692 => x"7f535753",
  2693 => x"83d53f80",
  2694 => x"08538008",
  2695 => x"ff2e81a0",
  2696 => x"3880ed98",
  2697 => x"08167080",
  2698 => x"ed980c74",
  2699 => x"7580edd4",
  2700 => x"0b88050c",
  2701 => x"74763118",
  2702 => x"70810751",
  2703 => x"5556587b",
  2704 => x"80edd42e",
  2705 => x"839c3879",
  2706 => x"8f2682cb",
  2707 => x"38810b84",
  2708 => x"150c8415",
  2709 => x"08fc0670",
  2710 => x"7a317a72",
  2711 => x"268f7225",
  2712 => x"07525553",
  2713 => x"72802efc",
  2714 => x"f93880db",
  2715 => x"3980089f",
  2716 => x"ff065372",
  2717 => x"feeb3877",
  2718 => x"80ed980c",
  2719 => x"80edd40b",
  2720 => x"8805087b",
  2721 => x"18810784",
  2722 => x"120c5580",
  2723 => x"edc40878",
  2724 => x"27863877",
  2725 => x"80edc40c",
  2726 => x"80edc008",
  2727 => x"7827fcac",
  2728 => x"387780ed",
  2729 => x"c00c8415",
  2730 => x"08fc0670",
  2731 => x"7a317a72",
  2732 => x"268f7225",
  2733 => x"07525553",
  2734 => x"72802efc",
  2735 => x"a5388839",
  2736 => x"80745456",
  2737 => x"fedb397d",
  2738 => x"51829f3f",
  2739 => x"800b800c",
  2740 => x"8f3d0d04",
  2741 => x"73538074",
  2742 => x"24a93872",
  2743 => x"822c8171",
  2744 => x"2b80edd8",
  2745 => x"08077080",
  2746 => x"edd40b84",
  2747 => x"050c5d53",
  2748 => x"778c180c",
  2749 => x"7488180c",
  2750 => x"7688190c",
  2751 => x"768c160c",
  2752 => x"f9b73983",
  2753 => x"1470822c",
  2754 => x"81712b80",
  2755 => x"edd80807",
  2756 => x"7080edd4",
  2757 => x"0b84050c",
  2758 => x"5e5153d4",
  2759 => x"397b7b06",
  2760 => x"5372fca3",
  2761 => x"38841a7b",
  2762 => x"105c5af1",
  2763 => x"39ff1a81",
  2764 => x"11515af7",
  2765 => x"b9397817",
  2766 => x"79810784",
  2767 => x"190c8c18",
  2768 => x"08881908",
  2769 => x"718c120c",
  2770 => x"88120c59",
  2771 => x"7080ede8",
  2772 => x"0c7080ed",
  2773 => x"e40c80ed",
  2774 => x"dc0b8c12",
  2775 => x"0c8c1108",
  2776 => x"88120c74",
  2777 => x"81078412",
  2778 => x"0c741175",
  2779 => x"710c5153",
  2780 => x"f9bd3975",
  2781 => x"17841108",
  2782 => x"81078412",
  2783 => x"0c538c17",
  2784 => x"08881808",
  2785 => x"718c120c",
  2786 => x"88120c58",
  2787 => x"7d5180da",
  2788 => x"3f881754",
  2789 => x"f5cf3972",
  2790 => x"84150cf4",
  2791 => x"1af80670",
  2792 => x"841e0881",
  2793 => x"0607841e",
  2794 => x"0c701d54",
  2795 => x"5b850b84",
  2796 => x"140c850b",
  2797 => x"88140c8f",
  2798 => x"7b27fdcf",
  2799 => x"38881c52",
  2800 => x"7d518290",
  2801 => x"3f80edd4",
  2802 => x"0b880508",
  2803 => x"80ed9808",
  2804 => x"5955fdb7",
  2805 => x"397780ed",
  2806 => x"980c7380",
  2807 => x"edc80cfc",
  2808 => x"91397284",
  2809 => x"150cfda3",
  2810 => x"390404fd",
  2811 => x"3d0d800b",
  2812 => x"80f68c0c",
  2813 => x"765186cc",
  2814 => x"3f800853",
  2815 => x"8008ff2e",
  2816 => x"88387280",
  2817 => x"0c853d0d",
  2818 => x"0480f68c",
  2819 => x"08547380",
  2820 => x"2ef03875",
  2821 => x"74710c52",
  2822 => x"72800c85",
  2823 => x"3d0d04fb",
  2824 => x"3d0d7770",
  2825 => x"5256c23f",
  2826 => x"80edd40b",
  2827 => x"88050884",
  2828 => x"1108fc06",
  2829 => x"707b319f",
  2830 => x"ef05e080",
  2831 => x"06e08005",
  2832 => x"565653a0",
  2833 => x"80742494",
  2834 => x"38805275",
  2835 => x"51ff9c3f",
  2836 => x"80eddc08",
  2837 => x"15537280",
  2838 => x"082e8f38",
  2839 => x"7551ff8a",
  2840 => x"3f805372",
  2841 => x"800c873d",
  2842 => x"0d047330",
  2843 => x"527551fe",
  2844 => x"fa3f8008",
  2845 => x"ff2ea838",
  2846 => x"80edd40b",
  2847 => x"88050875",
  2848 => x"75318107",
  2849 => x"84120c53",
  2850 => x"80ed9808",
  2851 => x"743180ed",
  2852 => x"980c7551",
  2853 => x"fed43f81",
  2854 => x"0b800c87",
  2855 => x"3d0d0480",
  2856 => x"527551fe",
  2857 => x"c63f80ed",
  2858 => x"d40b8805",
  2859 => x"08800871",
  2860 => x"3156538f",
  2861 => x"7525ffa4",
  2862 => x"38800880",
  2863 => x"edc80831",
  2864 => x"80ed980c",
  2865 => x"74810784",
  2866 => x"140c7551",
  2867 => x"fe9c3f80",
  2868 => x"53ff9039",
  2869 => x"f63d0d7c",
  2870 => x"7e545b72",
  2871 => x"802e8283",
  2872 => x"387a51fe",
  2873 => x"843ff813",
  2874 => x"84110870",
  2875 => x"fe067013",
  2876 => x"841108fc",
  2877 => x"065d5859",
  2878 => x"545880ed",
  2879 => x"dc08752e",
  2880 => x"82de3878",
  2881 => x"84160c80",
  2882 => x"73810654",
  2883 => x"5a727a2e",
  2884 => x"81d53878",
  2885 => x"15841108",
  2886 => x"81065153",
  2887 => x"72a03878",
  2888 => x"17577981",
  2889 => x"e6388815",
  2890 => x"08537280",
  2891 => x"eddc2e82",
  2892 => x"f9388c15",
  2893 => x"08708c15",
  2894 => x"0c738812",
  2895 => x"0c567681",
  2896 => x"0784190c",
  2897 => x"76187771",
  2898 => x"0c537981",
  2899 => x"913883ff",
  2900 => x"772781c8",
  2901 => x"3876892a",
  2902 => x"77832a56",
  2903 => x"5372802e",
  2904 => x"bf387686",
  2905 => x"2ab80555",
  2906 => x"847327b4",
  2907 => x"3880db13",
  2908 => x"55947327",
  2909 => x"ab38768c",
  2910 => x"2a80ee05",
  2911 => x"5580d473",
  2912 => x"279e3876",
  2913 => x"8f2a80f7",
  2914 => x"055582d4",
  2915 => x"73279138",
  2916 => x"76922a80",
  2917 => x"fc05558a",
  2918 => x"d4732784",
  2919 => x"3880fe55",
  2920 => x"74101010",
  2921 => x"80edd405",
  2922 => x"88110855",
  2923 => x"5673762e",
  2924 => x"82b33884",
  2925 => x"1408fc06",
  2926 => x"53767327",
  2927 => x"8d388814",
  2928 => x"08547376",
  2929 => x"2e098106",
  2930 => x"ea388c14",
  2931 => x"08708c1a",
  2932 => x"0c74881a",
  2933 => x"0c788812",
  2934 => x"0c56778c",
  2935 => x"150c7a51",
  2936 => x"fc883f8c",
  2937 => x"3d0d0477",
  2938 => x"08787131",
  2939 => x"59770588",
  2940 => x"19085457",
  2941 => x"7280eddc",
  2942 => x"2e80e038",
  2943 => x"8c180870",
  2944 => x"8c150c73",
  2945 => x"88120c56",
  2946 => x"fe893988",
  2947 => x"15088c16",
  2948 => x"08708c13",
  2949 => x"0c578817",
  2950 => x"0cfea339",
  2951 => x"76832a70",
  2952 => x"54558075",
  2953 => x"24819838",
  2954 => x"72822c81",
  2955 => x"712b80ed",
  2956 => x"d8080780",
  2957 => x"edd40b84",
  2958 => x"050c5374",
  2959 => x"10101080",
  2960 => x"edd40588",
  2961 => x"11085556",
  2962 => x"758c190c",
  2963 => x"7388190c",
  2964 => x"7788170c",
  2965 => x"778c150c",
  2966 => x"ff843981",
  2967 => x"5afdb439",
  2968 => x"78177381",
  2969 => x"06545772",
  2970 => x"98387708",
  2971 => x"78713159",
  2972 => x"77058c19",
  2973 => x"08881a08",
  2974 => x"718c120c",
  2975 => x"88120c57",
  2976 => x"57768107",
  2977 => x"84190c77",
  2978 => x"80edd40b",
  2979 => x"88050c80",
  2980 => x"edd00877",
  2981 => x"26fec738",
  2982 => x"80edcc08",
  2983 => x"527a51fa",
  2984 => x"fe3f7a51",
  2985 => x"fac43ffe",
  2986 => x"ba398178",
  2987 => x"8c150c78",
  2988 => x"88150c73",
  2989 => x"8c1a0c73",
  2990 => x"881a0c5a",
  2991 => x"fd803983",
  2992 => x"1570822c",
  2993 => x"81712b80",
  2994 => x"edd80807",
  2995 => x"80edd40b",
  2996 => x"84050c51",
  2997 => x"53741010",
  2998 => x"1080edd4",
  2999 => x"05881108",
  3000 => x"5556fee4",
  3001 => x"39745380",
  3002 => x"7524a738",
  3003 => x"72822c81",
  3004 => x"712b80ed",
  3005 => x"d8080780",
  3006 => x"edd40b84",
  3007 => x"050c5375",
  3008 => x"8c190c73",
  3009 => x"88190c77",
  3010 => x"88170c77",
  3011 => x"8c150cfd",
  3012 => x"cd398315",
  3013 => x"70822c81",
  3014 => x"712b80ed",
  3015 => x"d8080780",
  3016 => x"edd40b84",
  3017 => x"050c5153",
  3018 => x"d639810b",
  3019 => x"800c0480",
  3020 => x"3d0d7281",
  3021 => x"2e893880",
  3022 => x"0b800c82",
  3023 => x"3d0d0473",
  3024 => x"5180f83f",
  3025 => x"fe3d0d80",
  3026 => x"f6840851",
  3027 => x"708a3880",
  3028 => x"f6907080",
  3029 => x"f6840c51",
  3030 => x"70751252",
  3031 => x"52ff5370",
  3032 => x"87fb8080",
  3033 => x"26883870",
  3034 => x"80f6840c",
  3035 => x"71537280",
  3036 => x"0c843d0d",
  3037 => x"04fd3d0d",
  3038 => x"800b80e5",
  3039 => x"f8085454",
  3040 => x"72812e9c",
  3041 => x"387380f6",
  3042 => x"880cffa9",
  3043 => x"d33fffa8",
  3044 => x"ef3f80f5",
  3045 => x"dc528151",
  3046 => x"ddc73f80",
  3047 => x"0851a23f",
  3048 => x"7280f688",
  3049 => x"0cffa9b8",
  3050 => x"3fffa8d4",
  3051 => x"3f80f5dc",
  3052 => x"528151dd",
  3053 => x"ac3f8008",
  3054 => x"51873f00",
  3055 => x"ff3900ff",
  3056 => x"39f73d0d",
  3057 => x"7b80e698",
  3058 => x"0882c811",
  3059 => x"085a545a",
  3060 => x"77802e80",
  3061 => x"da388188",
  3062 => x"18841908",
  3063 => x"ff058171",
  3064 => x"2b595559",
  3065 => x"80742480",
  3066 => x"ea388074",
  3067 => x"24b53873",
  3068 => x"822b7811",
  3069 => x"88055656",
  3070 => x"81801908",
  3071 => x"77065372",
  3072 => x"802eb638",
  3073 => x"78167008",
  3074 => x"53537951",
  3075 => x"74085372",
  3076 => x"2dff14fc",
  3077 => x"17fc1779",
  3078 => x"812c5a57",
  3079 => x"57547380",
  3080 => x"25d63877",
  3081 => x"085877ff",
  3082 => x"ad3880e6",
  3083 => x"980853bc",
  3084 => x"1308a538",
  3085 => x"7951ff83",
  3086 => x"3f740853",
  3087 => x"722dff14",
  3088 => x"fc17fc17",
  3089 => x"79812c5a",
  3090 => x"57575473",
  3091 => x"8025ffa8",
  3092 => x"38d13980",
  3093 => x"57ff9339",
  3094 => x"7251bc13",
  3095 => x"0853722d",
  3096 => x"7951fed7",
  3097 => x"3fff3d0d",
  3098 => x"80f5e40b",
  3099 => x"fc057008",
  3100 => x"525270ff",
  3101 => x"2e913870",
  3102 => x"2dfc1270",
  3103 => x"08525270",
  3104 => x"ff2e0981",
  3105 => x"06f13883",
  3106 => x"3d0d0404",
  3107 => x"ffa8be3f",
  3108 => x"04000000",
  3109 => x"00000040",
  3110 => x"30782020",
  3111 => x"20202020",
  3112 => x"20200000",
  3113 => x"0a677265",
  3114 => x"74682072",
  3115 => x"65676973",
  3116 => x"74657273",
  3117 => x"3a000000",
  3118 => x"0a636f6e",
  3119 => x"74726f6c",
  3120 => x"3a202020",
  3121 => x"20202000",
  3122 => x"0a737461",
  3123 => x"7475733a",
  3124 => x"20202020",
  3125 => x"20202000",
  3126 => x"0a6d6163",
  3127 => x"5f6d7362",
  3128 => x"3a202020",
  3129 => x"20202000",
  3130 => x"0a6d6163",
  3131 => x"5f6c7362",
  3132 => x"3a202020",
  3133 => x"20202000",
  3134 => x"0a6d6469",
  3135 => x"6f5f636f",
  3136 => x"6e74726f",
  3137 => x"6c3a2000",
  3138 => x"0a74785f",
  3139 => x"706f696e",
  3140 => x"7465723a",
  3141 => x"20202000",
  3142 => x"0a72785f",
  3143 => x"706f696e",
  3144 => x"7465723a",
  3145 => x"20202000",
  3146 => x"0a656463",
  3147 => x"6c5f6970",
  3148 => x"3a202020",
  3149 => x"20202000",
  3150 => x"0a686173",
  3151 => x"685f6d73",
  3152 => x"623a2020",
  3153 => x"20202000",
  3154 => x"0a686173",
  3155 => x"685f6c73",
  3156 => x"623a2020",
  3157 => x"20202000",
  3158 => x"0a6d6469",
  3159 => x"6f207068",
  3160 => x"79207265",
  3161 => x"67697374",
  3162 => x"65727300",
  3163 => x"0a206d64",
  3164 => x"696f2070",
  3165 => x"68793a20",
  3166 => x"00000000",
  3167 => x"0a202072",
  3168 => x"65673a20",
  3169 => x"00000000",
  3170 => x"2d3e2000",
  3171 => x"0a677265",
  3172 => x"74682d3e",
  3173 => x"636f6e74",
  3174 => x"726f6c20",
  3175 => x"3a000000",
  3176 => x"0a677265",
  3177 => x"74682d3e",
  3178 => x"73746174",
  3179 => x"75732020",
  3180 => x"3a000000",
  3181 => x"0a646573",
  3182 => x"63722d3e",
  3183 => x"636f6e74",
  3184 => x"726f6c20",
  3185 => x"3a000000",
  3186 => x"0a0a0000",
  3187 => x"74657374",
  3188 => x"2e632000",
  3189 => x"286f6e20",
  3190 => x"73696d75",
  3191 => x"6c61746f",
  3192 => x"72290a00",
  3193 => x"636f6d70",
  3194 => x"696c6564",
  3195 => x"3a204175",
  3196 => x"67203138",
  3197 => x"20323031",
  3198 => x"30202031",
  3199 => x"343a3532",
  3200 => x"3a35340a",
  3201 => x"00000000",
  3202 => x"286f6e20",
  3203 => x"68617264",
  3204 => x"77617265",
  3205 => x"290a0000",
  3206 => x"000008b4",
  3207 => x"000008da",
  3208 => x"000008da",
  3209 => x"000008b4",
  3210 => x"000008da",
  3211 => x"000008da",
  3212 => x"000008da",
  3213 => x"000008da",
  3214 => x"000008da",
  3215 => x"000008da",
  3216 => x"000008da",
  3217 => x"000008da",
  3218 => x"000008da",
  3219 => x"000008da",
  3220 => x"000008da",
  3221 => x"000008da",
  3222 => x"000008da",
  3223 => x"000008da",
  3224 => x"000008da",
  3225 => x"000008da",
  3226 => x"000008da",
  3227 => x"000008da",
  3228 => x"000008da",
  3229 => x"000008da",
  3230 => x"000008da",
  3231 => x"000008da",
  3232 => x"000008da",
  3233 => x"000008da",
  3234 => x"000008da",
  3235 => x"000008da",
  3236 => x"000008da",
  3237 => x"000008da",
  3238 => x"000008da",
  3239 => x"000008da",
  3240 => x"000008da",
  3241 => x"000008da",
  3242 => x"000008da",
  3243 => x"000008da",
  3244 => x"00000986",
  3245 => x"0000097e",
  3246 => x"00000976",
  3247 => x"0000096e",
  3248 => x"00000966",
  3249 => x"0000095e",
  3250 => x"00000956",
  3251 => x"0000094d",
  3252 => x"00000944",
  3253 => x"43000000",
  3254 => x"64756d6d",
  3255 => x"792e6578",
  3256 => x"65000000",
  3257 => x"00ffffff",
  3258 => x"ff00ffff",
  3259 => x"ffff00ff",
  3260 => x"ffffff00",
  3261 => x"00000000",
  3262 => x"00000000",
  3263 => x"00000000",
  3264 => x"00003aec",
  3265 => x"80000c00",
  3266 => x"80000800",
  3267 => x"80000200",
  3268 => x"80000100",
  3269 => x"00000040",
  3270 => x"0000331c",
  3271 => x"00000000",
  3272 => x"00003584",
  3273 => x"000035e0",
  3274 => x"0000363c",
  3275 => x"00000000",
  3276 => x"00000000",
  3277 => x"00000000",
  3278 => x"00000000",
  3279 => x"00000000",
  3280 => x"00000000",
  3281 => x"00000000",
  3282 => x"00000000",
  3283 => x"00000000",
  3284 => x"000032d4",
  3285 => x"00000000",
  3286 => x"00000000",
  3287 => x"00000000",
  3288 => x"00000000",
  3289 => x"00000000",
  3290 => x"00000000",
  3291 => x"00000000",
  3292 => x"00000000",
  3293 => x"00000000",
  3294 => x"00000000",
  3295 => x"00000000",
  3296 => x"00000000",
  3297 => x"00000000",
  3298 => x"00000000",
  3299 => x"00000000",
  3300 => x"00000000",
  3301 => x"00000000",
  3302 => x"00000000",
  3303 => x"00000000",
  3304 => x"00000000",
  3305 => x"00000000",
  3306 => x"00000000",
  3307 => x"00000000",
  3308 => x"00000000",
  3309 => x"00000000",
  3310 => x"00000000",
  3311 => x"00000000",
  3312 => x"00000000",
  3313 => x"00000001",
  3314 => x"330eabcd",
  3315 => x"1234e66d",
  3316 => x"deec0005",
  3317 => x"000b0000",
  3318 => x"00000000",
  3319 => x"00000000",
  3320 => x"00000000",
  3321 => x"00000000",
  3322 => x"00000000",
  3323 => x"00000000",
  3324 => x"00000000",
  3325 => x"00000000",
  3326 => x"00000000",
  3327 => x"00000000",
  3328 => x"00000000",
  3329 => x"00000000",
  3330 => x"00000000",
  3331 => x"00000000",
  3332 => x"00000000",
  3333 => x"00000000",
  3334 => x"00000000",
  3335 => x"00000000",
  3336 => x"00000000",
  3337 => x"00000000",
  3338 => x"00000000",
  3339 => x"00000000",
  3340 => x"00000000",
  3341 => x"00000000",
  3342 => x"00000000",
  3343 => x"00000000",
  3344 => x"00000000",
  3345 => x"00000000",
  3346 => x"00000000",
  3347 => x"00000000",
  3348 => x"00000000",
  3349 => x"00000000",
  3350 => x"00000000",
  3351 => x"00000000",
  3352 => x"00000000",
  3353 => x"00000000",
  3354 => x"00000000",
  3355 => x"00000000",
  3356 => x"00000000",
  3357 => x"00000000",
  3358 => x"00000000",
  3359 => x"00000000",
  3360 => x"00000000",
  3361 => x"00000000",
  3362 => x"00000000",
  3363 => x"00000000",
  3364 => x"00000000",
  3365 => x"00000000",
  3366 => x"00000000",
  3367 => x"00000000",
  3368 => x"00000000",
  3369 => x"00000000",
  3370 => x"00000000",
  3371 => x"00000000",
  3372 => x"00000000",
  3373 => x"00000000",
  3374 => x"00000000",
  3375 => x"00000000",
  3376 => x"00000000",
  3377 => x"00000000",
  3378 => x"00000000",
  3379 => x"00000000",
  3380 => x"00000000",
  3381 => x"00000000",
  3382 => x"00000000",
  3383 => x"00000000",
  3384 => x"00000000",
  3385 => x"00000000",
  3386 => x"00000000",
  3387 => x"00000000",
  3388 => x"00000000",
  3389 => x"00000000",
  3390 => x"00000000",
  3391 => x"00000000",
  3392 => x"00000000",
  3393 => x"00000000",
  3394 => x"00000000",
  3395 => x"00000000",
  3396 => x"00000000",
  3397 => x"00000000",
  3398 => x"00000000",
  3399 => x"00000000",
  3400 => x"00000000",
  3401 => x"00000000",
  3402 => x"00000000",
  3403 => x"00000000",
  3404 => x"00000000",
  3405 => x"00000000",
  3406 => x"00000000",
  3407 => x"00000000",
  3408 => x"00000000",
  3409 => x"00000000",
  3410 => x"00000000",
  3411 => x"00000000",
  3412 => x"00000000",
  3413 => x"00000000",
  3414 => x"00000000",
  3415 => x"00000000",
  3416 => x"00000000",
  3417 => x"00000000",
  3418 => x"00000000",
  3419 => x"00000000",
  3420 => x"00000000",
  3421 => x"00000000",
  3422 => x"00000000",
  3423 => x"00000000",
  3424 => x"00000000",
  3425 => x"00000000",
  3426 => x"00000000",
  3427 => x"00000000",
  3428 => x"00000000",
  3429 => x"00000000",
  3430 => x"00000000",
  3431 => x"00000000",
  3432 => x"00000000",
  3433 => x"00000000",
  3434 => x"00000000",
  3435 => x"00000000",
  3436 => x"00000000",
  3437 => x"00000000",
  3438 => x"00000000",
  3439 => x"00000000",
  3440 => x"00000000",
  3441 => x"00000000",
  3442 => x"00000000",
  3443 => x"00000000",
  3444 => x"00000000",
  3445 => x"00000000",
  3446 => x"00000000",
  3447 => x"00000000",
  3448 => x"00000000",
  3449 => x"00000000",
  3450 => x"00000000",
  3451 => x"00000000",
  3452 => x"00000000",
  3453 => x"00000000",
  3454 => x"00000000",
  3455 => x"00000000",
  3456 => x"00000000",
  3457 => x"00000000",
  3458 => x"00000000",
  3459 => x"00000000",
  3460 => x"00000000",
  3461 => x"00000000",
  3462 => x"00000000",
  3463 => x"00000000",
  3464 => x"00000000",
  3465 => x"00000000",
  3466 => x"00000000",
  3467 => x"00000000",
  3468 => x"00000000",
  3469 => x"00000000",
  3470 => x"00000000",
  3471 => x"00000000",
  3472 => x"00000000",
  3473 => x"00000000",
  3474 => x"00000000",
  3475 => x"00000000",
  3476 => x"00000000",
  3477 => x"00000000",
  3478 => x"00000000",
  3479 => x"00000000",
  3480 => x"00000000",
  3481 => x"00000000",
  3482 => x"00000000",
  3483 => x"00000000",
  3484 => x"00000000",
  3485 => x"00000000",
  3486 => x"00000000",
  3487 => x"00000000",
  3488 => x"00000000",
  3489 => x"00000000",
  3490 => x"00000000",
  3491 => x"00000000",
  3492 => x"00000000",
  3493 => x"00000000",
  3494 => x"00000000",
  3495 => x"00000000",
  3496 => x"00000000",
  3497 => x"00000000",
  3498 => x"00000000",
  3499 => x"00000000",
  3500 => x"00000000",
  3501 => x"00000000",
  3502 => x"00000000",
  3503 => x"00000000",
  3504 => x"00000000",
  3505 => x"00000000",
  3506 => x"ffffffff",
  3507 => x"00000000",
  3508 => x"00020000",
  3509 => x"00000000",
  3510 => x"00000000",
  3511 => x"000036d4",
  3512 => x"000036d4",
  3513 => x"000036dc",
  3514 => x"000036dc",
  3515 => x"000036e4",
  3516 => x"000036e4",
  3517 => x"000036ec",
  3518 => x"000036ec",
  3519 => x"000036f4",
  3520 => x"000036f4",
  3521 => x"000036fc",
  3522 => x"000036fc",
  3523 => x"00003704",
  3524 => x"00003704",
  3525 => x"0000370c",
  3526 => x"0000370c",
  3527 => x"00003714",
  3528 => x"00003714",
  3529 => x"0000371c",
  3530 => x"0000371c",
  3531 => x"00003724",
  3532 => x"00003724",
  3533 => x"0000372c",
  3534 => x"0000372c",
  3535 => x"00003734",
  3536 => x"00003734",
  3537 => x"0000373c",
  3538 => x"0000373c",
  3539 => x"00003744",
  3540 => x"00003744",
  3541 => x"0000374c",
  3542 => x"0000374c",
  3543 => x"00003754",
  3544 => x"00003754",
  3545 => x"0000375c",
  3546 => x"0000375c",
  3547 => x"00003764",
  3548 => x"00003764",
  3549 => x"0000376c",
  3550 => x"0000376c",
  3551 => x"00003774",
  3552 => x"00003774",
  3553 => x"0000377c",
  3554 => x"0000377c",
  3555 => x"00003784",
  3556 => x"00003784",
  3557 => x"0000378c",
  3558 => x"0000378c",
  3559 => x"00003794",
  3560 => x"00003794",
  3561 => x"0000379c",
  3562 => x"0000379c",
  3563 => x"000037a4",
  3564 => x"000037a4",
  3565 => x"000037ac",
  3566 => x"000037ac",
  3567 => x"000037b4",
  3568 => x"000037b4",
  3569 => x"000037bc",
  3570 => x"000037bc",
  3571 => x"000037c4",
  3572 => x"000037c4",
  3573 => x"000037cc",
  3574 => x"000037cc",
  3575 => x"000037d4",
  3576 => x"000037d4",
  3577 => x"000037dc",
  3578 => x"000037dc",
  3579 => x"000037e4",
  3580 => x"000037e4",
  3581 => x"000037ec",
  3582 => x"000037ec",
  3583 => x"000037f4",
  3584 => x"000037f4",
  3585 => x"000037fc",
  3586 => x"000037fc",
  3587 => x"00003804",
  3588 => x"00003804",
  3589 => x"0000380c",
  3590 => x"0000380c",
  3591 => x"00003814",
  3592 => x"00003814",
  3593 => x"0000381c",
  3594 => x"0000381c",
  3595 => x"00003824",
  3596 => x"00003824",
  3597 => x"0000382c",
  3598 => x"0000382c",
  3599 => x"00003834",
  3600 => x"00003834",
  3601 => x"0000383c",
  3602 => x"0000383c",
  3603 => x"00003844",
  3604 => x"00003844",
  3605 => x"0000384c",
  3606 => x"0000384c",
  3607 => x"00003854",
  3608 => x"00003854",
  3609 => x"0000385c",
  3610 => x"0000385c",
  3611 => x"00003864",
  3612 => x"00003864",
  3613 => x"0000386c",
  3614 => x"0000386c",
  3615 => x"00003874",
  3616 => x"00003874",
  3617 => x"0000387c",
  3618 => x"0000387c",
  3619 => x"00003884",
  3620 => x"00003884",
  3621 => x"0000388c",
  3622 => x"0000388c",
  3623 => x"00003894",
  3624 => x"00003894",
  3625 => x"0000389c",
  3626 => x"0000389c",
  3627 => x"000038a4",
  3628 => x"000038a4",
  3629 => x"000038ac",
  3630 => x"000038ac",
  3631 => x"000038b4",
  3632 => x"000038b4",
  3633 => x"000038bc",
  3634 => x"000038bc",
  3635 => x"000038c4",
  3636 => x"000038c4",
  3637 => x"000038cc",
  3638 => x"000038cc",
  3639 => x"000038d4",
  3640 => x"000038d4",
  3641 => x"000038dc",
  3642 => x"000038dc",
  3643 => x"000038e4",
  3644 => x"000038e4",
  3645 => x"000038ec",
  3646 => x"000038ec",
  3647 => x"000038f4",
  3648 => x"000038f4",
  3649 => x"000038fc",
  3650 => x"000038fc",
  3651 => x"00003904",
  3652 => x"00003904",
  3653 => x"0000390c",
  3654 => x"0000390c",
  3655 => x"00003914",
  3656 => x"00003914",
  3657 => x"0000391c",
  3658 => x"0000391c",
  3659 => x"00003924",
  3660 => x"00003924",
  3661 => x"0000392c",
  3662 => x"0000392c",
  3663 => x"00003934",
  3664 => x"00003934",
  3665 => x"0000393c",
  3666 => x"0000393c",
  3667 => x"00003944",
  3668 => x"00003944",
  3669 => x"0000394c",
  3670 => x"0000394c",
  3671 => x"00003954",
  3672 => x"00003954",
  3673 => x"0000395c",
  3674 => x"0000395c",
  3675 => x"00003964",
  3676 => x"00003964",
  3677 => x"0000396c",
  3678 => x"0000396c",
  3679 => x"00003974",
  3680 => x"00003974",
  3681 => x"0000397c",
  3682 => x"0000397c",
  3683 => x"00003984",
  3684 => x"00003984",
  3685 => x"0000398c",
  3686 => x"0000398c",
  3687 => x"00003994",
  3688 => x"00003994",
  3689 => x"0000399c",
  3690 => x"0000399c",
  3691 => x"000039a4",
  3692 => x"000039a4",
  3693 => x"000039ac",
  3694 => x"000039ac",
  3695 => x"000039b4",
  3696 => x"000039b4",
  3697 => x"000039bc",
  3698 => x"000039bc",
  3699 => x"000039c4",
  3700 => x"000039c4",
  3701 => x"000039cc",
  3702 => x"000039cc",
  3703 => x"000039d4",
  3704 => x"000039d4",
  3705 => x"000039dc",
  3706 => x"000039dc",
  3707 => x"000039e4",
  3708 => x"000039e4",
  3709 => x"000039ec",
  3710 => x"000039ec",
  3711 => x"000039f4",
  3712 => x"000039f4",
  3713 => x"000039fc",
  3714 => x"000039fc",
  3715 => x"00003a04",
  3716 => x"00003a04",
  3717 => x"00003a0c",
  3718 => x"00003a0c",
  3719 => x"00003a14",
  3720 => x"00003a14",
  3721 => x"00003a1c",
  3722 => x"00003a1c",
  3723 => x"00003a24",
  3724 => x"00003a24",
  3725 => x"00003a2c",
  3726 => x"00003a2c",
  3727 => x"00003a34",
  3728 => x"00003a34",
  3729 => x"00003a3c",
  3730 => x"00003a3c",
  3731 => x"00003a44",
  3732 => x"00003a44",
  3733 => x"00003a4c",
  3734 => x"00003a4c",
  3735 => x"00003a54",
  3736 => x"00003a54",
  3737 => x"00003a5c",
  3738 => x"00003a5c",
  3739 => x"00003a64",
  3740 => x"00003a64",
  3741 => x"00003a6c",
  3742 => x"00003a6c",
  3743 => x"00003a74",
  3744 => x"00003a74",
  3745 => x"00003a7c",
  3746 => x"00003a7c",
  3747 => x"00003a84",
  3748 => x"00003a84",
  3749 => x"00003a8c",
  3750 => x"00003a8c",
  3751 => x"00003a94",
  3752 => x"00003a94",
  3753 => x"00003a9c",
  3754 => x"00003a9c",
  3755 => x"00003aa4",
  3756 => x"00003aa4",
  3757 => x"00003aac",
  3758 => x"00003aac",
  3759 => x"00003ab4",
  3760 => x"00003ab4",
  3761 => x"00003abc",
  3762 => x"00003abc",
  3763 => x"00003ac4",
  3764 => x"00003ac4",
  3765 => x"00003acc",
  3766 => x"00003acc",
  3767 => x"000032d8",
  3768 => x"ffffffff",
  3769 => x"00000000",
  3770 => x"ffffffff",
  3771 => x"00000000",
  3772 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
