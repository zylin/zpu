-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80ddc80c",
     3 => x"3a0b0b80",
     4 => x"d8990400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80d8e42d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80dd",
   162 => x"b4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0bbc",
   171 => x"fb2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bbe",
   179 => x"ad2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80ddc40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"d2853f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80ddc408",
   281 => x"802ea438",
   282 => x"80ddc808",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80e5",
   286 => x"800c82a0",
   287 => x"800b80e5",
   288 => x"840c8290",
   289 => x"800b80e5",
   290 => x"880c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"e5800cf8",
   294 => x"80808280",
   295 => x"0b80e584",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"e5880c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80e5800c",
   302 => x"80c0a880",
   303 => x"940b80e5",
   304 => x"840c0b0b",
   305 => x"80dab80b",
   306 => x"80e5880c",
   307 => x"04ff3d0d",
   308 => x"80e58c33",
   309 => x"5170a738",
   310 => x"80ddd008",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"ddd00c70",
   315 => x"2d80ddd0",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80e5",
   319 => x"8c34833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80e4fc08",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"e4fc510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404ff3d",
   333 => x"0d028f05",
   334 => x"33705252",
   335 => x"95ef3f71",
   336 => x"5196e53f",
   337 => x"71800c83",
   338 => x"3d0d04f6",
   339 => x"3d0d7c57",
   340 => x"80707179",
   341 => x"08700870",
   342 => x"9b2a8106",
   343 => x"8c1d0c70",
   344 => x"9f2a7094",
   345 => x"1e0c5859",
   346 => x"5b5d5b59",
   347 => x"72792e09",
   348 => x"81069138",
   349 => x"80c0780c",
   350 => x"77087086",
   351 => x"2a810657",
   352 => x"5575f538",
   353 => x"90187008",
   354 => x"708b2a9f",
   355 => x"06901a0c",
   356 => x"5556850a",
   357 => x"0b98180c",
   358 => x"850a0b9c",
   359 => x"180c9418",
   360 => x"53850a73",
   361 => x"0c981854",
   362 => x"850a740c",
   363 => x"800ba018",
   364 => x"0c800ba4",
   365 => x"180c800b",
   366 => x"a8180c80",
   367 => x"0bac180c",
   368 => x"80765555",
   369 => x"94170875",
   370 => x"2e098106",
   371 => x"84de3890",
   372 => x"17085475",
   373 => x"0870832a",
   374 => x"81065153",
   375 => x"72f53873",
   376 => x"8b2bf880",
   377 => x"80808107",
   378 => x"760c7508",
   379 => x"70832a81",
   380 => x"06555573",
   381 => x"f5389018",
   382 => x"56901708",
   383 => x"54750870",
   384 => x"832a8106",
   385 => x"515372f5",
   386 => x"38738b2b",
   387 => x"8207760c",
   388 => x"75087083",
   389 => x"2a810654",
   390 => x"5472f538",
   391 => x"73842a81",
   392 => x"0653ff54",
   393 => x"72883875",
   394 => x"0870902a",
   395 => x"5553738f",
   396 => x"2a810653",
   397 => x"72c33872",
   398 => x"748c2a81",
   399 => x"06575575",
   400 => x"802e859a",
   401 => x"38901708",
   402 => x"90195754",
   403 => x"75087083",
   404 => x"2a810651",
   405 => x"5b7af538",
   406 => x"738b2b80",
   407 => x"c207760c",
   408 => x"75087083",
   409 => x"2a81065c",
   410 => x"547af538",
   411 => x"73842a81",
   412 => x"065bff54",
   413 => x"7a883875",
   414 => x"0870902a",
   415 => x"555b7385",
   416 => x"2c810654",
   417 => x"73963881",
   418 => x"15558386",
   419 => x"d07525ff",
   420 => x"b43880da",
   421 => x"bc518fab",
   422 => x"3f760858",
   423 => x"800b9018",
   424 => x"08901a58",
   425 => x"555b7508",
   426 => x"70832a81",
   427 => x"06515574",
   428 => x"f538738b",
   429 => x"2b828207",
   430 => x"760c7508",
   431 => x"70832a81",
   432 => x"06565474",
   433 => x"f5387384",
   434 => x"2a810654",
   435 => x"ff557388",
   436 => x"38750870",
   437 => x"902a5653",
   438 => x"90170890",
   439 => x"19575475",
   440 => x"0870832a",
   441 => x"70810651",
   442 => x"515372f3",
   443 => x"38738b2b",
   444 => x"82c20776",
   445 => x"0c750870",
   446 => x"832a7081",
   447 => x"06515454",
   448 => x"72f33873",
   449 => x"842a7081",
   450 => x"065153ff",
   451 => x"54728838",
   452 => x"75087090",
   453 => x"2a555374",
   454 => x"882a8106",
   455 => x"5675802e",
   456 => x"90387388",
   457 => x"2a810656",
   458 => x"75802e85",
   459 => x"3881705b",
   460 => x"5974872a",
   461 => x"81065675",
   462 => x"802e9038",
   463 => x"73872a81",
   464 => x"06567580",
   465 => x"2e853881",
   466 => x"5a805974",
   467 => x"862a8106",
   468 => x"5574802e",
   469 => x"8e387386",
   470 => x"2a810654",
   471 => x"73802e83",
   472 => x"38815978",
   473 => x"842b7a87",
   474 => x"2b077b88",
   475 => x"2b07780c",
   476 => x"80dad851",
   477 => x"8dcd3f8c",
   478 => x"1708802e",
   479 => x"81c03880",
   480 => x"dae0518d",
   481 => x"be3f80da",
   482 => x"ec518db7",
   483 => x"3f760852",
   484 => x"a0518dd2",
   485 => x"3f80db84",
   486 => x"518da83f",
   487 => x"79802e81",
   488 => x"be3880db",
   489 => x"90518d9b",
   490 => x"3f80db94",
   491 => x"518d943f",
   492 => x"78802e81",
   493 => x"bc3880db",
   494 => x"9c518d87",
   495 => x"3f80dba4",
   496 => x"518d803f",
   497 => x"84175b81",
   498 => x"1b338518",
   499 => x"34821b33",
   500 => x"86183483",
   501 => x"1b338718",
   502 => x"34841b33",
   503 => x"88183485",
   504 => x"1b338918",
   505 => x"34760888",
   506 => x"117c3381",
   507 => x"1e337188",
   508 => x"2b07720c",
   509 => x"555b8c05",
   510 => x"821c3383",
   511 => x"1d337198",
   512 => x"2b71902b",
   513 => x"07841f33",
   514 => x"70882b72",
   515 => x"07608505",
   516 => x"33710776",
   517 => x"0c5e5c56",
   518 => x"59575a81",
   519 => x"0b800c8c",
   520 => x"3d0d0481",
   521 => x"15557482",
   522 => x"24fec538",
   523 => x"73087083",
   524 => x"2a810659",
   525 => x"5677802e",
   526 => x"ea388055",
   527 => x"ef3980db",
   528 => x"b0518bff",
   529 => x"3f80daec",
   530 => x"518bf83f",
   531 => x"760852a0",
   532 => x"518c933f",
   533 => x"80db8451",
   534 => x"8be93f79",
   535 => x"fec43880",
   536 => x"dbb8518b",
   537 => x"de3f80db",
   538 => x"94518bd7",
   539 => x"3f78fec6",
   540 => x"3880dbbc",
   541 => x"518bcc3f",
   542 => x"80dba451",
   543 => x"8bc53f84",
   544 => x"175b811b",
   545 => x"33851834",
   546 => x"821b3386",
   547 => x"1834831b",
   548 => x"33871834",
   549 => x"841b3388",
   550 => x"1834851b",
   551 => x"33891834",
   552 => x"76088811",
   553 => x"7c33811e",
   554 => x"3371882b",
   555 => x"07720c55",
   556 => x"5b8c0582",
   557 => x"1c33831d",
   558 => x"3371982b",
   559 => x"71902b07",
   560 => x"841f3370",
   561 => x"882b7207",
   562 => x"60850533",
   563 => x"7107760c",
   564 => x"5e5c5659",
   565 => x"575a810b",
   566 => x"800c8c3d",
   567 => x"0d049017",
   568 => x"08901957",
   569 => x"54750870",
   570 => x"832a8106",
   571 => x"5a5378f5",
   572 => x"38738b2b",
   573 => x"8207760c",
   574 => x"75087083",
   575 => x"2a810656",
   576 => x"5474f538",
   577 => x"73842a81",
   578 => x"0654ff55",
   579 => x"73883875",
   580 => x"0870902a",
   581 => x"5653748d",
   582 => x"2a548c17",
   583 => x"08802e92",
   584 => x"38738106",
   585 => x"56758b38",
   586 => x"74862a81",
   587 => x"06597880",
   588 => x"c9387381",
   589 => x"06567580",
   590 => x"2ea43874",
   591 => x"862a8106",
   592 => x"53729b38",
   593 => x"725b815a",
   594 => x"74882a81",
   595 => x"06597884",
   596 => x"2b7a872b",
   597 => x"077b882b",
   598 => x"07780cfc",
   599 => x"93397381",
   600 => x"065372e4",
   601 => x"3874862a",
   602 => x"81065372",
   603 => x"db387273",
   604 => x"76882a81",
   605 => x"065b5c5a",
   606 => x"d5398176",
   607 => x"76882a81",
   608 => x"065b5b5b",
   609 => x"c939ff3d",
   610 => x"0d739811",
   611 => x"085151bf",
   612 => x"5280710c",
   613 => x"ff128812",
   614 => x"52527180",
   615 => x"25f33883",
   616 => x"3d0d04fb",
   617 => x"3d0d777a",
   618 => x"981108a0",
   619 => x"12081010",
   620 => x"10117008",
   621 => x"708b2a81",
   622 => x"06515956",
   623 => x"54555680",
   624 => x"5174712e",
   625 => x"098106ad",
   626 => x"38788414",
   627 => x"0ca01408",
   628 => x"5170bf2e",
   629 => x"a7387010",
   630 => x"10101276",
   631 => x"90800771",
   632 => x"0c55a014",
   633 => x"088105a0",
   634 => x"150c7308",
   635 => x"70088107",
   636 => x"710c5681",
   637 => x"5170800c",
   638 => x"873d0d04",
   639 => x"83f81276",
   640 => x"b0800771",
   641 => x"0c5274a0",
   642 => x"150c7308",
   643 => x"70088107",
   644 => x"710c5681",
   645 => x"51df39e9",
   646 => x"3d0d80dd",
   647 => x"d8087008",
   648 => x"810a065c",
   649 => x"5781ff0b",
   650 => x"88180c8c",
   651 => x"d73f8bb6",
   652 => x"3f8be43f",
   653 => x"9c93567a",
   654 => x"84388ab2",
   655 => x"567580e5",
   656 => x"c00c80db",
   657 => x"c45187fb",
   658 => x"3f7a802e",
   659 => x"84ef3880",
   660 => x"dbd05187",
   661 => x"ee3ff880",
   662 => x"8098800b",
   663 => x"80e5900c",
   664 => x"800bfa80",
   665 => x"80858034",
   666 => x"9b0bfa80",
   667 => x"80858134",
   668 => x"a10bfa80",
   669 => x"80858234",
   670 => x"80e70bfa",
   671 => x"80808583",
   672 => x"34ffb80b",
   673 => x"fa808085",
   674 => x"8434ffb8",
   675 => x"0bfa8080",
   676 => x"858534de",
   677 => x"0bfa8080",
   678 => x"858634ff",
   679 => x"ad0bfa80",
   680 => x"80858734",
   681 => x"ffbe0bfa",
   682 => x"80808588",
   683 => x"34ef0bfa",
   684 => x"80808589",
   685 => x"34800bfa",
   686 => x"8080858a",
   687 => x"34a00bfa",
   688 => x"8080858b",
   689 => x"34850bfa",
   690 => x"8080858c",
   691 => x"34dc0bfa",
   692 => x"8080858d",
   693 => x"3480ddd8",
   694 => x"0858810b",
   695 => x"84190c86",
   696 => x"53fa8080",
   697 => x"85865280",
   698 => x"e5945180",
   699 => x"c1923f80",
   700 => x"ddd80856",
   701 => x"820b8417",
   702 => x"0c80598e",
   703 => x"5a7aab38",
   704 => x"fa808085",
   705 => x"801a5d79",
   706 => x"7d34811a",
   707 => x"7a71267a",
   708 => x"0570725d",
   709 => x"5b585876",
   710 => x"80268a38",
   711 => x"76e2388b",
   712 => x"e97827dc",
   713 => x"3880ddd8",
   714 => x"0856830b",
   715 => x"84170c80",
   716 => x"e59051f4",
   717 => x"963f80e5",
   718 => x"9051fcca",
   719 => x"3f80ddd8",
   720 => x"0859840b",
   721 => x"841a0c80",
   722 => x"dbdc5185",
   723 => x"f63f8059",
   724 => x"805afa80",
   725 => x"8085801a",
   726 => x"7033535e",
   727 => x"88518686",
   728 => x"3f788638",
   729 => x"79852e86",
   730 => x"38ba5185",
   731 => x"bc3f811a",
   732 => x"7a71267a",
   733 => x"0570725d",
   734 => x"5b585876",
   735 => x"80268938",
   736 => x"76d03885",
   737 => x"7827cb38",
   738 => x"8a51859d",
   739 => x"3f805d83",
   740 => x"5e7a8738",
   741 => x"805d9080",
   742 => x"0a5ea851",
   743 => x"858b3f7d",
   744 => x"5186e53f",
   745 => x"80dbfc51",
   746 => x"85993f80",
   747 => x"5b805c88",
   748 => x"a43f8008",
   749 => x"40888d3f",
   750 => x"80085f7c",
   751 => x"80268b38",
   752 => x"7c80cb38",
   753 => x"807e2780",
   754 => x"c53880e5",
   755 => x"b33380dd",
   756 => x"d8085b84",
   757 => x"1b0c80e5",
   758 => x"9053fa80",
   759 => x"80858052",
   760 => x"8bea51fb",
   761 => x"be3f8008",
   762 => x"9f2c8008",
   763 => x"1d7d7126",
   764 => x"5a5b7b05",
   765 => x"7805707b",
   766 => x"5e5c597c",
   767 => x"7926cb38",
   768 => x"7c792e09",
   769 => x"81068738",
   770 => x"7d7a26ff",
   771 => x"bd3887b4",
   772 => x"3f80085b",
   773 => x"87bf3f80",
   774 => x"ddd8085c",
   775 => x"81ff0b84",
   776 => x"1d0c7f80",
   777 => x"08317f7c",
   778 => x"31575880",
   779 => x"762482e4",
   780 => x"3880dc88",
   781 => x"51848c3f",
   782 => x"775185cc",
   783 => x"3fae5183",
   784 => x"e83f7551",
   785 => x"85c23f80",
   786 => x"dc905183",
   787 => x"f63f87e8",
   788 => x"527551a4",
   789 => x"a63f8008",
   790 => x"1852993d",
   791 => x"f805519d",
   792 => x"da3f805c",
   793 => x"807c5454",
   794 => x"825780f7",
   795 => x"0a775252",
   796 => x"8baf3f66",
   797 => x"685a5478",
   798 => x"55bbc0c2",
   799 => x"0a588078",
   800 => x"5353993d",
   801 => x"e005518d",
   802 => x"833f6062",
   803 => x"80dc9853",
   804 => x"5e5e83af",
   805 => x"3f7d517c",
   806 => x"529f9b3f",
   807 => x"80085680",
   808 => x"0b800824",
   809 => x"81d23875",
   810 => x"8a2c5184",
   811 => x"db3f80dc",
   812 => x"a451838f",
   813 => x"3f800b80",
   814 => x"0c993d0d",
   815 => x"0480dcac",
   816 => x"5183803f",
   817 => x"80dcbc51",
   818 => x"82f93ff8",
   819 => x"80809880",
   820 => x"0b80e590",
   821 => x"0c800bfa",
   822 => x"80808580",
   823 => x"349b0bfa",
   824 => x"80808581",
   825 => x"34a10bfa",
   826 => x"80808582",
   827 => x"3480e70b",
   828 => x"fa808085",
   829 => x"8334ffb8",
   830 => x"0bfa8080",
   831 => x"858434ff",
   832 => x"b80bfa80",
   833 => x"80858534",
   834 => x"de0bfa80",
   835 => x"80858634",
   836 => x"ffad0bfa",
   837 => x"80808587",
   838 => x"34ffbe0b",
   839 => x"fa808085",
   840 => x"8834ef0b",
   841 => x"fa808085",
   842 => x"8934800b",
   843 => x"fa808085",
   844 => x"8a34a00b",
   845 => x"fa808085",
   846 => x"8b34850b",
   847 => x"fa808085",
   848 => x"8c34dc0b",
   849 => x"fa808085",
   850 => x"8d3480dd",
   851 => x"d8085881",
   852 => x"0b84190c",
   853 => x"8653fa80",
   854 => x"80858652",
   855 => x"80e59451",
   856 => x"bc9e3f80",
   857 => x"ddd80856",
   858 => x"820b8417",
   859 => x"0c80598e",
   860 => x"5a7afbb6",
   861 => x"38fb8939",
   862 => x"800887ff",
   863 => x"05708a2c",
   864 => x"52568384",
   865 => x"3f80dca4",
   866 => x"5181b83f",
   867 => x"800b800c",
   868 => x"993d0d04",
   869 => x"87e81681",
   870 => x"1980dc88",
   871 => x"53595681",
   872 => x"a23f7751",
   873 => x"82e23fae",
   874 => x"5180fe3f",
   875 => x"755182d8",
   876 => x"3f80dc90",
   877 => x"51818c3f",
   878 => x"87e85275",
   879 => x"51a1bc3f",
   880 => x"80081852",
   881 => x"993df805",
   882 => x"519af03f",
   883 => x"805c807c",
   884 => x"54548257",
   885 => x"80f70a77",
   886 => x"525288c5",
   887 => x"3f66685a",
   888 => x"547855bb",
   889 => x"c0c20a58",
   890 => x"80785353",
   891 => x"993de005",
   892 => x"518a993f",
   893 => x"606280dc",
   894 => x"98535e5e",
   895 => x"80c53f7d",
   896 => x"517c529c",
   897 => x"b13f8008",
   898 => x"56800880",
   899 => x"25fd9838",
   900 => x"fee639ff",
   901 => x"3d0d028f",
   902 => x"053380dd",
   903 => x"d4085271",
   904 => x"0c800b80",
   905 => x"0c833d0d",
   906 => x"04ff3d0d",
   907 => x"028f0533",
   908 => x"5180e5c0",
   909 => x"0852712d",
   910 => x"800881ff",
   911 => x"06800c83",
   912 => x"3d0d04fe",
   913 => x"3d0d7470",
   914 => x"33535371",
   915 => x"802e9338",
   916 => x"81137252",
   917 => x"80e5c008",
   918 => x"5353712d",
   919 => x"72335271",
   920 => x"ef38843d",
   921 => x"0d04f43d",
   922 => x"0d7f0284",
   923 => x"05bb0533",
   924 => x"5557880b",
   925 => x"8c3d5a5a",
   926 => x"895380dd",
   927 => x"84527851",
   928 => x"b9fe3f73",
   929 => x"7a2e80fa",
   930 => x"38795673",
   931 => x"902e80e7",
   932 => x"3802a705",
   933 => x"58768f06",
   934 => x"54738926",
   935 => x"bf387518",
   936 => x"b0155555",
   937 => x"73753476",
   938 => x"842aff17",
   939 => x"7081ff06",
   940 => x"58555775",
   941 => x"e0387919",
   942 => x"55757534",
   943 => x"78703355",
   944 => x"5573802e",
   945 => x"93388115",
   946 => x"745280e5",
   947 => x"c0085755",
   948 => x"752d7433",
   949 => x"5473ef38",
   950 => x"8e3d0d04",
   951 => x"7518b715",
   952 => x"55557375",
   953 => x"3476842a",
   954 => x"ff177081",
   955 => x"ff065855",
   956 => x"5775ffa1",
   957 => x"38c03984",
   958 => x"70575a02",
   959 => x"a70558ff",
   960 => x"94398270",
   961 => x"575af439",
   962 => x"f23d0d60",
   963 => x"8c3d705b",
   964 => x"5b538073",
   965 => x"56577673",
   966 => x"2480f838",
   967 => x"7817548a",
   968 => x"5274519e",
   969 => x"b13f8008",
   970 => x"b0055372",
   971 => x"74348117",
   972 => x"578a5274",
   973 => x"519dfa3f",
   974 => x"80085580",
   975 => x"08de3880",
   976 => x"08779f2a",
   977 => x"1870812c",
   978 => x"5a565680",
   979 => x"78259e38",
   980 => x"7817ff05",
   981 => x"55751970",
   982 => x"33555374",
   983 => x"33733473",
   984 => x"75348116",
   985 => x"ff165656",
   986 => x"777624e9",
   987 => x"38761956",
   988 => x"80763479",
   989 => x"70335454",
   990 => x"72802e93",
   991 => x"38811473",
   992 => x"5280e5c0",
   993 => x"08585476",
   994 => x"2d733353",
   995 => x"72ef3890",
   996 => x"3d0d04ad",
   997 => x"7a3402a9",
   998 => x"05733071",
   999 => x"19565659",
  1000 => x"8a527451",
  1001 => x"9db03f80",
  1002 => x"08b00553",
  1003 => x"72743481",
  1004 => x"17578a52",
  1005 => x"74519cf9",
  1006 => x"3f800855",
  1007 => x"8008fedc",
  1008 => x"38fefc39",
  1009 => x"803d0d80",
  1010 => x"dde008a0",
  1011 => x"1108800c",
  1012 => x"51823d0d",
  1013 => x"04803d0d",
  1014 => x"80dde008",
  1015 => x"b0110880",
  1016 => x"0c51823d",
  1017 => x"0d04803d",
  1018 => x"0d80dde0",
  1019 => x"0851870b",
  1020 => x"84120cb0",
  1021 => x"ea0b9412",
  1022 => x"0c870b98",
  1023 => x"120c87e8",
  1024 => x"0ba4120c",
  1025 => x"a70ba812",
  1026 => x"0cff0bb4",
  1027 => x"120ca70b",
  1028 => x"b8120c82",
  1029 => x"3d0d0480",
  1030 => x"3d0d80dd",
  1031 => x"e40851b6",
  1032 => x"0b8c120c",
  1033 => x"830b8812",
  1034 => x"0c823d0d",
  1035 => x"04fe3d0d",
  1036 => x"02930533",
  1037 => x"53728a2e",
  1038 => x"9e3880dd",
  1039 => x"e4085284",
  1040 => x"12087082",
  1041 => x"2a708106",
  1042 => x"51515170",
  1043 => x"802ef038",
  1044 => x"72720c84",
  1045 => x"3d0d0480",
  1046 => x"dde40852",
  1047 => x"84120870",
  1048 => x"822a7081",
  1049 => x"06515151",
  1050 => x"70802ef0",
  1051 => x"388d720c",
  1052 => x"84120870",
  1053 => x"822a7081",
  1054 => x"06515151",
  1055 => x"70802eff",
  1056 => x"be38cd39",
  1057 => x"803d0d80",
  1058 => x"dddc0851",
  1059 => x"800b8412",
  1060 => x"0cfe800a",
  1061 => x"0b88120c",
  1062 => x"800b80e5",
  1063 => x"c434800b",
  1064 => x"80e5c834",
  1065 => x"823d0d04",
  1066 => x"fa3d0d02",
  1067 => x"a3053380",
  1068 => x"dddc0880",
  1069 => x"e5c43370",
  1070 => x"81ff0670",
  1071 => x"10101180",
  1072 => x"e5c83370",
  1073 => x"81ff0672",
  1074 => x"90291170",
  1075 => x"882b7807",
  1076 => x"770c535b",
  1077 => x"5b555559",
  1078 => x"5454738a",
  1079 => x"2e983874",
  1080 => x"80cf2e92",
  1081 => x"38738c2e",
  1082 => x"a4388116",
  1083 => x"537280e5",
  1084 => x"c834883d",
  1085 => x"0d0471a3",
  1086 => x"26a33881",
  1087 => x"17527180",
  1088 => x"e5c43480",
  1089 => x"0b80e5c8",
  1090 => x"34883d0d",
  1091 => x"04805271",
  1092 => x"882b730c",
  1093 => x"81125297",
  1094 => x"907226f3",
  1095 => x"38800b80",
  1096 => x"e5c43480",
  1097 => x"0b80e5c8",
  1098 => x"34df398c",
  1099 => x"08028c0c",
  1100 => x"f53d0d8c",
  1101 => x"08940508",
  1102 => x"9d388c08",
  1103 => x"8c05088c",
  1104 => x"08900508",
  1105 => x"8c088805",
  1106 => x"08585654",
  1107 => x"73760c74",
  1108 => x"84170c81",
  1109 => x"bf39800b",
  1110 => x"8c08f005",
  1111 => x"0c800b8c",
  1112 => x"08f4050c",
  1113 => x"8c088c05",
  1114 => x"088c0890",
  1115 => x"05085654",
  1116 => x"738c08f0",
  1117 => x"050c748c",
  1118 => x"08f4050c",
  1119 => x"8c08f805",
  1120 => x"8c08f005",
  1121 => x"56568870",
  1122 => x"54755376",
  1123 => x"5254b3f0",
  1124 => x"3fa00b8c",
  1125 => x"08940508",
  1126 => x"318c08ec",
  1127 => x"050c8c08",
  1128 => x"ec050880",
  1129 => x"249d3880",
  1130 => x"0b8c08f4",
  1131 => x"050c8c08",
  1132 => x"ec050830",
  1133 => x"8c08fc05",
  1134 => x"08712b8c",
  1135 => x"08f0050c",
  1136 => x"54b9398c",
  1137 => x"08fc0508",
  1138 => x"8c08ec05",
  1139 => x"082a8c08",
  1140 => x"e8050c8c",
  1141 => x"08fc0508",
  1142 => x"8c089405",
  1143 => x"082b8c08",
  1144 => x"f4050c8c",
  1145 => x"08f80508",
  1146 => x"8c089405",
  1147 => x"082b708c",
  1148 => x"08e80508",
  1149 => x"078c08f0",
  1150 => x"050c548c",
  1151 => x"08f00508",
  1152 => x"8c08f405",
  1153 => x"088c0888",
  1154 => x"05085856",
  1155 => x"5473760c",
  1156 => x"7484170c",
  1157 => x"8c088805",
  1158 => x"08800c8d",
  1159 => x"3d0d8c0c",
  1160 => x"048c0802",
  1161 => x"8c0cf43d",
  1162 => x"0d800b8c",
  1163 => x"08f0050c",
  1164 => x"800b8c08",
  1165 => x"f4050c8c",
  1166 => x"08880508",
  1167 => x"8c088c05",
  1168 => x"08565473",
  1169 => x"8c08f005",
  1170 => x"0c748c08",
  1171 => x"f4050c8c",
  1172 => x"08f8058c",
  1173 => x"08f00556",
  1174 => x"56887054",
  1175 => x"75537652",
  1176 => x"54b29d3f",
  1177 => x"800b8c08",
  1178 => x"e8050c80",
  1179 => x"0b8c08ec",
  1180 => x"050c8c08",
  1181 => x"9005088c",
  1182 => x"08940508",
  1183 => x"5654738c",
  1184 => x"08e8050c",
  1185 => x"748c08ec",
  1186 => x"050c8c08",
  1187 => x"f0058c08",
  1188 => x"e8055656",
  1189 => x"88705475",
  1190 => x"53765254",
  1191 => x"b1e23f8c",
  1192 => x"08f80508",
  1193 => x"8c08f005",
  1194 => x"08258b38",
  1195 => x"800b8c08",
  1196 => x"e4050c80",
  1197 => x"ca398c08",
  1198 => x"f005088c",
  1199 => x"08f80508",
  1200 => x"258a3882",
  1201 => x"0b8c08e4",
  1202 => x"050cb439",
  1203 => x"8c08fc05",
  1204 => x"088c08f4",
  1205 => x"0508278a",
  1206 => x"38800b8c",
  1207 => x"08e4050c",
  1208 => x"9e398c08",
  1209 => x"f405088c",
  1210 => x"08fc0508",
  1211 => x"278a3882",
  1212 => x"0b8c08e4",
  1213 => x"050c8839",
  1214 => x"810b8c08",
  1215 => x"e4050c8c",
  1216 => x"08e40508",
  1217 => x"800c8e3d",
  1218 => x"0d8c0c04",
  1219 => x"8c08028c",
  1220 => x"0cffbc3d",
  1221 => x"0d8c088c",
  1222 => x"05088c08",
  1223 => x"90050855",
  1224 => x"53728c08",
  1225 => x"cc050c73",
  1226 => x"8c08d005",
  1227 => x"0c8c0894",
  1228 => x"05088c08",
  1229 => x"98050855",
  1230 => x"53728c08",
  1231 => x"c4050c73",
  1232 => x"8c08c805",
  1233 => x"0c8c08ec",
  1234 => x"0570538c",
  1235 => x"08cc0570",
  1236 => x"535153ac",
  1237 => x"cd3f8c08",
  1238 => x"d8057053",
  1239 => x"8c08c405",
  1240 => x"70535153",
  1241 => x"acbc3f8c",
  1242 => x"08ec058c",
  1243 => x"08c0050c",
  1244 => x"8c08d805",
  1245 => x"8c08ffbc",
  1246 => x"050c8c08",
  1247 => x"c0050851",
  1248 => x"8efa3f80",
  1249 => x"08537280",
  1250 => x"2e8f388c",
  1251 => x"08c00508",
  1252 => x"8c08ffb8",
  1253 => x"050c8dbd",
  1254 => x"398c08ff",
  1255 => x"bc050851",
  1256 => x"8eda3f80",
  1257 => x"08537280",
  1258 => x"2e90388c",
  1259 => x"08ffbc05",
  1260 => x"088c08ff",
  1261 => x"b8050c8d",
  1262 => x"9c398c08",
  1263 => x"c005088c",
  1264 => x"08c00508",
  1265 => x"8c08ffbc",
  1266 => x"05088412",
  1267 => x"08841208",
  1268 => x"3284140c",
  1269 => x"8c08c005",
  1270 => x"08545555",
  1271 => x"558de93f",
  1272 => x"80085372",
  1273 => x"92388c08",
  1274 => x"c0050851",
  1275 => x"8da63f80",
  1276 => x"08537283",
  1277 => x"38b6398c",
  1278 => x"08c00508",
  1279 => x"8c08ffbc",
  1280 => x"05085454",
  1281 => x"73087308",
  1282 => x"2e098106",
  1283 => x"91388cef",
  1284 => x"3f800870",
  1285 => x"8c08ffb8",
  1286 => x"050c538c",
  1287 => x"b8398c08",
  1288 => x"c005088c",
  1289 => x"08ffb805",
  1290 => x"0c8caa39",
  1291 => x"8c08ffbc",
  1292 => x"0508518d",
  1293 => x"933f8008",
  1294 => x"5372802e",
  1295 => x"ac388c08",
  1296 => x"c0050853",
  1297 => x"80548055",
  1298 => x"738c140c",
  1299 => x"7490140c",
  1300 => x"8c08c005",
  1301 => x"0853800b",
  1302 => x"88140c8c",
  1303 => x"08c00508",
  1304 => x"8c08ffb8",
  1305 => x"050c8bed",
  1306 => x"398c08ff",
  1307 => x"bc050851",
  1308 => x"8ca23f80",
  1309 => x"08537280",
  1310 => x"2e98388c",
  1311 => x"08c00508",
  1312 => x"5384730c",
  1313 => x"8c08c005",
  1314 => x"088c08ff",
  1315 => x"b8050c8b",
  1316 => x"c4398c08",
  1317 => x"c005088c",
  1318 => x"08c00508",
  1319 => x"8c08ffbc",
  1320 => x"05088812",
  1321 => x"08881208",
  1322 => x"3188140c",
  1323 => x"8c08c005",
  1324 => x"08515555",
  1325 => x"55901308",
  1326 => x"8c140854",
  1327 => x"54728c08",
  1328 => x"ffa8050c",
  1329 => x"738c08ff",
  1330 => x"ac050c8c",
  1331 => x"08ffbc05",
  1332 => x"08539013",
  1333 => x"088c1408",
  1334 => x"5454728c",
  1335 => x"08ffa005",
  1336 => x"0c738c08",
  1337 => x"ffa4050c",
  1338 => x"8c08ffa0",
  1339 => x"05088c08",
  1340 => x"ffa80508",
  1341 => x"26a6388c",
  1342 => x"08ffa005",
  1343 => x"088c08ff",
  1344 => x"a805082e",
  1345 => x"09810681",
  1346 => x"de388c08",
  1347 => x"ffa40508",
  1348 => x"8c08ffac",
  1349 => x"05082684",
  1350 => x"3881cc39",
  1351 => x"8c08ffa8",
  1352 => x"05088c08",
  1353 => x"ffac0508",
  1354 => x"5553728c",
  1355 => x"08ff9005",
  1356 => x"0c738c08",
  1357 => x"ff94050c",
  1358 => x"8c08ff90",
  1359 => x"05088c08",
  1360 => x"ff940508",
  1361 => x"5553728c",
  1362 => x"08ff8805",
  1363 => x"0c738c08",
  1364 => x"ff8c050c",
  1365 => x"8c08ff8c",
  1366 => x"05088c08",
  1367 => x"ff940508",
  1368 => x"7012708c",
  1369 => x"08ff8405",
  1370 => x"0c525454",
  1371 => x"810b8c08",
  1372 => x"fefc050c",
  1373 => x"8c08ff84",
  1374 => x"05088c08",
  1375 => x"ff8c0508",
  1376 => x"54547274",
  1377 => x"26893880",
  1378 => x"0b8c08fe",
  1379 => x"fc050c8c",
  1380 => x"08ff8805",
  1381 => x"088c08ff",
  1382 => x"90050870",
  1383 => x"12708c08",
  1384 => x"ff80050c",
  1385 => x"8c08ff80",
  1386 => x"05088c08",
  1387 => x"fefc0508",
  1388 => x"11708c08",
  1389 => x"ff80050c",
  1390 => x"53515254",
  1391 => x"548c08ff",
  1392 => x"8005088c",
  1393 => x"08ff8405",
  1394 => x"08555372",
  1395 => x"8c08ffa8",
  1396 => x"050c738c",
  1397 => x"08ffac05",
  1398 => x"0c8c08c0",
  1399 => x"05088811",
  1400 => x"08ff0588",
  1401 => x"120c5388",
  1402 => x"0a538054",
  1403 => x"728c08ff",
  1404 => x"b0050c73",
  1405 => x"8c08ffb4",
  1406 => x"050c8053",
  1407 => x"8054728c",
  1408 => x"08ff9805",
  1409 => x"0c738c08",
  1410 => x"ff9c050c",
  1411 => x"8c08ffb0",
  1412 => x"0508708c",
  1413 => x"08ffb405",
  1414 => x"08075153",
  1415 => x"72802e84",
  1416 => x"8a388c08",
  1417 => x"ffa00508",
  1418 => x"8c08ffa8",
  1419 => x"05082682",
  1420 => x"8d388c08",
  1421 => x"ffa00508",
  1422 => x"8c08ffa8",
  1423 => x"05082e09",
  1424 => x"81069138",
  1425 => x"8c08ffa4",
  1426 => x"05088c08",
  1427 => x"ffac0508",
  1428 => x"2681eb38",
  1429 => x"8c08ff98",
  1430 => x"05088c08",
  1431 => x"ffb00508",
  1432 => x"078c08ff",
  1433 => x"9c05088c",
  1434 => x"08ffb405",
  1435 => x"08075553",
  1436 => x"728c08ff",
  1437 => x"98050c73",
  1438 => x"8c08ff9c",
  1439 => x"050c8c08",
  1440 => x"ffa80508",
  1441 => x"8c08ffac",
  1442 => x"05085553",
  1443 => x"728c08fe",
  1444 => x"f4050c73",
  1445 => x"8c08fef8",
  1446 => x"050c8c08",
  1447 => x"ffa00508",
  1448 => x"8c08ffa4",
  1449 => x"05085553",
  1450 => x"728c08fe",
  1451 => x"ec050c73",
  1452 => x"8c08fef0",
  1453 => x"050c8c08",
  1454 => x"fef80508",
  1455 => x"8c08fef0",
  1456 => x"05087171",
  1457 => x"31708c08",
  1458 => x"fee8050c",
  1459 => x"52545481",
  1460 => x"0b8c08fe",
  1461 => x"e0050c8c",
  1462 => x"08fee805",
  1463 => x"088c08fe",
  1464 => x"f8050854",
  1465 => x"54737326",
  1466 => x"8938800b",
  1467 => x"8c08fee0",
  1468 => x"050c8c08",
  1469 => x"fef40508",
  1470 => x"8c08feec",
  1471 => x"05087171",
  1472 => x"31708c08",
  1473 => x"fee4050c",
  1474 => x"8c08fee4",
  1475 => x"0508708c",
  1476 => x"08fee005",
  1477 => x"0831708c",
  1478 => x"08fee405",
  1479 => x"0c535152",
  1480 => x"54548c08",
  1481 => x"fee40508",
  1482 => x"8c08fee8",
  1483 => x"05085553",
  1484 => x"728c08ff",
  1485 => x"a8050c73",
  1486 => x"8c08ffac",
  1487 => x"050c8c08",
  1488 => x"ffb00508",
  1489 => x"9f2b8c08",
  1490 => x"ffb40508",
  1491 => x"812a7072",
  1492 => x"078c08ff",
  1493 => x"b0050881",
  1494 => x"2a565656",
  1495 => x"56728c08",
  1496 => x"ffb0050c",
  1497 => x"738c08ff",
  1498 => x"b4050c8c",
  1499 => x"08ffa805",
  1500 => x"088c08ff",
  1501 => x"ac050855",
  1502 => x"53728c08",
  1503 => x"fed8050c",
  1504 => x"738c08fe",
  1505 => x"dc050c8c",
  1506 => x"08fed805",
  1507 => x"088c08fe",
  1508 => x"dc050855",
  1509 => x"53728c08",
  1510 => x"fed0050c",
  1511 => x"738c08fe",
  1512 => x"d4050c8c",
  1513 => x"08fed405",
  1514 => x"088c08fe",
  1515 => x"dc050870",
  1516 => x"12708c08",
  1517 => x"fecc050c",
  1518 => x"52545481",
  1519 => x"0b8c08fe",
  1520 => x"c4050c8c",
  1521 => x"08fecc05",
  1522 => x"088c08fe",
  1523 => x"d4050854",
  1524 => x"54727426",
  1525 => x"8938800b",
  1526 => x"8c08fec4",
  1527 => x"050c8c08",
  1528 => x"fed00508",
  1529 => x"8c08fed8",
  1530 => x"05087012",
  1531 => x"708c08fe",
  1532 => x"c8050c8c",
  1533 => x"08fec805",
  1534 => x"088c08fe",
  1535 => x"c4050811",
  1536 => x"708c08fe",
  1537 => x"c8050c53",
  1538 => x"51525454",
  1539 => x"8c08fec8",
  1540 => x"05088c08",
  1541 => x"fecc0508",
  1542 => x"5553728c",
  1543 => x"08ffa805",
  1544 => x"0c738c08",
  1545 => x"ffac050c",
  1546 => x"fbe2398c",
  1547 => x"08ff9805",
  1548 => x"08800670",
  1549 => x"8c08febc",
  1550 => x"050c8c08",
  1551 => x"ff9c0508",
  1552 => x"81ff0670",
  1553 => x"8c08fec0",
  1554 => x"050c5454",
  1555 => x"8c08febc",
  1556 => x"05088c08",
  1557 => x"fec00508",
  1558 => x"5553728c",
  1559 => x"08febc05",
  1560 => x"0c738c08",
  1561 => x"fec0050c",
  1562 => x"8c08febc",
  1563 => x"05085473",
  1564 => x"83bc388c",
  1565 => x"08fec005",
  1566 => x"08537281",
  1567 => x"802e0981",
  1568 => x"0683ab38",
  1569 => x"8c08ff98",
  1570 => x"0508982b",
  1571 => x"8c08ff9c",
  1572 => x"0508882a",
  1573 => x"7072078c",
  1574 => x"08ff9805",
  1575 => x"08882a71",
  1576 => x"81065156",
  1577 => x"56565672",
  1578 => x"802e81b8",
  1579 => x"388c08ff",
  1580 => x"9805088c",
  1581 => x"08ff9c05",
  1582 => x"08555372",
  1583 => x"8c08feb4",
  1584 => x"050c738c",
  1585 => x"08feb805",
  1586 => x"0c805381",
  1587 => x"8054728c",
  1588 => x"08feac05",
  1589 => x"0c738c08",
  1590 => x"feb0050c",
  1591 => x"8c08feb8",
  1592 => x"05088c08",
  1593 => x"feb00508",
  1594 => x"7012708c",
  1595 => x"08fea805",
  1596 => x"0c525454",
  1597 => x"810b8c08",
  1598 => x"fea0050c",
  1599 => x"8c08fea8",
  1600 => x"05088c08",
  1601 => x"feb80508",
  1602 => x"54547274",
  1603 => x"26893880",
  1604 => x"0b8c08fe",
  1605 => x"a0050c8c",
  1606 => x"08feb405",
  1607 => x"088c08fe",
  1608 => x"ac050870",
  1609 => x"12708c08",
  1610 => x"fea4050c",
  1611 => x"8c08fea4",
  1612 => x"05088c08",
  1613 => x"fea00508",
  1614 => x"11708c08",
  1615 => x"fea4050c",
  1616 => x"53515254",
  1617 => x"548c08fe",
  1618 => x"a405088c",
  1619 => x"08fea805",
  1620 => x"08555372",
  1621 => x"8c08ff98",
  1622 => x"050c738c",
  1623 => x"08ff9c05",
  1624 => x"0c81cb39",
  1625 => x"8c08ffa8",
  1626 => x"0508708c",
  1627 => x"08ffac05",
  1628 => x"08075153",
  1629 => x"72802e81",
  1630 => x"b5388c08",
  1631 => x"ff980508",
  1632 => x"8c08ff9c",
  1633 => x"05085553",
  1634 => x"728c08fe",
  1635 => x"98050c73",
  1636 => x"8c08fe9c",
  1637 => x"050c8053",
  1638 => x"81805472",
  1639 => x"8c08fe90",
  1640 => x"050c738c",
  1641 => x"08fe9405",
  1642 => x"0c8c08fe",
  1643 => x"9c05088c",
  1644 => x"08fe9405",
  1645 => x"08701270",
  1646 => x"8c08fe8c",
  1647 => x"050c5254",
  1648 => x"54810b8c",
  1649 => x"08fe8405",
  1650 => x"0c8c08fe",
  1651 => x"8c05088c",
  1652 => x"08fe9c05",
  1653 => x"08545472",
  1654 => x"74268938",
  1655 => x"800b8c08",
  1656 => x"fe84050c",
  1657 => x"8c08fe98",
  1658 => x"05088c08",
  1659 => x"fe900508",
  1660 => x"7012708c",
  1661 => x"08fe8805",
  1662 => x"0c8c08fe",
  1663 => x"8805088c",
  1664 => x"08fe8405",
  1665 => x"0811708c",
  1666 => x"08fe8805",
  1667 => x"0c535152",
  1668 => x"54548c08",
  1669 => x"fe880508",
  1670 => x"8c08fe8c",
  1671 => x"05085553",
  1672 => x"728c08ff",
  1673 => x"98050c73",
  1674 => x"8c08ff9c",
  1675 => x"050c8c08",
  1676 => x"c0050855",
  1677 => x"8c08ff98",
  1678 => x"05088c08",
  1679 => x"ff9c0508",
  1680 => x"5553728c",
  1681 => x"160c7390",
  1682 => x"160c8c08",
  1683 => x"c005088c",
  1684 => x"08ffb805",
  1685 => x"0c8c08ff",
  1686 => x"b8050870",
  1687 => x"8c08d405",
  1688 => x"0c8c08d4",
  1689 => x"0508538c",
  1690 => x"08880508",
  1691 => x"52538dfd",
  1692 => x"3f8c0888",
  1693 => x"0508800c",
  1694 => x"80c63d0d",
  1695 => x"8c0c048c",
  1696 => x"08028c0c",
  1697 => x"803d0d80",
  1698 => x"dd907080",
  1699 => x"0c51823d",
  1700 => x"0d8c0c04",
  1701 => x"8c08028c",
  1702 => x"0cff3d0d",
  1703 => x"800b8c08",
  1704 => x"fc050c8c",
  1705 => x"08880508",
  1706 => x"51700882",
  1707 => x"2e098106",
  1708 => x"8838810b",
  1709 => x"8c08fc05",
  1710 => x"0c8c08fc",
  1711 => x"05087080",
  1712 => x"0c51833d",
  1713 => x"0d8c0c04",
  1714 => x"8c08028c",
  1715 => x"0cff3d0d",
  1716 => x"800b8c08",
  1717 => x"fc050c8c",
  1718 => x"08880508",
  1719 => x"51700884",
  1720 => x"2e098106",
  1721 => x"8838810b",
  1722 => x"8c08fc05",
  1723 => x"0c8c08fc",
  1724 => x"05087080",
  1725 => x"0c51833d",
  1726 => x"0d8c0c04",
  1727 => x"8c08028c",
  1728 => x"0cff3d0d",
  1729 => x"800b8c08",
  1730 => x"fc050c8c",
  1731 => x"08880508",
  1732 => x"51700880",
  1733 => x"2e8f388c",
  1734 => x"08880508",
  1735 => x"51700881",
  1736 => x"2e833888",
  1737 => x"39810b8c",
  1738 => x"08fc050c",
  1739 => x"8c08fc05",
  1740 => x"0870800c",
  1741 => x"51833d0d",
  1742 => x"8c0c048c",
  1743 => x"08028c0c",
  1744 => x"f63d0d83",
  1745 => x"0b8c08ec",
  1746 => x"050c800b",
  1747 => x"8c08e805",
  1748 => x"0c8c088c",
  1749 => x"05088025",
  1750 => x"8838810b",
  1751 => x"8c08e805",
  1752 => x"0c8c08e8",
  1753 => x"05088c08",
  1754 => x"f0050c8c",
  1755 => x"088c0508",
  1756 => x"8b38820b",
  1757 => x"8c08ec05",
  1758 => x"0c819e39",
  1759 => x"bc0b8c08",
  1760 => x"f4050c8c",
  1761 => x"08f00508",
  1762 => x"802ebe38",
  1763 => x"8c088c05",
  1764 => x"08810a2e",
  1765 => x"09810698",
  1766 => x"388f830a",
  1767 => x"53800b8c",
  1768 => x"08880508",
  1769 => x"56547275",
  1770 => x"0c738416",
  1771 => x"0c80fa39",
  1772 => x"8c088c05",
  1773 => x"0830708c",
  1774 => x"08fc050c",
  1775 => x"709f2c70",
  1776 => x"8c08f805",
  1777 => x"0c515397",
  1778 => x"398c088c",
  1779 => x"0508708c",
  1780 => x"08fc050c",
  1781 => x"709f2c70",
  1782 => x"8c08f805",
  1783 => x"0c51538c",
  1784 => x"08f80508",
  1785 => x"f00a26b1",
  1786 => x"388c08fc",
  1787 => x"05089f2a",
  1788 => x"8c08f805",
  1789 => x"08107072",
  1790 => x"078c08f8",
  1791 => x"050c8c08",
  1792 => x"fc050810",
  1793 => x"8c08fc05",
  1794 => x"0c8c08f4",
  1795 => x"0508ff05",
  1796 => x"8c08f405",
  1797 => x"0c5454c7",
  1798 => x"398c08ec",
  1799 => x"0570538c",
  1800 => x"08880508",
  1801 => x"52538ac5",
  1802 => x"3f8c0888",
  1803 => x"0508800c",
  1804 => x"8c3d0d8c",
  1805 => x"0c048c08",
  1806 => x"028c0cec",
  1807 => x"3d0d8c08",
  1808 => x"8805088c",
  1809 => x"088c0508",
  1810 => x"5755748c",
  1811 => x"08e0050c",
  1812 => x"758c08e4",
  1813 => x"050c8c08",
  1814 => x"ec057053",
  1815 => x"8c08e005",
  1816 => x"70535155",
  1817 => x"9abc3f8c",
  1818 => x"08ec0570",
  1819 => x"5255838d",
  1820 => x"3f800855",
  1821 => x"74802e8b",
  1822 => x"38800b8c",
  1823 => x"08d4050c",
  1824 => x"81fb398c",
  1825 => x"08ec0570",
  1826 => x"525582b2",
  1827 => x"3f800855",
  1828 => x"74802e8b",
  1829 => x"38800b8c",
  1830 => x"08d4050c",
  1831 => x"81df398c",
  1832 => x"08ec0570",
  1833 => x"525581e2",
  1834 => x"3f800855",
  1835 => x"74802ea9",
  1836 => x"388c08f0",
  1837 => x"0508802e",
  1838 => x"8b38810a",
  1839 => x"0b8c08d0",
  1840 => x"050c8939",
  1841 => x"fe0a0b8c",
  1842 => x"08d0050c",
  1843 => x"8c08d005",
  1844 => x"088c08d4",
  1845 => x"050c81a5",
  1846 => x"398c08f4",
  1847 => x"05088025",
  1848 => x"8b38800b",
  1849 => x"8c08d405",
  1850 => x"0c819239",
  1851 => x"9e0b8c08",
  1852 => x"f4050825",
  1853 => x"a9388c08",
  1854 => x"f0050880",
  1855 => x"2e8b3881",
  1856 => x"0a0b8c08",
  1857 => x"cc050c89",
  1858 => x"39fe0a0b",
  1859 => x"8c08cc05",
  1860 => x"0c8c08cc",
  1861 => x"05088c08",
  1862 => x"d4050c80",
  1863 => x"e039bc0b",
  1864 => x"8c08f405",
  1865 => x"08318c08",
  1866 => x"d8057156",
  1867 => x"58558c08",
  1868 => x"f805088c",
  1869 => x"08fc0508",
  1870 => x"57557452",
  1871 => x"75537651",
  1872 => x"86b53f8c",
  1873 => x"08d80508",
  1874 => x"8c08dc05",
  1875 => x"08708c08",
  1876 => x"e8050c8c",
  1877 => x"08e80508",
  1878 => x"8c08c805",
  1879 => x"0c57558c",
  1880 => x"08f00508",
  1881 => x"802e8c38",
  1882 => x"8c08c805",
  1883 => x"08308c08",
  1884 => x"c8050c8c",
  1885 => x"08c80508",
  1886 => x"8c08d405",
  1887 => x"0c8c08d4",
  1888 => x"0508800c",
  1889 => x"963d0d8c",
  1890 => x"0c048c08",
  1891 => x"028c0cff",
  1892 => x"3d0d800b",
  1893 => x"8c08fc05",
  1894 => x"0c8c0888",
  1895 => x"05085170",
  1896 => x"08842e09",
  1897 => x"81068838",
  1898 => x"810b8c08",
  1899 => x"fc050c8c",
  1900 => x"08fc0508",
  1901 => x"70800c51",
  1902 => x"833d0d8c",
  1903 => x"0c048c08",
  1904 => x"028c0cff",
  1905 => x"3d0d800b",
  1906 => x"8c08fc05",
  1907 => x"0c8c0888",
  1908 => x"05085170",
  1909 => x"08802e8f",
  1910 => x"388c0888",
  1911 => x"05085170",
  1912 => x"08812e83",
  1913 => x"38883981",
  1914 => x"0b8c08fc",
  1915 => x"050c8c08",
  1916 => x"fc050870",
  1917 => x"800c5183",
  1918 => x"3d0d8c0c",
  1919 => x"048c0802",
  1920 => x"8c0cff3d",
  1921 => x"0d800b8c",
  1922 => x"08fc050c",
  1923 => x"8c088805",
  1924 => x"08517008",
  1925 => x"822e0981",
  1926 => x"06883881",
  1927 => x"0b8c08fc",
  1928 => x"050c8c08",
  1929 => x"fc050870",
  1930 => x"800c5183",
  1931 => x"3d0d8c0c",
  1932 => x"048c0802",
  1933 => x"8c0cfd3d",
  1934 => x"0d80538c",
  1935 => x"088c0508",
  1936 => x"528c0888",
  1937 => x"05085182",
  1938 => x"de3f8008",
  1939 => x"70800c54",
  1940 => x"853d0d8c",
  1941 => x"0c048c08",
  1942 => x"028c0cfd",
  1943 => x"3d0d8153",
  1944 => x"8c088c05",
  1945 => x"08528c08",
  1946 => x"88050851",
  1947 => x"82b93f80",
  1948 => x"0870800c",
  1949 => x"54853d0d",
  1950 => x"8c0c048c",
  1951 => x"08028c0c",
  1952 => x"f93d0d80",
  1953 => x"0b8c08fc",
  1954 => x"050c8c08",
  1955 => x"88050880",
  1956 => x"25ab388c",
  1957 => x"08880508",
  1958 => x"308c0888",
  1959 => x"050c800b",
  1960 => x"8c08f405",
  1961 => x"0c8c08fc",
  1962 => x"05088838",
  1963 => x"810b8c08",
  1964 => x"f4050c8c",
  1965 => x"08f40508",
  1966 => x"8c08fc05",
  1967 => x"0c8c088c",
  1968 => x"05088025",
  1969 => x"ab388c08",
  1970 => x"8c050830",
  1971 => x"8c088c05",
  1972 => x"0c800b8c",
  1973 => x"08f0050c",
  1974 => x"8c08fc05",
  1975 => x"08883881",
  1976 => x"0b8c08f0",
  1977 => x"050c8c08",
  1978 => x"f005088c",
  1979 => x"08fc050c",
  1980 => x"80538c08",
  1981 => x"8c050852",
  1982 => x"8c088805",
  1983 => x"085181a7",
  1984 => x"3f800870",
  1985 => x"8c08f805",
  1986 => x"0c548c08",
  1987 => x"fc050880",
  1988 => x"2e8c388c",
  1989 => x"08f80508",
  1990 => x"308c08f8",
  1991 => x"050c8c08",
  1992 => x"f8050870",
  1993 => x"800c5489",
  1994 => x"3d0d8c0c",
  1995 => x"048c0802",
  1996 => x"8c0cfb3d",
  1997 => x"0d800b8c",
  1998 => x"08fc050c",
  1999 => x"8c088805",
  2000 => x"08802593",
  2001 => x"388c0888",
  2002 => x"0508308c",
  2003 => x"0888050c",
  2004 => x"810b8c08",
  2005 => x"fc050c8c",
  2006 => x"088c0508",
  2007 => x"80258c38",
  2008 => x"8c088c05",
  2009 => x"08308c08",
  2010 => x"8c050c81",
  2011 => x"538c088c",
  2012 => x"0508528c",
  2013 => x"08880508",
  2014 => x"51ad3f80",
  2015 => x"08708c08",
  2016 => x"f8050c54",
  2017 => x"8c08fc05",
  2018 => x"08802e8c",
  2019 => x"388c08f8",
  2020 => x"0508308c",
  2021 => x"08f8050c",
  2022 => x"8c08f805",
  2023 => x"0870800c",
  2024 => x"54873d0d",
  2025 => x"8c0c048c",
  2026 => x"08028c0c",
  2027 => x"fd3d0d81",
  2028 => x"0b8c08fc",
  2029 => x"050c800b",
  2030 => x"8c08f805",
  2031 => x"0c8c088c",
  2032 => x"05088c08",
  2033 => x"88050827",
  2034 => x"ac388c08",
  2035 => x"fc050880",
  2036 => x"2ea33880",
  2037 => x"0b8c088c",
  2038 => x"05082499",
  2039 => x"388c088c",
  2040 => x"0508108c",
  2041 => x"088c050c",
  2042 => x"8c08fc05",
  2043 => x"08108c08",
  2044 => x"fc050cc9",
  2045 => x"398c08fc",
  2046 => x"0508802e",
  2047 => x"80c9388c",
  2048 => x"088c0508",
  2049 => x"8c088805",
  2050 => x"0826a138",
  2051 => x"8c088805",
  2052 => x"088c088c",
  2053 => x"0508318c",
  2054 => x"0888050c",
  2055 => x"8c08f805",
  2056 => x"088c08fc",
  2057 => x"0508078c",
  2058 => x"08f8050c",
  2059 => x"8c08fc05",
  2060 => x"08812a8c",
  2061 => x"08fc050c",
  2062 => x"8c088c05",
  2063 => x"08812a8c",
  2064 => x"088c050c",
  2065 => x"ffaf398c",
  2066 => x"08900508",
  2067 => x"802e8f38",
  2068 => x"8c088805",
  2069 => x"08708c08",
  2070 => x"f4050c51",
  2071 => x"8d398c08",
  2072 => x"f8050870",
  2073 => x"8c08f405",
  2074 => x"0c518c08",
  2075 => x"f4050880",
  2076 => x"0c853d0d",
  2077 => x"8c0c048c",
  2078 => x"08028c0c",
  2079 => x"f53d0d8c",
  2080 => x"08940508",
  2081 => x"9d388c08",
  2082 => x"8c05088c",
  2083 => x"08900508",
  2084 => x"8c088805",
  2085 => x"08585654",
  2086 => x"73760c74",
  2087 => x"84170c81",
  2088 => x"bf39800b",
  2089 => x"8c08f005",
  2090 => x"0c800b8c",
  2091 => x"08f4050c",
  2092 => x"8c088c05",
  2093 => x"088c0890",
  2094 => x"05085654",
  2095 => x"738c08f0",
  2096 => x"050c748c",
  2097 => x"08f4050c",
  2098 => x"8c08f805",
  2099 => x"8c08f005",
  2100 => x"56568870",
  2101 => x"54755376",
  2102 => x"525495a4",
  2103 => x"3fa00b8c",
  2104 => x"08940508",
  2105 => x"318c08ec",
  2106 => x"050c8c08",
  2107 => x"ec050880",
  2108 => x"249d3880",
  2109 => x"0b8c08f0",
  2110 => x"050c8c08",
  2111 => x"ec050830",
  2112 => x"8c08f805",
  2113 => x"08712a8c",
  2114 => x"08f4050c",
  2115 => x"54b9398c",
  2116 => x"08f80508",
  2117 => x"8c08ec05",
  2118 => x"082b8c08",
  2119 => x"e8050c8c",
  2120 => x"08f80508",
  2121 => x"8c089405",
  2122 => x"082a8c08",
  2123 => x"f0050c8c",
  2124 => x"08fc0508",
  2125 => x"8c089405",
  2126 => x"082a708c",
  2127 => x"08e80508",
  2128 => x"078c08f4",
  2129 => x"050c548c",
  2130 => x"08f00508",
  2131 => x"8c08f405",
  2132 => x"088c0888",
  2133 => x"05085856",
  2134 => x"5473760c",
  2135 => x"7484170c",
  2136 => x"8c088805",
  2137 => x"08800c8d",
  2138 => x"3d0d8c0c",
  2139 => x"048c0802",
  2140 => x"8c0cc73d",
  2141 => x"0d8c088c",
  2142 => x"05085590",
  2143 => x"15088c16",
  2144 => x"08565674",
  2145 => x"8c08f005",
  2146 => x"0c758c08",
  2147 => x"f4050c8c",
  2148 => x"088c0508",
  2149 => x"8411088c",
  2150 => x"08ec050c",
  2151 => x"55800b8c",
  2152 => x"08e8050c",
  2153 => x"8c088c05",
  2154 => x"08518fb7",
  2155 => x"3f800855",
  2156 => x"74802eaa",
  2157 => x"388fff0b",
  2158 => x"8c08e805",
  2159 => x"0c8c08f0",
  2160 => x"0508a080",
  2161 => x"80078c08",
  2162 => x"f4050880",
  2163 => x"07575574",
  2164 => x"8c08f005",
  2165 => x"0c758c08",
  2166 => x"f4050c8c",
  2167 => x"ff398c08",
  2168 => x"8c050851",
  2169 => x"8ec93f80",
  2170 => x"08557480",
  2171 => x"2e9c388f",
  2172 => x"ff0b8c08",
  2173 => x"e8050c80",
  2174 => x"55805674",
  2175 => x"8c08f005",
  2176 => x"0c758c08",
  2177 => x"f4050c8c",
  2178 => x"d3398c08",
  2179 => x"8c050851",
  2180 => x"8de93f80",
  2181 => x"08557480",
  2182 => x"2e9b3880",
  2183 => x"0b8c08e8",
  2184 => x"050c8055",
  2185 => x"8056748c",
  2186 => x"08f0050c",
  2187 => x"758c08f4",
  2188 => x"050c8ca8",
  2189 => x"398c08f0",
  2190 => x"0508708c",
  2191 => x"08f40508",
  2192 => x"07515574",
  2193 => x"8b38800b",
  2194 => x"8c08e805",
  2195 => x"0c8c8d39",
  2196 => x"8c088c05",
  2197 => x"08558815",
  2198 => x"08f88225",
  2199 => x"86fb388c",
  2200 => x"088c0508",
  2201 => x"f8820b88",
  2202 => x"1208318c",
  2203 => x"08e4050c",
  2204 => x"55800b8c",
  2205 => x"08e8050c",
  2206 => x"b80b8c08",
  2207 => x"e4050825",
  2208 => x"94388055",
  2209 => x"8056748c",
  2210 => x"08f0050c",
  2211 => x"758c08f4",
  2212 => x"050c82a2",
  2213 => x"39800b8c",
  2214 => x"08e0050c",
  2215 => x"8c08d805",
  2216 => x"57805581",
  2217 => x"0b8c08e4",
  2218 => x"05085556",
  2219 => x"74527553",
  2220 => x"7651dcf7",
  2221 => x"3f8c08d8",
  2222 => x"05088c08",
  2223 => x"dc050857",
  2224 => x"55748c08",
  2225 => x"d0050c75",
  2226 => x"8c08d405",
  2227 => x"0cff56ff",
  2228 => x"57758c08",
  2229 => x"c8050c76",
  2230 => x"8c08cc05",
  2231 => x"0c8c08d4",
  2232 => x"05088c08",
  2233 => x"cc050870",
  2234 => x"12708c08",
  2235 => x"c4050c52",
  2236 => x"5657810b",
  2237 => x"8c08ffbc",
  2238 => x"050c8c08",
  2239 => x"c405088c",
  2240 => x"08d40508",
  2241 => x"58567676",
  2242 => x"26893880",
  2243 => x"0b8c08ff",
  2244 => x"bc050c8c",
  2245 => x"08d00508",
  2246 => x"8c08c805",
  2247 => x"08701270",
  2248 => x"8c08c005",
  2249 => x"0c8c08c0",
  2250 => x"05088c08",
  2251 => x"ffbc0508",
  2252 => x"11708c08",
  2253 => x"c0050c8c",
  2254 => x"08c00508",
  2255 => x"708c08f0",
  2256 => x"0508068c",
  2257 => x"08c40508",
  2258 => x"708c08f4",
  2259 => x"05080672",
  2260 => x"70720751",
  2261 => x"52575252",
  2262 => x"52525a52",
  2263 => x"57557680",
  2264 => x"2e883881",
  2265 => x"0b8c08e0",
  2266 => x"050c8c08",
  2267 => x"d8058c08",
  2268 => x"e4050855",
  2269 => x"578c08f0",
  2270 => x"05088c08",
  2271 => x"f4050857",
  2272 => x"55745275",
  2273 => x"537651f9",
  2274 => x"ee3f8c08",
  2275 => x"d805088c",
  2276 => x"08dc0508",
  2277 => x"8c08e005",
  2278 => x"089f2c8c",
  2279 => x"08e00508",
  2280 => x"71707507",
  2281 => x"8c08f005",
  2282 => x"0c737207",
  2283 => x"8c08f405",
  2284 => x"0c59595b",
  2285 => x"59578c08",
  2286 => x"f0050880",
  2287 => x"06708c08",
  2288 => x"ffb4050c",
  2289 => x"8c08f405",
  2290 => x"0881ff06",
  2291 => x"708c08ff",
  2292 => x"b8050c57",
  2293 => x"558c08ff",
  2294 => x"b405088c",
  2295 => x"08ffb805",
  2296 => x"08575574",
  2297 => x"8c08ffb4",
  2298 => x"050c758c",
  2299 => x"08ffb805",
  2300 => x"0c8c08ff",
  2301 => x"b4050856",
  2302 => x"7581eb38",
  2303 => x"8c08ffb8",
  2304 => x"05085776",
  2305 => x"81802e09",
  2306 => x"810681da",
  2307 => x"388c08f0",
  2308 => x"0508982b",
  2309 => x"8c08f405",
  2310 => x"08882a70",
  2311 => x"72078c08",
  2312 => x"f0050888",
  2313 => x"2a718106",
  2314 => x"51585858",
  2315 => x"5874802e",
  2316 => x"82e4388c",
  2317 => x"08f00508",
  2318 => x"8c08f405",
  2319 => x"08575574",
  2320 => x"8c08ffac",
  2321 => x"050c758c",
  2322 => x"08ffb005",
  2323 => x"0c805681",
  2324 => x"8057758c",
  2325 => x"08ffa405",
  2326 => x"0c768c08",
  2327 => x"ffa8050c",
  2328 => x"8c08ffb0",
  2329 => x"05088c08",
  2330 => x"ffa80508",
  2331 => x"7012708c",
  2332 => x"08ffa005",
  2333 => x"0c525657",
  2334 => x"810b8c08",
  2335 => x"ff98050c",
  2336 => x"8c08ffa0",
  2337 => x"05088c08",
  2338 => x"ffb00508",
  2339 => x"58567676",
  2340 => x"26893880",
  2341 => x"0b8c08ff",
  2342 => x"98050c8c",
  2343 => x"08ffac05",
  2344 => x"088c08ff",
  2345 => x"a4050870",
  2346 => x"12708c08",
  2347 => x"ff9c050c",
  2348 => x"8c08ff9c",
  2349 => x"05088c08",
  2350 => x"ff980508",
  2351 => x"11708c08",
  2352 => x"ff9c050c",
  2353 => x"525a5257",
  2354 => x"558c08ff",
  2355 => x"9c05088c",
  2356 => x"08ffa005",
  2357 => x"08575574",
  2358 => x"8c08f005",
  2359 => x"0c758c08",
  2360 => x"f4050c81",
  2361 => x"b1398c08",
  2362 => x"f005088c",
  2363 => x"08f40508",
  2364 => x"5856758c",
  2365 => x"08ff9005",
  2366 => x"0c768c08",
  2367 => x"ff94050c",
  2368 => x"805580ff",
  2369 => x"56748c08",
  2370 => x"ff88050c",
  2371 => x"758c08ff",
  2372 => x"8c050c8c",
  2373 => x"08ff9405",
  2374 => x"088c08ff",
  2375 => x"8c050870",
  2376 => x"12708c08",
  2377 => x"ff84050c",
  2378 => x"52585681",
  2379 => x"0b8c08fe",
  2380 => x"fc050c8c",
  2381 => x"08ff8405",
  2382 => x"088c08ff",
  2383 => x"94050857",
  2384 => x"55757526",
  2385 => x"8938800b",
  2386 => x"8c08fefc",
  2387 => x"050c8c08",
  2388 => x"ff900508",
  2389 => x"8c08ff88",
  2390 => x"05087012",
  2391 => x"708c08ff",
  2392 => x"80050c8c",
  2393 => x"08ff8005",
  2394 => x"088c08fe",
  2395 => x"fc050811",
  2396 => x"708c08ff",
  2397 => x"80050c53",
  2398 => x"59525657",
  2399 => x"8c08ff80",
  2400 => x"05088c08",
  2401 => x"ff840508",
  2402 => x"5755748c",
  2403 => x"08f0050c",
  2404 => x"758c08f4",
  2405 => x"050c8c08",
  2406 => x"f00508f0",
  2407 => x"0a268338",
  2408 => x"8d398c08",
  2409 => x"e8050881",
  2410 => x"058c08e8",
  2411 => x"050c8c08",
  2412 => x"f0050898",
  2413 => x"2b8c08f4",
  2414 => x"0508882a",
  2415 => x"7072078c",
  2416 => x"08f00508",
  2417 => x"882a5858",
  2418 => x"5858748c",
  2419 => x"08f0050c",
  2420 => x"758c08f4",
  2421 => x"050c8584",
  2422 => x"398c088c",
  2423 => x"05085587",
  2424 => x"ff0b8816",
  2425 => x"08259c38",
  2426 => x"8fff0b8c",
  2427 => x"08e8050c",
  2428 => x"80558056",
  2429 => x"748c08f0",
  2430 => x"050c758c",
  2431 => x"08f4050c",
  2432 => x"84da398c",
  2433 => x"088c0508",
  2434 => x"88110887",
  2435 => x"ff058c08",
  2436 => x"e8050c8c",
  2437 => x"08f00508",
  2438 => x"8006708c",
  2439 => x"08fef405",
  2440 => x"0c8c08f4",
  2441 => x"050881ff",
  2442 => x"06708c08",
  2443 => x"fef8050c",
  2444 => x"5957558c",
  2445 => x"08fef405",
  2446 => x"088c08fe",
  2447 => x"f8050857",
  2448 => x"55748c08",
  2449 => x"fef4050c",
  2450 => x"758c08fe",
  2451 => x"f8050c8c",
  2452 => x"08fef405",
  2453 => x"08567581",
  2454 => x"eb388c08",
  2455 => x"fef80508",
  2456 => x"57768180",
  2457 => x"2e098106",
  2458 => x"81da388c",
  2459 => x"08f00508",
  2460 => x"982b8c08",
  2461 => x"f4050888",
  2462 => x"2a707207",
  2463 => x"8c08f005",
  2464 => x"08882a71",
  2465 => x"81065158",
  2466 => x"58585874",
  2467 => x"802e82e4",
  2468 => x"388c08f0",
  2469 => x"05088c08",
  2470 => x"f4050857",
  2471 => x"55748c08",
  2472 => x"feec050c",
  2473 => x"758c08fe",
  2474 => x"f0050c80",
  2475 => x"56818057",
  2476 => x"758c08fe",
  2477 => x"e4050c76",
  2478 => x"8c08fee8",
  2479 => x"050c8c08",
  2480 => x"fef00508",
  2481 => x"8c08fee8",
  2482 => x"05087012",
  2483 => x"708c08fe",
  2484 => x"e0050c52",
  2485 => x"5657810b",
  2486 => x"8c08fed8",
  2487 => x"050c8c08",
  2488 => x"fee00508",
  2489 => x"8c08fef0",
  2490 => x"05085856",
  2491 => x"76762689",
  2492 => x"38800b8c",
  2493 => x"08fed805",
  2494 => x"0c8c08fe",
  2495 => x"ec05088c",
  2496 => x"08fee405",
  2497 => x"08701270",
  2498 => x"8c08fedc",
  2499 => x"050c8c08",
  2500 => x"fedc0508",
  2501 => x"8c08fed8",
  2502 => x"05081170",
  2503 => x"8c08fedc",
  2504 => x"050c525a",
  2505 => x"5257558c",
  2506 => x"08fedc05",
  2507 => x"088c08fe",
  2508 => x"e0050857",
  2509 => x"55748c08",
  2510 => x"f0050c75",
  2511 => x"8c08f405",
  2512 => x"0c81b139",
  2513 => x"8c08f005",
  2514 => x"088c08f4",
  2515 => x"05085856",
  2516 => x"758c08fe",
  2517 => x"d0050c76",
  2518 => x"8c08fed4",
  2519 => x"050c8055",
  2520 => x"80ff5674",
  2521 => x"8c08fec8",
  2522 => x"050c758c",
  2523 => x"08fecc05",
  2524 => x"0c8c08fe",
  2525 => x"d405088c",
  2526 => x"08fecc05",
  2527 => x"08701270",
  2528 => x"8c08fec4",
  2529 => x"050c5258",
  2530 => x"56810b8c",
  2531 => x"08febc05",
  2532 => x"0c8c08fe",
  2533 => x"c405088c",
  2534 => x"08fed405",
  2535 => x"08575575",
  2536 => x"75268938",
  2537 => x"800b8c08",
  2538 => x"febc050c",
  2539 => x"8c08fed0",
  2540 => x"05088c08",
  2541 => x"fec80508",
  2542 => x"7012708c",
  2543 => x"08fec005",
  2544 => x"0c8c08fe",
  2545 => x"c005088c",
  2546 => x"08febc05",
  2547 => x"0811708c",
  2548 => x"08fec005",
  2549 => x"0c535952",
  2550 => x"56578c08",
  2551 => x"fec00508",
  2552 => x"8c08fec4",
  2553 => x"05085755",
  2554 => x"748c08f0",
  2555 => x"050c758c",
  2556 => x"08f4050c",
  2557 => x"8c08f005",
  2558 => x"08f80a26",
  2559 => x"8338b539",
  2560 => x"8c08f005",
  2561 => x"089f2b8c",
  2562 => x"08f40508",
  2563 => x"812a7072",
  2564 => x"078c08f0",
  2565 => x"0508812a",
  2566 => x"58585858",
  2567 => x"748c08f0",
  2568 => x"050c758c",
  2569 => x"08f4050c",
  2570 => x"8c08e805",
  2571 => x"0881058c",
  2572 => x"08e8050c",
  2573 => x"8c08f005",
  2574 => x"08982b8c",
  2575 => x"08f40508",
  2576 => x"882a7072",
  2577 => x"078c08f0",
  2578 => x"0508882a",
  2579 => x"58585858",
  2580 => x"748c08f0",
  2581 => x"050c758c",
  2582 => x"08f4050c",
  2583 => x"8c08f005",
  2584 => x"08bfffff",
  2585 => x"068c08f8",
  2586 => x"050c8c08",
  2587 => x"f40508ff",
  2588 => x"068c08fc",
  2589 => x"050c8c08",
  2590 => x"e8050856",
  2591 => x"80708006",
  2592 => x"778fff06",
  2593 => x"70942b53",
  2594 => x"5a585580",
  2595 => x"0b8c08f8",
  2596 => x"05087607",
  2597 => x"8c08f805",
  2598 => x"0c708c08",
  2599 => x"fc050807",
  2600 => x"8c08fc05",
  2601 => x"0c8c08ec",
  2602 => x"05085156",
  2603 => x"80708006",
  2604 => x"77810670",
  2605 => x"9f2b535a",
  2606 => x"5855800b",
  2607 => x"8c08f805",
  2608 => x"0876078c",
  2609 => x"08f8050c",
  2610 => x"708c08fc",
  2611 => x"0508078c",
  2612 => x"08fc050c",
  2613 => x"568c08f8",
  2614 => x"05088c08",
  2615 => x"fc05088c",
  2616 => x"08880508",
  2617 => x"59575574",
  2618 => x"770c7584",
  2619 => x"180c8c08",
  2620 => x"88050880",
  2621 => x"0cbb3d0d",
  2622 => x"8c0c048c",
  2623 => x"08028c0c",
  2624 => x"ff3d0d80",
  2625 => x"0b8c08fc",
  2626 => x"050c8c08",
  2627 => x"88050851",
  2628 => x"7008822e",
  2629 => x"09810688",
  2630 => x"38810b8c",
  2631 => x"08fc050c",
  2632 => x"8c08fc05",
  2633 => x"0870800c",
  2634 => x"51833d0d",
  2635 => x"8c0c048c",
  2636 => x"08028c0c",
  2637 => x"ff3d0d80",
  2638 => x"0b8c08fc",
  2639 => x"050c8c08",
  2640 => x"88050851",
  2641 => x"7008842e",
  2642 => x"09810688",
  2643 => x"38810b8c",
  2644 => x"08fc050c",
  2645 => x"8c08fc05",
  2646 => x"0870800c",
  2647 => x"51833d0d",
  2648 => x"8c0c048c",
  2649 => x"08028c0c",
  2650 => x"ff3d0d80",
  2651 => x"0b8c08fc",
  2652 => x"050c8c08",
  2653 => x"88050851",
  2654 => x"7008802e",
  2655 => x"8f388c08",
  2656 => x"88050851",
  2657 => x"7008812e",
  2658 => x"83388839",
  2659 => x"810b8c08",
  2660 => x"fc050c8c",
  2661 => x"08fc0508",
  2662 => x"70800c51",
  2663 => x"833d0d8c",
  2664 => x"0c048c08",
  2665 => x"028c0cf8",
  2666 => x"3d0d8c08",
  2667 => x"88050870",
  2668 => x"08bfffff",
  2669 => x"068c08f8",
  2670 => x"050c8411",
  2671 => x"08ff068c",
  2672 => x"08fc050c",
  2673 => x"8c088805",
  2674 => x"08700894",
  2675 => x"2a545451",
  2676 => x"80728fff",
  2677 => x"068c08f4",
  2678 => x"050c8c08",
  2679 => x"88050870",
  2680 => x"089f2a54",
  2681 => x"54518072",
  2682 => x"81068c08",
  2683 => x"f0050c8c",
  2684 => x"088c0508",
  2685 => x"8c08f005",
  2686 => x"0884120c",
  2687 => x"51518c08",
  2688 => x"f4050881",
  2689 => x"bd388c08",
  2690 => x"f8050870",
  2691 => x"8c08fc05",
  2692 => x"08075151",
  2693 => x"708d388c",
  2694 => x"088c0508",
  2695 => x"5182710c",
  2696 => x"82d8398c",
  2697 => x"088c0508",
  2698 => x"8c08f405",
  2699 => x"08f88205",
  2700 => x"88120c8c",
  2701 => x"08fc0508",
  2702 => x"982a8c08",
  2703 => x"f8050888",
  2704 => x"2b707207",
  2705 => x"8c08fc05",
  2706 => x"08882b56",
  2707 => x"53555551",
  2708 => x"708c08f8",
  2709 => x"050c718c",
  2710 => x"08fc050c",
  2711 => x"8c088c05",
  2712 => x"08518371",
  2713 => x"0c8c08f8",
  2714 => x"0508f00a",
  2715 => x"26b7388c",
  2716 => x"08fc0508",
  2717 => x"9f2a8c08",
  2718 => x"f8050810",
  2719 => x"7072078c",
  2720 => x"08fc0508",
  2721 => x"10555354",
  2722 => x"54708c08",
  2723 => x"f8050c71",
  2724 => x"8c08fc05",
  2725 => x"0c8c088c",
  2726 => x"05088811",
  2727 => x"08ff0588",
  2728 => x"120c51c1",
  2729 => x"398c088c",
  2730 => x"0508538c",
  2731 => x"08f80508",
  2732 => x"8c08fc05",
  2733 => x"08535170",
  2734 => x"8c140c71",
  2735 => x"90140c81",
  2736 => x"b9398c08",
  2737 => x"f405088f",
  2738 => x"ff2e0981",
  2739 => x"0680e238",
  2740 => x"8c08f805",
  2741 => x"08708c08",
  2742 => x"fc050807",
  2743 => x"5151708d",
  2744 => x"388c088c",
  2745 => x"05085184",
  2746 => x"710c818e",
  2747 => x"398c08f8",
  2748 => x"0508932a",
  2749 => x"52807281",
  2750 => x"06515170",
  2751 => x"802e8c38",
  2752 => x"8c088c05",
  2753 => x"08518171",
  2754 => x"0c8a398c",
  2755 => x"088c0508",
  2756 => x"5180710c",
  2757 => x"8c088c05",
  2758 => x"08538c08",
  2759 => x"f805088c",
  2760 => x"08fc0508",
  2761 => x"5351708c",
  2762 => x"140c7190",
  2763 => x"140c80ca",
  2764 => x"398c088c",
  2765 => x"05088c08",
  2766 => x"f40508f8",
  2767 => x"81058812",
  2768 => x"0c8c088c",
  2769 => x"05085151",
  2770 => x"83710c8c",
  2771 => x"088c0508",
  2772 => x"8c08fc05",
  2773 => x"08982a8c",
  2774 => x"08f80508",
  2775 => x"882b7072",
  2776 => x"078c08fc",
  2777 => x"0508882b",
  2778 => x"71880a07",
  2779 => x"8c160c70",
  2780 => x"80079016",
  2781 => x"0c565455",
  2782 => x"55558a3d",
  2783 => x"0d8c0c04",
  2784 => x"fc3d0d76",
  2785 => x"70797b55",
  2786 => x"5555558f",
  2787 => x"72278c38",
  2788 => x"72750783",
  2789 => x"06517080",
  2790 => x"2ea738ff",
  2791 => x"125271ff",
  2792 => x"2e983872",
  2793 => x"70810554",
  2794 => x"33747081",
  2795 => x"055634ff",
  2796 => x"125271ff",
  2797 => x"2e098106",
  2798 => x"ea387480",
  2799 => x"0c863d0d",
  2800 => x"04745172",
  2801 => x"70840554",
  2802 => x"08717084",
  2803 => x"05530c72",
  2804 => x"70840554",
  2805 => x"08717084",
  2806 => x"05530c72",
  2807 => x"70840554",
  2808 => x"08717084",
  2809 => x"05530c72",
  2810 => x"70840554",
  2811 => x"08717084",
  2812 => x"05530cf0",
  2813 => x"1252718f",
  2814 => x"26c93883",
  2815 => x"72279538",
  2816 => x"72708405",
  2817 => x"54087170",
  2818 => x"8405530c",
  2819 => x"fc125271",
  2820 => x"8326ed38",
  2821 => x"7054ff83",
  2822 => x"39fd3d0d",
  2823 => x"800b80dd",
  2824 => x"c8085454",
  2825 => x"72812e9d",
  2826 => x"387380e5",
  2827 => x"cc0cffb0",
  2828 => x"af3fffaf",
  2829 => x"cb3f80dd",
  2830 => x"e8528151",
  2831 => x"ffbbd83f",
  2832 => x"800851a3",
  2833 => x"3f7280e5",
  2834 => x"cc0cffb0",
  2835 => x"933fffaf",
  2836 => x"af3f80dd",
  2837 => x"e8528151",
  2838 => x"ffbbbc3f",
  2839 => x"80085187",
  2840 => x"3f00ff39",
  2841 => x"00ff39f7",
  2842 => x"3d0d7b80",
  2843 => x"ddec0882",
  2844 => x"c811085a",
  2845 => x"545a7780",
  2846 => x"2e80da38",
  2847 => x"81881884",
  2848 => x"1908ff05",
  2849 => x"81712b59",
  2850 => x"55598074",
  2851 => x"2480ea38",
  2852 => x"807424b5",
  2853 => x"3873822b",
  2854 => x"78118805",
  2855 => x"56568180",
  2856 => x"19087706",
  2857 => x"5372802e",
  2858 => x"b6387816",
  2859 => x"70085353",
  2860 => x"79517408",
  2861 => x"53722dff",
  2862 => x"14fc17fc",
  2863 => x"1779812c",
  2864 => x"5a575754",
  2865 => x"738025d6",
  2866 => x"38770858",
  2867 => x"77ffad38",
  2868 => x"80ddec08",
  2869 => x"53bc1308",
  2870 => x"a5387951",
  2871 => x"ff833f74",
  2872 => x"0853722d",
  2873 => x"ff14fc17",
  2874 => x"fc177981",
  2875 => x"2c5a5757",
  2876 => x"54738025",
  2877 => x"ffa838d1",
  2878 => x"398057ff",
  2879 => x"93397251",
  2880 => x"bc130853",
  2881 => x"722d7951",
  2882 => x"fed73fff",
  2883 => x"3d0d80e4",
  2884 => x"f00bfc05",
  2885 => x"70085252",
  2886 => x"70ff2e91",
  2887 => x"38702dfc",
  2888 => x"12700852",
  2889 => x"5270ff2e",
  2890 => x"098106f1",
  2891 => x"38833d0d",
  2892 => x"0404ffaf",
  2893 => x"983f0400",
  2894 => x"00000040",
  2895 => x"4175746f",
  2896 => x"2d6e6567",
  2897 => x"6f746961",
  2898 => x"74696f6e",
  2899 => x"20666169",
  2900 => x"6c65640a",
  2901 => x"00000000",
  2902 => x"47524554",
  2903 => x"48280000",
  2904 => x"31302f31",
  2905 => x"30302f31",
  2906 => x"30303000",
  2907 => x"29204574",
  2908 => x"6865726e",
  2909 => x"6574204d",
  2910 => x"41432061",
  2911 => x"74205b30",
  2912 => x"78000000",
  2913 => x"5d2e2052",
  2914 => x"756e6e69",
  2915 => x"6e672000",
  2916 => x"31303000",
  2917 => x"204d6270",
  2918 => x"73200000",
  2919 => x"66756c6c",
  2920 => x"00000000",
  2921 => x"20647570",
  2922 => x"6c65780a",
  2923 => x"00000000",
  2924 => x"31302f31",
  2925 => x"30300000",
  2926 => x"31300000",
  2927 => x"68616c66",
  2928 => x"00000000",
  2929 => x"0c677265",
  2930 => x"74682e63",
  2931 => x"00000000",
  2932 => x"20286f6e",
  2933 => x"2073696d",
  2934 => x"290a0000",
  2935 => x"0a53656e",
  2936 => x"64696e67",
  2937 => x"20313530",
  2938 => x"30204d62",
  2939 => x"79746520",
  2940 => x"6f662064",
  2941 => x"61746120",
  2942 => x"746f2000",
  2943 => x"20706163",
  2944 => x"6b657473",
  2945 => x"290a0000",
  2946 => x"0a54696d",
  2947 => x"653a2000",
  2948 => x"20736563",
  2949 => x"0a000000",
  2950 => x"42697472",
  2951 => x"6174653a",
  2952 => x"20000000",
  2953 => x"206b6270",
  2954 => x"730a0000",
  2955 => x"20286f6e",
  2956 => x"20686172",
  2957 => x"64776172",
  2958 => x"65290a00",
  2959 => x"636f6d70",
  2960 => x"696c6564",
  2961 => x"3a204465",
  2962 => x"63202032",
  2963 => x"20323031",
  2964 => x"30202031",
  2965 => x"363a3034",
  2966 => x"3a34330a",
  2967 => x"00000000",
  2968 => x"30622020",
  2969 => x"20202020",
  2970 => x"20202020",
  2971 => x"20202020",
  2972 => x"20202020",
  2973 => x"20202020",
  2974 => x"20202020",
  2975 => x"20202020",
  2976 => x"20200000",
  2977 => x"20202020",
  2978 => x"20202020",
  2979 => x"00000000",
  2980 => x"00000000",
  2981 => x"00000000",
  2982 => x"00000000",
  2983 => x"00000000",
  2984 => x"00000000",
  2985 => x"64756d6d",
  2986 => x"792e6578",
  2987 => x"65000000",
  2988 => x"43000000",
  2989 => x"00ffffff",
  2990 => x"ff00ffff",
  2991 => x"ffff00ff",
  2992 => x"ffffff00",
  2993 => x"00000000",
  2994 => x"00000000",
  2995 => x"00000000",
  2996 => x"00003278",
  2997 => x"80000d00",
  2998 => x"80000800",
  2999 => x"80000600",
  3000 => x"80000200",
  3001 => x"80000100",
  3002 => x"00002ea4",
  3003 => x"00002ef0",
  3004 => x"00000000",
  3005 => x"00003158",
  3006 => x"000031b4",
  3007 => x"00003210",
  3008 => x"00000000",
  3009 => x"00000000",
  3010 => x"00000000",
  3011 => x"00000000",
  3012 => x"00000000",
  3013 => x"00000000",
  3014 => x"00000000",
  3015 => x"00000000",
  3016 => x"00000000",
  3017 => x"00002eb0",
  3018 => x"00000000",
  3019 => x"00000000",
  3020 => x"00000000",
  3021 => x"00000000",
  3022 => x"00000000",
  3023 => x"00000000",
  3024 => x"00000000",
  3025 => x"00000000",
  3026 => x"00000000",
  3027 => x"00000000",
  3028 => x"00000000",
  3029 => x"00000000",
  3030 => x"00000000",
  3031 => x"00000000",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"00000000",
  3041 => x"00000000",
  3042 => x"00000000",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000000",
  3046 => x"00000001",
  3047 => x"330eabcd",
  3048 => x"1234e66d",
  3049 => x"deec0005",
  3050 => x"000b0000",
  3051 => x"00000000",
  3052 => x"00000000",
  3053 => x"00000000",
  3054 => x"00000000",
  3055 => x"00000000",
  3056 => x"00000000",
  3057 => x"00000000",
  3058 => x"00000000",
  3059 => x"00000000",
  3060 => x"00000000",
  3061 => x"00000000",
  3062 => x"00000000",
  3063 => x"00000000",
  3064 => x"00000000",
  3065 => x"00000000",
  3066 => x"00000000",
  3067 => x"00000000",
  3068 => x"00000000",
  3069 => x"00000000",
  3070 => x"00000000",
  3071 => x"00000000",
  3072 => x"00000000",
  3073 => x"00000000",
  3074 => x"00000000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000000",
  3084 => x"00000000",
  3085 => x"00000000",
  3086 => x"00000000",
  3087 => x"00000000",
  3088 => x"00000000",
  3089 => x"00000000",
  3090 => x"00000000",
  3091 => x"00000000",
  3092 => x"00000000",
  3093 => x"00000000",
  3094 => x"00000000",
  3095 => x"00000000",
  3096 => x"00000000",
  3097 => x"00000000",
  3098 => x"00000000",
  3099 => x"00000000",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00000000",
  3103 => x"00000000",
  3104 => x"00000000",
  3105 => x"00000000",
  3106 => x"00000000",
  3107 => x"00000000",
  3108 => x"00000000",
  3109 => x"00000000",
  3110 => x"00000000",
  3111 => x"00000000",
  3112 => x"00000000",
  3113 => x"00000000",
  3114 => x"00000000",
  3115 => x"00000000",
  3116 => x"00000000",
  3117 => x"00000000",
  3118 => x"00000000",
  3119 => x"00000000",
  3120 => x"00000000",
  3121 => x"00000000",
  3122 => x"00000000",
  3123 => x"00000000",
  3124 => x"00000000",
  3125 => x"00000000",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000000",
  3151 => x"00000000",
  3152 => x"00000000",
  3153 => x"00000000",
  3154 => x"00000000",
  3155 => x"00000000",
  3156 => x"00000000",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"00000000",
  3161 => x"00000000",
  3162 => x"00000000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"00000000",
  3166 => x"00000000",
  3167 => x"00000000",
  3168 => x"00000000",
  3169 => x"00000000",
  3170 => x"00000000",
  3171 => x"00000000",
  3172 => x"00000000",
  3173 => x"00000000",
  3174 => x"00000000",
  3175 => x"00000000",
  3176 => x"00000000",
  3177 => x"00000000",
  3178 => x"00000000",
  3179 => x"00000000",
  3180 => x"00000000",
  3181 => x"00000000",
  3182 => x"00000000",
  3183 => x"00000000",
  3184 => x"00000000",
  3185 => x"00000000",
  3186 => x"00000000",
  3187 => x"00000000",
  3188 => x"00000000",
  3189 => x"00000000",
  3190 => x"00000000",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00000000",
  3195 => x"00000000",
  3196 => x"00000000",
  3197 => x"00000000",
  3198 => x"00000000",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"ffffffff",
  3228 => x"00000000",
  3229 => x"ffffffff",
  3230 => x"00000000",
  3231 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
