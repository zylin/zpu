-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0bbedc0c",
     3 => x"3a0b0b0b",
     4 => x"b1d50400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0bb2972d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bbe",
   162 => x"c8738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0bac",
   171 => x"c02d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bad",
   179 => x"f22d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bbed80c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81fb3fab",
   257 => x"b73f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104be",
   280 => x"d808802e",
   281 => x"a338bedc",
   282 => x"08822ebd",
   283 => x"38838080",
   284 => x"0b0b0b80",
   285 => x"c6980c82",
   286 => x"a0800b80",
   287 => x"c69c0c82",
   288 => x"90800b80",
   289 => x"c6a00c04",
   290 => x"f8808080",
   291 => x"a40b0b0b",
   292 => x"80c6980c",
   293 => x"f8808082",
   294 => x"800b80c6",
   295 => x"9c0cf880",
   296 => x"8084800b",
   297 => x"80c6a00c",
   298 => x"0480c0a8",
   299 => x"808c0b0b",
   300 => x"0b80c698",
   301 => x"0c80c0a8",
   302 => x"80940b80",
   303 => x"c69c0c0b",
   304 => x"0b0bb3e8",
   305 => x"0b80c6a0",
   306 => x"0c04ff3d",
   307 => x"0d80c6a4",
   308 => x"335170a4",
   309 => x"38bee408",
   310 => x"70085252",
   311 => x"70802e92",
   312 => x"388412be",
   313 => x"e40c702d",
   314 => x"bee40870",
   315 => x"08525270",
   316 => x"f038810b",
   317 => x"80c6a434",
   318 => x"833d0d04",
   319 => x"04803d0d",
   320 => x"0b0b80c6",
   321 => x"9408802e",
   322 => x"8e380b0b",
   323 => x"0b0b800b",
   324 => x"802e0981",
   325 => x"06853882",
   326 => x"3d0d040b",
   327 => x"0b80c694",
   328 => x"510b0b0b",
   329 => x"f5da3f82",
   330 => x"3d0d0404",
   331 => x"fb3d0d77",
   332 => x"70713370",
   333 => x"81ff0654",
   334 => x"55555570",
   335 => x"802eb038",
   336 => x"befc0852",
   337 => x"7281ff06",
   338 => x"81155553",
   339 => x"728a2e80",
   340 => x"e7388412",
   341 => x"0870822a",
   342 => x"81065151",
   343 => x"70802ef2",
   344 => x"3872720c",
   345 => x"73337081",
   346 => x"ff065753",
   347 => x"75d63874",
   348 => x"75335253",
   349 => x"70802ebc",
   350 => x"3870bef4",
   351 => x"08555281",
   352 => x"1353718a",
   353 => x"2e80d638",
   354 => x"80c6ac33",
   355 => x"70101011",
   356 => x"80c6b033",
   357 => x"71902905",
   358 => x"70882b75",
   359 => x"07770c80",
   360 => x"c6b03381",
   361 => x"05595152",
   362 => x"557580c6",
   363 => x"b0347233",
   364 => x"5271cc38",
   365 => x"873d0d04",
   366 => x"84120870",
   367 => x"822a8106",
   368 => x"51567580",
   369 => x"2ef2388d",
   370 => x"720c8412",
   371 => x"0870822a",
   372 => x"81065151",
   373 => x"70802efe",
   374 => x"f938ff85",
   375 => x"3980c6ac",
   376 => x"337081ff",
   377 => x"06565274",
   378 => x"a3269938",
   379 => x"81125170",
   380 => x"80c6ac34",
   381 => x"800b80c6",
   382 => x"b0347233",
   383 => x"5271feff",
   384 => x"38ffb139",
   385 => x"800b80c6",
   386 => x"ac34800b",
   387 => x"80c6b034",
   388 => x"e939f53d",
   389 => x"0d7e0284",
   390 => x"05b70533",
   391 => x"8c3d5b55",
   392 => x"578b53b3",
   393 => x"ec527851",
   394 => x"a4923f82",
   395 => x"5673882e",
   396 => x"96388456",
   397 => x"73902e8f",
   398 => x"38885673",
   399 => x"a02e8838",
   400 => x"74567480",
   401 => x"2ea73802",
   402 => x"a5055876",
   403 => x"8f065473",
   404 => x"89268193",
   405 => x"387518b0",
   406 => x"15555573",
   407 => x"75347684",
   408 => x"2aff1770",
   409 => x"81ff0658",
   410 => x"555775df",
   411 => x"38787933",
   412 => x"55577380",
   413 => x"2ea83873",
   414 => x"befc0856",
   415 => x"56811757",
   416 => x"758a2e80",
   417 => x"fe388415",
   418 => x"0870822a",
   419 => x"81065154",
   420 => x"73802ef2",
   421 => x"3875750c",
   422 => x"76335675",
   423 => x"e0387879",
   424 => x"33555673",
   425 => x"802ebc38",
   426 => x"73bef408",
   427 => x"58558116",
   428 => x"56748a2e",
   429 => x"80f23880",
   430 => x"c6ac3370",
   431 => x"10101180",
   432 => x"c6b03371",
   433 => x"90290570",
   434 => x"882b7807",
   435 => x"7a0c80c6",
   436 => x"b0338105",
   437 => x"52525558",
   438 => x"7380c6b0",
   439 => x"34753355",
   440 => x"74cc388d",
   441 => x"3d0d0475",
   442 => x"18b71555",
   443 => x"55737534",
   444 => x"76842aff",
   445 => x"177081ff",
   446 => x"06585557",
   447 => x"75fecc38",
   448 => x"feeb3984",
   449 => x"15087082",
   450 => x"2a810651",
   451 => x"5877802e",
   452 => x"f2388d75",
   453 => x"0c841508",
   454 => x"70822a81",
   455 => x"06515473",
   456 => x"802efee2",
   457 => x"38feee39",
   458 => x"80c6ac33",
   459 => x"7081ff06",
   460 => x"5a5578a3",
   461 => x"26993881",
   462 => x"15587780",
   463 => x"c6ac3480",
   464 => x"0b80c6b0",
   465 => x"34753355",
   466 => x"74fee338",
   467 => x"ff953980",
   468 => x"0b80c6ac",
   469 => x"34800b80",
   470 => x"c6b034e9",
   471 => x"39fd3d0d",
   472 => x"bef00854",
   473 => x"80d50b84",
   474 => x"150cbefc",
   475 => x"08528412",
   476 => x"08810651",
   477 => x"70802ef6",
   478 => x"38710870",
   479 => x"81ff06f6",
   480 => x"11525451",
   481 => x"70ae268b",
   482 => x"38701010",
   483 => x"bcc80551",
   484 => x"70080484",
   485 => x"12087082",
   486 => x"2a708106",
   487 => x"51515170",
   488 => x"802ef038",
   489 => x"ab720c72",
   490 => x"8a2eaa38",
   491 => x"84120870",
   492 => x"822a7081",
   493 => x"06515151",
   494 => x"70802ef0",
   495 => x"3872720c",
   496 => x"84120870",
   497 => x"822a8106",
   498 => x"51537280",
   499 => x"2ef238ad",
   500 => x"720cff9a",
   501 => x"39841208",
   502 => x"70822a70",
   503 => x"81065151",
   504 => x"5170802e",
   505 => x"f0388d72",
   506 => x"0c841208",
   507 => x"70822a70",
   508 => x"81065151",
   509 => x"5170802e",
   510 => x"ffb238c1",
   511 => x"3981ff0b",
   512 => x"84150cfe",
   513 => x"e93980ff",
   514 => x"0b84150c",
   515 => x"fee039bf",
   516 => x"0b84150c",
   517 => x"fed8399f",
   518 => x"0b84150c",
   519 => x"fed0398f",
   520 => x"0b84150c",
   521 => x"fec83987",
   522 => x"0b84150c",
   523 => x"fec03983",
   524 => x"0b84150c",
   525 => x"feb83981",
   526 => x"0b84150c",
   527 => x"feb03980",
   528 => x"0b84150c",
   529 => x"fea839fc",
   530 => x"3d0d890a",
   531 => x"0bb69c52",
   532 => x"54f9d93f",
   533 => x"7352a051",
   534 => x"fbb83fb6",
   535 => x"ac51f9cc",
   536 => x"3f9452a0",
   537 => x"51fbab3f",
   538 => x"b6b851f9",
   539 => x"bf3f8053",
   540 => x"72747084",
   541 => x"05560c81",
   542 => x"13539473",
   543 => x"26f23889",
   544 => x"0a558054",
   545 => x"74085380",
   546 => x"c6a80880",
   547 => x"c938b6bc",
   548 => x"51f9993f",
   549 => x"7452a051",
   550 => x"faf83fb6",
   551 => x"cc51f98c",
   552 => x"3f7352a0",
   553 => x"51faeb3f",
   554 => x"b6d851f8",
   555 => x"ff3f7252",
   556 => x"a051fade",
   557 => x"3f73732e",
   558 => x"be38b6e0",
   559 => x"51f8ed3f",
   560 => x"b6e851f8",
   561 => x"e73f8415",
   562 => x"81155555",
   563 => x"947426ff",
   564 => x"b338863d",
   565 => x"0d04b6d8",
   566 => x"51f8d13f",
   567 => x"7252a051",
   568 => x"fab03fb6",
   569 => x"e851f8c4",
   570 => x"3f841581",
   571 => x"15555594",
   572 => x"7426ff90",
   573 => x"38dc39b6",
   574 => x"ec51f8b0",
   575 => x"3fc239f1",
   576 => x"3d0db6f0",
   577 => x"51f8a53f",
   578 => x"bee80870",
   579 => x"08b78053",
   580 => x"5b53f898",
   581 => x"3f7981ff",
   582 => x"ff068d3d",
   583 => x"705b5c53",
   584 => x"80735657",
   585 => x"76732487",
   586 => x"ba387817",
   587 => x"548a5274",
   588 => x"5199e83f",
   589 => x"8008b005",
   590 => x"56757434",
   591 => x"8117578a",
   592 => x"52745199",
   593 => x"b13f8008",
   594 => x"558008de",
   595 => x"38800877",
   596 => x"9f2a1870",
   597 => x"812c5a56",
   598 => x"56807825",
   599 => x"9e387817",
   600 => x"ff055575",
   601 => x"19703355",
   602 => x"53743373",
   603 => x"34737534",
   604 => x"8116ff16",
   605 => x"56567776",
   606 => x"24e93876",
   607 => x"19568076",
   608 => x"347a51f7",
   609 => x"a73fb794",
   610 => x"51f7a13f",
   611 => x"798f2a81",
   612 => x"06528851",
   613 => x"f8fc3fb7",
   614 => x"a851f790",
   615 => x"3f79902a",
   616 => x"81065288",
   617 => x"51f8eb3f",
   618 => x"b7bc51f6",
   619 => x"ff3f7995",
   620 => x"2a830653",
   621 => x"72812e90",
   622 => x"b2388173",
   623 => x"26909b38",
   624 => x"72822e90",
   625 => x"b8387283",
   626 => x"2e8fdf38",
   627 => x"b7d051f6",
   628 => x"db3f7997",
   629 => x"2a870683",
   630 => x"0581712b",
   631 => x"7c5b5455",
   632 => x"80735657",
   633 => x"76732488",
   634 => x"a0387817",
   635 => x"588a5274",
   636 => x"5198a83f",
   637 => x"8008b005",
   638 => x"53727834",
   639 => x"8117578a",
   640 => x"52745197",
   641 => x"f13f8008",
   642 => x"558008de",
   643 => x"38800877",
   644 => x"9f2a1870",
   645 => x"812c5a56",
   646 => x"56807825",
   647 => x"9e387817",
   648 => x"ff055575",
   649 => x"19703355",
   650 => x"53743373",
   651 => x"34737534",
   652 => x"8116ff16",
   653 => x"56567776",
   654 => x"24e93876",
   655 => x"19568076",
   656 => x"347a51f5",
   657 => x"e73fb7e4",
   658 => x"51f5e13f",
   659 => x"b7ec51f5",
   660 => x"db3f799a",
   661 => x"2a810681",
   662 => x"057b5a53",
   663 => x"80735657",
   664 => x"76732486",
   665 => x"f3387817",
   666 => x"588a5274",
   667 => x"5197ac3f",
   668 => x"8008b005",
   669 => x"54737834",
   670 => x"8117578a",
   671 => x"52745196",
   672 => x"f53f8008",
   673 => x"558008de",
   674 => x"38800877",
   675 => x"9f2a1870",
   676 => x"812c5a56",
   677 => x"56807825",
   678 => x"9e387817",
   679 => x"ff055575",
   680 => x"19703355",
   681 => x"53743373",
   682 => x"34737534",
   683 => x"8116ff16",
   684 => x"56567776",
   685 => x"24e93876",
   686 => x"19568076",
   687 => x"347a51f4",
   688 => x"eb3fb880",
   689 => x"51f4e53f",
   690 => x"799b2a87",
   691 => x"0683057b",
   692 => x"5a538073",
   693 => x"56577673",
   694 => x"2485cc38",
   695 => x"7817588a",
   696 => x"52745196",
   697 => x"b63f8008",
   698 => x"b0055473",
   699 => x"78348117",
   700 => x"578a5274",
   701 => x"5195ff3f",
   702 => x"80085580",
   703 => x"08de3880",
   704 => x"08779f2a",
   705 => x"1870812c",
   706 => x"5a565680",
   707 => x"78259e38",
   708 => x"7817ff05",
   709 => x"55751970",
   710 => x"33555374",
   711 => x"33733473",
   712 => x"75348116",
   713 => x"ff165656",
   714 => x"777624e9",
   715 => x"38761956",
   716 => x"8076347a",
   717 => x"51f3f53f",
   718 => x"b89451f3",
   719 => x"ef3f799e",
   720 => x"2a82077b",
   721 => x"5a538073",
   722 => x"56577673",
   723 => x"2484a738",
   724 => x"7817588a",
   725 => x"52745195",
   726 => x"c23f8008",
   727 => x"b0055473",
   728 => x"78348117",
   729 => x"578a5274",
   730 => x"51958b3f",
   731 => x"80085580",
   732 => x"08de3880",
   733 => x"08779f2a",
   734 => x"1870812c",
   735 => x"5a565680",
   736 => x"78259e38",
   737 => x"7817ff05",
   738 => x"55751970",
   739 => x"33555374",
   740 => x"33733473",
   741 => x"75348116",
   742 => x"ff165656",
   743 => x"777624e9",
   744 => x"38761956",
   745 => x"8076347a",
   746 => x"51f3813f",
   747 => x"b8a851f2",
   748 => x"fb3f799f",
   749 => x"2a528851",
   750 => x"f4d83fbe",
   751 => x"e8088411",
   752 => x"08b8bc53",
   753 => x"5b57f2e4",
   754 => x"3f799fff",
   755 => x"067b5a53",
   756 => x"80735657",
   757 => x"76732482",
   758 => x"ec387817",
   759 => x"588a5274",
   760 => x"5194b83f",
   761 => x"8008b005",
   762 => x"54737834",
   763 => x"8117578a",
   764 => x"52745194",
   765 => x"813f8008",
   766 => x"558008de",
   767 => x"38800877",
   768 => x"9f2a1870",
   769 => x"812c5a56",
   770 => x"56807825",
   771 => x"9e387817",
   772 => x"ff055575",
   773 => x"19703355",
   774 => x"53743373",
   775 => x"34737534",
   776 => x"8116ff16",
   777 => x"56567776",
   778 => x"24e93876",
   779 => x"19568076",
   780 => x"347a51f1",
   781 => x"f73fb8d0",
   782 => x"51f1f13f",
   783 => x"798c2a87",
   784 => x"06830581",
   785 => x"712b7c52",
   786 => x"54598073",
   787 => x"56577673",
   788 => x"2481c138",
   789 => x"7817588a",
   790 => x"52745193",
   791 => x"be3f8008",
   792 => x"b0055473",
   793 => x"78348117",
   794 => x"578a5274",
   795 => x"5193873f",
   796 => x"80085580",
   797 => x"08de3880",
   798 => x"08779f2a",
   799 => x"1870812c",
   800 => x"5a565680",
   801 => x"78259e38",
   802 => x"7817ff05",
   803 => x"55751970",
   804 => x"33555374",
   805 => x"33733473",
   806 => x"75348116",
   807 => x"ff165656",
   808 => x"777624e9",
   809 => x"38761956",
   810 => x"8076347a",
   811 => x"51f0fd3f",
   812 => x"b8e451f0",
   813 => x"f73f798f",
   814 => x"2a810652",
   815 => x"8851f2d2",
   816 => x"3fbee808",
   817 => x"881108b8",
   818 => x"f8535b59",
   819 => x"f0de3f79",
   820 => x"87065372",
   821 => x"862682e2",
   822 => x"38721010",
   823 => x"be840558",
   824 => x"770804ad",
   825 => x"7b3402ad",
   826 => x"05733071",
   827 => x"19565659",
   828 => x"8a527451",
   829 => x"92a53f80",
   830 => x"08b00556",
   831 => x"75743481",
   832 => x"17578a52",
   833 => x"745191ee",
   834 => x"3f800855",
   835 => x"8008f89a",
   836 => x"38f8ba39",
   837 => x"ad7b3402",
   838 => x"ad057330",
   839 => x"71195a56",
   840 => x"598a5274",
   841 => x"5191f43f",
   842 => x"8008b005",
   843 => x"54737834",
   844 => x"8117578a",
   845 => x"52745191",
   846 => x"bd3f8008",
   847 => x"558008fe",
   848 => x"9338feb3",
   849 => x"39ad7b34",
   850 => x"02ad0573",
   851 => x"3071195a",
   852 => x"56598a52",
   853 => x"745191c3",
   854 => x"3f8008b0",
   855 => x"05547378",
   856 => x"34811757",
   857 => x"8a527451",
   858 => x"918c3f80",
   859 => x"08558008",
   860 => x"fce838fd",
   861 => x"8839ad7b",
   862 => x"3402ad05",
   863 => x"73307119",
   864 => x"5a56598a",
   865 => x"52745191",
   866 => x"923f8008",
   867 => x"b0055473",
   868 => x"78348117",
   869 => x"578a5274",
   870 => x"5190db3f",
   871 => x"80085580",
   872 => x"08fbad38",
   873 => x"fbcd39ad",
   874 => x"7b3402ad",
   875 => x"05733071",
   876 => x"195a5659",
   877 => x"8a527451",
   878 => x"90e13f80",
   879 => x"08b00554",
   880 => x"73783481",
   881 => x"17578a52",
   882 => x"745190aa",
   883 => x"3f800855",
   884 => x"8008fa88",
   885 => x"38faa839",
   886 => x"ad7b3402",
   887 => x"ad057330",
   888 => x"71195a56",
   889 => x"598a5274",
   890 => x"5190b03f",
   891 => x"8008b005",
   892 => x"54737834",
   893 => x"8117578a",
   894 => x"5274518f",
   895 => x"f93f8008",
   896 => x"558008f8",
   897 => x"e138f981",
   898 => x"39ad7b34",
   899 => x"02ad0573",
   900 => x"3071195a",
   901 => x"56598a52",
   902 => x"74518fff",
   903 => x"3f8008b0",
   904 => x"05537278",
   905 => x"34811757",
   906 => x"8a527451",
   907 => x"8fc83f80",
   908 => x"08558008",
   909 => x"f7b438f7",
   910 => x"d439b98c",
   911 => x"51eded3f",
   912 => x"b99451ed",
   913 => x"e73fb99c",
   914 => x"51ede13f",
   915 => x"79832a83",
   916 => x"06537281",
   917 => x"2e879d38",
   918 => x"81732687",
   919 => x"85387282",
   920 => x"2e87ac38",
   921 => x"72832e86",
   922 => x"9738b9b0",
   923 => x"51edbd3f",
   924 => x"b9b451ed",
   925 => x"b73f7985",
   926 => x"2a870653",
   927 => x"72812e86",
   928 => x"a0388173",
   929 => x"2686ca38",
   930 => x"72822e86",
   931 => x"f9387283",
   932 => x"2e85e438",
   933 => x"b9c851ed",
   934 => x"933f7990",
   935 => x"2a708706",
   936 => x"51537285",
   937 => x"268b3872",
   938 => x"1010bea0",
   939 => x"05597808",
   940 => x"04b98c51",
   941 => x"ecf63fb9",
   942 => x"dc51ecf0",
   943 => x"3f79932a",
   944 => x"83068207",
   945 => x"7b5a5380",
   946 => x"73565776",
   947 => x"732484f6",
   948 => x"38781756",
   949 => x"8a527451",
   950 => x"8ec13f80",
   951 => x"08b00558",
   952 => x"77763481",
   953 => x"17578a52",
   954 => x"74518e8a",
   955 => x"3f800855",
   956 => x"8008de38",
   957 => x"8008779f",
   958 => x"2a187081",
   959 => x"2c5a5656",
   960 => x"8078259e",
   961 => x"387817ff",
   962 => x"05557519",
   963 => x"70335553",
   964 => x"74337334",
   965 => x"73753481",
   966 => x"16ff1656",
   967 => x"56777624",
   968 => x"e9387619",
   969 => x"56807634",
   970 => x"7a51ec80",
   971 => x"3fb9f051",
   972 => x"ebfa3f79",
   973 => x"942a8f06",
   974 => x"7b5a5380",
   975 => x"73565776",
   976 => x"732483d1",
   977 => x"38781758",
   978 => x"8a527451",
   979 => x"8dcd3f80",
   980 => x"08b00554",
   981 => x"73783481",
   982 => x"17578a52",
   983 => x"74518d96",
   984 => x"3f800855",
   985 => x"8008de38",
   986 => x"8008779f",
   987 => x"2a187081",
   988 => x"2c5a5656",
   989 => x"8078259e",
   990 => x"387817ff",
   991 => x"05557519",
   992 => x"70335553",
   993 => x"74337334",
   994 => x"73753481",
   995 => x"16ff1656",
   996 => x"56777624",
   997 => x"e9387619",
   998 => x"56807634",
   999 => x"7a51eb8c",
  1000 => x"3fba8451",
  1001 => x"eb863f79",
  1002 => x"982a8106",
  1003 => x"81057b5a",
  1004 => x"53807356",
  1005 => x"57767324",
  1006 => x"82aa3878",
  1007 => x"17588a52",
  1008 => x"74518cd7",
  1009 => x"3f8008b0",
  1010 => x"05547378",
  1011 => x"34811757",
  1012 => x"8a527451",
  1013 => x"8ca03f80",
  1014 => x"08558008",
  1015 => x"de388008",
  1016 => x"779f2a18",
  1017 => x"70812c5a",
  1018 => x"56568078",
  1019 => x"259e3878",
  1020 => x"17ff0555",
  1021 => x"75197033",
  1022 => x"55537433",
  1023 => x"73347375",
  1024 => x"348116ff",
  1025 => x"16565677",
  1026 => x"7624e938",
  1027 => x"76195680",
  1028 => x"76347a51",
  1029 => x"ea963fba",
  1030 => x"9851ea90",
  1031 => x"3f799e2a",
  1032 => x"82077b5a",
  1033 => x"53807356",
  1034 => x"57767324",
  1035 => x"81853878",
  1036 => x"17588a52",
  1037 => x"74518be3",
  1038 => x"3f8008b0",
  1039 => x"05547378",
  1040 => x"34811757",
  1041 => x"8a527451",
  1042 => x"8bac3f80",
  1043 => x"08558008",
  1044 => x"de388008",
  1045 => x"779f2a18",
  1046 => x"70812c5a",
  1047 => x"56568078",
  1048 => x"259e3878",
  1049 => x"17ff0555",
  1050 => x"75197033",
  1051 => x"55537433",
  1052 => x"73347375",
  1053 => x"348116ff",
  1054 => x"16565677",
  1055 => x"7624e938",
  1056 => x"76195680",
  1057 => x"76347a51",
  1058 => x"e9a23fba",
  1059 => x"ac51e99c",
  1060 => x"3f799f2a",
  1061 => x"528851ea",
  1062 => x"f93fbee8",
  1063 => x"08901108",
  1064 => x"bac0535b",
  1065 => x"5be9853f",
  1066 => x"7952a051",
  1067 => x"eae43f91",
  1068 => x"3d0d04ad",
  1069 => x"7b3402ad",
  1070 => x"05733071",
  1071 => x"195a5659",
  1072 => x"8a527451",
  1073 => x"8ad53f80",
  1074 => x"08b00554",
  1075 => x"73783481",
  1076 => x"17578a52",
  1077 => x"74518a9e",
  1078 => x"3f800855",
  1079 => x"8008fecf",
  1080 => x"38feef39",
  1081 => x"ad7b3402",
  1082 => x"ad057330",
  1083 => x"71195a56",
  1084 => x"598a5274",
  1085 => x"518aa43f",
  1086 => x"8008b005",
  1087 => x"54737834",
  1088 => x"8117578a",
  1089 => x"52745189",
  1090 => x"ed3f8008",
  1091 => x"558008fd",
  1092 => x"aa38fdca",
  1093 => x"39ad7b34",
  1094 => x"02ad0573",
  1095 => x"3071195a",
  1096 => x"56598a52",
  1097 => x"745189f3",
  1098 => x"3f8008b0",
  1099 => x"05547378",
  1100 => x"34811757",
  1101 => x"8a527451",
  1102 => x"89bc3f80",
  1103 => x"08558008",
  1104 => x"fc8338fc",
  1105 => x"a339ad7b",
  1106 => x"3402ad05",
  1107 => x"73307119",
  1108 => x"5856598a",
  1109 => x"52745189",
  1110 => x"c23f8008",
  1111 => x"b0055877",
  1112 => x"76348117",
  1113 => x"578a5274",
  1114 => x"51898b3f",
  1115 => x"80085580",
  1116 => x"08fade38",
  1117 => x"fafe39ba",
  1118 => x"d451e7b0",
  1119 => x"3ffa9539",
  1120 => x"bad851e7",
  1121 => x"a73fb9b0",
  1122 => x"51e7a13f",
  1123 => x"b9b451e7",
  1124 => x"9b3f7985",
  1125 => x"2a870653",
  1126 => x"72812e09",
  1127 => x"8106f9e2",
  1128 => x"38badc51",
  1129 => x"e7863ff9",
  1130 => x"eb39bae4",
  1131 => x"51e6fd3f",
  1132 => x"b7d051e6",
  1133 => x"f73f7997",
  1134 => x"2a870683",
  1135 => x"0581712b",
  1136 => x"7c5b5455",
  1137 => x"80735657",
  1138 => x"727725f0",
  1139 => x"9d38f8b9",
  1140 => x"39baec51",
  1141 => x"e6d63ff9",
  1142 => x"bb39baf4",
  1143 => x"51e6cd3f",
  1144 => x"cf39bafc",
  1145 => x"51e6c53f",
  1146 => x"ff9c39bb",
  1147 => x"8051e6bc",
  1148 => x"3fffbd39",
  1149 => x"bb8851e6",
  1150 => x"b33fff8a",
  1151 => x"39bb8c51",
  1152 => x"e6aa3fff",
  1153 => x"ab39bb94",
  1154 => x"51e6a13f",
  1155 => x"f98639bb",
  1156 => x"9851e698",
  1157 => x"3ffeef39",
  1158 => x"bb9c51f8",
  1159 => x"a039bb94",
  1160 => x"51f89a39",
  1161 => x"bba051f8",
  1162 => x"9439bba4",
  1163 => x"51f88e39",
  1164 => x"bba851e5",
  1165 => x"f73fb9dc",
  1166 => x"51e5f13f",
  1167 => x"79932a83",
  1168 => x"0682077b",
  1169 => x"5a538073",
  1170 => x"56577277",
  1171 => x"25f98238",
  1172 => x"fdf439bb",
  1173 => x"b851e5d4",
  1174 => x"3fb9dc51",
  1175 => x"e5ce3f79",
  1176 => x"932a8306",
  1177 => x"82077b5a",
  1178 => x"53807356",
  1179 => x"57727725",
  1180 => x"f8df38fd",
  1181 => x"d139bbc4",
  1182 => x"51e5b13f",
  1183 => x"b9dc51e5",
  1184 => x"ab3f7993",
  1185 => x"2a830682",
  1186 => x"077b5a53",
  1187 => x"80735657",
  1188 => x"727725f8",
  1189 => x"bc38fdae",
  1190 => x"39bbd451",
  1191 => x"e58e3fb9",
  1192 => x"dc51e588",
  1193 => x"3f79932a",
  1194 => x"83068207",
  1195 => x"7b5a5380",
  1196 => x"73565772",
  1197 => x"7725f899",
  1198 => x"38fd8b39",
  1199 => x"bbe051e4",
  1200 => x"eb3fb9dc",
  1201 => x"51e4e53f",
  1202 => x"79932a83",
  1203 => x"0682077b",
  1204 => x"5a538073",
  1205 => x"56577277",
  1206 => x"25f7f638",
  1207 => x"fce839fc",
  1208 => x"3d0dbef0",
  1209 => x"08700881",
  1210 => x"0a0680c6",
  1211 => x"a80cbef8",
  1212 => x"08545487",
  1213 => x"0b84140c",
  1214 => x"bef40855",
  1215 => x"800b8416",
  1216 => x"0c83ffff",
  1217 => x"0b88160c",
  1218 => x"800b80c6",
  1219 => x"ac34800b",
  1220 => x"80c6b034",
  1221 => x"befc0853",
  1222 => x"b60b8c14",
  1223 => x"0c830b88",
  1224 => x"140c81ff",
  1225 => x"0b88150c",
  1226 => x"beec0854",
  1227 => x"ff0b8415",
  1228 => x"0cfc9480",
  1229 => x"0b88150c",
  1230 => x"82d0affd",
  1231 => x"fb0b8c15",
  1232 => x"0c80c074",
  1233 => x"0c730870",
  1234 => x"862a8106",
  1235 => x"515372f5",
  1236 => x"38901408",
  1237 => x"70832a81",
  1238 => x"06515574",
  1239 => x"f43881fc",
  1240 => x"80810b90",
  1241 => x"150c9014",
  1242 => x"0870832a",
  1243 => x"81065153",
  1244 => x"72f43880",
  1245 => x"fdc0810b",
  1246 => x"90150cb6",
  1247 => x"b851e3ac",
  1248 => x"3fbbfc51",
  1249 => x"e3a63f80",
  1250 => x"c6a80880",
  1251 => x"2e84e138",
  1252 => x"bc8451e3",
  1253 => x"973fbc94",
  1254 => x"51e3913f",
  1255 => x"c0808053",
  1256 => x"bbe851e3",
  1257 => x"873f7252",
  1258 => x"a051e4e6",
  1259 => x"3fbbf451",
  1260 => x"e2fa3f72",
  1261 => x"70840554",
  1262 => x"0852a051",
  1263 => x"e4d43fb6",
  1264 => x"e851e2e8",
  1265 => x"3fc08098",
  1266 => x"7327d538",
  1267 => x"800bbef8",
  1268 => x"085555bf",
  1269 => x"a9bc0b94",
  1270 => x"150c850b",
  1271 => x"98150c98",
  1272 => x"14087081",
  1273 => x"06515372",
  1274 => x"f638bfa9",
  1275 => x"bc0b9415",
  1276 => x"0c850b98",
  1277 => x"150c9814",
  1278 => x"08708106",
  1279 => x"515372f6",
  1280 => x"38bfa9bc",
  1281 => x"0b94150c",
  1282 => x"850b9815",
  1283 => x"0c981408",
  1284 => x"70810651",
  1285 => x"5372f638",
  1286 => x"bfa9bc0b",
  1287 => x"94150c85",
  1288 => x"0b98150c",
  1289 => x"98140870",
  1290 => x"81065153",
  1291 => x"72f638bf",
  1292 => x"a9bc0b94",
  1293 => x"150c850b",
  1294 => x"98150c98",
  1295 => x"14087081",
  1296 => x"06515372",
  1297 => x"f638bfa9",
  1298 => x"bc0b9415",
  1299 => x"0c850b98",
  1300 => x"150c9814",
  1301 => x"08708106",
  1302 => x"515372f6",
  1303 => x"38811555",
  1304 => x"8a7526fe",
  1305 => x"ee38800b",
  1306 => x"bef40856",
  1307 => x"5473882b",
  1308 => x"750c8114",
  1309 => x"54979074",
  1310 => x"26f33880",
  1311 => x"0b80c6ac",
  1312 => x"34800b80",
  1313 => x"c6b034e7",
  1314 => x"be3f800b",
  1315 => x"bef80855",
  1316 => x"55bfa9bc",
  1317 => x"0b94150c",
  1318 => x"850b9815",
  1319 => x"0c981408",
  1320 => x"70810651",
  1321 => x"5372f638",
  1322 => x"bfa9bc0b",
  1323 => x"94150c85",
  1324 => x"0b98150c",
  1325 => x"98140870",
  1326 => x"81065153",
  1327 => x"72f638bf",
  1328 => x"a9bc0b94",
  1329 => x"150c850b",
  1330 => x"98150c98",
  1331 => x"14087081",
  1332 => x"06515372",
  1333 => x"f638bfa9",
  1334 => x"bc0b9415",
  1335 => x"0c850b98",
  1336 => x"150c9814",
  1337 => x"08708106",
  1338 => x"515372f6",
  1339 => x"38bfa9bc",
  1340 => x"0b94150c",
  1341 => x"850b9815",
  1342 => x"0c981408",
  1343 => x"70810651",
  1344 => x"5372f638",
  1345 => x"bfa9bc0b",
  1346 => x"94150c85",
  1347 => x"0b98150c",
  1348 => x"98140870",
  1349 => x"81065153",
  1350 => x"72f63881",
  1351 => x"15558575",
  1352 => x"26feee38",
  1353 => x"72bef408",
  1354 => x"56547388",
  1355 => x"2b750c81",
  1356 => x"14549790",
  1357 => x"7426f338",
  1358 => x"800b80c6",
  1359 => x"ac34800b",
  1360 => x"80c6b034",
  1361 => x"e7b93f80",
  1362 => x"0bbef808",
  1363 => x"5555bfa9",
  1364 => x"bc0b9415",
  1365 => x"0c850b98",
  1366 => x"150c9814",
  1367 => x"08708106",
  1368 => x"515372f6",
  1369 => x"38bfa9bc",
  1370 => x"0b94150c",
  1371 => x"850b9815",
  1372 => x"0c981408",
  1373 => x"70810651",
  1374 => x"5372f638",
  1375 => x"bfa9bc0b",
  1376 => x"94150c85",
  1377 => x"0b98150c",
  1378 => x"98140870",
  1379 => x"81065153",
  1380 => x"72f638bf",
  1381 => x"a9bc0b94",
  1382 => x"150c850b",
  1383 => x"98150c98",
  1384 => x"14087081",
  1385 => x"06515372",
  1386 => x"f638bfa9",
  1387 => x"bc0b9415",
  1388 => x"0c850b98",
  1389 => x"150c9814",
  1390 => x"08708106",
  1391 => x"515372f6",
  1392 => x"38bfa9bc",
  1393 => x"0b94150c",
  1394 => x"850b9815",
  1395 => x"0c981408",
  1396 => x"70810651",
  1397 => x"5372f638",
  1398 => x"81155574",
  1399 => x"8527fd86",
  1400 => x"38bfa9bc",
  1401 => x"0b94150c",
  1402 => x"850b9815",
  1403 => x"0cfeeb39",
  1404 => x"bcb851fb",
  1405 => x"9e398c08",
  1406 => x"028c0cfd",
  1407 => x"3d0d8053",
  1408 => x"8c088c05",
  1409 => x"08528c08",
  1410 => x"88050851",
  1411 => x"82de3f80",
  1412 => x"0870800c",
  1413 => x"54853d0d",
  1414 => x"8c0c048c",
  1415 => x"08028c0c",
  1416 => x"fd3d0d81",
  1417 => x"538c088c",
  1418 => x"0508528c",
  1419 => x"08880508",
  1420 => x"5182b93f",
  1421 => x"80087080",
  1422 => x"0c54853d",
  1423 => x"0d8c0c04",
  1424 => x"8c08028c",
  1425 => x"0cf93d0d",
  1426 => x"800b8c08",
  1427 => x"fc050c8c",
  1428 => x"08880508",
  1429 => x"8025ab38",
  1430 => x"8c088805",
  1431 => x"08308c08",
  1432 => x"88050c80",
  1433 => x"0b8c08f4",
  1434 => x"050c8c08",
  1435 => x"fc050888",
  1436 => x"38810b8c",
  1437 => x"08f4050c",
  1438 => x"8c08f405",
  1439 => x"088c08fc",
  1440 => x"050c8c08",
  1441 => x"8c050880",
  1442 => x"25ab388c",
  1443 => x"088c0508",
  1444 => x"308c088c",
  1445 => x"050c800b",
  1446 => x"8c08f005",
  1447 => x"0c8c08fc",
  1448 => x"05088838",
  1449 => x"810b8c08",
  1450 => x"f0050c8c",
  1451 => x"08f00508",
  1452 => x"8c08fc05",
  1453 => x"0c80538c",
  1454 => x"088c0508",
  1455 => x"528c0888",
  1456 => x"05085181",
  1457 => x"a73f8008",
  1458 => x"708c08f8",
  1459 => x"050c548c",
  1460 => x"08fc0508",
  1461 => x"802e8c38",
  1462 => x"8c08f805",
  1463 => x"08308c08",
  1464 => x"f8050c8c",
  1465 => x"08f80508",
  1466 => x"70800c54",
  1467 => x"893d0d8c",
  1468 => x"0c048c08",
  1469 => x"028c0cfb",
  1470 => x"3d0d800b",
  1471 => x"8c08fc05",
  1472 => x"0c8c0888",
  1473 => x"05088025",
  1474 => x"93388c08",
  1475 => x"88050830",
  1476 => x"8c088805",
  1477 => x"0c810b8c",
  1478 => x"08fc050c",
  1479 => x"8c088c05",
  1480 => x"0880258c",
  1481 => x"388c088c",
  1482 => x"0508308c",
  1483 => x"088c050c",
  1484 => x"81538c08",
  1485 => x"8c050852",
  1486 => x"8c088805",
  1487 => x"0851ad3f",
  1488 => x"8008708c",
  1489 => x"08f8050c",
  1490 => x"548c08fc",
  1491 => x"0508802e",
  1492 => x"8c388c08",
  1493 => x"f8050830",
  1494 => x"8c08f805",
  1495 => x"0c8c08f8",
  1496 => x"05087080",
  1497 => x"0c54873d",
  1498 => x"0d8c0c04",
  1499 => x"8c08028c",
  1500 => x"0cfd3d0d",
  1501 => x"810b8c08",
  1502 => x"fc050c80",
  1503 => x"0b8c08f8",
  1504 => x"050c8c08",
  1505 => x"8c05088c",
  1506 => x"08880508",
  1507 => x"27ac388c",
  1508 => x"08fc0508",
  1509 => x"802ea338",
  1510 => x"800b8c08",
  1511 => x"8c050824",
  1512 => x"99388c08",
  1513 => x"8c050810",
  1514 => x"8c088c05",
  1515 => x"0c8c08fc",
  1516 => x"0508108c",
  1517 => x"08fc050c",
  1518 => x"c9398c08",
  1519 => x"fc050880",
  1520 => x"2e80c938",
  1521 => x"8c088c05",
  1522 => x"088c0888",
  1523 => x"050826a1",
  1524 => x"388c0888",
  1525 => x"05088c08",
  1526 => x"8c050831",
  1527 => x"8c088805",
  1528 => x"0c8c08f8",
  1529 => x"05088c08",
  1530 => x"fc050807",
  1531 => x"8c08f805",
  1532 => x"0c8c08fc",
  1533 => x"0508812a",
  1534 => x"8c08fc05",
  1535 => x"0c8c088c",
  1536 => x"0508812a",
  1537 => x"8c088c05",
  1538 => x"0cffaf39",
  1539 => x"8c089005",
  1540 => x"08802e8f",
  1541 => x"388c0888",
  1542 => x"0508708c",
  1543 => x"08f4050c",
  1544 => x"518d398c",
  1545 => x"08f80508",
  1546 => x"708c08f4",
  1547 => x"050c518c",
  1548 => x"08f40508",
  1549 => x"800c853d",
  1550 => x"0d8c0c04",
  1551 => x"fc3d0d76",
  1552 => x"70797b55",
  1553 => x"5555558f",
  1554 => x"72278c38",
  1555 => x"72750783",
  1556 => x"06517080",
  1557 => x"2ea738ff",
  1558 => x"125271ff",
  1559 => x"2e983872",
  1560 => x"70810554",
  1561 => x"33747081",
  1562 => x"055634ff",
  1563 => x"125271ff",
  1564 => x"2e098106",
  1565 => x"ea387480",
  1566 => x"0c863d0d",
  1567 => x"04745172",
  1568 => x"70840554",
  1569 => x"08717084",
  1570 => x"05530c72",
  1571 => x"70840554",
  1572 => x"08717084",
  1573 => x"05530c72",
  1574 => x"70840554",
  1575 => x"08717084",
  1576 => x"05530c72",
  1577 => x"70840554",
  1578 => x"08717084",
  1579 => x"05530cf0",
  1580 => x"1252718f",
  1581 => x"26c93883",
  1582 => x"72279538",
  1583 => x"72708405",
  1584 => x"54087170",
  1585 => x"8405530c",
  1586 => x"fc125271",
  1587 => x"8326ed38",
  1588 => x"7054ff83",
  1589 => x"39fd3d0d",
  1590 => x"800bbedc",
  1591 => x"08545472",
  1592 => x"812e9938",
  1593 => x"7380c6b4",
  1594 => x"0cd6f43f",
  1595 => x"d6923fbf",
  1596 => x"80528151",
  1597 => x"f3e93f80",
  1598 => x"08519f3f",
  1599 => x"7280c6b4",
  1600 => x"0cd6dc3f",
  1601 => x"d5fa3fbf",
  1602 => x"80528151",
  1603 => x"f3d13f80",
  1604 => x"0851873f",
  1605 => x"00ff3900",
  1606 => x"ff39f73d",
  1607 => x"0d7bbf84",
  1608 => x"0882c811",
  1609 => x"085a545a",
  1610 => x"77802e80",
  1611 => x"d9388188",
  1612 => x"18841908",
  1613 => x"ff058171",
  1614 => x"2b595559",
  1615 => x"80742480",
  1616 => x"e9388074",
  1617 => x"24b53873",
  1618 => x"822b7811",
  1619 => x"88055656",
  1620 => x"81801908",
  1621 => x"77065372",
  1622 => x"802eb538",
  1623 => x"78167008",
  1624 => x"53537951",
  1625 => x"74085372",
  1626 => x"2dff14fc",
  1627 => x"17fc1779",
  1628 => x"812c5a57",
  1629 => x"57547380",
  1630 => x"25d63877",
  1631 => x"085877ff",
  1632 => x"ad38bf84",
  1633 => x"0853bc13",
  1634 => x"08a53879",
  1635 => x"51ff853f",
  1636 => x"74085372",
  1637 => x"2dff14fc",
  1638 => x"17fc1779",
  1639 => x"812c5a57",
  1640 => x"57547380",
  1641 => x"25ffa938",
  1642 => x"d2398057",
  1643 => x"ff943972",
  1644 => x"51bc1308",
  1645 => x"53722d79",
  1646 => x"51fed93f",
  1647 => x"ff3d0d80",
  1648 => x"c6880bfc",
  1649 => x"05700852",
  1650 => x"5270ff2e",
  1651 => x"9138702d",
  1652 => x"fc127008",
  1653 => x"525270ff",
  1654 => x"2e098106",
  1655 => x"f138833d",
  1656 => x"0d0404d5",
  1657 => x"e53f0400",
  1658 => x"00000040",
  1659 => x"30782020",
  1660 => x"20202020",
  1661 => x"20200000",
  1662 => x"0a677265",
  1663 => x"74682072",
  1664 => x"65676973",
  1665 => x"74657273",
  1666 => x"3a000000",
  1667 => x"0a636f6e",
  1668 => x"74726f6c",
  1669 => x"3a202020",
  1670 => x"20202000",
  1671 => x"0a737461",
  1672 => x"7475733a",
  1673 => x"20202020",
  1674 => x"20202000",
  1675 => x"0a6d6163",
  1676 => x"5f6d7362",
  1677 => x"3a202020",
  1678 => x"20202000",
  1679 => x"0a6d6163",
  1680 => x"5f6c7362",
  1681 => x"3a202020",
  1682 => x"20202000",
  1683 => x"0a6d6469",
  1684 => x"6f5f636f",
  1685 => x"6e74726f",
  1686 => x"6c3a2000",
  1687 => x"0a74785f",
  1688 => x"706f696e",
  1689 => x"7465723a",
  1690 => x"20202000",
  1691 => x"0a72785f",
  1692 => x"706f696e",
  1693 => x"7465723a",
  1694 => x"20202000",
  1695 => x"0a656463",
  1696 => x"6c5f6970",
  1697 => x"3a202020",
  1698 => x"20202000",
  1699 => x"0a686173",
  1700 => x"685f6d73",
  1701 => x"623a2020",
  1702 => x"20202000",
  1703 => x"0a686173",
  1704 => x"685f6c73",
  1705 => x"623a2020",
  1706 => x"20202000",
  1707 => x"0a6d6469",
  1708 => x"6f207068",
  1709 => x"79207265",
  1710 => x"67697374",
  1711 => x"65727300",
  1712 => x"0a206d64",
  1713 => x"696f2070",
  1714 => x"68793a20",
  1715 => x"00000000",
  1716 => x"0a202072",
  1717 => x"65673a20",
  1718 => x"00000000",
  1719 => x"2d3e2000",
  1720 => x"0a677265",
  1721 => x"74682d3e",
  1722 => x"636f6e74",
  1723 => x"726f6c20",
  1724 => x"3a000000",
  1725 => x"0a677265",
  1726 => x"74682d3e",
  1727 => x"73746174",
  1728 => x"75732020",
  1729 => x"3a000000",
  1730 => x"0a646573",
  1731 => x"63722d3e",
  1732 => x"636f6e74",
  1733 => x"726f6c20",
  1734 => x"3a000000",
  1735 => x"77726974",
  1736 => x"65206164",
  1737 => x"64726573",
  1738 => x"733a2000",
  1739 => x"20206c65",
  1740 => x"6e677468",
  1741 => x"3a200000",
  1742 => x"0a0a0000",
  1743 => x"72656164",
  1744 => x"20206164",
  1745 => x"64726573",
  1746 => x"733a2000",
  1747 => x"20206578",
  1748 => x"70656374",
  1749 => x"3a200000",
  1750 => x"2020676f",
  1751 => x"743a2000",
  1752 => x"20657272",
  1753 => x"6f720000",
  1754 => x"0a000000",
  1755 => x"206f6b00",
  1756 => x"44445220",
  1757 => x"6d656d6f",
  1758 => x"72792069",
  1759 => x"6e666f00",
  1760 => x"0a617574",
  1761 => x"6f20745f",
  1762 => x"52455245",
  1763 => x"5348203a",
  1764 => x"00000000",
  1765 => x"0a636c6f",
  1766 => x"636b2065",
  1767 => x"6e61626c",
  1768 => x"6520203a",
  1769 => x"00000000",
  1770 => x"0a696e69",
  1771 => x"74616c69",
  1772 => x"7a652020",
  1773 => x"2020203a",
  1774 => x"00000000",
  1775 => x"0a636f6c",
  1776 => x"756d6e20",
  1777 => x"73697a65",
  1778 => x"2020203a",
  1779 => x"00000000",
  1780 => x"0a62616e",
  1781 => x"6b73697a",
  1782 => x"65202020",
  1783 => x"2020203a",
  1784 => x"00000000",
  1785 => x"4d627974",
  1786 => x"65000000",
  1787 => x"0a745f52",
  1788 => x"43442020",
  1789 => x"20202020",
  1790 => x"2020203a",
  1791 => x"00000000",
  1792 => x"0a745f52",
  1793 => x"46432020",
  1794 => x"20202020",
  1795 => x"2020203a",
  1796 => x"00000000",
  1797 => x"0a745f52",
  1798 => x"50202020",
  1799 => x"20202020",
  1800 => x"2020203a",
  1801 => x"00000000",
  1802 => x"0a726566",
  1803 => x"72657368",
  1804 => x"20656e2e",
  1805 => x"2020203a",
  1806 => x"00000000",
  1807 => x"0a444452",
  1808 => x"20667265",
  1809 => x"7175656e",
  1810 => x"6379203a",
  1811 => x"00000000",
  1812 => x"0a444452",
  1813 => x"20646174",
  1814 => x"61207769",
  1815 => x"6474683a",
  1816 => x"00000000",
  1817 => x"0a6d6f62",
  1818 => x"696c6520",
  1819 => x"73757070",
  1820 => x"6f72743a",
  1821 => x"00000000",
  1822 => x"0a73656c",
  1823 => x"66207265",
  1824 => x"66726573",
  1825 => x"6820203a",
  1826 => x"00000000",
  1827 => x"756e6b6e",
  1828 => x"6f776e00",
  1829 => x"20617272",
  1830 => x"61790000",
  1831 => x"0a74656d",
  1832 => x"702d636f",
  1833 => x"6d702072",
  1834 => x"6566723a",
  1835 => x"00000000",
  1836 => x"c2b04300",
  1837 => x"0a647269",
  1838 => x"76652073",
  1839 => x"7472656e",
  1840 => x"6774683a",
  1841 => x"00000000",
  1842 => x"0a706f77",
  1843 => x"65722073",
  1844 => x"6176696e",
  1845 => x"6720203a",
  1846 => x"00000000",
  1847 => x"0a745f58",
  1848 => x"50202020",
  1849 => x"20202020",
  1850 => x"2020203a",
  1851 => x"00000000",
  1852 => x"0a745f58",
  1853 => x"53522020",
  1854 => x"20202020",
  1855 => x"2020203a",
  1856 => x"00000000",
  1857 => x"0a745f43",
  1858 => x"4b452020",
  1859 => x"20202020",
  1860 => x"2020203a",
  1861 => x"00000000",
  1862 => x"0a434153",
  1863 => x"206c6174",
  1864 => x"656e6379",
  1865 => x"2020203a",
  1866 => x"00000000",
  1867 => x"0a6d6f62",
  1868 => x"696c6520",
  1869 => x"656e6162",
  1870 => x"6c65643a",
  1871 => x"00000000",
  1872 => x"0a737461",
  1873 => x"74757320",
  1874 => x"72656164",
  1875 => x"2020203a",
  1876 => x"00000000",
  1877 => x"332f3400",
  1878 => x"38350000",
  1879 => x"68616c66",
  1880 => x"00000000",
  1881 => x"34303639",
  1882 => x"00000000",
  1883 => x"66756c6c",
  1884 => x"00000000",
  1885 => x"20353132",
  1886 => x"00000000",
  1887 => x"37300000",
  1888 => x"31303234",
  1889 => x"00000000",
  1890 => x"34350000",
  1891 => x"32303438",
  1892 => x"00000000",
  1893 => x"312f3400",
  1894 => x"31350000",
  1895 => x"312f3800",
  1896 => x"312f3200",
  1897 => x"312f3100",
  1898 => x"64656570",
  1899 => x"20706f77",
  1900 => x"65722064",
  1901 => x"6f776e00",
  1902 => x"636c6f63",
  1903 => x"6b207374",
  1904 => x"6f700000",
  1905 => x"73656c66",
  1906 => x"20726566",
  1907 => x"72657368",
  1908 => x"00000000",
  1909 => x"706f7765",
  1910 => x"7220646f",
  1911 => x"776e0000",
  1912 => x"6e6f6e65",
  1913 => x"00000000",
  1914 => x"61646472",
  1915 => x"6573733a",
  1916 => x"20000000",
  1917 => x"20646174",
  1918 => x"613a2000",
  1919 => x"74657374",
  1920 => x"2e632000",
  1921 => x"286f6e20",
  1922 => x"73696d75",
  1923 => x"6c61746f",
  1924 => x"72290a00",
  1925 => x"636f6d70",
  1926 => x"696c6564",
  1927 => x"3a204175",
  1928 => x"67203233",
  1929 => x"20323031",
  1930 => x"30202031",
  1931 => x"373a3030",
  1932 => x"3a31390a",
  1933 => x"00000000",
  1934 => x"286f6e20",
  1935 => x"68617264",
  1936 => x"77617265",
  1937 => x"290a0000",
  1938 => x"0000076e",
  1939 => x"00000793",
  1940 => x"00000793",
  1941 => x"0000076e",
  1942 => x"00000793",
  1943 => x"00000793",
  1944 => x"00000793",
  1945 => x"00000793",
  1946 => x"00000793",
  1947 => x"00000793",
  1948 => x"00000793",
  1949 => x"00000793",
  1950 => x"00000793",
  1951 => x"00000793",
  1952 => x"00000793",
  1953 => x"00000793",
  1954 => x"00000793",
  1955 => x"00000793",
  1956 => x"00000793",
  1957 => x"00000793",
  1958 => x"00000793",
  1959 => x"00000793",
  1960 => x"00000793",
  1961 => x"00000793",
  1962 => x"00000793",
  1963 => x"00000793",
  1964 => x"00000793",
  1965 => x"00000793",
  1966 => x"00000793",
  1967 => x"00000793",
  1968 => x"00000793",
  1969 => x"00000793",
  1970 => x"00000793",
  1971 => x"00000793",
  1972 => x"00000793",
  1973 => x"00000793",
  1974 => x"00000793",
  1975 => x"00000793",
  1976 => x"0000083f",
  1977 => x"00000837",
  1978 => x"0000082f",
  1979 => x"00000827",
  1980 => x"0000081f",
  1981 => x"00000817",
  1982 => x"0000080f",
  1983 => x"00000806",
  1984 => x"000007fd",
  1985 => x"0000122a",
  1986 => x"00001224",
  1987 => x"0000121e",
  1988 => x"00000e3a",
  1989 => x"00000e3a",
  1990 => x"00001218",
  1991 => x"00001218",
  1992 => x"000012bc",
  1993 => x"00001299",
  1994 => x"00001276",
  1995 => x"00000eb1",
  1996 => x"00001253",
  1997 => x"00001230",
  1998 => x"64756d6d",
  1999 => x"792e6578",
  2000 => x"65000000",
  2001 => x"43000000",
  2002 => x"00ffffff",
  2003 => x"ff00ffff",
  2004 => x"ffff00ff",
  2005 => x"ffffff00",
  2006 => x"00000000",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00002310",
  2010 => x"fff00000",
  2011 => x"80000c00",
  2012 => x"80000800",
  2013 => x"80000600",
  2014 => x"80000200",
  2015 => x"80000100",
  2016 => x"00001f38",
  2017 => x"00001f88",
  2018 => x"00000000",
  2019 => x"000021f0",
  2020 => x"0000224c",
  2021 => x"000022a8",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00000000",
  2026 => x"00000000",
  2027 => x"00000000",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000000",
  2031 => x"00001f44",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"00000000",
  2049 => x"00000000",
  2050 => x"00000000",
  2051 => x"00000000",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000001",
  2061 => x"330eabcd",
  2062 => x"1234e66d",
  2063 => x"deec0005",
  2064 => x"000b0000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"00000000",
  2102 => x"00000000",
  2103 => x"00000000",
  2104 => x"00000000",
  2105 => x"00000000",
  2106 => x"00000000",
  2107 => x"00000000",
  2108 => x"00000000",
  2109 => x"00000000",
  2110 => x"00000000",
  2111 => x"00000000",
  2112 => x"00000000",
  2113 => x"00000000",
  2114 => x"00000000",
  2115 => x"00000000",
  2116 => x"00000000",
  2117 => x"00000000",
  2118 => x"00000000",
  2119 => x"00000000",
  2120 => x"00000000",
  2121 => x"00000000",
  2122 => x"00000000",
  2123 => x"00000000",
  2124 => x"00000000",
  2125 => x"00000000",
  2126 => x"00000000",
  2127 => x"00000000",
  2128 => x"00000000",
  2129 => x"00000000",
  2130 => x"00000000",
  2131 => x"00000000",
  2132 => x"00000000",
  2133 => x"00000000",
  2134 => x"00000000",
  2135 => x"00000000",
  2136 => x"00000000",
  2137 => x"00000000",
  2138 => x"00000000",
  2139 => x"00000000",
  2140 => x"00000000",
  2141 => x"00000000",
  2142 => x"00000000",
  2143 => x"00000000",
  2144 => x"00000000",
  2145 => x"00000000",
  2146 => x"00000000",
  2147 => x"00000000",
  2148 => x"00000000",
  2149 => x"00000000",
  2150 => x"00000000",
  2151 => x"00000000",
  2152 => x"00000000",
  2153 => x"00000000",
  2154 => x"00000000",
  2155 => x"00000000",
  2156 => x"00000000",
  2157 => x"00000000",
  2158 => x"00000000",
  2159 => x"00000000",
  2160 => x"00000000",
  2161 => x"00000000",
  2162 => x"00000000",
  2163 => x"00000000",
  2164 => x"00000000",
  2165 => x"00000000",
  2166 => x"00000000",
  2167 => x"00000000",
  2168 => x"00000000",
  2169 => x"00000000",
  2170 => x"00000000",
  2171 => x"00000000",
  2172 => x"00000000",
  2173 => x"00000000",
  2174 => x"00000000",
  2175 => x"00000000",
  2176 => x"00000000",
  2177 => x"00000000",
  2178 => x"00000000",
  2179 => x"00000000",
  2180 => x"00000000",
  2181 => x"00000000",
  2182 => x"00000000",
  2183 => x"00000000",
  2184 => x"00000000",
  2185 => x"00000000",
  2186 => x"00000000",
  2187 => x"00000000",
  2188 => x"00000000",
  2189 => x"00000000",
  2190 => x"00000000",
  2191 => x"00000000",
  2192 => x"00000000",
  2193 => x"00000000",
  2194 => x"00000000",
  2195 => x"00000000",
  2196 => x"00000000",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"00000000",
  2203 => x"00000000",
  2204 => x"00000000",
  2205 => x"00000000",
  2206 => x"00000000",
  2207 => x"00000000",
  2208 => x"00000000",
  2209 => x"00000000",
  2210 => x"00000000",
  2211 => x"00000000",
  2212 => x"00000000",
  2213 => x"00000000",
  2214 => x"00000000",
  2215 => x"00000000",
  2216 => x"00000000",
  2217 => x"00000000",
  2218 => x"00000000",
  2219 => x"00000000",
  2220 => x"00000000",
  2221 => x"00000000",
  2222 => x"00000000",
  2223 => x"00000000",
  2224 => x"00000000",
  2225 => x"00000000",
  2226 => x"00000000",
  2227 => x"00000000",
  2228 => x"00000000",
  2229 => x"00000000",
  2230 => x"00000000",
  2231 => x"00000000",
  2232 => x"00000000",
  2233 => x"00000000",
  2234 => x"00000000",
  2235 => x"00000000",
  2236 => x"00000000",
  2237 => x"00000000",
  2238 => x"00000000",
  2239 => x"00000000",
  2240 => x"00000000",
  2241 => x"ffffffff",
  2242 => x"00000000",
  2243 => x"ffffffff",
  2244 => x"00000000",
  2245 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
