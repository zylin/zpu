-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0b9ad40c",
     3 => x"3a0b0b0b",
     4 => x"97bb0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b97fb2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b9a",
   162 => x"c0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b93",
   171 => x"bf2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b94",
   179 => x"f12d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0b9ad00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f91",
   257 => x"9b3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"5351049a",
   280 => x"d008802e",
   281 => x"a1389ad4",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"a2840c82",
   286 => x"a0800ba2",
   287 => x"880c8290",
   288 => x"800ba28c",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0ba2",
   292 => x"840cf880",
   293 => x"8082800b",
   294 => x"a2880cf8",
   295 => x"80808480",
   296 => x"0ba28c0c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0ba284",
   300 => x"0c80c0a8",
   301 => x"80940ba2",
   302 => x"880c0b0b",
   303 => x"0b99cc0b",
   304 => x"a28c0c04",
   305 => x"ff3d0da2",
   306 => x"90335170",
   307 => x"a3389adc",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"9adc0c70",
   312 => x"2d9adc08",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0ba29034",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0ba2",
   319 => x"8008802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0ba280",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"fd3d0d9a",
   330 => x"e40876b0",
   331 => x"ea299412",
   332 => x"0c54850b",
   333 => x"98150c98",
   334 => x"14087081",
   335 => x"06515372",
   336 => x"f638853d",
   337 => x"0d04ff3d",
   338 => x"0d9ae408",
   339 => x"74101075",
   340 => x"10059412",
   341 => x"0c52850b",
   342 => x"98130c98",
   343 => x"12087081",
   344 => x"06515170",
   345 => x"f638833d",
   346 => x"0d04803d",
   347 => x"0d725180",
   348 => x"71278738",
   349 => x"ff115170",
   350 => x"fb38823d",
   351 => x"0d04803d",
   352 => x"0d9ae408",
   353 => x"51870b84",
   354 => x"120c823d",
   355 => x"0d04803d",
   356 => x"0d9ae808",
   357 => x"51b60b8c",
   358 => x"120c830b",
   359 => x"88120c82",
   360 => x"3d0d04ff",
   361 => x"3d0d9ae8",
   362 => x"08528412",
   363 => x"08708106",
   364 => x"51517080",
   365 => x"2ef43871",
   366 => x"087081ff",
   367 => x"06800c51",
   368 => x"833d0d04",
   369 => x"fe3d0d02",
   370 => x"9305339a",
   371 => x"e8085353",
   372 => x"84120870",
   373 => x"892a7081",
   374 => x"06515151",
   375 => x"70f23872",
   376 => x"720c843d",
   377 => x"0d04fe3d",
   378 => x"0d029305",
   379 => x"3353728a",
   380 => x"2e9b389a",
   381 => x"e8085284",
   382 => x"12087089",
   383 => x"2a708106",
   384 => x"51515170",
   385 => x"f2387272",
   386 => x"0c843d0d",
   387 => x"049ae808",
   388 => x"52841208",
   389 => x"70892a70",
   390 => x"81065151",
   391 => x"5170f238",
   392 => x"8d720c84",
   393 => x"12087089",
   394 => x"2a708106",
   395 => x"51515170",
   396 => x"c638d339",
   397 => x"fd3d0d75",
   398 => x"70335254",
   399 => x"70802ea7",
   400 => x"38709ae8",
   401 => x"08535381",
   402 => x"1454728a",
   403 => x"2e9d3884",
   404 => x"12087089",
   405 => x"2a708106",
   406 => x"51515170",
   407 => x"f2387272",
   408 => x"0c733353",
   409 => x"72e13885",
   410 => x"3d0d0484",
   411 => x"12087089",
   412 => x"2a708106",
   413 => x"51515170",
   414 => x"f2388d72",
   415 => x"0c841208",
   416 => x"70892a70",
   417 => x"81065151",
   418 => x"5170c438",
   419 => x"d139803d",
   420 => x"0d9ae008",
   421 => x"5181ff0b",
   422 => x"88120c82",
   423 => x"3d0d04fb",
   424 => x"3d0d8880",
   425 => x"e0870b9a",
   426 => x"e0089ae4",
   427 => x"08728413",
   428 => x"0c565755",
   429 => x"afd7c20b",
   430 => x"94150c85",
   431 => x"0b98150c",
   432 => x"98140870",
   433 => x"81065153",
   434 => x"72f63874",
   435 => x"9f2a7510",
   436 => x"07708418",
   437 => x"0c55afd7",
   438 => x"c20b9415",
   439 => x"0c850b98",
   440 => x"150cdd39",
   441 => x"fe3d0d9a",
   442 => x"e8085284",
   443 => x"12088106",
   444 => x"5170802e",
   445 => x"f6387108",
   446 => x"7081ff06",
   447 => x"54518412",
   448 => x"0870892a",
   449 => x"70810651",
   450 => x"515170f2",
   451 => x"38ab720c",
   452 => x"728a2ea6",
   453 => x"38841208",
   454 => x"70892a70",
   455 => x"81065151",
   456 => x"5170f238",
   457 => x"72720c84",
   458 => x"12087089",
   459 => x"2a810651",
   460 => x"5372f438",
   461 => x"ad720cff",
   462 => x"b2398412",
   463 => x"0870892a",
   464 => x"70810651",
   465 => x"515170f2",
   466 => x"388d720c",
   467 => x"84120870",
   468 => x"892a7081",
   469 => x"06515151",
   470 => x"70ffba38",
   471 => x"c739ff3d",
   472 => x"0d9ae008",
   473 => x"52710870",
   474 => x"8f067071",
   475 => x"842b0784",
   476 => x"150c5151",
   477 => x"7108708f",
   478 => x"06707184",
   479 => x"2b078415",
   480 => x"0c5151e1",
   481 => x"39fa3d0d",
   482 => x"9ae00870",
   483 => x"08810a06",
   484 => x"9ae40855",
   485 => x"5855870b",
   486 => x"84140c9a",
   487 => x"e80854b6",
   488 => x"0b8c150c",
   489 => x"830b8815",
   490 => x"0c99d00b",
   491 => x"99d03354",
   492 => x"5672802e",
   493 => x"a4387255",
   494 => x"81165674",
   495 => x"8a2e81f7",
   496 => x"38841408",
   497 => x"70892a70",
   498 => x"81065151",
   499 => x"5372f238",
   500 => x"74740c75",
   501 => x"335574e0",
   502 => x"3899d40b",
   503 => x"99d43354",
   504 => x"5672802e",
   505 => x"a4387255",
   506 => x"81165674",
   507 => x"8a2e81ec",
   508 => x"38841408",
   509 => x"70892a70",
   510 => x"81065151",
   511 => x"5372f238",
   512 => x"74740c75",
   513 => x"335574e0",
   514 => x"3876802e",
   515 => x"82b53899",
   516 => x"ec0b99ec",
   517 => x"33545672",
   518 => x"802ea238",
   519 => x"72558116",
   520 => x"56748a2e",
   521 => x"81db3884",
   522 => x"14087089",
   523 => x"2a810651",
   524 => x"5372f438",
   525 => x"74740c75",
   526 => x"335574e2",
   527 => x"3899fc0b",
   528 => x"99fc3354",
   529 => x"5672802e",
   530 => x"a2387255",
   531 => x"81165674",
   532 => x"8a2e81ce",
   533 => x"38841408",
   534 => x"70892a81",
   535 => x"06515372",
   536 => x"f4387474",
   537 => x"0c753355",
   538 => x"74e23884",
   539 => x"14088106",
   540 => x"5675802e",
   541 => x"f6387308",
   542 => x"7081ff06",
   543 => x"56578414",
   544 => x"0870892a",
   545 => x"81065457",
   546 => x"72f438ab",
   547 => x"740c748a",
   548 => x"2e828b38",
   549 => x"84140870",
   550 => x"892a8106",
   551 => x"545772f4",
   552 => x"3874740c",
   553 => x"84140870",
   554 => x"892a8106",
   555 => x"565674f4",
   556 => x"38ad740c",
   557 => x"ffb53984",
   558 => x"14087089",
   559 => x"2a708106",
   560 => x"51515372",
   561 => x"f2388d74",
   562 => x"0c841408",
   563 => x"70892a70",
   564 => x"81065151",
   565 => x"5372fde9",
   566 => x"38fdf539",
   567 => x"84140870",
   568 => x"892a7081",
   569 => x"06515153",
   570 => x"72f2388d",
   571 => x"740c8414",
   572 => x"0870892a",
   573 => x"70810651",
   574 => x"515372fd",
   575 => x"f438fe80",
   576 => x"39841408",
   577 => x"70892a81",
   578 => x"06515776",
   579 => x"f4388d74",
   580 => x"0c841408",
   581 => x"70892a81",
   582 => x"06515372",
   583 => x"fe8938fe",
   584 => x"93398414",
   585 => x"0870892a",
   586 => x"81065157",
   587 => x"76f4388d",
   588 => x"740c8414",
   589 => x"0870892a",
   590 => x"81065153",
   591 => x"72fe9638",
   592 => x"fea0399a",
   593 => x"a00b9aa0",
   594 => x"33545672",
   595 => x"802efded",
   596 => x"38728117",
   597 => x"5755748a",
   598 => x"2ea53884",
   599 => x"14087089",
   600 => x"2a810651",
   601 => x"5372f438",
   602 => x"74740c75",
   603 => x"33557480",
   604 => x"2efdca38",
   605 => x"81165674",
   606 => x"8a2e0981",
   607 => x"06dd3884",
   608 => x"14087089",
   609 => x"2a810651",
   610 => x"5776f438",
   611 => x"8d740c84",
   612 => x"14087089",
   613 => x"2a810651",
   614 => x"5372c038",
   615 => x"cb398414",
   616 => x"0870892a",
   617 => x"81065457",
   618 => x"72f4388d",
   619 => x"740c8414",
   620 => x"0870892a",
   621 => x"81065457",
   622 => x"72fdd938",
   623 => x"fde3398c",
   624 => x"08028c0c",
   625 => x"f93d0d80",
   626 => x"0b8c08fc",
   627 => x"050c8c08",
   628 => x"88050880",
   629 => x"25ab388c",
   630 => x"08880508",
   631 => x"308c0888",
   632 => x"050c800b",
   633 => x"8c08f405",
   634 => x"0c8c08fc",
   635 => x"05088838",
   636 => x"810b8c08",
   637 => x"f4050c8c",
   638 => x"08f40508",
   639 => x"8c08fc05",
   640 => x"0c8c088c",
   641 => x"05088025",
   642 => x"ab388c08",
   643 => x"8c050830",
   644 => x"8c088c05",
   645 => x"0c800b8c",
   646 => x"08f0050c",
   647 => x"8c08fc05",
   648 => x"08883881",
   649 => x"0b8c08f0",
   650 => x"050c8c08",
   651 => x"f005088c",
   652 => x"08fc050c",
   653 => x"80538c08",
   654 => x"8c050852",
   655 => x"8c088805",
   656 => x"085181a7",
   657 => x"3f800870",
   658 => x"8c08f805",
   659 => x"0c548c08",
   660 => x"fc050880",
   661 => x"2e8c388c",
   662 => x"08f80508",
   663 => x"308c08f8",
   664 => x"050c8c08",
   665 => x"f8050870",
   666 => x"800c5489",
   667 => x"3d0d8c0c",
   668 => x"048c0802",
   669 => x"8c0cfb3d",
   670 => x"0d800b8c",
   671 => x"08fc050c",
   672 => x"8c088805",
   673 => x"08802593",
   674 => x"388c0888",
   675 => x"0508308c",
   676 => x"0888050c",
   677 => x"810b8c08",
   678 => x"fc050c8c",
   679 => x"088c0508",
   680 => x"80258c38",
   681 => x"8c088c05",
   682 => x"08308c08",
   683 => x"8c050c81",
   684 => x"538c088c",
   685 => x"0508528c",
   686 => x"08880508",
   687 => x"51ad3f80",
   688 => x"08708c08",
   689 => x"f8050c54",
   690 => x"8c08fc05",
   691 => x"08802e8c",
   692 => x"388c08f8",
   693 => x"0508308c",
   694 => x"08f8050c",
   695 => x"8c08f805",
   696 => x"0870800c",
   697 => x"54873d0d",
   698 => x"8c0c048c",
   699 => x"08028c0c",
   700 => x"fd3d0d81",
   701 => x"0b8c08fc",
   702 => x"050c800b",
   703 => x"8c08f805",
   704 => x"0c8c088c",
   705 => x"05088c08",
   706 => x"88050827",
   707 => x"ac388c08",
   708 => x"fc050880",
   709 => x"2ea33880",
   710 => x"0b8c088c",
   711 => x"05082499",
   712 => x"388c088c",
   713 => x"0508108c",
   714 => x"088c050c",
   715 => x"8c08fc05",
   716 => x"08108c08",
   717 => x"fc050cc9",
   718 => x"398c08fc",
   719 => x"0508802e",
   720 => x"80c9388c",
   721 => x"088c0508",
   722 => x"8c088805",
   723 => x"0826a138",
   724 => x"8c088805",
   725 => x"088c088c",
   726 => x"0508318c",
   727 => x"0888050c",
   728 => x"8c08f805",
   729 => x"088c08fc",
   730 => x"0508078c",
   731 => x"08f8050c",
   732 => x"8c08fc05",
   733 => x"08812a8c",
   734 => x"08fc050c",
   735 => x"8c088c05",
   736 => x"08812a8c",
   737 => x"088c050c",
   738 => x"ffaf398c",
   739 => x"08900508",
   740 => x"802e8f38",
   741 => x"8c088805",
   742 => x"08708c08",
   743 => x"f4050c51",
   744 => x"8d398c08",
   745 => x"f8050870",
   746 => x"8c08f405",
   747 => x"0c518c08",
   748 => x"f4050880",
   749 => x"0c853d0d",
   750 => x"8c0c04fd",
   751 => x"3d0d800b",
   752 => x"9ad40854",
   753 => x"5472812e",
   754 => x"983873a2",
   755 => x"940cf18f",
   756 => x"3ff0ad3f",
   757 => x"9aec5281",
   758 => x"51f7aa3f",
   759 => x"8008519e",
   760 => x"3f72a294",
   761 => x"0cf0f83f",
   762 => x"f0963f9a",
   763 => x"ec528151",
   764 => x"f7933f80",
   765 => x"0851873f",
   766 => x"00ff3900",
   767 => x"ff39f73d",
   768 => x"0d7b9af0",
   769 => x"0882c811",
   770 => x"085a545a",
   771 => x"77802e80",
   772 => x"d9388188",
   773 => x"18841908",
   774 => x"ff058171",
   775 => x"2b595559",
   776 => x"80742480",
   777 => x"e9388074",
   778 => x"24b53873",
   779 => x"822b7811",
   780 => x"88055656",
   781 => x"81801908",
   782 => x"77065372",
   783 => x"802eb538",
   784 => x"78167008",
   785 => x"53537951",
   786 => x"74085372",
   787 => x"2dff14fc",
   788 => x"17fc1779",
   789 => x"812c5a57",
   790 => x"57547380",
   791 => x"25d63877",
   792 => x"085877ff",
   793 => x"ad389af0",
   794 => x"0853bc13",
   795 => x"08a53879",
   796 => x"51ff853f",
   797 => x"74085372",
   798 => x"2dff14fc",
   799 => x"17fc1779",
   800 => x"812c5a57",
   801 => x"57547380",
   802 => x"25ffa938",
   803 => x"d2398057",
   804 => x"ff943972",
   805 => x"51bc1308",
   806 => x"53722d79",
   807 => x"51fed93f",
   808 => x"ff3d0da1",
   809 => x"f40bfc05",
   810 => x"70085252",
   811 => x"70ff2e91",
   812 => x"38702dfc",
   813 => x"12700852",
   814 => x"5270ff2e",
   815 => x"098106f1",
   816 => x"38833d0d",
   817 => x"0404effc",
   818 => x"3f040000",
   819 => x"00000040",
   820 => x"0a0a0000",
   821 => x"536f432c",
   822 => x"205a5055",
   823 => x"20746573",
   824 => x"74207072",
   825 => x"6f677261",
   826 => x"6d200000",
   827 => x"286f6e20",
   828 => x"73696d75",
   829 => x"6c61746f",
   830 => x"72290a00",
   831 => x"636f6d70",
   832 => x"696c6564",
   833 => x"3a204175",
   834 => x"67202035",
   835 => x"20323031",
   836 => x"30202020",
   837 => x"31343a31",
   838 => x"343a3337",
   839 => x"0a000000",
   840 => x"286f6e20",
   841 => x"68617264",
   842 => x"77617265",
   843 => x"290a0000",
   844 => x"64756d6d",
   845 => x"792e6578",
   846 => x"65000000",
   847 => x"43000000",
   848 => x"00ffffff",
   849 => x"ff00ffff",
   850 => x"ffff00ff",
   851 => x"ffffff00",
   852 => x"00000000",
   853 => x"00000000",
   854 => x"00000000",
   855 => x"000010fc",
   856 => x"80000800",
   857 => x"80000200",
   858 => x"80000100",
   859 => x"00000d30",
   860 => x"00000d74",
   861 => x"00000000",
   862 => x"00000fdc",
   863 => x"00001038",
   864 => x"00001094",
   865 => x"00000000",
   866 => x"00000000",
   867 => x"00000000",
   868 => x"00000000",
   869 => x"00000000",
   870 => x"00000000",
   871 => x"00000000",
   872 => x"00000000",
   873 => x"00000000",
   874 => x"00000d3c",
   875 => x"00000000",
   876 => x"00000000",
   877 => x"00000000",
   878 => x"00000000",
   879 => x"00000000",
   880 => x"00000000",
   881 => x"00000000",
   882 => x"00000000",
   883 => x"00000000",
   884 => x"00000000",
   885 => x"00000000",
   886 => x"00000000",
   887 => x"00000000",
   888 => x"00000000",
   889 => x"00000000",
   890 => x"00000000",
   891 => x"00000000",
   892 => x"00000000",
   893 => x"00000000",
   894 => x"00000000",
   895 => x"00000000",
   896 => x"00000000",
   897 => x"00000000",
   898 => x"00000000",
   899 => x"00000000",
   900 => x"00000000",
   901 => x"00000000",
   902 => x"00000000",
   903 => x"00000001",
   904 => x"330eabcd",
   905 => x"1234e66d",
   906 => x"deec0005",
   907 => x"000b0000",
   908 => x"00000000",
   909 => x"00000000",
   910 => x"00000000",
   911 => x"00000000",
   912 => x"00000000",
   913 => x"00000000",
   914 => x"00000000",
   915 => x"00000000",
   916 => x"00000000",
   917 => x"00000000",
   918 => x"00000000",
   919 => x"00000000",
   920 => x"00000000",
   921 => x"00000000",
   922 => x"00000000",
   923 => x"00000000",
   924 => x"00000000",
   925 => x"00000000",
   926 => x"00000000",
   927 => x"00000000",
   928 => x"00000000",
   929 => x"00000000",
   930 => x"00000000",
   931 => x"00000000",
   932 => x"00000000",
   933 => x"00000000",
   934 => x"00000000",
   935 => x"00000000",
   936 => x"00000000",
   937 => x"00000000",
   938 => x"00000000",
   939 => x"00000000",
   940 => x"00000000",
   941 => x"00000000",
   942 => x"00000000",
   943 => x"00000000",
   944 => x"00000000",
   945 => x"00000000",
   946 => x"00000000",
   947 => x"00000000",
   948 => x"00000000",
   949 => x"00000000",
   950 => x"00000000",
   951 => x"00000000",
   952 => x"00000000",
   953 => x"00000000",
   954 => x"00000000",
   955 => x"00000000",
   956 => x"00000000",
   957 => x"00000000",
   958 => x"00000000",
   959 => x"00000000",
   960 => x"00000000",
   961 => x"00000000",
   962 => x"00000000",
   963 => x"00000000",
   964 => x"00000000",
   965 => x"00000000",
   966 => x"00000000",
   967 => x"00000000",
   968 => x"00000000",
   969 => x"00000000",
   970 => x"00000000",
   971 => x"00000000",
   972 => x"00000000",
   973 => x"00000000",
   974 => x"00000000",
   975 => x"00000000",
   976 => x"00000000",
   977 => x"00000000",
   978 => x"00000000",
   979 => x"00000000",
   980 => x"00000000",
   981 => x"00000000",
   982 => x"00000000",
   983 => x"00000000",
   984 => x"00000000",
   985 => x"00000000",
   986 => x"00000000",
   987 => x"00000000",
   988 => x"00000000",
   989 => x"00000000",
   990 => x"00000000",
   991 => x"00000000",
   992 => x"00000000",
   993 => x"00000000",
   994 => x"00000000",
   995 => x"00000000",
   996 => x"00000000",
   997 => x"00000000",
   998 => x"00000000",
   999 => x"00000000",
  1000 => x"00000000",
  1001 => x"00000000",
  1002 => x"00000000",
  1003 => x"00000000",
  1004 => x"00000000",
  1005 => x"00000000",
  1006 => x"00000000",
  1007 => x"00000000",
  1008 => x"00000000",
  1009 => x"00000000",
  1010 => x"00000000",
  1011 => x"00000000",
  1012 => x"00000000",
  1013 => x"00000000",
  1014 => x"00000000",
  1015 => x"00000000",
  1016 => x"00000000",
  1017 => x"00000000",
  1018 => x"00000000",
  1019 => x"00000000",
  1020 => x"00000000",
  1021 => x"00000000",
  1022 => x"00000000",
  1023 => x"00000000",
  1024 => x"00000000",
  1025 => x"00000000",
  1026 => x"00000000",
  1027 => x"00000000",
  1028 => x"00000000",
  1029 => x"00000000",
  1030 => x"00000000",
  1031 => x"00000000",
  1032 => x"00000000",
  1033 => x"00000000",
  1034 => x"00000000",
  1035 => x"00000000",
  1036 => x"00000000",
  1037 => x"00000000",
  1038 => x"00000000",
  1039 => x"00000000",
  1040 => x"00000000",
  1041 => x"00000000",
  1042 => x"00000000",
  1043 => x"00000000",
  1044 => x"00000000",
  1045 => x"00000000",
  1046 => x"00000000",
  1047 => x"00000000",
  1048 => x"00000000",
  1049 => x"00000000",
  1050 => x"00000000",
  1051 => x"00000000",
  1052 => x"00000000",
  1053 => x"00000000",
  1054 => x"00000000",
  1055 => x"00000000",
  1056 => x"00000000",
  1057 => x"00000000",
  1058 => x"00000000",
  1059 => x"00000000",
  1060 => x"00000000",
  1061 => x"00000000",
  1062 => x"00000000",
  1063 => x"00000000",
  1064 => x"00000000",
  1065 => x"00000000",
  1066 => x"00000000",
  1067 => x"00000000",
  1068 => x"00000000",
  1069 => x"00000000",
  1070 => x"00000000",
  1071 => x"00000000",
  1072 => x"00000000",
  1073 => x"00000000",
  1074 => x"00000000",
  1075 => x"00000000",
  1076 => x"00000000",
  1077 => x"00000000",
  1078 => x"00000000",
  1079 => x"00000000",
  1080 => x"00000000",
  1081 => x"00000000",
  1082 => x"00000000",
  1083 => x"00000000",
  1084 => x"ffffffff",
  1085 => x"00000000",
  1086 => x"ffffffff",
  1087 => x"00000000",
  1088 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
