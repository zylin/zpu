------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2003 - 2008, Gaisler Research
--  Copyright (C) 2008 - 2010, Aeroflex Gaisler
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 
-----------------------------------------------------------------------------
-- Entity:      charrom
-- File:        charrom.vhd
-- Author:      Marcus Hellqvist
-- Description: Character ROM for video controller
-----------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;
library grlib;
use grlib.stdlib.all;

entity charrom is
  port(
    clk         : in std_ulogic;
    addr        : in std_logic_vector(11 downto 0);
    data        : out std_logic_vector(7 downto 0)
    );
end entity;

architecture rtl of charrom is

    type rom_t is array (0 to 2**12-1) of std_logic_vector (data'range);

    signal rom : rom_t:= 
    (
        16#000# => X"00", -- 
        16#100# => X"00", -- 
        16#200# => X"00", -- 
        16#300# => X"00", -- 
        16#400# => X"00", -- 
        16#500# => X"00", -- 
        16#600# => X"00", -- 
        16#700# => X"00", -- 
        16#800# => X"00", -- 
        16#900# => X"00", -- 
        16#a00# => X"00", -- 
        16#b00# => X"00", -- 
        16#c00# => X"00", -- 
        16#020# => X"00", --  
        16#120# => X"00", --  
        16#220# => X"00", --  
        16#320# => X"00", --  
        16#420# => X"00", --  
        16#520# => X"00", --  
        16#620# => X"00", --  
        16#720# => X"00", --  
        16#820# => X"00", --  
        16#920# => X"00", --  
        16#a20# => X"00", --  
        16#b20# => X"00", --  
        16#c20# => X"00", --  
        16#021# => X"00", -- !
        16#121# => X"00", -- !
        16#221# => X"10", -- !
        16#321# => X"10", -- !
        16#421# => X"10", -- !
        16#521# => X"10", -- !
        16#621# => X"10", -- !
        16#721# => X"10", -- !
        16#821# => X"10", -- !
        16#921# => X"00", -- !
        16#a21# => X"10", -- !
        16#b21# => X"00", -- !
        16#c21# => X"00", -- !
        16#022# => X"00", -- "
        16#122# => X"00", -- "
        16#222# => X"24", -- "
        16#322# => X"24", -- "
        16#422# => X"24", -- "
        16#522# => X"00", -- "
        16#622# => X"00", -- "
        16#722# => X"00", -- "
        16#822# => X"00", -- "
        16#922# => X"00", -- "
        16#a22# => X"00", -- "
        16#b22# => X"00", -- "
        16#c22# => X"00", -- "
        16#023# => X"00", -- #
        16#123# => X"00", -- #
        16#223# => X"00", -- #
        16#323# => X"24", -- #
        16#423# => X"24", -- #
        16#523# => X"7e", -- #
        16#623# => X"24", -- #
        16#723# => X"7e", -- #
        16#823# => X"24", -- #
        16#923# => X"24", -- #
        16#a23# => X"00", -- #
        16#b23# => X"00", -- #
        16#c23# => X"00", -- #
        16#024# => X"00", -- $
        16#124# => X"00", -- $
        16#224# => X"10", -- $
        16#324# => X"3c", -- $
        16#424# => X"50", -- $
        16#524# => X"50", -- $
        16#624# => X"38", -- $
        16#724# => X"14", -- $
        16#824# => X"14", -- $
        16#924# => X"78", -- $
        16#a24# => X"10", -- $
        16#b24# => X"00", -- $
        16#c24# => X"00", -- $
        16#025# => X"00", -- %
        16#125# => X"00", -- %
        16#225# => X"22", -- %
        16#325# => X"52", -- %
        16#425# => X"24", -- %
        16#525# => X"08", -- %
        16#625# => X"08", -- %
        16#725# => X"10", -- %
        16#825# => X"24", -- %
        16#925# => X"2a", -- %
        16#a25# => X"44", -- %
        16#b25# => X"00", -- %
        16#c25# => X"00", -- %
        16#026# => X"00", -- &
        16#126# => X"00", -- &
        16#226# => X"00", -- &
        16#326# => X"00", -- &
        16#426# => X"30", -- &
        16#526# => X"48", -- &
        16#626# => X"48", -- &
        16#726# => X"30", -- &
        16#826# => X"4a", -- &
        16#926# => X"44", -- &
        16#a26# => X"3a", -- &
        16#b26# => X"00", -- &
        16#c26# => X"00", -- &
        16#027# => X"00", -- '
        16#127# => X"00", -- '
        16#227# => X"10", -- '
        16#327# => X"10", -- '
        16#427# => X"10", -- '
        16#527# => X"00", -- '
        16#627# => X"00", -- '
        16#727# => X"00", -- '
        16#827# => X"00", -- '
        16#927# => X"00", -- '
        16#a27# => X"00", -- '
        16#b27# => X"00", -- '
        16#c27# => X"00", -- '
        16#028# => X"00", -- (
        16#128# => X"00", -- (
        16#228# => X"04", -- (
        16#328# => X"08", -- (
        16#428# => X"08", -- (
        16#528# => X"10", -- (
        16#628# => X"10", -- (
        16#728# => X"10", -- (
        16#828# => X"08", -- (
        16#928# => X"08", -- (
        16#a28# => X"04", -- (
        16#b28# => X"00", -- (
        16#c28# => X"00", -- (
        16#029# => X"00", -- )
        16#129# => X"00", -- )
        16#229# => X"20", -- )
        16#329# => X"10", -- )
        16#429# => X"10", -- )
        16#529# => X"08", -- )
        16#629# => X"08", -- )
        16#729# => X"08", -- )
        16#829# => X"10", -- )
        16#929# => X"10", -- )
        16#a29# => X"20", -- )
        16#b29# => X"00", -- )
        16#c29# => X"00", -- )
        16#02a# => X"00", -- *
        16#12a# => X"00", -- *
        16#22a# => X"24", -- *
        16#32a# => X"18", -- *
        16#42a# => X"7e", -- *
        16#52a# => X"18", -- *
        16#62a# => X"24", -- *
        16#72a# => X"00", -- *
        16#82a# => X"00", -- *
        16#92a# => X"00", -- *
        16#a2a# => X"00", -- *
        16#b2a# => X"00", -- *
        16#c2a# => X"00", -- *
        16#02b# => X"00", -- +
        16#12b# => X"00", -- +
        16#22b# => X"00", -- +
        16#32b# => X"00", -- +
        16#42b# => X"10", -- +
        16#52b# => X"10", -- +
        16#62b# => X"7c", -- +
        16#72b# => X"10", -- +
        16#82b# => X"10", -- +
        16#92b# => X"00", -- +
        16#a2b# => X"00", -- +
        16#b2b# => X"00", -- +
        16#c2b# => X"00", -- +
        16#02c# => X"00", -- ,
        16#12c# => X"00", -- ,
        16#22c# => X"00", -- ,
        16#32c# => X"00", -- ,
        16#42c# => X"00", -- ,
        16#52c# => X"00", -- ,
        16#62c# => X"00", -- ,
        16#72c# => X"00", -- ,
        16#82c# => X"00", -- ,
        16#92c# => X"38", -- ,
        16#a2c# => X"30", -- ,
        16#b2c# => X"40", -- ,
        16#c2c# => X"00", -- ,
        16#02d# => X"00", -- -
        16#12d# => X"00", -- -
        16#22d# => X"00", -- -
        16#32d# => X"00", -- -
        16#42d# => X"00", -- -
        16#52d# => X"00", -- -
        16#62d# => X"7c", -- -
        16#72d# => X"00", -- -
        16#82d# => X"00", -- -
        16#92d# => X"00", -- -
        16#a2d# => X"00", -- -
        16#b2d# => X"00", -- -
        16#c2d# => X"00", -- -
        16#02e# => X"00", -- .
        16#12e# => X"00", -- .
        16#22e# => X"00", -- .
        16#32e# => X"00", -- .
        16#42e# => X"00", -- .
        16#52e# => X"00", -- .
        16#62e# => X"00", -- .
        16#72e# => X"00", -- .
        16#82e# => X"00", -- .
        16#92e# => X"10", -- .
        16#a2e# => X"38", -- .
        16#b2e# => X"10", -- .
        16#c2e# => X"00", -- .
        16#02f# => X"00", -- /
        16#12f# => X"00", -- /
        16#22f# => X"02", -- /
        16#32f# => X"02", -- /
        16#42f# => X"04", -- /
        16#52f# => X"08", -- /
        16#62f# => X"10", -- /
        16#72f# => X"20", -- /
        16#82f# => X"40", -- /
        16#92f# => X"80", -- /
        16#a2f# => X"80", -- /
        16#b2f# => X"00", -- /
        16#c2f# => X"00", -- /
        16#030# => X"00", -- 0
        16#130# => X"00", -- 0
        16#230# => X"18", -- 0
        16#330# => X"24", -- 0
        16#430# => X"42", -- 0
        16#530# => X"42", -- 0
        16#630# => X"42", -- 0
        16#730# => X"42", -- 0
        16#830# => X"42", -- 0
        16#930# => X"24", -- 0
        16#a30# => X"18", -- 0
        16#b30# => X"00", -- 0
        16#c30# => X"00", -- 0
        16#031# => X"00", -- 1
        16#131# => X"00", -- 1
        16#231# => X"10", -- 1
        16#331# => X"30", -- 1
        16#431# => X"50", -- 1
        16#531# => X"10", -- 1
        16#631# => X"10", -- 1
        16#731# => X"10", -- 1
        16#831# => X"10", -- 1
        16#931# => X"10", -- 1
        16#a31# => X"7c", -- 1
        16#b31# => X"00", -- 1
        16#c31# => X"00", -- 1
        16#032# => X"00", -- 2
        16#132# => X"00", -- 2
        16#232# => X"3c", -- 2
        16#332# => X"42", -- 2
        16#432# => X"42", -- 2
        16#532# => X"02", -- 2
        16#632# => X"04", -- 2
        16#732# => X"18", -- 2
        16#832# => X"20", -- 2
        16#932# => X"40", -- 2
        16#a32# => X"7e", -- 2
        16#b32# => X"00", -- 2
        16#c32# => X"00", -- 2
        16#033# => X"00", -- 3
        16#133# => X"00", -- 3
        16#233# => X"7e", -- 3
        16#333# => X"02", -- 3
        16#433# => X"04", -- 3
        16#533# => X"08", -- 3
        16#633# => X"1c", -- 3
        16#733# => X"02", -- 3
        16#833# => X"02", -- 3
        16#933# => X"42", -- 3
        16#a33# => X"3c", -- 3
        16#b33# => X"00", -- 3
        16#c33# => X"00", -- 3
        16#034# => X"00", -- 4
        16#134# => X"00", -- 4
        16#234# => X"04", -- 4
        16#334# => X"0c", -- 4
        16#434# => X"14", -- 4
        16#534# => X"24", -- 4
        16#634# => X"44", -- 4
        16#734# => X"44", -- 4
        16#834# => X"7e", -- 4
        16#934# => X"04", -- 4
        16#a34# => X"04", -- 4
        16#b34# => X"00", -- 4
        16#c34# => X"00", -- 4
        16#035# => X"00", -- 5
        16#135# => X"00", -- 5
        16#235# => X"7e", -- 5
        16#335# => X"40", -- 5
        16#435# => X"40", -- 5
        16#535# => X"5c", -- 5
        16#635# => X"62", -- 5
        16#735# => X"02", -- 5
        16#835# => X"02", -- 5
        16#935# => X"42", -- 5
        16#a35# => X"3c", -- 5
        16#b35# => X"00", -- 5
        16#c35# => X"00", -- 5
        16#036# => X"00", -- 6
        16#136# => X"00", -- 6
        16#236# => X"1c", -- 6
        16#336# => X"20", -- 6
        16#436# => X"40", -- 6
        16#536# => X"40", -- 6
        16#636# => X"5c", -- 6
        16#736# => X"62", -- 6
        16#836# => X"42", -- 6
        16#936# => X"42", -- 6
        16#a36# => X"3c", -- 6
        16#b36# => X"00", -- 6
        16#c36# => X"00", -- 6
        16#037# => X"00", -- 7
        16#137# => X"00", -- 7
        16#237# => X"7e", -- 7
        16#337# => X"02", -- 7
        16#437# => X"04", -- 7
        16#537# => X"08", -- 7
        16#637# => X"08", -- 7
        16#737# => X"10", -- 7
        16#837# => X"10", -- 7
        16#937# => X"20", -- 7
        16#a37# => X"20", -- 7
        16#b37# => X"00", -- 7
        16#c37# => X"00", -- 7
        16#038# => X"00", -- 8
        16#138# => X"00", -- 8
        16#238# => X"3c", -- 8
        16#338# => X"42", -- 8
        16#438# => X"42", -- 8
        16#538# => X"42", -- 8
        16#638# => X"3c", -- 8
        16#738# => X"42", -- 8
        16#838# => X"42", -- 8
        16#938# => X"42", -- 8
        16#a38# => X"3c", -- 8
        16#b38# => X"00", -- 8
        16#c38# => X"00", -- 8
        16#039# => X"00", -- 9
        16#139# => X"00", -- 9
        16#239# => X"3c", -- 9
        16#339# => X"42", -- 9
        16#439# => X"42", -- 9
        16#539# => X"46", -- 9
        16#639# => X"3a", -- 9
        16#739# => X"02", -- 9
        16#839# => X"02", -- 9
        16#939# => X"04", -- 9
        16#a39# => X"38", -- 9
        16#b39# => X"00", -- 9
        16#c39# => X"00", -- 9
        16#03a# => X"00", -- :
        16#13a# => X"00", -- :
        16#23a# => X"00", -- :
        16#33a# => X"00", -- :
        16#43a# => X"10", -- :
        16#53a# => X"38", -- :
        16#63a# => X"10", -- :
        16#73a# => X"00", -- :
        16#83a# => X"00", -- :
        16#93a# => X"10", -- :
        16#a3a# => X"38", -- :
        16#b3a# => X"10", -- :
        16#c3a# => X"00", -- :
        16#03b# => X"00", -- ;
        16#13b# => X"00", -- ;
        16#23b# => X"00", -- ;
        16#33b# => X"00", -- ;
        16#43b# => X"10", -- ;
        16#53b# => X"38", -- ;
        16#63b# => X"10", -- ;
        16#73b# => X"00", -- ;
        16#83b# => X"00", -- ;
        16#93b# => X"38", -- ;
        16#a3b# => X"30", -- ;
        16#b3b# => X"40", -- ;
        16#c3b# => X"00", -- ;
        16#03c# => X"00", -- <
        16#13c# => X"00", -- <
        16#23c# => X"02", -- <
        16#33c# => X"04", -- <
        16#43c# => X"08", -- <
        16#53c# => X"10", -- <
        16#63c# => X"20", -- <
        16#73c# => X"10", -- <
        16#83c# => X"08", -- <
        16#93c# => X"04", -- <
        16#a3c# => X"02", -- <
        16#b3c# => X"00", -- <
        16#c3c# => X"00", -- <
        16#03d# => X"00", -- =
        16#13d# => X"00", -- =
        16#23d# => X"00", -- =
        16#33d# => X"00", -- =
        16#43d# => X"00", -- =
        16#53d# => X"7e", -- =
        16#63d# => X"00", -- =
        16#73d# => X"00", -- =
        16#83d# => X"7e", -- =
        16#93d# => X"00", -- =
        16#a3d# => X"00", -- =
        16#b3d# => X"00", -- =
        16#c3d# => X"00", -- =
        16#03e# => X"00", -- >
        16#13e# => X"00", -- >
        16#23e# => X"40", -- >
        16#33e# => X"20", -- >
        16#43e# => X"10", -- >
        16#53e# => X"08", -- >
        16#63e# => X"04", -- >
        16#73e# => X"08", -- >
        16#83e# => X"10", -- >
        16#93e# => X"20", -- >
        16#a3e# => X"40", -- >
        16#b3e# => X"00", -- >
        16#c3e# => X"00", -- >
        16#03f# => X"00", -- ?
        16#13f# => X"00", -- ?
        16#23f# => X"3c", -- ?
        16#33f# => X"42", -- ?
        16#43f# => X"42", -- ?
        16#53f# => X"02", -- ?
        16#63f# => X"04", -- ?
        16#73f# => X"08", -- ?
        16#83f# => X"08", -- ?
        16#93f# => X"00", -- ?
        16#a3f# => X"08", -- ?
        16#b3f# => X"00", -- ?
        16#c3f# => X"00", -- ?
        16#040# => X"00", -- @
        16#140# => X"00", -- @
        16#240# => X"3c", -- @
        16#340# => X"42", -- @
        16#440# => X"42", -- @
        16#540# => X"4e", -- @
        16#640# => X"52", -- @
        16#740# => X"56", -- @
        16#840# => X"4a", -- @
        16#940# => X"40", -- @
        16#a40# => X"3c", -- @
        16#b40# => X"00", -- @
        16#c40# => X"00", -- @
        16#041# => X"00", -- A
        16#141# => X"00", -- A
        16#241# => X"18", -- A
        16#341# => X"24", -- A
        16#441# => X"42", -- A
        16#541# => X"42", -- A
        16#641# => X"42", -- A
        16#741# => X"7e", -- A
        16#841# => X"42", -- A
        16#941# => X"42", -- A
        16#a41# => X"42", -- A
        16#b41# => X"00", -- A
        16#c41# => X"00", -- A
        16#042# => X"00", -- B
        16#142# => X"00", -- B
        16#242# => X"78", -- B
        16#342# => X"44", -- B
        16#442# => X"42", -- B
        16#542# => X"44", -- B
        16#642# => X"78", -- B
        16#742# => X"44", -- B
        16#842# => X"42", -- B
        16#942# => X"44", -- B
        16#a42# => X"78", -- B
        16#b42# => X"00", -- B
        16#c42# => X"00", -- B
        16#043# => X"00", -- C
        16#143# => X"00", -- C
        16#243# => X"3c", -- C
        16#343# => X"42", -- C
        16#443# => X"40", -- C
        16#543# => X"40", -- C
        16#643# => X"40", -- C
        16#743# => X"40", -- C
        16#843# => X"40", -- C
        16#943# => X"42", -- C
        16#a43# => X"3c", -- C
        16#b43# => X"00", -- C
        16#c43# => X"00", -- C
        16#044# => X"00", -- D
        16#144# => X"00", -- D
        16#244# => X"78", -- D
        16#344# => X"44", -- D
        16#444# => X"42", -- D
        16#544# => X"42", -- D
        16#644# => X"42", -- D
        16#744# => X"42", -- D
        16#844# => X"42", -- D
        16#944# => X"44", -- D
        16#a44# => X"78", -- D
        16#b44# => X"00", -- D
        16#c44# => X"00", -- D
        16#045# => X"00", -- E
        16#145# => X"00", -- E
        16#245# => X"7e", -- E
        16#345# => X"40", -- E
        16#445# => X"40", -- E
        16#545# => X"40", -- E
        16#645# => X"78", -- E
        16#745# => X"40", -- E
        16#845# => X"40", -- E
        16#945# => X"40", -- E
        16#a45# => X"7e", -- E
        16#b45# => X"00", -- E
        16#c45# => X"00", -- E
        16#046# => X"00", -- F
        16#146# => X"00", -- F
        16#246# => X"7e", -- F
        16#346# => X"40", -- F
        16#446# => X"40", -- F
        16#546# => X"40", -- F
        16#646# => X"78", -- F
        16#746# => X"40", -- F
        16#846# => X"40", -- F
        16#946# => X"40", -- F
        16#a46# => X"40", -- F
        16#b46# => X"00", -- F
        16#c46# => X"00", -- F
        16#047# => X"00", -- G
        16#147# => X"00", -- G
        16#247# => X"3c", -- G
        16#347# => X"42", -- G
        16#447# => X"40", -- G
        16#547# => X"40", -- G
        16#647# => X"40", -- G
        16#747# => X"4e", -- G
        16#847# => X"42", -- G
        16#947# => X"46", -- G
        16#a47# => X"3a", -- G
        16#b47# => X"00", -- G
        16#c47# => X"00", -- G
        16#048# => X"00", -- H
        16#148# => X"00", -- H
        16#248# => X"42", -- H
        16#348# => X"42", -- H
        16#448# => X"42", -- H
        16#548# => X"42", -- H
        16#648# => X"7e", -- H
        16#748# => X"42", -- H
        16#848# => X"42", -- H
        16#948# => X"42", -- H
        16#a48# => X"42", -- H
        16#b48# => X"00", -- H
        16#c48# => X"00", -- H
        16#049# => X"00", -- I
        16#149# => X"00", -- I
        16#249# => X"7c", -- I
        16#349# => X"10", -- I
        16#449# => X"10", -- I
        16#549# => X"10", -- I
        16#649# => X"10", -- I
        16#749# => X"10", -- I
        16#849# => X"10", -- I
        16#949# => X"10", -- I
        16#a49# => X"7c", -- I
        16#b49# => X"00", -- I
        16#c49# => X"00", -- I
        16#04a# => X"00", -- J
        16#14a# => X"00", -- J
        16#24a# => X"1f", -- J
        16#34a# => X"04", -- J
        16#44a# => X"04", -- J
        16#54a# => X"04", -- J
        16#64a# => X"04", -- J
        16#74a# => X"04", -- J
        16#84a# => X"04", -- J
        16#94a# => X"44", -- J
        16#a4a# => X"38", -- J
        16#b4a# => X"00", -- J
        16#c4a# => X"00", -- J
        16#04b# => X"00", -- K
        16#14b# => X"00", -- K
        16#24b# => X"42", -- K
        16#34b# => X"44", -- K
        16#44b# => X"48", -- K
        16#54b# => X"50", -- K
        16#64b# => X"60", -- K
        16#74b# => X"50", -- K
        16#84b# => X"48", -- K
        16#94b# => X"44", -- K
        16#a4b# => X"42", -- K
        16#b4b# => X"00", -- K
        16#c4b# => X"00", -- K
        16#04c# => X"00", -- L
        16#14c# => X"00", -- L
        16#24c# => X"40", -- L
        16#34c# => X"40", -- L
        16#44c# => X"40", -- L
        16#54c# => X"40", -- L
        16#64c# => X"40", -- L
        16#74c# => X"40", -- L
        16#84c# => X"40", -- L
        16#94c# => X"40", -- L
        16#a4c# => X"7e", -- L
        16#b4c# => X"00", -- L
        16#c4c# => X"00", -- L
        16#04d# => X"00", -- M
        16#14d# => X"00", -- M
        16#24d# => X"82", -- M
        16#34d# => X"82", -- M
        16#44d# => X"c6", -- M
        16#54d# => X"aa", -- M
        16#64d# => X"92", -- M
        16#74d# => X"92", -- M
        16#84d# => X"82", -- M
        16#94d# => X"82", -- M
        16#a4d# => X"82", -- M
        16#b4d# => X"00", -- M
        16#c4d# => X"00", -- M
        16#04e# => X"00", -- N
        16#14e# => X"00", -- N
        16#24e# => X"42", -- N
        16#34e# => X"42", -- N
        16#44e# => X"62", -- N
        16#54e# => X"52", -- N
        16#64e# => X"4a", -- N
        16#74e# => X"46", -- N
        16#84e# => X"42", -- N
        16#94e# => X"42", -- N
        16#a4e# => X"42", -- N
        16#b4e# => X"00", -- N
        16#c4e# => X"00", -- N
        16#04f# => X"00", -- O
        16#14f# => X"00", -- O
        16#24f# => X"3c", -- O
        16#34f# => X"42", -- O
        16#44f# => X"42", -- O
        16#54f# => X"42", -- O
        16#64f# => X"42", -- O
        16#74f# => X"42", -- O
        16#84f# => X"42", -- O
        16#94f# => X"42", -- O
        16#a4f# => X"3c", -- O
        16#b4f# => X"00", -- O
        16#c4f# => X"00", -- O
        16#050# => X"00", -- P
        16#150# => X"00", -- P
        16#250# => X"7c", -- P
        16#350# => X"42", -- P
        16#450# => X"42", -- P
        16#550# => X"42", -- P
        16#650# => X"7c", -- P
        16#750# => X"40", -- P
        16#850# => X"40", -- P
        16#950# => X"40", -- P
        16#a50# => X"40", -- P
        16#b50# => X"00", -- P
        16#c50# => X"00", -- P
        16#051# => X"00", -- Q
        16#151# => X"00", -- Q
        16#251# => X"3c", -- Q
        16#351# => X"42", -- Q
        16#451# => X"42", -- Q
        16#551# => X"42", -- Q
        16#651# => X"42", -- Q
        16#751# => X"42", -- Q
        16#851# => X"52", -- Q
        16#951# => X"4a", -- Q
        16#a51# => X"3c", -- Q
        16#b51# => X"02", -- Q
        16#c51# => X"00", -- Q
        16#052# => X"00", -- R
        16#152# => X"00", -- R
        16#252# => X"7c", -- R
        16#352# => X"42", -- R
        16#452# => X"42", -- R
        16#552# => X"42", -- R
        16#652# => X"7c", -- R
        16#752# => X"50", -- R
        16#852# => X"48", -- R
        16#952# => X"44", -- R
        16#a52# => X"42", -- R
        16#b52# => X"00", -- R
        16#c52# => X"00", -- R
        16#053# => X"00", -- S
        16#153# => X"00", -- S
        16#253# => X"3c", -- S
        16#353# => X"42", -- S
        16#453# => X"40", -- S
        16#553# => X"40", -- S
        16#653# => X"3c", -- S
        16#753# => X"02", -- S
        16#853# => X"02", -- S
        16#953# => X"42", -- S
        16#a53# => X"3c", -- S
        16#b53# => X"00", -- S
        16#c53# => X"00", -- S
        16#054# => X"00", -- T
        16#154# => X"00", -- T
        16#254# => X"fe", -- T
        16#354# => X"10", -- T
        16#454# => X"10", -- T
        16#554# => X"10", -- T
        16#654# => X"10", -- T
        16#754# => X"10", -- T
        16#854# => X"10", -- T
        16#954# => X"10", -- T
        16#a54# => X"10", -- T
        16#b54# => X"00", -- T
        16#c54# => X"00", -- T
        16#055# => X"00", -- U
        16#155# => X"00", -- U
        16#255# => X"42", -- U
        16#355# => X"42", -- U
        16#455# => X"42", -- U
        16#555# => X"42", -- U
        16#655# => X"42", -- U
        16#755# => X"42", -- U
        16#855# => X"42", -- U
        16#955# => X"42", -- U
        16#a55# => X"3c", -- U
        16#b55# => X"00", -- U
        16#c55# => X"00", -- U
        16#056# => X"00", -- V
        16#156# => X"00", -- V
        16#256# => X"82", -- V
        16#356# => X"82", -- V
        16#456# => X"44", -- V
        16#556# => X"44", -- V
        16#656# => X"44", -- V
        16#756# => X"28", -- V
        16#856# => X"28", -- V
        16#956# => X"28", -- V
        16#a56# => X"10", -- V
        16#b56# => X"00", -- V
        16#c56# => X"00", -- V
        16#057# => X"00", -- W
        16#157# => X"00", -- W
        16#257# => X"82", -- W
        16#357# => X"82", -- W
        16#457# => X"82", -- W
        16#557# => X"82", -- W
        16#657# => X"92", -- W
        16#757# => X"92", -- W
        16#857# => X"92", -- W
        16#957# => X"aa", -- W
        16#a57# => X"44", -- W
        16#b57# => X"00", -- W
        16#c57# => X"00", -- W
        16#058# => X"00", -- X
        16#158# => X"00", -- X
        16#258# => X"82", -- X
        16#358# => X"82", -- X
        16#458# => X"44", -- X
        16#558# => X"28", -- X
        16#658# => X"10", -- X
        16#758# => X"28", -- X
        16#858# => X"44", -- X
        16#958# => X"82", -- X
        16#a58# => X"82", -- X
        16#b58# => X"00", -- X
        16#c58# => X"00", -- X
        16#059# => X"00", -- Y
        16#159# => X"00", -- Y
        16#259# => X"82", -- Y
        16#359# => X"82", -- Y
        16#459# => X"44", -- Y
        16#559# => X"28", -- Y
        16#659# => X"10", -- Y
        16#759# => X"10", -- Y
        16#859# => X"10", -- Y
        16#959# => X"10", -- Y
        16#a59# => X"10", -- Y
        16#b59# => X"00", -- Y
        16#c59# => X"00", -- Y
        16#05a# => X"00", -- Z
        16#15a# => X"00", -- Z
        16#25a# => X"7e", -- Z
        16#35a# => X"02", -- Z
        16#45a# => X"04", -- Z
        16#55a# => X"08", -- Z
        16#65a# => X"10", -- Z
        16#75a# => X"20", -- Z
        16#85a# => X"40", -- Z
        16#95a# => X"40", -- Z
        16#a5a# => X"7e", -- Z
        16#b5a# => X"00", -- Z
        16#c5a# => X"00", -- Z
        16#05b# => X"00", -- [
        16#15b# => X"00", -- [
        16#25b# => X"3c", -- [
        16#35b# => X"20", -- [
        16#45b# => X"20", -- [
        16#55b# => X"20", -- [
        16#65b# => X"20", -- [
        16#75b# => X"20", -- [
        16#85b# => X"20", -- [
        16#95b# => X"20", -- [
        16#a5b# => X"3c", -- [
        16#b5b# => X"00", -- [
        16#c5b# => X"00", -- [
        16#05c# => X"00", -- \
        16#15c# => X"00", -- \
        16#25c# => X"80", -- \
        16#35c# => X"80", -- \
        16#45c# => X"40", -- \
        16#55c# => X"20", -- \
        16#65c# => X"10", -- \
        16#75c# => X"08", -- \
        16#85c# => X"04", -- \
        16#95c# => X"02", -- \
        16#a5c# => X"02", -- \
        16#b5c# => X"00", -- \
        16#c5c# => X"00", -- \
        16#05d# => X"00", -- ]
        16#15d# => X"00", -- ]
        16#25d# => X"78", -- ]
        16#35d# => X"08", -- ]
        16#45d# => X"08", -- ]
        16#55d# => X"08", -- ]
        16#65d# => X"08", -- ]
        16#75d# => X"08", -- ]
        16#85d# => X"08", -- ]
        16#95d# => X"08", -- ]
        16#a5d# => X"78", -- ]
        16#b5d# => X"00", -- ]
        16#c5d# => X"00", -- ]
        16#05e# => X"00", -- ^
        16#15e# => X"00", -- ^
        16#25e# => X"10", -- ^
        16#35e# => X"28", -- ^
        16#45e# => X"44", -- ^
        16#55e# => X"00", -- ^
        16#65e# => X"00", -- ^
        16#75e# => X"00", -- ^
        16#85e# => X"00", -- ^
        16#95e# => X"00", -- ^
        16#a5e# => X"00", -- ^
        16#b5e# => X"00", -- ^
        16#c5e# => X"00", -- ^
        16#05f# => X"00", -- _
        16#15f# => X"00", -- _
        16#25f# => X"00", -- _
        16#35f# => X"00", -- _
        16#45f# => X"00", -- _
        16#55f# => X"00", -- _
        16#65f# => X"00", -- _
        16#75f# => X"00", -- _
        16#85f# => X"00", -- _
        16#95f# => X"00", -- _
        16#a5f# => X"00", -- _
        16#b5f# => X"fe", -- _
        16#c5f# => X"00", -- _
        16#060# => X"00", -- `
        16#160# => X"10", -- `
        16#260# => X"08", -- `
        16#360# => X"00", -- `
        16#460# => X"00", -- `
        16#560# => X"00", -- `
        16#660# => X"00", -- `
        16#760# => X"00", -- `
        16#860# => X"00", -- `
        16#960# => X"00", -- `
        16#a60# => X"00", -- `
        16#b60# => X"00", -- `
        16#c60# => X"00", -- `
        16#061# => X"00", -- a
        16#161# => X"00", -- a
        16#261# => X"00", -- a
        16#361# => X"00", -- a
        16#461# => X"00", -- a
        16#561# => X"3c", -- a
        16#661# => X"02", -- a
        16#761# => X"3e", -- a
        16#861# => X"42", -- a
        16#961# => X"46", -- a
        16#a61# => X"3a", -- a
        16#b61# => X"00", -- a
        16#c61# => X"00", -- a
        16#062# => X"00", -- b
        16#162# => X"00", -- b
        16#262# => X"40", -- b
        16#362# => X"40", -- b
        16#462# => X"40", -- b
        16#562# => X"5c", -- b
        16#662# => X"62", -- b
        16#762# => X"42", -- b
        16#862# => X"42", -- b
        16#962# => X"62", -- b
        16#a62# => X"5c", -- b
        16#b62# => X"00", -- b
        16#c62# => X"00", -- b
        16#063# => X"00", -- c
        16#163# => X"00", -- c
        16#263# => X"00", -- c
        16#363# => X"00", -- c
        16#463# => X"00", -- c
        16#563# => X"3c", -- c
        16#663# => X"42", -- c
        16#763# => X"40", -- c
        16#863# => X"40", -- c
        16#963# => X"42", -- c
        16#a63# => X"3c", -- c
        16#b63# => X"00", -- c
        16#c63# => X"00", -- c
        16#064# => X"00", -- d
        16#164# => X"00", -- d
        16#264# => X"02", -- d
        16#364# => X"02", -- d
        16#464# => X"02", -- d
        16#564# => X"3a", -- d
        16#664# => X"46", -- d
        16#764# => X"42", -- d
        16#864# => X"42", -- d
        16#964# => X"46", -- d
        16#a64# => X"3a", -- d
        16#b64# => X"00", -- d
        16#c64# => X"00", -- d
        16#065# => X"00", -- e
        16#165# => X"00", -- e
        16#265# => X"00", -- e
        16#365# => X"00", -- e
        16#465# => X"00", -- e
        16#565# => X"3c", -- e
        16#665# => X"42", -- e
        16#765# => X"7e", -- e
        16#865# => X"40", -- e
        16#965# => X"42", -- e
        16#a65# => X"3c", -- e
        16#b65# => X"00", -- e
        16#c65# => X"00", -- e
        16#066# => X"00", -- f
        16#166# => X"00", -- f
        16#266# => X"1c", -- f
        16#366# => X"22", -- f
        16#466# => X"20", -- f
        16#566# => X"20", -- f
        16#666# => X"7c", -- f
        16#766# => X"20", -- f
        16#866# => X"20", -- f
        16#966# => X"20", -- f
        16#a66# => X"20", -- f
        16#b66# => X"00", -- f
        16#c66# => X"00", -- f
        16#067# => X"00", -- g
        16#167# => X"00", -- g
        16#267# => X"00", -- g
        16#367# => X"00", -- g
        16#467# => X"00", -- g
        16#567# => X"3a", -- g
        16#667# => X"44", -- g
        16#767# => X"44", -- g
        16#867# => X"38", -- g
        16#967# => X"40", -- g
        16#a67# => X"3c", -- g
        16#b67# => X"42", -- g
        16#c67# => X"3c", -- g
        16#068# => X"00", -- h
        16#168# => X"00", -- h
        16#268# => X"40", -- h
        16#368# => X"40", -- h
        16#468# => X"40", -- h
        16#568# => X"5c", -- h
        16#668# => X"62", -- h
        16#768# => X"42", -- h
        16#868# => X"42", -- h
        16#968# => X"42", -- h
        16#a68# => X"42", -- h
        16#b68# => X"00", -- h
        16#c68# => X"00", -- h
        16#069# => X"00", -- i
        16#169# => X"00", -- i
        16#269# => X"00", -- i
        16#369# => X"10", -- i
        16#469# => X"00", -- i
        16#569# => X"30", -- i
        16#669# => X"10", -- i
        16#769# => X"10", -- i
        16#869# => X"10", -- i
        16#969# => X"10", -- i
        16#a69# => X"7c", -- i
        16#b69# => X"00", -- i
        16#c69# => X"00", -- i
        16#06a# => X"00", -- j
        16#16a# => X"00", -- j
        16#26a# => X"00", -- j
        16#36a# => X"04", -- j
        16#46a# => X"00", -- j
        16#56a# => X"0c", -- j
        16#66a# => X"04", -- j
        16#76a# => X"04", -- j
        16#86a# => X"04", -- j
        16#96a# => X"04", -- j
        16#a6a# => X"44", -- j
        16#b6a# => X"44", -- j
        16#c6a# => X"38", -- j
        16#06b# => X"00", -- k
        16#16b# => X"00", -- k
        16#26b# => X"40", -- k
        16#36b# => X"40", -- k
        16#46b# => X"40", -- k
        16#56b# => X"44", -- k
        16#66b# => X"48", -- k
        16#76b# => X"70", -- k
        16#86b# => X"48", -- k
        16#96b# => X"44", -- k
        16#a6b# => X"42", -- k
        16#b6b# => X"00", -- k
        16#c6b# => X"00", -- k
        16#06c# => X"00", -- l
        16#16c# => X"00", -- l
        16#26c# => X"30", -- l
        16#36c# => X"10", -- l
        16#46c# => X"10", -- l
        16#56c# => X"10", -- l
        16#66c# => X"10", -- l
        16#76c# => X"10", -- l
        16#86c# => X"10", -- l
        16#96c# => X"10", -- l
        16#a6c# => X"7c", -- l
        16#b6c# => X"00", -- l
        16#c6c# => X"00", -- l
        16#06d# => X"00", -- m
        16#16d# => X"00", -- m
        16#26d# => X"00", -- m
        16#36d# => X"00", -- m
        16#46d# => X"00", -- m
        16#56d# => X"ec", -- m
        16#66d# => X"92", -- m
        16#76d# => X"92", -- m
        16#86d# => X"92", -- m
        16#96d# => X"92", -- m
        16#a6d# => X"82", -- m
        16#b6d# => X"00", -- m
        16#c6d# => X"00", -- m
        16#06e# => X"00", -- n
        16#16e# => X"00", -- n
        16#26e# => X"00", -- n
        16#36e# => X"00", -- n
        16#46e# => X"00", -- n
        16#56e# => X"5c", -- n
        16#66e# => X"62", -- n
        16#76e# => X"42", -- n
        16#86e# => X"42", -- n
        16#96e# => X"42", -- n
        16#a6e# => X"42", -- n
        16#b6e# => X"00", -- n
        16#c6e# => X"00", -- n
        16#06f# => X"00", -- o
        16#16f# => X"00", -- o
        16#26f# => X"00", -- o
        16#36f# => X"00", -- o
        16#46f# => X"00", -- o
        16#56f# => X"3c", -- o
        16#66f# => X"42", -- o
        16#76f# => X"42", -- o
        16#86f# => X"42", -- o
        16#96f# => X"42", -- o
        16#a6f# => X"3c", -- o
        16#b6f# => X"00", -- o
        16#c6f# => X"00", -- o
        16#070# => X"00", -- p
        16#170# => X"00", -- p
        16#270# => X"00", -- p
        16#370# => X"00", -- p
        16#470# => X"00", -- p
        16#570# => X"5c", -- p
        16#670# => X"62", -- p
        16#770# => X"42", -- p
        16#870# => X"62", -- p
        16#970# => X"5c", -- p
        16#a70# => X"40", -- p
        16#b70# => X"40", -- p
        16#c70# => X"40", -- p
        16#071# => X"00", -- q
        16#171# => X"00", -- q
        16#271# => X"00", -- q
        16#371# => X"00", -- q
        16#471# => X"00", -- q
        16#571# => X"3a", -- q
        16#671# => X"46", -- q
        16#771# => X"42", -- q
        16#871# => X"46", -- q
        16#971# => X"3a", -- q
        16#a71# => X"02", -- q
        16#b71# => X"02", -- q
        16#c71# => X"02", -- q
        16#072# => X"00", -- r
        16#172# => X"00", -- r
        16#272# => X"00", -- r
        16#372# => X"00", -- r
        16#472# => X"00", -- r
        16#572# => X"5c", -- r
        16#672# => X"22", -- r
        16#772# => X"20", -- r
        16#872# => X"20", -- r
        16#972# => X"20", -- r
        16#a72# => X"20", -- r
        16#b72# => X"00", -- r
        16#c72# => X"00", -- r
        16#073# => X"00", -- s
        16#173# => X"00", -- s
        16#273# => X"00", -- s
        16#373# => X"00", -- s
        16#473# => X"00", -- s
        16#573# => X"3c", -- s
        16#673# => X"42", -- s
        16#773# => X"30", -- s
        16#873# => X"0c", -- s
        16#973# => X"42", -- s
        16#a73# => X"3c", -- s
        16#b73# => X"00", -- s
        16#c73# => X"00", -- s
        16#074# => X"00", -- t
        16#174# => X"00", -- t
        16#274# => X"00", -- t
        16#374# => X"20", -- t
        16#474# => X"20", -- t
        16#574# => X"7c", -- t
        16#674# => X"20", -- t
        16#774# => X"20", -- t
        16#874# => X"20", -- t
        16#974# => X"22", -- t
        16#a74# => X"1c", -- t
        16#b74# => X"00", -- t
        16#c74# => X"00", -- t
        16#075# => X"00", -- u
        16#175# => X"00", -- u
        16#275# => X"00", -- u
        16#375# => X"00", -- u
        16#475# => X"00", -- u
        16#575# => X"44", -- u
        16#675# => X"44", -- u
        16#775# => X"44", -- u
        16#875# => X"44", -- u
        16#975# => X"44", -- u
        16#a75# => X"3a", -- u
        16#b75# => X"00", -- u
        16#c75# => X"00", -- u
        16#076# => X"00", -- v
        16#176# => X"00", -- v
        16#276# => X"00", -- v
        16#376# => X"00", -- v
        16#476# => X"00", -- v
        16#576# => X"44", -- v
        16#676# => X"44", -- v
        16#776# => X"44", -- v
        16#876# => X"28", -- v
        16#976# => X"28", -- v
        16#a76# => X"10", -- v
        16#b76# => X"00", -- v
        16#c76# => X"00", -- v
        16#077# => X"00", -- w
        16#177# => X"00", -- w
        16#277# => X"00", -- w
        16#377# => X"00", -- w
        16#477# => X"00", -- w
        16#577# => X"82", -- w
        16#677# => X"82", -- w
        16#777# => X"92", -- w
        16#877# => X"92", -- w
        16#977# => X"aa", -- w
        16#a77# => X"44", -- w
        16#b77# => X"00", -- w
        16#c77# => X"00", -- w
        16#078# => X"00", -- x
        16#178# => X"00", -- x
        16#278# => X"00", -- x
        16#378# => X"00", -- x
        16#478# => X"00", -- x
        16#578# => X"42", -- x
        16#678# => X"24", -- x
        16#778# => X"18", -- x
        16#878# => X"18", -- x
        16#978# => X"24", -- x
        16#a78# => X"42", -- x
        16#b78# => X"00", -- x
        16#c78# => X"00", -- x
        16#079# => X"00", -- y
        16#179# => X"00", -- y
        16#279# => X"00", -- y
        16#379# => X"00", -- y
        16#479# => X"00", -- y
        16#579# => X"42", -- y
        16#679# => X"42", -- y
        16#779# => X"42", -- y
        16#879# => X"46", -- y
        16#979# => X"3a", -- y
        16#a79# => X"02", -- y
        16#b79# => X"42", -- y
        16#c79# => X"3c", -- y
        16#07a# => X"00", -- z
        16#17a# => X"00", -- z
        16#27a# => X"00", -- z
        16#37a# => X"00", -- z
        16#47a# => X"00", -- z
        16#57a# => X"7e", -- z
        16#67a# => X"04", -- z
        16#77a# => X"08", -- z
        16#87a# => X"10", -- z
        16#97a# => X"20", -- z
        16#a7a# => X"7e", -- z
        16#b7a# => X"00", -- z
        16#c7a# => X"00", -- z
        16#07b# => X"00", -- {
        16#17b# => X"00", -- {
        16#27b# => X"0e", -- {
        16#37b# => X"10", -- {
        16#47b# => X"10", -- {
        16#57b# => X"08", -- {
        16#67b# => X"30", -- {
        16#77b# => X"08", -- {
        16#87b# => X"10", -- {
        16#97b# => X"10", -- {
        16#a7b# => X"0e", -- {
        16#b7b# => X"00", -- {
        16#c7b# => X"00", -- {
        16#07c# => X"00", -- |
        16#17c# => X"00", -- |
        16#27c# => X"10", -- |
        16#37c# => X"10", -- |
        16#47c# => X"10", -- |
        16#57c# => X"10", -- |
        16#67c# => X"10", -- |
        16#77c# => X"10", -- |
        16#87c# => X"10", -- |
        16#97c# => X"10", -- |
        16#a7c# => X"10", -- |
        16#b7c# => X"00", -- |
        16#c7c# => X"00", -- |
        16#07d# => X"00", -- }
        16#17d# => X"00", -- }
        16#27d# => X"70", -- }
        16#37d# => X"08", -- }
        16#47d# => X"08", -- }
        16#57d# => X"10", -- }
        16#67d# => X"0c", -- }
        16#77d# => X"10", -- }
        16#87d# => X"08", -- }
        16#97d# => X"08", -- }
        16#a7d# => X"70", -- }
        16#b7d# => X"00", -- }
        16#c7d# => X"00", -- }
        16#07e# => X"00", -- ~
        16#17e# => X"00", -- ~
        16#27e# => X"24", -- ~
        16#37e# => X"54", -- ~
        16#47e# => X"48", -- ~
        16#57e# => X"00", -- ~
        16#67e# => X"00", -- ~
        16#77e# => X"00", -- ~
        16#87e# => X"00", -- ~
        16#97e# => X"00", -- ~
        16#a7e# => X"00", -- ~
        16#b7e# => X"00", -- ~
        16#c7e# => X"00", -- ~
        16#0a0# => X"00", -- �
        16#1a0# => X"00", -- �
        16#2a0# => X"00", -- �
        16#3a0# => X"00", -- �
        16#4a0# => X"00", -- �
        16#5a0# => X"00", -- �
        16#6a0# => X"00", -- �
        16#7a0# => X"00", -- �
        16#8a0# => X"00", -- �
        16#9a0# => X"00", -- �
        16#aa0# => X"00", -- �
        16#ba0# => X"00", -- �
        16#ca0# => X"00", -- �
        16#0a1# => X"00", -- �
        16#1a1# => X"00", -- �
        16#2a1# => X"10", -- �
        16#3a1# => X"00", -- �
        16#4a1# => X"10", -- �
        16#5a1# => X"10", -- �
        16#6a1# => X"10", -- �
        16#7a1# => X"10", -- �
        16#8a1# => X"10", -- �
        16#9a1# => X"10", -- �
        16#aa1# => X"10", -- �
        16#ba1# => X"00", -- �
        16#ca1# => X"00", -- �
        16#0a2# => X"00", -- �
        16#1a2# => X"00", -- �
        16#2a2# => X"10", -- �
        16#3a2# => X"38", -- �
        16#4a2# => X"54", -- �
        16#5a2# => X"50", -- �
        16#6a2# => X"50", -- �
        16#7a2# => X"54", -- �
        16#8a2# => X"38", -- �
        16#9a2# => X"10", -- �
        16#aa2# => X"00", -- �
        16#ba2# => X"00", -- �
        16#ca2# => X"00", -- �
        16#0a3# => X"00", -- �
        16#1a3# => X"00", -- �
        16#2a3# => X"1c", -- �
        16#3a3# => X"22", -- �
        16#4a3# => X"20", -- �
        16#5a3# => X"70", -- �
        16#6a3# => X"20", -- �
        16#7a3# => X"20", -- �
        16#8a3# => X"20", -- �
        16#9a3# => X"62", -- �
        16#aa3# => X"dc", -- �
        16#ba3# => X"00", -- �
        16#ca3# => X"00", -- �
        16#0a4# => X"00", -- �
        16#1a4# => X"00", -- �
        16#2a4# => X"00", -- �
        16#3a4# => X"00", -- �
        16#4a4# => X"42", -- �
        16#5a4# => X"3c", -- �
        16#6a4# => X"24", -- �
        16#7a4# => X"24", -- �
        16#8a4# => X"3c", -- �
        16#9a4# => X"42", -- �
        16#aa4# => X"00", -- �
        16#ba4# => X"00", -- �
        16#ca4# => X"00", -- �
        16#0a5# => X"00", -- �
        16#1a5# => X"00", -- �
        16#2a5# => X"82", -- �
        16#3a5# => X"82", -- �
        16#4a5# => X"44", -- �
        16#5a5# => X"28", -- �
        16#6a5# => X"7c", -- �
        16#7a5# => X"10", -- �
        16#8a5# => X"7c", -- �
        16#9a5# => X"10", -- �
        16#aa5# => X"10", -- �
        16#ba5# => X"00", -- �
        16#ca5# => X"00", -- �
        16#0a6# => X"00", -- �
        16#1a6# => X"00", -- �
        16#2a6# => X"10", -- �
        16#3a6# => X"10", -- �
        16#4a6# => X"10", -- �
        16#5a6# => X"10", -- �
        16#6a6# => X"00", -- �
        16#7a6# => X"10", -- �
        16#8a6# => X"10", -- �
        16#9a6# => X"10", -- �
        16#aa6# => X"10", -- �
        16#ba6# => X"00", -- �
        16#ca6# => X"00", -- �
        16#0a7# => X"00", -- �
        16#1a7# => X"18", -- �
        16#2a7# => X"24", -- �
        16#3a7# => X"20", -- �
        16#4a7# => X"18", -- �
        16#5a7# => X"24", -- �
        16#6a7# => X"24", -- �
        16#7a7# => X"18", -- �
        16#8a7# => X"04", -- �
        16#9a7# => X"24", -- �
        16#aa7# => X"18", -- �
        16#ba7# => X"00", -- �
        16#ca7# => X"00", -- �
        16#0a8# => X"00", -- �
        16#1a8# => X"24", -- �
        16#2a8# => X"24", -- �
        16#3a8# => X"00", -- �
        16#4a8# => X"00", -- �
        16#5a8# => X"00", -- �
        16#6a8# => X"00", -- �
        16#7a8# => X"00", -- �
        16#8a8# => X"00", -- �
        16#9a8# => X"00", -- �
        16#aa8# => X"00", -- �
        16#ba8# => X"00", -- �
        16#ca8# => X"00", -- �
        16#0a9# => X"00", -- �
        16#1a9# => X"38", -- �
        16#2a9# => X"44", -- �
        16#3a9# => X"92", -- �
        16#4a9# => X"aa", -- �
        16#5a9# => X"a2", -- �
        16#6a9# => X"aa", -- �
        16#7a9# => X"92", -- �
        16#8a9# => X"44", -- �
        16#9a9# => X"38", -- �
        16#aa9# => X"00", -- �
        16#ba9# => X"00", -- �
        16#ca9# => X"00", -- �
        16#0aa# => X"00", -- �
        16#1aa# => X"00", -- �
        16#2aa# => X"38", -- �
        16#3aa# => X"04", -- �
        16#4aa# => X"3c", -- �
        16#5aa# => X"44", -- �
        16#6aa# => X"3c", -- �
        16#7aa# => X"00", -- �
        16#8aa# => X"7c", -- �
        16#9aa# => X"00", -- �
        16#aaa# => X"00", -- �
        16#baa# => X"00", -- �
        16#caa# => X"00", -- �
        16#0ab# => X"00", -- �
        16#1ab# => X"00", -- �
        16#2ab# => X"00", -- �
        16#3ab# => X"12", -- �
        16#4ab# => X"24", -- �
        16#5ab# => X"48", -- �
        16#6ab# => X"90", -- �
        16#7ab# => X"48", -- �
        16#8ab# => X"24", -- �
        16#9ab# => X"12", -- �
        16#aab# => X"00", -- �
        16#bab# => X"00", -- �
        16#cab# => X"00", -- �
        16#0ac# => X"00", -- �
        16#1ac# => X"00", -- �
        16#2ac# => X"00", -- �
        16#3ac# => X"00", -- �
        16#4ac# => X"00", -- �
        16#5ac# => X"00", -- �
        16#6ac# => X"7e", -- �
        16#7ac# => X"02", -- �
        16#8ac# => X"02", -- �
        16#9ac# => X"02", -- �
        16#aac# => X"00", -- �
        16#bac# => X"00", -- �
        16#cac# => X"00", -- �
        16#0ad# => X"00", -- �
        16#1ad# => X"00", -- �
        16#2ad# => X"00", -- �
        16#3ad# => X"00", -- �
        16#4ad# => X"00", -- �
        16#5ad# => X"00", -- �
        16#6ad# => X"3c", -- �
        16#7ad# => X"00", -- �
        16#8ad# => X"00", -- �
        16#9ad# => X"00", -- �
        16#aad# => X"00", -- �
        16#bad# => X"00", -- �
        16#cad# => X"00", -- �
        16#0ae# => X"00", -- �
        16#1ae# => X"38", -- �
        16#2ae# => X"44", -- �
        16#3ae# => X"92", -- �
        16#4ae# => X"aa", -- �
        16#5ae# => X"aa", -- �
        16#6ae# => X"b2", -- �
        16#7ae# => X"aa", -- �
        16#8ae# => X"44", -- �
        16#9ae# => X"38", -- �
        16#aae# => X"00", -- �
        16#bae# => X"00", -- �
        16#cae# => X"00", -- �
        16#0af# => X"00", -- �
        16#1af# => X"00", -- �
        16#2af# => X"7e", -- �
        16#3af# => X"00", -- �
        16#4af# => X"00", -- �
        16#5af# => X"00", -- �
        16#6af# => X"00", -- �
        16#7af# => X"00", -- �
        16#8af# => X"00", -- �
        16#9af# => X"00", -- �
        16#aaf# => X"00", -- �
        16#baf# => X"00", -- �
        16#caf# => X"00", -- �
        16#0b0# => X"00", -- �
        16#1b0# => X"00", -- �
        16#2b0# => X"18", -- �
        16#3b0# => X"24", -- �
        16#4b0# => X"24", -- �
        16#5b0# => X"18", -- �
        16#6b0# => X"00", -- �
        16#7b0# => X"00", -- �
        16#8b0# => X"00", -- �
        16#9b0# => X"00", -- �
        16#ab0# => X"00", -- �
        16#bb0# => X"00", -- �
        16#cb0# => X"00", -- �
        16#0b1# => X"00", -- �
        16#1b1# => X"00", -- �
        16#2b1# => X"00", -- �
        16#3b1# => X"10", -- �
        16#4b1# => X"10", -- �
        16#5b1# => X"7c", -- �
        16#6b1# => X"10", -- �
        16#7b1# => X"10", -- �
        16#8b1# => X"00", -- �
        16#9b1# => X"7c", -- �
        16#ab1# => X"00", -- �
        16#bb1# => X"00", -- �
        16#cb1# => X"00", -- �
        16#0b2# => X"00", -- �
        16#1b2# => X"30", -- �
        16#2b2# => X"48", -- �
        16#3b2# => X"08", -- �
        16#4b2# => X"30", -- �
        16#5b2# => X"40", -- �
        16#6b2# => X"78", -- �
        16#7b2# => X"00", -- �
        16#8b2# => X"00", -- �
        16#9b2# => X"00", -- �
        16#ab2# => X"00", -- �
        16#bb2# => X"00", -- �
        16#cb2# => X"00", -- �
        16#0b3# => X"00", -- �
        16#1b3# => X"30", -- �
        16#2b3# => X"48", -- �
        16#3b3# => X"10", -- �
        16#4b3# => X"08", -- �
        16#5b3# => X"48", -- �
        16#6b3# => X"30", -- �
        16#7b3# => X"00", -- �
        16#8b3# => X"00", -- �
        16#9b3# => X"00", -- �
        16#ab3# => X"00", -- �
        16#bb3# => X"00", -- �
        16#cb3# => X"00", -- �
        16#0b4# => X"00", -- �
        16#1b4# => X"08", -- �
        16#2b4# => X"10", -- �
        16#3b4# => X"00", -- �
        16#4b4# => X"00", -- �
        16#5b4# => X"00", -- �
        16#6b4# => X"00", -- �
        16#7b4# => X"00", -- �
        16#8b4# => X"00", -- �
        16#9b4# => X"00", -- �
        16#ab4# => X"00", -- �
        16#bb4# => X"00", -- �
        16#cb4# => X"00", -- �
        16#0b5# => X"00", -- �
        16#1b5# => X"00", -- �
        16#2b5# => X"00", -- �
        16#3b5# => X"00", -- �
        16#4b5# => X"00", -- �
        16#5b5# => X"42", -- �
        16#6b5# => X"42", -- �
        16#7b5# => X"42", -- �
        16#8b5# => X"42", -- �
        16#9b5# => X"66", -- �
        16#ab5# => X"5a", -- �
        16#bb5# => X"40", -- �
        16#cb5# => X"00", -- �
        16#0b6# => X"00", -- �
        16#1b6# => X"00", -- �
        16#2b6# => X"3e", -- �
        16#3b6# => X"74", -- �
        16#4b6# => X"74", -- �
        16#5b6# => X"74", -- �
        16#6b6# => X"34", -- �
        16#7b6# => X"14", -- �
        16#8b6# => X"14", -- �
        16#9b6# => X"14", -- �
        16#ab6# => X"14", -- �
        16#bb6# => X"00", -- �
        16#cb6# => X"00", -- �
        16#0b7# => X"00", -- �
        16#1b7# => X"00", -- �
        16#2b7# => X"00", -- �
        16#3b7# => X"00", -- �
        16#4b7# => X"00", -- �
        16#5b7# => X"00", -- �
        16#6b7# => X"18", -- �
        16#7b7# => X"00", -- �
        16#8b7# => X"00", -- �
        16#9b7# => X"00", -- �
        16#ab7# => X"00", -- �
        16#bb7# => X"00", -- �
        16#cb7# => X"00", -- �
        16#0b8# => X"00", -- �
        16#1b8# => X"00", -- �
        16#2b8# => X"00", -- �
        16#3b8# => X"00", -- �
        16#4b8# => X"00", -- �
        16#5b8# => X"00", -- �
        16#6b8# => X"00", -- �
        16#7b8# => X"00", -- �
        16#8b8# => X"00", -- �
        16#9b8# => X"00", -- �
        16#ab8# => X"00", -- �
        16#bb8# => X"08", -- �
        16#cb8# => X"18", -- �
        16#0b9# => X"00", -- �
        16#1b9# => X"20", -- �
        16#2b9# => X"60", -- �
        16#3b9# => X"20", -- �
        16#4b9# => X"20", -- �
        16#5b9# => X"20", -- �
        16#6b9# => X"70", -- �
        16#7b9# => X"00", -- �
        16#8b9# => X"00", -- �
        16#9b9# => X"00", -- �
        16#ab9# => X"00", -- �
        16#bb9# => X"00", -- �
        16#cb9# => X"00", -- �
        16#0ba# => X"00", -- �
        16#1ba# => X"00", -- �
        16#2ba# => X"30", -- �
        16#3ba# => X"48", -- �
        16#4ba# => X"48", -- �
        16#5ba# => X"30", -- �
        16#6ba# => X"00", -- �
        16#7ba# => X"78", -- �
        16#8ba# => X"00", -- �
        16#9ba# => X"00", -- �
        16#aba# => X"00", -- �
        16#bba# => X"00", -- �
        16#cba# => X"00", -- �
        16#0bb# => X"00", -- �
        16#1bb# => X"00", -- �
        16#2bb# => X"00", -- �
        16#3bb# => X"90", -- �
        16#4bb# => X"48", -- �
        16#5bb# => X"24", -- �
        16#6bb# => X"12", -- �
        16#7bb# => X"24", -- �
        16#8bb# => X"48", -- �
        16#9bb# => X"90", -- �
        16#abb# => X"00", -- �
        16#bbb# => X"00", -- �
        16#cbb# => X"00", -- �
        16#0bc# => X"00", -- �
        16#1bc# => X"40", -- �
        16#2bc# => X"c0", -- �
        16#3bc# => X"40", -- �
        16#4bc# => X"40", -- �
        16#5bc# => X"42", -- �
        16#6bc# => X"e6", -- �
        16#7bc# => X"0a", -- �
        16#8bc# => X"12", -- �
        16#9bc# => X"1a", -- �
        16#abc# => X"06", -- �
        16#bbc# => X"00", -- �
        16#cbc# => X"00", -- �
        16#0bd# => X"00", -- �
        16#1bd# => X"40", -- �
        16#2bd# => X"c0", -- �
        16#3bd# => X"40", -- �
        16#4bd# => X"40", -- �
        16#5bd# => X"4c", -- �
        16#6bd# => X"f2", -- �
        16#7bd# => X"02", -- �
        16#8bd# => X"0c", -- �
        16#9bd# => X"10", -- �
        16#abd# => X"1e", -- �
        16#bbd# => X"00", -- �
        16#cbd# => X"00", -- �
        16#0be# => X"00", -- �
        16#1be# => X"60", -- �
        16#2be# => X"90", -- �
        16#3be# => X"20", -- �
        16#4be# => X"10", -- �
        16#5be# => X"92", -- �
        16#6be# => X"66", -- �
        16#7be# => X"0a", -- �
        16#8be# => X"12", -- �
        16#9be# => X"1a", -- �
        16#abe# => X"06", -- �
        16#bbe# => X"00", -- �
        16#cbe# => X"00", -- �
        16#0bf# => X"00", -- �
        16#1bf# => X"00", -- �
        16#2bf# => X"10", -- �
        16#3bf# => X"00", -- �
        16#4bf# => X"10", -- �
        16#5bf# => X"10", -- �
        16#6bf# => X"20", -- �
        16#7bf# => X"40", -- �
        16#8bf# => X"42", -- �
        16#9bf# => X"42", -- �
        16#abf# => X"3c", -- �
        16#bbf# => X"00", -- �
        16#cbf# => X"00", -- �
        16#0c0# => X"00", -- �
        16#1c0# => X"10", -- �
        16#2c0# => X"08", -- �
        16#3c0# => X"00", -- �
        16#4c0# => X"18", -- �
        16#5c0# => X"24", -- �
        16#6c0# => X"42", -- �
        16#7c0# => X"42", -- �
        16#8c0# => X"7e", -- �
        16#9c0# => X"42", -- �
        16#ac0# => X"42", -- �
        16#bc0# => X"00", -- �
        16#cc0# => X"00", -- �
        16#0c1# => X"00", -- �
        16#1c1# => X"08", -- �
        16#2c1# => X"10", -- �
        16#3c1# => X"00", -- �
        16#4c1# => X"18", -- �
        16#5c1# => X"24", -- �
        16#6c1# => X"42", -- �
        16#7c1# => X"42", -- �
        16#8c1# => X"7e", -- �
        16#9c1# => X"42", -- �
        16#ac1# => X"42", -- �
        16#bc1# => X"00", -- �
        16#cc1# => X"00", -- �
        16#0c2# => X"00", -- �
        16#1c2# => X"18", -- �
        16#2c2# => X"24", -- �
        16#3c2# => X"00", -- �
        16#4c2# => X"18", -- �
        16#5c2# => X"24", -- �
        16#6c2# => X"42", -- �
        16#7c2# => X"42", -- �
        16#8c2# => X"7e", -- �
        16#9c2# => X"42", -- �
        16#ac2# => X"42", -- �
        16#bc2# => X"00", -- �
        16#cc2# => X"00", -- �
        16#0c3# => X"00", -- �
        16#1c3# => X"32", -- �
        16#2c3# => X"4c", -- �
        16#3c3# => X"00", -- �
        16#4c3# => X"18", -- �
        16#5c3# => X"24", -- �
        16#6c3# => X"42", -- �
        16#7c3# => X"42", -- �
        16#8c3# => X"7e", -- �
        16#9c3# => X"42", -- �
        16#ac3# => X"42", -- �
        16#bc3# => X"00", -- �
        16#cc3# => X"00", -- �
        16#0c4# => X"00", -- �
        16#1c4# => X"24", -- �
        16#2c4# => X"24", -- �
        16#3c4# => X"00", -- �
        16#4c4# => X"18", -- �
        16#5c4# => X"24", -- �
        16#6c4# => X"42", -- �
        16#7c4# => X"42", -- �
        16#8c4# => X"7e", -- �
        16#9c4# => X"42", -- �
        16#ac4# => X"42", -- �
        16#bc4# => X"00", -- �
        16#cc4# => X"00", -- �
        16#0c5# => X"00", -- �
        16#1c5# => X"18", -- �
        16#2c5# => X"24", -- �
        16#3c5# => X"18", -- �
        16#4c5# => X"18", -- �
        16#5c5# => X"24", -- �
        16#6c5# => X"42", -- �
        16#7c5# => X"42", -- �
        16#8c5# => X"7e", -- �
        16#9c5# => X"42", -- �
        16#ac5# => X"42", -- �
        16#bc5# => X"00", -- �
        16#cc5# => X"00", -- �
        16#0c6# => X"00", -- �
        16#1c6# => X"00", -- �
        16#2c6# => X"6e", -- �
        16#3c6# => X"90", -- �
        16#4c6# => X"90", -- �
        16#5c6# => X"90", -- �
        16#6c6# => X"9c", -- �
        16#7c6# => X"f0", -- �
        16#8c6# => X"90", -- �
        16#9c6# => X"90", -- �
        16#ac6# => X"9e", -- �
        16#bc6# => X"00", -- �
        16#cc6# => X"00", -- �
        16#0c7# => X"00", -- �
        16#1c7# => X"00", -- �
        16#2c7# => X"3c", -- �
        16#3c7# => X"42", -- �
        16#4c7# => X"40", -- �
        16#5c7# => X"40", -- �
        16#6c7# => X"40", -- �
        16#7c7# => X"40", -- �
        16#8c7# => X"40", -- �
        16#9c7# => X"42", -- �
        16#ac7# => X"3c", -- �
        16#bc7# => X"08", -- �
        16#cc7# => X"10", -- �
        16#0c8# => X"00", -- �
        16#1c8# => X"10", -- �
        16#2c8# => X"08", -- �
        16#3c8# => X"00", -- �
        16#4c8# => X"7e", -- �
        16#5c8# => X"40", -- �
        16#6c8# => X"40", -- �
        16#7c8# => X"78", -- �
        16#8c8# => X"40", -- �
        16#9c8# => X"40", -- �
        16#ac8# => X"7e", -- �
        16#bc8# => X"00", -- �
        16#cc8# => X"00", -- �
        16#0c9# => X"00", -- �
        16#1c9# => X"08", -- �
        16#2c9# => X"10", -- �
        16#3c9# => X"00", -- �
        16#4c9# => X"7e", -- �
        16#5c9# => X"40", -- �
        16#6c9# => X"40", -- �
        16#7c9# => X"78", -- �
        16#8c9# => X"40", -- �
        16#9c9# => X"40", -- �
        16#ac9# => X"7e", -- �
        16#bc9# => X"00", -- �
        16#cc9# => X"00", -- �
        16#0ca# => X"00", -- �
        16#1ca# => X"18", -- �
        16#2ca# => X"24", -- �
        16#3ca# => X"00", -- �
        16#4ca# => X"7e", -- �
        16#5ca# => X"40", -- �
        16#6ca# => X"40", -- �
        16#7ca# => X"78", -- �
        16#8ca# => X"40", -- �
        16#9ca# => X"40", -- �
        16#aca# => X"7e", -- �
        16#bca# => X"00", -- �
        16#cca# => X"00", -- �
        16#0cb# => X"00", -- �
        16#1cb# => X"24", -- �
        16#2cb# => X"24", -- �
        16#3cb# => X"00", -- �
        16#4cb# => X"7e", -- �
        16#5cb# => X"40", -- �
        16#6cb# => X"40", -- �
        16#7cb# => X"78", -- �
        16#8cb# => X"40", -- �
        16#9cb# => X"40", -- �
        16#acb# => X"7e", -- �
        16#bcb# => X"00", -- �
        16#ccb# => X"00", -- �
        16#0cc# => X"00", -- �
        16#1cc# => X"20", -- �
        16#2cc# => X"10", -- �
        16#3cc# => X"00", -- �
        16#4cc# => X"7c", -- �
        16#5cc# => X"10", -- �
        16#6cc# => X"10", -- �
        16#7cc# => X"10", -- �
        16#8cc# => X"10", -- �
        16#9cc# => X"10", -- �
        16#acc# => X"7c", -- �
        16#bcc# => X"00", -- �
        16#ccc# => X"00", -- �
        16#0cd# => X"00", -- �
        16#1cd# => X"08", -- �
        16#2cd# => X"10", -- �
        16#3cd# => X"00", -- �
        16#4cd# => X"7c", -- �
        16#5cd# => X"10", -- �
        16#6cd# => X"10", -- �
        16#7cd# => X"10", -- �
        16#8cd# => X"10", -- �
        16#9cd# => X"10", -- �
        16#acd# => X"7c", -- �
        16#bcd# => X"00", -- �
        16#ccd# => X"00", -- �
        16#0ce# => X"00", -- �
        16#1ce# => X"18", -- �
        16#2ce# => X"24", -- �
        16#3ce# => X"00", -- �
        16#4ce# => X"7c", -- �
        16#5ce# => X"10", -- �
        16#6ce# => X"10", -- �
        16#7ce# => X"10", -- �
        16#8ce# => X"10", -- �
        16#9ce# => X"10", -- �
        16#ace# => X"7c", -- �
        16#bce# => X"00", -- �
        16#cce# => X"00", -- �
        16#0cf# => X"00", -- �
        16#1cf# => X"44", -- �
        16#2cf# => X"44", -- �
        16#3cf# => X"00", -- �
        16#4cf# => X"7c", -- �
        16#5cf# => X"10", -- �
        16#6cf# => X"10", -- �
        16#7cf# => X"10", -- �
        16#8cf# => X"10", -- �
        16#9cf# => X"10", -- �
        16#acf# => X"7c", -- �
        16#bcf# => X"00", -- �
        16#ccf# => X"00", -- �
        16#0d0# => X"00", -- �
        16#1d0# => X"00", -- �
        16#2d0# => X"78", -- �
        16#3d0# => X"44", -- �
        16#4d0# => X"42", -- �
        16#5d0# => X"42", -- �
        16#6d0# => X"e2", -- �
        16#7d0# => X"42", -- �
        16#8d0# => X"42", -- �
        16#9d0# => X"44", -- �
        16#ad0# => X"78", -- �
        16#bd0# => X"00", -- �
        16#cd0# => X"00", -- �
        16#0d1# => X"00", -- �
        16#1d1# => X"64", -- �
        16#2d1# => X"98", -- �
        16#3d1# => X"00", -- �
        16#4d1# => X"82", -- �
        16#5d1# => X"c2", -- �
        16#6d1# => X"a2", -- �
        16#7d1# => X"92", -- �
        16#8d1# => X"8a", -- �
        16#9d1# => X"86", -- �
        16#ad1# => X"82", -- �
        16#bd1# => X"00", -- �
        16#cd1# => X"00", -- �
        16#0d2# => X"00", -- �
        16#1d2# => X"20", -- �
        16#2d2# => X"10", -- �
        16#3d2# => X"00", -- �
        16#4d2# => X"7c", -- �
        16#5d2# => X"82", -- �
        16#6d2# => X"82", -- �
        16#7d2# => X"82", -- �
        16#8d2# => X"82", -- �
        16#9d2# => X"82", -- �
        16#ad2# => X"7c", -- �
        16#bd2# => X"00", -- �
        16#cd2# => X"00", -- �
        16#0d3# => X"00", -- �
        16#1d3# => X"08", -- �
        16#2d3# => X"10", -- �
        16#3d3# => X"00", -- �
        16#4d3# => X"7c", -- �
        16#5d3# => X"82", -- �
        16#6d3# => X"82", -- �
        16#7d3# => X"82", -- �
        16#8d3# => X"82", -- �
        16#9d3# => X"82", -- �
        16#ad3# => X"7c", -- �
        16#bd3# => X"00", -- �
        16#cd3# => X"00", -- �
        16#0d4# => X"00", -- �
        16#1d4# => X"18", -- �
        16#2d4# => X"24", -- �
        16#3d4# => X"00", -- �
        16#4d4# => X"7c", -- �
        16#5d4# => X"82", -- �
        16#6d4# => X"82", -- �
        16#7d4# => X"82", -- �
        16#8d4# => X"82", -- �
        16#9d4# => X"82", -- �
        16#ad4# => X"7c", -- �
        16#bd4# => X"00", -- �
        16#cd4# => X"00", -- �
        16#0d5# => X"00", -- �
        16#1d5# => X"64", -- �
        16#2d5# => X"98", -- �
        16#3d5# => X"00", -- �
        16#4d5# => X"7c", -- �
        16#5d5# => X"82", -- �
        16#6d5# => X"82", -- �
        16#7d5# => X"82", -- �
        16#8d5# => X"82", -- �
        16#9d5# => X"82", -- �
        16#ad5# => X"7c", -- �
        16#bd5# => X"00", -- �
        16#cd5# => X"00", -- �
        16#0d6# => X"00", -- �
        16#1d6# => X"44", -- �
        16#2d6# => X"44", -- �
        16#3d6# => X"00", -- �
        16#4d6# => X"7c", -- �
        16#5d6# => X"82", -- �
        16#6d6# => X"82", -- �
        16#7d6# => X"82", -- �
        16#8d6# => X"82", -- �
        16#9d6# => X"82", -- �
        16#ad6# => X"7c", -- �
        16#bd6# => X"00", -- �
        16#cd6# => X"00", -- �
        16#0d7# => X"00", -- �
        16#1d7# => X"00", -- �
        16#2d7# => X"00", -- �
        16#3d7# => X"00", -- �
        16#4d7# => X"42", -- �
        16#5d7# => X"24", -- �
        16#6d7# => X"18", -- �
        16#7d7# => X"18", -- �
        16#8d7# => X"24", -- �
        16#9d7# => X"42", -- �
        16#ad7# => X"00", -- �
        16#bd7# => X"00", -- �
        16#cd7# => X"00", -- �
        16#0d8# => X"00", -- �
        16#1d8# => X"02", -- �
        16#2d8# => X"3c", -- �
        16#3d8# => X"46", -- �
        16#4d8# => X"4a", -- �
        16#5d8# => X"4a", -- �
        16#6d8# => X"52", -- �
        16#7d8# => X"52", -- �
        16#8d8# => X"52", -- �
        16#9d8# => X"62", -- �
        16#ad8# => X"3c", -- �
        16#bd8# => X"40", -- �
        16#cd8# => X"00", -- �
        16#0d9# => X"00", -- �
        16#1d9# => X"20", -- �
        16#2d9# => X"10", -- �
        16#3d9# => X"00", -- �
        16#4d9# => X"42", -- �
        16#5d9# => X"42", -- �
        16#6d9# => X"42", -- �
        16#7d9# => X"42", -- �
        16#8d9# => X"42", -- �
        16#9d9# => X"42", -- �
        16#ad9# => X"3c", -- �
        16#bd9# => X"00", -- �
        16#cd9# => X"00", -- �
        16#0da# => X"00", -- �
        16#1da# => X"08", -- �
        16#2da# => X"10", -- �
        16#3da# => X"00", -- �
        16#4da# => X"42", -- �
        16#5da# => X"42", -- �
        16#6da# => X"42", -- �
        16#7da# => X"42", -- �
        16#8da# => X"42", -- �
        16#9da# => X"42", -- �
        16#ada# => X"3c", -- �
        16#bda# => X"00", -- �
        16#cda# => X"00", -- �
        16#0db# => X"00", -- �
        16#1db# => X"18", -- �
        16#2db# => X"24", -- �
        16#3db# => X"00", -- �
        16#4db# => X"42", -- �
        16#5db# => X"42", -- �
        16#6db# => X"42", -- �
        16#7db# => X"42", -- �
        16#8db# => X"42", -- �
        16#9db# => X"42", -- �
        16#adb# => X"3c", -- �
        16#bdb# => X"00", -- �
        16#cdb# => X"00", -- �
        16#0dc# => X"00", -- �
        16#1dc# => X"24", -- �
        16#2dc# => X"24", -- �
        16#3dc# => X"00", -- �
        16#4dc# => X"42", -- �
        16#5dc# => X"42", -- �
        16#6dc# => X"42", -- �
        16#7dc# => X"42", -- �
        16#8dc# => X"42", -- �
        16#9dc# => X"42", -- �
        16#adc# => X"3c", -- �
        16#bdc# => X"00", -- �
        16#cdc# => X"00", -- �
        16#0dd# => X"00", -- �
        16#1dd# => X"08", -- �
        16#2dd# => X"10", -- �
        16#3dd# => X"00", -- �
        16#4dd# => X"44", -- �
        16#5dd# => X"44", -- �
        16#6dd# => X"28", -- �
        16#7dd# => X"10", -- �
        16#8dd# => X"10", -- �
        16#9dd# => X"10", -- �
        16#add# => X"10", -- �
        16#bdd# => X"00", -- �
        16#cdd# => X"00", -- �
        16#0de# => X"00", -- �
        16#1de# => X"00", -- �
        16#2de# => X"40", -- �
        16#3de# => X"7c", -- �
        16#4de# => X"42", -- �
        16#5de# => X"42", -- �
        16#6de# => X"42", -- �
        16#7de# => X"7c", -- �
        16#8de# => X"40", -- �
        16#9de# => X"40", -- �
        16#ade# => X"40", -- �
        16#bde# => X"00", -- �
        16#cde# => X"00", -- �
        16#0df# => X"00", -- �
        16#1df# => X"00", -- �
        16#2df# => X"38", -- �
        16#3df# => X"44", -- �
        16#4df# => X"44", -- �
        16#5df# => X"48", -- �
        16#6df# => X"50", -- �
        16#7df# => X"4c", -- �
        16#8df# => X"42", -- �
        16#9df# => X"42", -- �
        16#adf# => X"5c", -- �
        16#bdf# => X"00", -- �
        16#cdf# => X"00", -- �
        16#0e0# => X"00", -- �
        16#1e0# => X"00", -- �
        16#2e0# => X"10", -- �
        16#3e0# => X"08", -- �
        16#4e0# => X"00", -- �
        16#5e0# => X"3c", -- �
        16#6e0# => X"02", -- �
        16#7e0# => X"3e", -- �
        16#8e0# => X"42", -- �
        16#9e0# => X"46", -- �
        16#ae0# => X"3a", -- �
        16#be0# => X"00", -- �
        16#ce0# => X"00", -- �
        16#0e1# => X"00", -- �
        16#1e1# => X"00", -- �
        16#2e1# => X"04", -- �
        16#3e1# => X"08", -- �
        16#4e1# => X"00", -- �
        16#5e1# => X"3c", -- �
        16#6e1# => X"02", -- �
        16#7e1# => X"3e", -- �
        16#8e1# => X"42", -- �
        16#9e1# => X"46", -- �
        16#ae1# => X"3a", -- �
        16#be1# => X"00", -- �
        16#ce1# => X"00", -- �
        16#0e2# => X"00", -- �
        16#1e2# => X"00", -- �
        16#2e2# => X"18", -- �
        16#3e2# => X"24", -- �
        16#4e2# => X"00", -- �
        16#5e2# => X"3c", -- �
        16#6e2# => X"02", -- �
        16#7e2# => X"3e", -- �
        16#8e2# => X"42", -- �
        16#9e2# => X"46", -- �
        16#ae2# => X"3a", -- �
        16#be2# => X"00", -- �
        16#ce2# => X"00", -- �
        16#0e3# => X"00", -- �
        16#1e3# => X"00", -- �
        16#2e3# => X"32", -- �
        16#3e3# => X"4c", -- �
        16#4e3# => X"00", -- �
        16#5e3# => X"3c", -- �
        16#6e3# => X"02", -- �
        16#7e3# => X"3e", -- �
        16#8e3# => X"42", -- �
        16#9e3# => X"46", -- �
        16#ae3# => X"3a", -- �
        16#be3# => X"00", -- �
        16#ce3# => X"00", -- �
        16#0e4# => X"00", -- �
        16#1e4# => X"00", -- �
        16#2e4# => X"24", -- �
        16#3e4# => X"24", -- �
        16#4e4# => X"00", -- �
        16#5e4# => X"3c", -- �
        16#6e4# => X"02", -- �
        16#7e4# => X"3e", -- �
        16#8e4# => X"42", -- �
        16#9e4# => X"46", -- �
        16#ae4# => X"3a", -- �
        16#be4# => X"00", -- �
        16#ce4# => X"00", -- �
        16#0e5# => X"00", -- �
        16#1e5# => X"18", -- �
        16#2e5# => X"24", -- �
        16#3e5# => X"18", -- �
        16#4e5# => X"00", -- �
        16#5e5# => X"3c", -- �
        16#6e5# => X"02", -- �
        16#7e5# => X"3e", -- �
        16#8e5# => X"42", -- �
        16#9e5# => X"46", -- �
        16#ae5# => X"3a", -- �
        16#be5# => X"00", -- �
        16#ce5# => X"00", -- �
        16#0e6# => X"00", -- �
        16#1e6# => X"00", -- �
        16#2e6# => X"00", -- �
        16#3e6# => X"00", -- �
        16#4e6# => X"00", -- �
        16#5e6# => X"6c", -- �
        16#6e6# => X"12", -- �
        16#7e6# => X"7c", -- �
        16#8e6# => X"90", -- �
        16#9e6# => X"92", -- �
        16#ae6# => X"6c", -- �
        16#be6# => X"00", -- �
        16#ce6# => X"00", -- �
        16#0e7# => X"00", -- �
        16#1e7# => X"00", -- �
        16#2e7# => X"00", -- �
        16#3e7# => X"00", -- �
        16#4e7# => X"00", -- �
        16#5e7# => X"3c", -- �
        16#6e7# => X"42", -- �
        16#7e7# => X"40", -- �
        16#8e7# => X"40", -- �
        16#9e7# => X"42", -- �
        16#ae7# => X"3c", -- �
        16#be7# => X"08", -- �
        16#ce7# => X"10", -- �
        16#0e8# => X"00", -- �
        16#1e8# => X"00", -- �
        16#2e8# => X"10", -- �
        16#3e8# => X"08", -- �
        16#4e8# => X"00", -- �
        16#5e8# => X"3c", -- �
        16#6e8# => X"42", -- �
        16#7e8# => X"7e", -- �
        16#8e8# => X"40", -- �
        16#9e8# => X"42", -- �
        16#ae8# => X"3c", -- �
        16#be8# => X"00", -- �
        16#ce8# => X"00", -- �
        16#0e9# => X"00", -- �
        16#1e9# => X"00", -- �
        16#2e9# => X"08", -- �
        16#3e9# => X"10", -- �
        16#4e9# => X"00", -- �
        16#5e9# => X"3c", -- �
        16#6e9# => X"42", -- �
        16#7e9# => X"7e", -- �
        16#8e9# => X"40", -- �
        16#9e9# => X"42", -- �
        16#ae9# => X"3c", -- �
        16#be9# => X"00", -- �
        16#ce9# => X"00", -- �
        16#0ea# => X"00", -- �
        16#1ea# => X"00", -- �
        16#2ea# => X"18", -- �
        16#3ea# => X"24", -- �
        16#4ea# => X"00", -- �
        16#5ea# => X"3c", -- �
        16#6ea# => X"42", -- �
        16#7ea# => X"7e", -- �
        16#8ea# => X"40", -- �
        16#9ea# => X"42", -- �
        16#aea# => X"3c", -- �
        16#bea# => X"00", -- �
        16#cea# => X"00", -- �
        16#0eb# => X"00", -- �
        16#1eb# => X"00", -- �
        16#2eb# => X"24", -- �
        16#3eb# => X"24", -- �
        16#4eb# => X"00", -- �
        16#5eb# => X"3c", -- �
        16#6eb# => X"42", -- �
        16#7eb# => X"7e", -- �
        16#8eb# => X"40", -- �
        16#9eb# => X"42", -- �
        16#aeb# => X"3c", -- �
        16#beb# => X"00", -- �
        16#ceb# => X"00", -- �
        16#0ec# => X"00", -- �
        16#1ec# => X"00", -- �
        16#2ec# => X"20", -- �
        16#3ec# => X"10", -- �
        16#4ec# => X"00", -- �
        16#5ec# => X"30", -- �
        16#6ec# => X"10", -- �
        16#7ec# => X"10", -- �
        16#8ec# => X"10", -- �
        16#9ec# => X"10", -- �
        16#aec# => X"7c", -- �
        16#bec# => X"00", -- �
        16#cec# => X"00", -- �
        16#0ed# => X"00", -- �
        16#1ed# => X"00", -- �
        16#2ed# => X"10", -- �
        16#3ed# => X"20", -- �
        16#4ed# => X"00", -- �
        16#5ed# => X"30", -- �
        16#6ed# => X"10", -- �
        16#7ed# => X"10", -- �
        16#8ed# => X"10", -- �
        16#9ed# => X"10", -- �
        16#aed# => X"7c", -- �
        16#bed# => X"00", -- �
        16#ced# => X"00", -- �
        16#0ee# => X"00", -- �
        16#1ee# => X"00", -- �
        16#2ee# => X"30", -- �
        16#3ee# => X"48", -- �
        16#4ee# => X"00", -- �
        16#5ee# => X"30", -- �
        16#6ee# => X"10", -- �
        16#7ee# => X"10", -- �
        16#8ee# => X"10", -- �
        16#9ee# => X"10", -- �
        16#aee# => X"7c", -- �
        16#bee# => X"00", -- �
        16#cee# => X"00", -- �
        16#0ef# => X"00", -- �
        16#1ef# => X"00", -- �
        16#2ef# => X"48", -- �
        16#3ef# => X"48", -- �
        16#4ef# => X"00", -- �
        16#5ef# => X"30", -- �
        16#6ef# => X"10", -- �
        16#7ef# => X"10", -- �
        16#8ef# => X"10", -- �
        16#9ef# => X"10", -- �
        16#aef# => X"7c", -- �
        16#bef# => X"00", -- �
        16#cef# => X"00", -- �
        16#0f0# => X"00", -- �
        16#1f0# => X"24", -- �
        16#2f0# => X"18", -- �
        16#3f0# => X"28", -- �
        16#4f0# => X"04", -- �
        16#5f0# => X"3c", -- �
        16#6f0# => X"42", -- �
        16#7f0# => X"42", -- �
        16#8f0# => X"42", -- �
        16#9f0# => X"42", -- �
        16#af0# => X"3c", -- �
        16#bf0# => X"00", -- �
        16#cf0# => X"00", -- �
        16#0f1# => X"00", -- �
        16#1f1# => X"00", -- �
        16#2f1# => X"32", -- �
        16#3f1# => X"4c", -- �
        16#4f1# => X"00", -- �
        16#5f1# => X"5c", -- �
        16#6f1# => X"62", -- �
        16#7f1# => X"42", -- �
        16#8f1# => X"42", -- �
        16#9f1# => X"42", -- �
        16#af1# => X"42", -- �
        16#bf1# => X"00", -- �
        16#cf1# => X"00", -- �
        16#0f2# => X"00", -- �
        16#1f2# => X"00", -- �
        16#2f2# => X"20", -- �
        16#3f2# => X"10", -- �
        16#4f2# => X"00", -- �
        16#5f2# => X"3c", -- �
        16#6f2# => X"42", -- �
        16#7f2# => X"42", -- �
        16#8f2# => X"42", -- �
        16#9f2# => X"42", -- �
        16#af2# => X"3c", -- �
        16#bf2# => X"00", -- �
        16#cf2# => X"00", -- �
        16#0f3# => X"00", -- �
        16#1f3# => X"00", -- �
        16#2f3# => X"08", -- �
        16#3f3# => X"10", -- �
        16#4f3# => X"00", -- �
        16#5f3# => X"3c", -- �
        16#6f3# => X"42", -- �
        16#7f3# => X"42", -- �
        16#8f3# => X"42", -- �
        16#9f3# => X"42", -- �
        16#af3# => X"3c", -- �
        16#bf3# => X"00", -- �
        16#cf3# => X"00", -- �
        16#0f4# => X"00", -- �
        16#1f4# => X"00", -- �
        16#2f4# => X"18", -- �
        16#3f4# => X"24", -- �
        16#4f4# => X"00", -- �
        16#5f4# => X"3c", -- �
        16#6f4# => X"42", -- �
        16#7f4# => X"42", -- �
        16#8f4# => X"42", -- �
        16#9f4# => X"42", -- �
        16#af4# => X"3c", -- �
        16#bf4# => X"00", -- �
        16#cf4# => X"00", -- �
        16#0f5# => X"00", -- �
        16#1f5# => X"00", -- �
        16#2f5# => X"32", -- �
        16#3f5# => X"4c", -- �
        16#4f5# => X"00", -- �
        16#5f5# => X"3c", -- �
        16#6f5# => X"42", -- �
        16#7f5# => X"42", -- �
        16#8f5# => X"42", -- �
        16#9f5# => X"42", -- �
        16#af5# => X"3c", -- �
        16#bf5# => X"00", -- �
        16#cf5# => X"00", -- �
        16#0f6# => X"00", -- �
        16#1f6# => X"00", -- �
        16#2f6# => X"24", -- �
        16#3f6# => X"24", -- �
        16#4f6# => X"00", -- �
        16#5f6# => X"3c", -- �
        16#6f6# => X"42", -- �
        16#7f6# => X"42", -- �
        16#8f6# => X"42", -- �
        16#9f6# => X"42", -- �
        16#af6# => X"3c", -- �
        16#bf6# => X"00", -- �
        16#cf6# => X"00", -- �
        16#0f7# => X"00", -- �
        16#1f7# => X"00", -- �
        16#2f7# => X"00", -- �
        16#3f7# => X"10", -- �
        16#4f7# => X"10", -- �
        16#5f7# => X"00", -- �
        16#6f7# => X"7c", -- �
        16#7f7# => X"00", -- �
        16#8f7# => X"10", -- �
        16#9f7# => X"10", -- �
        16#af7# => X"00", -- �
        16#bf7# => X"00", -- �
        16#cf7# => X"00", -- �
        16#0f8# => X"00", -- �
        16#1f8# => X"00", -- �
        16#2f8# => X"00", -- �
        16#3f8# => X"00", -- �
        16#4f8# => X"02", -- �
        16#5f8# => X"3c", -- �
        16#6f8# => X"46", -- �
        16#7f8# => X"4a", -- �
        16#8f8# => X"52", -- �
        16#9f8# => X"62", -- �
        16#af8# => X"3c", -- �
        16#bf8# => X"40", -- �
        16#cf8# => X"00", -- �
        16#0f9# => X"00", -- �
        16#1f9# => X"00", -- �
        16#2f9# => X"20", -- �
        16#3f9# => X"10", -- �
        16#4f9# => X"00", -- �
        16#5f9# => X"44", -- �
        16#6f9# => X"44", -- �
        16#7f9# => X"44", -- �
        16#8f9# => X"44", -- �
        16#9f9# => X"44", -- �
        16#af9# => X"3a", -- �
        16#bf9# => X"00", -- �
        16#cf9# => X"00", -- �
        16#0fa# => X"00", -- �
        16#1fa# => X"00", -- �
        16#2fa# => X"08", -- �
        16#3fa# => X"10", -- �
        16#4fa# => X"00", -- �
        16#5fa# => X"44", -- �
        16#6fa# => X"44", -- �
        16#7fa# => X"44", -- �
        16#8fa# => X"44", -- �
        16#9fa# => X"44", -- �
        16#afa# => X"3a", -- �
        16#bfa# => X"00", -- �
        16#cfa# => X"00", -- �
        16#0fb# => X"00", -- �
        16#1fb# => X"00", -- �
        16#2fb# => X"18", -- �
        16#3fb# => X"24", -- �
        16#4fb# => X"00", -- �
        16#5fb# => X"44", -- �
        16#6fb# => X"44", -- �
        16#7fb# => X"44", -- �
        16#8fb# => X"44", -- �
        16#9fb# => X"44", -- �
        16#afb# => X"3a", -- �
        16#bfb# => X"00", -- �
        16#cfb# => X"00", -- �
        16#0fc# => X"00", -- �
        16#1fc# => X"00", -- �
        16#2fc# => X"28", -- �
        16#3fc# => X"28", -- �
        16#4fc# => X"00", -- �
        16#5fc# => X"44", -- �
        16#6fc# => X"44", -- �
        16#7fc# => X"44", -- �
        16#8fc# => X"44", -- �
        16#9fc# => X"44", -- �
        16#afc# => X"3a", -- �
        16#bfc# => X"00", -- �
        16#cfc# => X"00", -- �
        16#0fd# => X"00", -- �
        16#1fd# => X"00", -- �
        16#2fd# => X"08", -- �
        16#3fd# => X"10", -- �
        16#4fd# => X"00", -- �
        16#5fd# => X"42", -- �
        16#6fd# => X"42", -- �
        16#7fd# => X"42", -- �
        16#8fd# => X"46", -- �
        16#9fd# => X"3a", -- �
        16#afd# => X"02", -- �
        16#bfd# => X"42", -- �
        16#cfd# => X"3c", -- �
        16#0fe# => X"00", -- �
        16#1fe# => X"00", -- �
        16#2fe# => X"00", -- �
        16#3fe# => X"40", -- �
        16#4fe# => X"40", -- �
        16#5fe# => X"5c", -- �
        16#6fe# => X"62", -- �
        16#7fe# => X"42", -- �
        16#8fe# => X"42", -- �
        16#9fe# => X"62", -- �
        16#afe# => X"5c", -- �
        16#bfe# => X"40", -- �
        16#cfe# => X"40", -- �
        16#0ff# => X"00", -- �
        16#1ff# => X"00", -- �
        16#2ff# => X"24", -- �
        16#3ff# => X"24", -- �
        16#4ff# => X"00", -- �
        16#5ff# => X"42", -- �
        16#6ff# => X"42", -- �
        16#7ff# => X"42", -- �
        16#8ff# => X"46", -- �
        16#9ff# => X"3a", -- �
        16#aff# => X"02", -- �
        16#bff# => X"42", -- �
        16#cff# => X"3c", -- �
        others  => x"00"
    );

begin
    process
    begin
        wait until rising_edge( clk);
        if not is_x( addr) then -- avoid simulation warnings
            data <= rom( to_integer( unsigned( addr)));
        end if;
    end process;
end rtl;

