-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0b98b00c",
     3 => x"3a0b0b0b",
     4 => x"95bc0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0b95fc2d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0b98",
   162 => x"9c738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0b91",
   171 => x"c02d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0b92",
   179 => x"f22d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0b98ac0c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81f33f8f",
   257 => x"9c3f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"53510498",
   280 => x"ac08802e",
   281 => x"a13898b0",
   282 => x"08822eb9",
   283 => x"38838080",
   284 => x"0b0b0b0b",
   285 => x"9fe00c82",
   286 => x"a0800b9f",
   287 => x"e40c8290",
   288 => x"800b9fe8",
   289 => x"0c04f880",
   290 => x"8080a40b",
   291 => x"0b0b0b9f",
   292 => x"e00cf880",
   293 => x"8082800b",
   294 => x"9fe40cf8",
   295 => x"80808480",
   296 => x"0b9fe80c",
   297 => x"0480c0a8",
   298 => x"808c0b0b",
   299 => x"0b0b9fe0",
   300 => x"0c80c0a8",
   301 => x"80940b9f",
   302 => x"e40c0b0b",
   303 => x"0b97cc0b",
   304 => x"9fe80c04",
   305 => x"ff3d0d9f",
   306 => x"ec335170",
   307 => x"a33898b8",
   308 => x"08700852",
   309 => x"5270802e",
   310 => x"92388412",
   311 => x"98b80c70",
   312 => x"2d98b808",
   313 => x"70085252",
   314 => x"70f03881",
   315 => x"0b9fec34",
   316 => x"833d0d04",
   317 => x"04803d0d",
   318 => x"0b0b0b9f",
   319 => x"dc08802e",
   320 => x"8e380b0b",
   321 => x"0b0b800b",
   322 => x"802e0981",
   323 => x"06853882",
   324 => x"3d0d040b",
   325 => x"0b0b9fdc",
   326 => x"510b0b0b",
   327 => x"f5e23f82",
   328 => x"3d0d0404",
   329 => x"fd3d0d98",
   330 => x"c00876b0",
   331 => x"ea299412",
   332 => x"0c54850b",
   333 => x"98150c98",
   334 => x"14087081",
   335 => x"06515372",
   336 => x"f638853d",
   337 => x"0d04ff3d",
   338 => x"0d98c008",
   339 => x"74101075",
   340 => x"10059412",
   341 => x"0c52850b",
   342 => x"98130c98",
   343 => x"12087081",
   344 => x"06515170",
   345 => x"f638833d",
   346 => x"0d04803d",
   347 => x"0d725180",
   348 => x"71278738",
   349 => x"ff115170",
   350 => x"fb38823d",
   351 => x"0d04803d",
   352 => x"0d98c008",
   353 => x"51870b84",
   354 => x"120c823d",
   355 => x"0d04803d",
   356 => x"0d98c408",
   357 => x"51b60b8c",
   358 => x"120c830b",
   359 => x"88120c82",
   360 => x"3d0d04ff",
   361 => x"3d0d98c4",
   362 => x"08528412",
   363 => x"08708106",
   364 => x"51517080",
   365 => x"2ef43871",
   366 => x"087081ff",
   367 => x"06800c51",
   368 => x"833d0d04",
   369 => x"fe3d0d02",
   370 => x"93053398",
   371 => x"c4085353",
   372 => x"84120870",
   373 => x"892a7081",
   374 => x"06515151",
   375 => x"70f23872",
   376 => x"720c843d",
   377 => x"0d04fe3d",
   378 => x"0d029305",
   379 => x"3353728a",
   380 => x"2e9b3898",
   381 => x"c4085284",
   382 => x"12087089",
   383 => x"2a708106",
   384 => x"51515170",
   385 => x"f2387272",
   386 => x"0c843d0d",
   387 => x"0498c408",
   388 => x"52841208",
   389 => x"70892a70",
   390 => x"81065151",
   391 => x"5170f238",
   392 => x"8d720c84",
   393 => x"12087089",
   394 => x"2a708106",
   395 => x"51515170",
   396 => x"c638d339",
   397 => x"fd3d0d75",
   398 => x"70335254",
   399 => x"70802ea7",
   400 => x"387098c4",
   401 => x"08535381",
   402 => x"1454728a",
   403 => x"2e9d3884",
   404 => x"12087089",
   405 => x"2a708106",
   406 => x"51515170",
   407 => x"f2387272",
   408 => x"0c733353",
   409 => x"72e13885",
   410 => x"3d0d0484",
   411 => x"12087089",
   412 => x"2a708106",
   413 => x"51515170",
   414 => x"f2388d72",
   415 => x"0c841208",
   416 => x"70892a70",
   417 => x"81065151",
   418 => x"5170c438",
   419 => x"d139803d",
   420 => x"0d98bc08",
   421 => x"5181ff0b",
   422 => x"88120c82",
   423 => x"3d0d04fb",
   424 => x"3d0d8880",
   425 => x"e0870b98",
   426 => x"bc0898c0",
   427 => x"08728413",
   428 => x"0c565755",
   429 => x"afd7c20b",
   430 => x"94150c85",
   431 => x"0b98150c",
   432 => x"98140870",
   433 => x"81065153",
   434 => x"72f63874",
   435 => x"9f2a7510",
   436 => x"07708418",
   437 => x"0c55afd7",
   438 => x"c20b9415",
   439 => x"0c850b98",
   440 => x"150cdd39",
   441 => x"fe3d0d98",
   442 => x"c4085284",
   443 => x"12088106",
   444 => x"5170802e",
   445 => x"f6387108",
   446 => x"7081ff06",
   447 => x"54518412",
   448 => x"0870892a",
   449 => x"70810651",
   450 => x"515170f2",
   451 => x"38ab720c",
   452 => x"728a2ea6",
   453 => x"38841208",
   454 => x"70892a70",
   455 => x"81065151",
   456 => x"5170f238",
   457 => x"72720c84",
   458 => x"12087089",
   459 => x"2a810651",
   460 => x"5372f438",
   461 => x"ad720cff",
   462 => x"b2398412",
   463 => x"0870892a",
   464 => x"70810651",
   465 => x"515170f2",
   466 => x"388d720c",
   467 => x"84120870",
   468 => x"892a7081",
   469 => x"06515151",
   470 => x"70ffba38",
   471 => x"c739ff3d",
   472 => x"0d98bc08",
   473 => x"52710870",
   474 => x"8f067071",
   475 => x"842b0784",
   476 => x"150c5151",
   477 => x"7108708f",
   478 => x"06707184",
   479 => x"2b078415",
   480 => x"0c5151e1",
   481 => x"39fb3d0d",
   482 => x"98c00853",
   483 => x"870b8414",
   484 => x"0c98c408",
   485 => x"54b60b8c",
   486 => x"150c830b",
   487 => x"88150c97",
   488 => x"d00b97d0",
   489 => x"33545672",
   490 => x"802ea438",
   491 => x"72558116",
   492 => x"56748a2e",
   493 => x"819f3884",
   494 => x"14087089",
   495 => x"2a708106",
   496 => x"51515372",
   497 => x"f2387474",
   498 => x"0c753355",
   499 => x"74e03897",
   500 => x"e80b97e8",
   501 => x"33545672",
   502 => x"802ea438",
   503 => x"72558116",
   504 => x"56748a2e",
   505 => x"81943884",
   506 => x"14087089",
   507 => x"2a708106",
   508 => x"51515372",
   509 => x"f2387474",
   510 => x"0c753355",
   511 => x"74e03898",
   512 => x"bc085581",
   513 => x"ff0b8816",
   514 => x"0c841408",
   515 => x"81065675",
   516 => x"802ef638",
   517 => x"73087081",
   518 => x"ff065656",
   519 => x"84140870",
   520 => x"892a8106",
   521 => x"515372f4",
   522 => x"38ab740c",
   523 => x"748a2e80",
   524 => x"ee388414",
   525 => x"0870892a",
   526 => x"81065153",
   527 => x"72f43874",
   528 => x"740c8414",
   529 => x"0870892a",
   530 => x"81065653",
   531 => x"74f438ad",
   532 => x"740cffb5",
   533 => x"39841408",
   534 => x"70892a70",
   535 => x"81065151",
   536 => x"5372f238",
   537 => x"8d740c84",
   538 => x"14087089",
   539 => x"2a708106",
   540 => x"51515372",
   541 => x"fec138fe",
   542 => x"cd398414",
   543 => x"0870892a",
   544 => x"70810651",
   545 => x"515372f2",
   546 => x"388d740c",
   547 => x"84140870",
   548 => x"892a7081",
   549 => x"06515153",
   550 => x"72fecc38",
   551 => x"fed83984",
   552 => x"14087089",
   553 => x"2a810651",
   554 => x"5675f438",
   555 => x"8d740c84",
   556 => x"14087089",
   557 => x"2a810651",
   558 => x"5372fef6",
   559 => x"38ff8039",
   560 => x"8c08028c",
   561 => x"0cf93d0d",
   562 => x"800b8c08",
   563 => x"fc050c8c",
   564 => x"08880508",
   565 => x"8025ab38",
   566 => x"8c088805",
   567 => x"08308c08",
   568 => x"88050c80",
   569 => x"0b8c08f4",
   570 => x"050c8c08",
   571 => x"fc050888",
   572 => x"38810b8c",
   573 => x"08f4050c",
   574 => x"8c08f405",
   575 => x"088c08fc",
   576 => x"050c8c08",
   577 => x"8c050880",
   578 => x"25ab388c",
   579 => x"088c0508",
   580 => x"308c088c",
   581 => x"050c800b",
   582 => x"8c08f005",
   583 => x"0c8c08fc",
   584 => x"05088838",
   585 => x"810b8c08",
   586 => x"f0050c8c",
   587 => x"08f00508",
   588 => x"8c08fc05",
   589 => x"0c80538c",
   590 => x"088c0508",
   591 => x"528c0888",
   592 => x"05085181",
   593 => x"a73f8008",
   594 => x"708c08f8",
   595 => x"050c548c",
   596 => x"08fc0508",
   597 => x"802e8c38",
   598 => x"8c08f805",
   599 => x"08308c08",
   600 => x"f8050c8c",
   601 => x"08f80508",
   602 => x"70800c54",
   603 => x"893d0d8c",
   604 => x"0c048c08",
   605 => x"028c0cfb",
   606 => x"3d0d800b",
   607 => x"8c08fc05",
   608 => x"0c8c0888",
   609 => x"05088025",
   610 => x"93388c08",
   611 => x"88050830",
   612 => x"8c088805",
   613 => x"0c810b8c",
   614 => x"08fc050c",
   615 => x"8c088c05",
   616 => x"0880258c",
   617 => x"388c088c",
   618 => x"0508308c",
   619 => x"088c050c",
   620 => x"81538c08",
   621 => x"8c050852",
   622 => x"8c088805",
   623 => x"0851ad3f",
   624 => x"8008708c",
   625 => x"08f8050c",
   626 => x"548c08fc",
   627 => x"0508802e",
   628 => x"8c388c08",
   629 => x"f8050830",
   630 => x"8c08f805",
   631 => x"0c8c08f8",
   632 => x"05087080",
   633 => x"0c54873d",
   634 => x"0d8c0c04",
   635 => x"8c08028c",
   636 => x"0cfd3d0d",
   637 => x"810b8c08",
   638 => x"fc050c80",
   639 => x"0b8c08f8",
   640 => x"050c8c08",
   641 => x"8c05088c",
   642 => x"08880508",
   643 => x"27ac388c",
   644 => x"08fc0508",
   645 => x"802ea338",
   646 => x"800b8c08",
   647 => x"8c050824",
   648 => x"99388c08",
   649 => x"8c050810",
   650 => x"8c088c05",
   651 => x"0c8c08fc",
   652 => x"0508108c",
   653 => x"08fc050c",
   654 => x"c9398c08",
   655 => x"fc050880",
   656 => x"2e80c938",
   657 => x"8c088c05",
   658 => x"088c0888",
   659 => x"050826a1",
   660 => x"388c0888",
   661 => x"05088c08",
   662 => x"8c050831",
   663 => x"8c088805",
   664 => x"0c8c08f8",
   665 => x"05088c08",
   666 => x"fc050807",
   667 => x"8c08f805",
   668 => x"0c8c08fc",
   669 => x"0508812a",
   670 => x"8c08fc05",
   671 => x"0c8c088c",
   672 => x"0508812a",
   673 => x"8c088c05",
   674 => x"0cffaf39",
   675 => x"8c089005",
   676 => x"08802e8f",
   677 => x"388c0888",
   678 => x"0508708c",
   679 => x"08f4050c",
   680 => x"518d398c",
   681 => x"08f80508",
   682 => x"708c08f4",
   683 => x"050c518c",
   684 => x"08f40508",
   685 => x"800c853d",
   686 => x"0d8c0c04",
   687 => x"fd3d0d80",
   688 => x"0b98b008",
   689 => x"54547281",
   690 => x"2e983873",
   691 => x"9ff00cf3",
   692 => x"8e3ff2ac",
   693 => x"3f98c852",
   694 => x"8151f9a9",
   695 => x"3f800851",
   696 => x"9e3f729f",
   697 => x"f00cf2f7",
   698 => x"3ff2953f",
   699 => x"98c85281",
   700 => x"51f9923f",
   701 => x"80085187",
   702 => x"3f00ff39",
   703 => x"00ff39f7",
   704 => x"3d0d7b98",
   705 => x"cc0882c8",
   706 => x"11085a54",
   707 => x"5a77802e",
   708 => x"80d93881",
   709 => x"88188419",
   710 => x"08ff0581",
   711 => x"712b5955",
   712 => x"59807424",
   713 => x"80e93880",
   714 => x"7424b538",
   715 => x"73822b78",
   716 => x"11880556",
   717 => x"56818019",
   718 => x"08770653",
   719 => x"72802eb5",
   720 => x"38781670",
   721 => x"08535379",
   722 => x"51740853",
   723 => x"722dff14",
   724 => x"fc17fc17",
   725 => x"79812c5a",
   726 => x"57575473",
   727 => x"8025d638",
   728 => x"77085877",
   729 => x"ffad3898",
   730 => x"cc0853bc",
   731 => x"1308a538",
   732 => x"7951ff85",
   733 => x"3f740853",
   734 => x"722dff14",
   735 => x"fc17fc17",
   736 => x"79812c5a",
   737 => x"57575473",
   738 => x"8025ffa9",
   739 => x"38d23980",
   740 => x"57ff9439",
   741 => x"7251bc13",
   742 => x"0853722d",
   743 => x"7951fed9",
   744 => x"3fff3d0d",
   745 => x"9fd00bfc",
   746 => x"05700852",
   747 => x"5270ff2e",
   748 => x"9138702d",
   749 => x"fc127008",
   750 => x"525270ff",
   751 => x"2e098106",
   752 => x"f138833d",
   753 => x"0d0404f1",
   754 => x"fb3f0400",
   755 => x"00000040",
   756 => x"536f432c",
   757 => x"205a5055",
   758 => x"20746573",
   759 => x"74207072",
   760 => x"6f677261",
   761 => x"6d0a0000",
   762 => x"636f6d70",
   763 => x"696c6564",
   764 => x"3a204175",
   765 => x"67202035",
   766 => x"20323031",
   767 => x"30202020",
   768 => x"31313a30",
   769 => x"393a3436",
   770 => x"0a000000",
   771 => x"64756d6d",
   772 => x"792e6578",
   773 => x"65000000",
   774 => x"43000000",
   775 => x"00ffffff",
   776 => x"ff00ffff",
   777 => x"ffff00ff",
   778 => x"ffffff00",
   779 => x"00000000",
   780 => x"00000000",
   781 => x"00000000",
   782 => x"00000fd8",
   783 => x"80000800",
   784 => x"80000200",
   785 => x"80000100",
   786 => x"00000c0c",
   787 => x"00000c50",
   788 => x"00000000",
   789 => x"00000eb8",
   790 => x"00000f14",
   791 => x"00000f70",
   792 => x"00000000",
   793 => x"00000000",
   794 => x"00000000",
   795 => x"00000000",
   796 => x"00000000",
   797 => x"00000000",
   798 => x"00000000",
   799 => x"00000000",
   800 => x"00000000",
   801 => x"00000c18",
   802 => x"00000000",
   803 => x"00000000",
   804 => x"00000000",
   805 => x"00000000",
   806 => x"00000000",
   807 => x"00000000",
   808 => x"00000000",
   809 => x"00000000",
   810 => x"00000000",
   811 => x"00000000",
   812 => x"00000000",
   813 => x"00000000",
   814 => x"00000000",
   815 => x"00000000",
   816 => x"00000000",
   817 => x"00000000",
   818 => x"00000000",
   819 => x"00000000",
   820 => x"00000000",
   821 => x"00000000",
   822 => x"00000000",
   823 => x"00000000",
   824 => x"00000000",
   825 => x"00000000",
   826 => x"00000000",
   827 => x"00000000",
   828 => x"00000000",
   829 => x"00000000",
   830 => x"00000001",
   831 => x"330eabcd",
   832 => x"1234e66d",
   833 => x"deec0005",
   834 => x"000b0000",
   835 => x"00000000",
   836 => x"00000000",
   837 => x"00000000",
   838 => x"00000000",
   839 => x"00000000",
   840 => x"00000000",
   841 => x"00000000",
   842 => x"00000000",
   843 => x"00000000",
   844 => x"00000000",
   845 => x"00000000",
   846 => x"00000000",
   847 => x"00000000",
   848 => x"00000000",
   849 => x"00000000",
   850 => x"00000000",
   851 => x"00000000",
   852 => x"00000000",
   853 => x"00000000",
   854 => x"00000000",
   855 => x"00000000",
   856 => x"00000000",
   857 => x"00000000",
   858 => x"00000000",
   859 => x"00000000",
   860 => x"00000000",
   861 => x"00000000",
   862 => x"00000000",
   863 => x"00000000",
   864 => x"00000000",
   865 => x"00000000",
   866 => x"00000000",
   867 => x"00000000",
   868 => x"00000000",
   869 => x"00000000",
   870 => x"00000000",
   871 => x"00000000",
   872 => x"00000000",
   873 => x"00000000",
   874 => x"00000000",
   875 => x"00000000",
   876 => x"00000000",
   877 => x"00000000",
   878 => x"00000000",
   879 => x"00000000",
   880 => x"00000000",
   881 => x"00000000",
   882 => x"00000000",
   883 => x"00000000",
   884 => x"00000000",
   885 => x"00000000",
   886 => x"00000000",
   887 => x"00000000",
   888 => x"00000000",
   889 => x"00000000",
   890 => x"00000000",
   891 => x"00000000",
   892 => x"00000000",
   893 => x"00000000",
   894 => x"00000000",
   895 => x"00000000",
   896 => x"00000000",
   897 => x"00000000",
   898 => x"00000000",
   899 => x"00000000",
   900 => x"00000000",
   901 => x"00000000",
   902 => x"00000000",
   903 => x"00000000",
   904 => x"00000000",
   905 => x"00000000",
   906 => x"00000000",
   907 => x"00000000",
   908 => x"00000000",
   909 => x"00000000",
   910 => x"00000000",
   911 => x"00000000",
   912 => x"00000000",
   913 => x"00000000",
   914 => x"00000000",
   915 => x"00000000",
   916 => x"00000000",
   917 => x"00000000",
   918 => x"00000000",
   919 => x"00000000",
   920 => x"00000000",
   921 => x"00000000",
   922 => x"00000000",
   923 => x"00000000",
   924 => x"00000000",
   925 => x"00000000",
   926 => x"00000000",
   927 => x"00000000",
   928 => x"00000000",
   929 => x"00000000",
   930 => x"00000000",
   931 => x"00000000",
   932 => x"00000000",
   933 => x"00000000",
   934 => x"00000000",
   935 => x"00000000",
   936 => x"00000000",
   937 => x"00000000",
   938 => x"00000000",
   939 => x"00000000",
   940 => x"00000000",
   941 => x"00000000",
   942 => x"00000000",
   943 => x"00000000",
   944 => x"00000000",
   945 => x"00000000",
   946 => x"00000000",
   947 => x"00000000",
   948 => x"00000000",
   949 => x"00000000",
   950 => x"00000000",
   951 => x"00000000",
   952 => x"00000000",
   953 => x"00000000",
   954 => x"00000000",
   955 => x"00000000",
   956 => x"00000000",
   957 => x"00000000",
   958 => x"00000000",
   959 => x"00000000",
   960 => x"00000000",
   961 => x"00000000",
   962 => x"00000000",
   963 => x"00000000",
   964 => x"00000000",
   965 => x"00000000",
   966 => x"00000000",
   967 => x"00000000",
   968 => x"00000000",
   969 => x"00000000",
   970 => x"00000000",
   971 => x"00000000",
   972 => x"00000000",
   973 => x"00000000",
   974 => x"00000000",
   975 => x"00000000",
   976 => x"00000000",
   977 => x"00000000",
   978 => x"00000000",
   979 => x"00000000",
   980 => x"00000000",
   981 => x"00000000",
   982 => x"00000000",
   983 => x"00000000",
   984 => x"00000000",
   985 => x"00000000",
   986 => x"00000000",
   987 => x"00000000",
   988 => x"00000000",
   989 => x"00000000",
   990 => x"00000000",
   991 => x"00000000",
   992 => x"00000000",
   993 => x"00000000",
   994 => x"00000000",
   995 => x"00000000",
   996 => x"00000000",
   997 => x"00000000",
   998 => x"00000000",
   999 => x"00000000",
  1000 => x"00000000",
  1001 => x"00000000",
  1002 => x"00000000",
  1003 => x"00000000",
  1004 => x"00000000",
  1005 => x"00000000",
  1006 => x"00000000",
  1007 => x"00000000",
  1008 => x"00000000",
  1009 => x"00000000",
  1010 => x"00000000",
  1011 => x"ffffffff",
  1012 => x"00000000",
  1013 => x"ffffffff",
  1014 => x"00000000",
  1015 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
