
----------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2010 Aeroflex Gaisler
----------------------------------------------------------------------------
-- Entity: 	ahbrom
-- File:	ahbrom.vhd
-- Author:	Jiri Gaisler - Gaisler Research
-- Description:	AHB rom. 0/1-waitstate read
----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
library grlib;
use grlib.amba.all;
use grlib.stdlib.all;
use grlib.devices.all;

entity ahbrom is
  generic (
    hindex  : integer := 0;
    haddr   : integer := 0;
    hmask   : integer := 16#fff#;
    pipe    : integer := 0;
    tech    : integer := 0;
    kbytes  : integer := 1);
  port (
    rst     : in  std_ulogic;
    clk     : in  std_ulogic;
    ahbsi   : in  ahb_slv_in_type;
    ahbso   : out ahb_slv_out_type
  );
end;

architecture rtl of ahbrom is
constant abits : integer := 15;
constant bytes : integer := 16436;

constant hconfig : ahb_config_type := (
  0 => ahb_device_reg ( VENDOR_GAISLER, GAISLER_AHBROM, 0, 0, 0),
  4 => ahb_membar(haddr, '1', '1', hmask), others => zero32);

signal romdata : std_logic_vector(31 downto 0);
signal addr : std_logic_vector(abits-1 downto 2);
signal hsel, hready : std_ulogic;

begin

  ahbso.hresp   <= "00"; 
  ahbso.hsplit  <= (others => '0'); 
  ahbso.hirq    <= (others => '0');
  ahbso.hcache  <= '1';
  ahbso.hconfig <= hconfig;
  ahbso.hindex  <= hindex;

  reg : process (clk)
  begin
    if rising_edge(clk) then 
      addr <= ahbsi.haddr(abits-1 downto 2);
    end if;
  end process;

  p0 : if pipe = 0 generate
    ahbso.hrdata  <= romdata;
    ahbso.hready  <= '1';
  end generate;

  p1 : if pipe = 1 generate
    reg2 : process (clk)
    begin
      if rising_edge(clk) then
	hsel <= ahbsi.hsel(hindex) and ahbsi.htrans(1);
	hready <= ahbsi.hready;
	ahbso.hready <=  (not rst) or (hsel and hready) or
	  (ahbsi.hsel(hindex) and not ahbsi.htrans(1) and ahbsi.hready);
	ahbso.hrdata  <= romdata;
      end if;
    end process;
  end generate;

  comb : process (addr)
  begin
    case conv_integer(addr) is
    when 16#00000# => romdata <= X"0B0B0B0B";
    when 16#00001# => romdata <= X"82700B0B";
    when 16#00002# => romdata <= X"80F0AC0C";
    when 16#00003# => romdata <= X"3A0B0B80";
    when 16#00004# => romdata <= X"E2D80400";
    when 16#00005# => romdata <= X"00000000";
    when 16#00006# => romdata <= X"00000000";
    when 16#00007# => romdata <= X"00000000";
    when 16#00008# => romdata <= X"0B0B0B89";
    when 16#00009# => romdata <= X"92040000";
    when 16#0000A# => romdata <= X"00000000";
    when 16#0000B# => romdata <= X"00000000";
    when 16#0000C# => romdata <= X"00000000";
    when 16#0000D# => romdata <= X"00000000";
    when 16#0000E# => romdata <= X"00000000";
    when 16#0000F# => romdata <= X"00000000";
    when 16#00010# => romdata <= X"71FD0608";
    when 16#00011# => romdata <= X"72830609";
    when 16#00012# => romdata <= X"81058205";
    when 16#00013# => romdata <= X"832B2A83";
    when 16#00014# => romdata <= X"FFFF0652";
    when 16#00015# => romdata <= X"04000000";
    when 16#00016# => romdata <= X"00000000";
    when 16#00017# => romdata <= X"00000000";
    when 16#00018# => romdata <= X"71FD0608";
    when 16#00019# => romdata <= X"83FFFF73";
    when 16#0001A# => romdata <= X"83060981";
    when 16#0001B# => romdata <= X"05820583";
    when 16#0001C# => romdata <= X"2B2B0906";
    when 16#0001D# => romdata <= X"7383FFFF";
    when 16#0001E# => romdata <= X"0B0B0B0B";
    when 16#0001F# => romdata <= X"83A70400";
    when 16#00020# => romdata <= X"72098105";
    when 16#00021# => romdata <= X"72057373";
    when 16#00022# => romdata <= X"09060906";
    when 16#00023# => romdata <= X"73097306";
    when 16#00024# => romdata <= X"070A8106";
    when 16#00025# => romdata <= X"53510400";
    when 16#00026# => romdata <= X"00000000";
    when 16#00027# => romdata <= X"00000000";
    when 16#00028# => romdata <= X"72722473";
    when 16#00029# => romdata <= X"732E0753";
    when 16#0002A# => romdata <= X"51040000";
    when 16#0002B# => romdata <= X"00000000";
    when 16#0002C# => romdata <= X"00000000";
    when 16#0002D# => romdata <= X"00000000";
    when 16#0002E# => romdata <= X"00000000";
    when 16#0002F# => romdata <= X"00000000";
    when 16#00030# => romdata <= X"71737109";
    when 16#00031# => romdata <= X"71068106";
    when 16#00032# => romdata <= X"30720A10";
    when 16#00033# => romdata <= X"0A720A10";
    when 16#00034# => romdata <= X"0A31050A";
    when 16#00035# => romdata <= X"81065151";
    when 16#00036# => romdata <= X"53510400";
    when 16#00037# => romdata <= X"00000000";
    when 16#00038# => romdata <= X"72722673";
    when 16#00039# => romdata <= X"732E0753";
    when 16#0003A# => romdata <= X"51040000";
    when 16#0003B# => romdata <= X"00000000";
    when 16#0003C# => romdata <= X"00000000";
    when 16#0003D# => romdata <= X"00000000";
    when 16#0003E# => romdata <= X"00000000";
    when 16#0003F# => romdata <= X"00000000";
    when 16#00040# => romdata <= X"00000000";
    when 16#00041# => romdata <= X"00000000";
    when 16#00042# => romdata <= X"00000000";
    when 16#00043# => romdata <= X"00000000";
    when 16#00044# => romdata <= X"00000000";
    when 16#00045# => romdata <= X"00000000";
    when 16#00046# => romdata <= X"00000000";
    when 16#00047# => romdata <= X"00000000";
    when 16#00048# => romdata <= X"0B0B0B88";
    when 16#00049# => romdata <= X"C4040000";
    when 16#0004A# => romdata <= X"00000000";
    when 16#0004B# => romdata <= X"00000000";
    when 16#0004C# => romdata <= X"00000000";
    when 16#0004D# => romdata <= X"00000000";
    when 16#0004E# => romdata <= X"00000000";
    when 16#0004F# => romdata <= X"00000000";
    when 16#00050# => romdata <= X"720A722B";
    when 16#00051# => romdata <= X"0A535104";
    when 16#00052# => romdata <= X"00000000";
    when 16#00053# => romdata <= X"00000000";
    when 16#00054# => romdata <= X"00000000";
    when 16#00055# => romdata <= X"00000000";
    when 16#00056# => romdata <= X"00000000";
    when 16#00057# => romdata <= X"00000000";
    when 16#00058# => romdata <= X"72729F06";
    when 16#00059# => romdata <= X"0981050B";
    when 16#0005A# => romdata <= X"0B0B88A7";
    when 16#0005B# => romdata <= X"05040000";
    when 16#0005C# => romdata <= X"00000000";
    when 16#0005D# => romdata <= X"00000000";
    when 16#0005E# => romdata <= X"00000000";
    when 16#0005F# => romdata <= X"00000000";
    when 16#00060# => romdata <= X"72722AFF";
    when 16#00061# => romdata <= X"739F062A";
    when 16#00062# => romdata <= X"0974090A";
    when 16#00063# => romdata <= X"8106FF05";
    when 16#00064# => romdata <= X"06075351";
    when 16#00065# => romdata <= X"04000000";
    when 16#00066# => romdata <= X"00000000";
    when 16#00067# => romdata <= X"00000000";
    when 16#00068# => romdata <= X"71715351";
    when 16#00069# => romdata <= X"020D0406";
    when 16#0006A# => romdata <= X"73830609";
    when 16#0006B# => romdata <= X"81058205";
    when 16#0006C# => romdata <= X"832B0B2B";
    when 16#0006D# => romdata <= X"0772FC06";
    when 16#0006E# => romdata <= X"0C515104";
    when 16#0006F# => romdata <= X"00000000";
    when 16#00070# => romdata <= X"72098105";
    when 16#00071# => romdata <= X"72050970";
    when 16#00072# => romdata <= X"81050906";
    when 16#00073# => romdata <= X"0A810653";
    when 16#00074# => romdata <= X"51040000";
    when 16#00075# => romdata <= X"00000000";
    when 16#00076# => romdata <= X"00000000";
    when 16#00077# => romdata <= X"00000000";
    when 16#00078# => romdata <= X"72098105";
    when 16#00079# => romdata <= X"72050970";
    when 16#0007A# => romdata <= X"81050906";
    when 16#0007B# => romdata <= X"0A098106";
    when 16#0007C# => romdata <= X"53510400";
    when 16#0007D# => romdata <= X"00000000";
    when 16#0007E# => romdata <= X"00000000";
    when 16#0007F# => romdata <= X"00000000";
    when 16#00080# => romdata <= X"71098105";
    when 16#00081# => romdata <= X"52040000";
    when 16#00082# => romdata <= X"00000000";
    when 16#00083# => romdata <= X"00000000";
    when 16#00084# => romdata <= X"00000000";
    when 16#00085# => romdata <= X"00000000";
    when 16#00086# => romdata <= X"00000000";
    when 16#00087# => romdata <= X"00000000";
    when 16#00088# => romdata <= X"72720981";
    when 16#00089# => romdata <= X"05055351";
    when 16#0008A# => romdata <= X"04000000";
    when 16#0008B# => romdata <= X"00000000";
    when 16#0008C# => romdata <= X"00000000";
    when 16#0008D# => romdata <= X"00000000";
    when 16#0008E# => romdata <= X"00000000";
    when 16#0008F# => romdata <= X"00000000";
    when 16#00090# => romdata <= X"72097206";
    when 16#00091# => romdata <= X"73730906";
    when 16#00092# => romdata <= X"07535104";
    when 16#00093# => romdata <= X"00000000";
    when 16#00094# => romdata <= X"00000000";
    when 16#00095# => romdata <= X"00000000";
    when 16#00096# => romdata <= X"00000000";
    when 16#00097# => romdata <= X"00000000";
    when 16#00098# => romdata <= X"71FC0608";
    when 16#00099# => romdata <= X"72830609";
    when 16#0009A# => romdata <= X"81058305";
    when 16#0009B# => romdata <= X"1010102A";
    when 16#0009C# => romdata <= X"81FF0652";
    when 16#0009D# => romdata <= X"04000000";
    when 16#0009E# => romdata <= X"00000000";
    when 16#0009F# => romdata <= X"00000000";
    when 16#000A0# => romdata <= X"71FC0608";
    when 16#000A1# => romdata <= X"0B0B80F0";
    when 16#000A2# => romdata <= X"98738306";
    when 16#000A3# => romdata <= X"10100508";
    when 16#000A4# => romdata <= X"060B0B0B";
    when 16#000A5# => romdata <= X"88AA0400";
    when 16#000A6# => romdata <= X"00000000";
    when 16#000A7# => romdata <= X"00000000";
    when 16#000A8# => romdata <= X"0B0B0B88";
    when 16#000A9# => romdata <= X"F9040000";
    when 16#000AA# => romdata <= X"00000000";
    when 16#000AB# => romdata <= X"00000000";
    when 16#000AC# => romdata <= X"00000000";
    when 16#000AD# => romdata <= X"00000000";
    when 16#000AE# => romdata <= X"00000000";
    when 16#000AF# => romdata <= X"00000000";
    when 16#000B0# => romdata <= X"0B0B0B88";
    when 16#000B1# => romdata <= X"E0040000";
    when 16#000B2# => romdata <= X"00000000";
    when 16#000B3# => romdata <= X"00000000";
    when 16#000B4# => romdata <= X"00000000";
    when 16#000B5# => romdata <= X"00000000";
    when 16#000B6# => romdata <= X"00000000";
    when 16#000B7# => romdata <= X"00000000";
    when 16#000B8# => romdata <= X"72097081";
    when 16#000B9# => romdata <= X"0509060A";
    when 16#000BA# => romdata <= X"8106FF05";
    when 16#000BB# => romdata <= X"70547106";
    when 16#000BC# => romdata <= X"73097274";
    when 16#000BD# => romdata <= X"05FF0506";
    when 16#000BE# => romdata <= X"07515151";
    when 16#000BF# => romdata <= X"04000000";
    when 16#000C0# => romdata <= X"72097081";
    when 16#000C1# => romdata <= X"0509060A";
    when 16#000C2# => romdata <= X"098106FF";
    when 16#000C3# => romdata <= X"05705471";
    when 16#000C4# => romdata <= X"06730972";
    when 16#000C5# => romdata <= X"7405FF05";
    when 16#000C6# => romdata <= X"06075151";
    when 16#000C7# => romdata <= X"51040000";
    when 16#000C8# => romdata <= X"05FF0504";
    when 16#000C9# => romdata <= X"00000000";
    when 16#000CA# => romdata <= X"00000000";
    when 16#000CB# => romdata <= X"00000000";
    when 16#000CC# => romdata <= X"00000000";
    when 16#000CD# => romdata <= X"00000000";
    when 16#000CE# => romdata <= X"00000000";
    when 16#000CF# => romdata <= X"00000000";
    when 16#000D0# => romdata <= X"810B0B0B";
    when 16#000D1# => romdata <= X"80F0A80C";
    when 16#000D2# => romdata <= X"51040000";
    when 16#000D3# => romdata <= X"00000000";
    when 16#000D4# => romdata <= X"00000000";
    when 16#000D5# => romdata <= X"00000000";
    when 16#000D6# => romdata <= X"00000000";
    when 16#000D7# => romdata <= X"00000000";
    when 16#000D8# => romdata <= X"71810552";
    when 16#000D9# => romdata <= X"04000000";
    when 16#000DA# => romdata <= X"00000000";
    when 16#000DB# => romdata <= X"00000000";
    when 16#000DC# => romdata <= X"00000000";
    when 16#000DD# => romdata <= X"00000000";
    when 16#000DE# => romdata <= X"00000000";
    when 16#000DF# => romdata <= X"00000000";
    when 16#000E0# => romdata <= X"00000000";
    when 16#000E1# => romdata <= X"00000000";
    when 16#000E2# => romdata <= X"00000000";
    when 16#000E3# => romdata <= X"00000000";
    when 16#000E4# => romdata <= X"00000000";
    when 16#000E5# => romdata <= X"00000000";
    when 16#000E6# => romdata <= X"00000000";
    when 16#000E7# => romdata <= X"00000000";
    when 16#000E8# => romdata <= X"02840572";
    when 16#000E9# => romdata <= X"10100552";
    when 16#000EA# => romdata <= X"04000000";
    when 16#000EB# => romdata <= X"00000000";
    when 16#000EC# => romdata <= X"00000000";
    when 16#000ED# => romdata <= X"00000000";
    when 16#000EE# => romdata <= X"00000000";
    when 16#000EF# => romdata <= X"00000000";
    when 16#000F0# => romdata <= X"00000000";
    when 16#000F1# => romdata <= X"00000000";
    when 16#000F2# => romdata <= X"00000000";
    when 16#000F3# => romdata <= X"00000000";
    when 16#000F4# => romdata <= X"00000000";
    when 16#000F5# => romdata <= X"00000000";
    when 16#000F6# => romdata <= X"00000000";
    when 16#000F7# => romdata <= X"00000000";
    when 16#000F8# => romdata <= X"717105FF";
    when 16#000F9# => romdata <= X"05715351";
    when 16#000FA# => romdata <= X"020D0400";
    when 16#000FB# => romdata <= X"00000000";
    when 16#000FC# => romdata <= X"00000000";
    when 16#000FD# => romdata <= X"00000000";
    when 16#000FE# => romdata <= X"00000000";
    when 16#000FF# => romdata <= X"00000000";
    when 16#00100# => romdata <= X"82C43F80";
    when 16#00101# => romdata <= X"DCC23F04";
    when 16#00102# => romdata <= X"10101010";
    when 16#00103# => romdata <= X"10101010";
    when 16#00104# => romdata <= X"10101010";
    when 16#00105# => romdata <= X"10101010";
    when 16#00106# => romdata <= X"10101010";
    when 16#00107# => romdata <= X"10101010";
    when 16#00108# => romdata <= X"10101010";
    when 16#00109# => romdata <= X"10101053";
    when 16#0010A# => romdata <= X"51047381";
    when 16#0010B# => romdata <= X"FF067383";
    when 16#0010C# => romdata <= X"06098105";
    when 16#0010D# => romdata <= X"83051010";
    when 16#0010E# => romdata <= X"102B0772";
    when 16#0010F# => romdata <= X"FC060C51";
    when 16#00110# => romdata <= X"51043C04";
    when 16#00111# => romdata <= X"72728072";
    when 16#00112# => romdata <= X"8106FF05";
    when 16#00113# => romdata <= X"09720605";
    when 16#00114# => romdata <= X"71105272";
    when 16#00115# => romdata <= X"0A100A53";
    when 16#00116# => romdata <= X"72ED3851";
    when 16#00117# => romdata <= X"51535104";
    when 16#00118# => romdata <= X"80088408";
    when 16#00119# => romdata <= X"88087575";
    when 16#0011A# => romdata <= X"80C1C12D";
    when 16#0011B# => romdata <= X"50508008";
    when 16#0011C# => romdata <= X"56880C84";
    when 16#0011D# => romdata <= X"0C800C51";
    when 16#0011E# => romdata <= X"04800884";
    when 16#0011F# => romdata <= X"08880875";
    when 16#00120# => romdata <= X"7580C08F";
    when 16#00121# => romdata <= X"2D505080";
    when 16#00122# => romdata <= X"0856880C";
    when 16#00123# => romdata <= X"840C800C";
    when 16#00124# => romdata <= X"51048008";
    when 16#00125# => romdata <= X"84088808";
    when 16#00126# => romdata <= X"80E3A12D";
    when 16#00127# => romdata <= X"880C840C";
    when 16#00128# => romdata <= X"800C0480";
    when 16#00129# => romdata <= X"F0A80880";
    when 16#0012A# => romdata <= X"2EA43880";
    when 16#0012B# => romdata <= X"F0AC0882";
    when 16#0012C# => romdata <= X"2EBD3883";
    when 16#0012D# => romdata <= X"80800B0B";
    when 16#0012E# => romdata <= X"0B8180B4";
    when 16#0012F# => romdata <= X"0C82A080";
    when 16#00130# => romdata <= X"0B8180B8";
    when 16#00131# => romdata <= X"0C829080";
    when 16#00132# => romdata <= X"0B8180BC";
    when 16#00133# => romdata <= X"0C04F880";
    when 16#00134# => romdata <= X"8080A40B";
    when 16#00135# => romdata <= X"0B0B8180";
    when 16#00136# => romdata <= X"B40CF880";
    when 16#00137# => romdata <= X"8082800B";
    when 16#00138# => romdata <= X"8180B80C";
    when 16#00139# => romdata <= X"F8808084";
    when 16#0013A# => romdata <= X"800B8180";
    when 16#0013B# => romdata <= X"BC0C0480";
    when 16#0013C# => romdata <= X"C0A8808C";
    when 16#0013D# => romdata <= X"0B0B0B81";
    when 16#0013E# => romdata <= X"80B40C80";
    when 16#0013F# => romdata <= X"C0A88094";
    when 16#00140# => romdata <= X"0B8180B8";
    when 16#00141# => romdata <= X"0C0B0B80";
    when 16#00142# => romdata <= X"E4F40B81";
    when 16#00143# => romdata <= X"80BC0C04";
    when 16#00144# => romdata <= X"FF3D0D81";
    when 16#00145# => romdata <= X"80C03351";
    when 16#00146# => romdata <= X"70A73880";
    when 16#00147# => romdata <= X"F0B40870";
    when 16#00148# => romdata <= X"08525270";
    when 16#00149# => romdata <= X"802E9438";
    when 16#0014A# => romdata <= X"841280F0";
    when 16#0014B# => romdata <= X"B40C702D";
    when 16#0014C# => romdata <= X"80F0B408";
    when 16#0014D# => romdata <= X"70085252";
    when 16#0014E# => romdata <= X"70EE3881";
    when 16#0014F# => romdata <= X"0B8180C0";
    when 16#00150# => romdata <= X"34833D0D";
    when 16#00151# => romdata <= X"0404803D";
    when 16#00152# => romdata <= X"0D0B0B81";
    when 16#00153# => romdata <= X"80B00880";
    when 16#00154# => romdata <= X"2E8E380B";
    when 16#00155# => romdata <= X"0B0B0B80";
    when 16#00156# => romdata <= X"0B802E09";
    when 16#00157# => romdata <= X"81068538";
    when 16#00158# => romdata <= X"823D0D04";
    when 16#00159# => romdata <= X"0B0B8180";
    when 16#0015A# => romdata <= X"B0510B0B";
    when 16#0015B# => romdata <= X"0BF5913F";
    when 16#0015C# => romdata <= X"823D0D04";
    when 16#0015D# => romdata <= X"04FF3D0D";
    when 16#0015E# => romdata <= X"028F0533";
    when 16#0015F# => romdata <= X"705252B2";
    when 16#00160# => romdata <= X"CD3F7151";
    when 16#00161# => romdata <= X"B3BC3F71";
    when 16#00162# => romdata <= X"800C833D";
    when 16#00163# => romdata <= X"0D04FA3D";
    when 16#00164# => romdata <= X"0D02A305";
    when 16#00165# => romdata <= X"3356758D";
    when 16#00166# => romdata <= X"2E80F438";
    when 16#00167# => romdata <= X"75883270";
    when 16#00168# => romdata <= X"307780FF";
    when 16#00169# => romdata <= X"32703072";
    when 16#0016A# => romdata <= X"80257180";
    when 16#0016B# => romdata <= X"25075451";
    when 16#0016C# => romdata <= X"56585574";
    when 16#0016D# => romdata <= X"95389F76";
    when 16#0016E# => romdata <= X"278C3881";
    when 16#0016F# => romdata <= X"8ABC3355";
    when 16#00170# => romdata <= X"80CE7527";
    when 16#00171# => romdata <= X"AE38883D";
    when 16#00172# => romdata <= X"0D04818A";
    when 16#00173# => romdata <= X"BC335675";
    when 16#00174# => romdata <= X"802EF338";
    when 16#00175# => romdata <= X"8851ADB4";
    when 16#00176# => romdata <= X"3FA051AD";
    when 16#00177# => romdata <= X"AF3F8851";
    when 16#00178# => romdata <= X"ADAA3F81";
    when 16#00179# => romdata <= X"8ABC33FF";
    when 16#0017A# => romdata <= X"05577681";
    when 16#0017B# => romdata <= X"8ABC3488";
    when 16#0017C# => romdata <= X"3D0D0475";
    when 16#0017D# => romdata <= X"51AD953F";
    when 16#0017E# => romdata <= X"818ABC33";
    when 16#0017F# => romdata <= X"81115557";
    when 16#00180# => romdata <= X"73818ABC";
    when 16#00181# => romdata <= X"34758189";
    when 16#00182# => romdata <= X"E8183488";
    when 16#00183# => romdata <= X"3D0D048A";
    when 16#00184# => romdata <= X"51ACF93F";
    when 16#00185# => romdata <= X"818ABC33";
    when 16#00186# => romdata <= X"81115654";
    when 16#00187# => romdata <= X"74818ABC";
    when 16#00188# => romdata <= X"34800B81";
    when 16#00189# => romdata <= X"89E81534";
    when 16#0018A# => romdata <= X"8056800B";
    when 16#0018B# => romdata <= X"8189E817";
    when 16#0018C# => romdata <= X"33565474";
    when 16#0018D# => romdata <= X"A02E8338";
    when 16#0018E# => romdata <= X"81547480";
    when 16#0018F# => romdata <= X"2E903873";
    when 16#00190# => romdata <= X"802E8B38";
    when 16#00191# => romdata <= X"81167081";
    when 16#00192# => romdata <= X"FF065757";
    when 16#00193# => romdata <= X"DD397580";
    when 16#00194# => romdata <= X"2EBF3880";
    when 16#00195# => romdata <= X"0B818AB8";
    when 16#00196# => romdata <= X"33555574";
    when 16#00197# => romdata <= X"7427AB38";
    when 16#00198# => romdata <= X"73577410";
    when 16#00199# => romdata <= X"10107510";
    when 16#0019A# => romdata <= X"05765481";
    when 16#0019B# => romdata <= X"89E85381";
    when 16#0019C# => romdata <= X"80C80551";
    when 16#0019D# => romdata <= X"BDFC3F80";
    when 16#0019E# => romdata <= X"08802EA6";
    when 16#0019F# => romdata <= X"38811570";
    when 16#001A0# => romdata <= X"81FF0656";
    when 16#001A1# => romdata <= X"54767526";
    when 16#001A2# => romdata <= X"D93880E5";
    when 16#001A3# => romdata <= X"8451AC96";
    when 16#001A4# => romdata <= X"3F80E580";
    when 16#001A5# => romdata <= X"51AC8F3F";
    when 16#001A6# => romdata <= X"800B818A";
    when 16#001A7# => romdata <= X"BC34883D";
    when 16#001A8# => romdata <= X"0D047410";
    when 16#001A9# => romdata <= X"108189A8";
    when 16#001AA# => romdata <= X"05700881";
    when 16#001AB# => romdata <= X"8AC00C56";
    when 16#001AC# => romdata <= X"800B818A";
    when 16#001AD# => romdata <= X"BC34E739";
    when 16#001AE# => romdata <= X"800B818A";
    when 16#001AF# => romdata <= X"C43404FC";
    when 16#001B0# => romdata <= X"3D0D8A51";
    when 16#001B1# => romdata <= X"ABC63F80";
    when 16#001B2# => romdata <= X"E59851AB";
    when 16#001B3# => romdata <= X"D93F800B";
    when 16#001B4# => romdata <= X"818AB833";
    when 16#001B5# => romdata <= X"53537272";
    when 16#001B6# => romdata <= X"2780F538";
    when 16#001B7# => romdata <= X"72101010";
    when 16#001B8# => romdata <= X"73100581";
    when 16#001B9# => romdata <= X"80C80570";
    when 16#001BA# => romdata <= X"5254ABBA";
    when 16#001BB# => romdata <= X"3F72842B";
    when 16#001BC# => romdata <= X"70743182";
    when 16#001BD# => romdata <= X"2B8181E8";
    when 16#001BE# => romdata <= X"11335153";
    when 16#001BF# => romdata <= X"5571802E";
    when 16#001C0# => romdata <= X"B7387351";
    when 16#001C1# => romdata <= X"BC8D3F80";
    when 16#001C2# => romdata <= X"0881FF06";
    when 16#001C3# => romdata <= X"52718926";
    when 16#001C4# => romdata <= X"9338A051";
    when 16#001C5# => romdata <= X"AAF63F81";
    when 16#001C6# => romdata <= X"127081FF";
    when 16#001C7# => romdata <= X"06535489";
    when 16#001C8# => romdata <= X"7227EF38";
    when 16#001C9# => romdata <= X"80E5B051";
    when 16#001CA# => romdata <= X"AAFC3F74";
    when 16#001CB# => romdata <= X"7331822B";
    when 16#001CC# => romdata <= X"8181E805";
    when 16#001CD# => romdata <= X"51AAEF3F";
    when 16#001CE# => romdata <= X"8A51AAD0";
    when 16#001CF# => romdata <= X"3F811370";
    when 16#001D0# => romdata <= X"81FF0681";
    when 16#001D1# => romdata <= X"8AB83354";
    when 16#001D2# => romdata <= X"54557173";
    when 16#001D3# => romdata <= X"26FF8D38";
    when 16#001D4# => romdata <= X"8A51AAB8";
    when 16#001D5# => romdata <= X"3F863D0D";
    when 16#001D6# => romdata <= X"04FC3D0D";
    when 16#001D7# => romdata <= X"8A51AAAC";
    when 16#001D8# => romdata <= X"3F800B81";
    when 16#001D9# => romdata <= X"8ABC3480";
    when 16#001DA# => romdata <= X"0B818AB8";
    when 16#001DB# => romdata <= X"34800B81";
    when 16#001DC# => romdata <= X"8AC00C80";
    when 16#001DD# => romdata <= X"E5B45281";
    when 16#001DE# => romdata <= X"80C851BA";
    when 16#001DF# => romdata <= X"A93F80E5";
    when 16#001E0# => romdata <= X"B852818A";
    when 16#001E1# => romdata <= X"B8337090";
    when 16#001E2# => romdata <= X"29713170";
    when 16#001E3# => romdata <= X"10108181";
    when 16#001E4# => romdata <= X"E8055356";
    when 16#001E5# => romdata <= X"54BA8F3F";
    when 16#001E6# => romdata <= X"818AB833";
    when 16#001E7# => romdata <= X"70101081";
    when 16#001E8# => romdata <= X"89A805AB";
    when 16#001E9# => romdata <= X"94710C54";
    when 16#001EA# => romdata <= X"81115155";
    when 16#001EB# => romdata <= X"74818AB8";
    when 16#001EC# => romdata <= X"3480E5CC";
    when 16#001ED# => romdata <= X"527481FF";
    when 16#001EE# => romdata <= X"06708A29";
    when 16#001EF# => romdata <= X"8180C805";
    when 16#001F0# => romdata <= X"5253B9E2";
    when 16#001F1# => romdata <= X"3F80E5D4";
    when 16#001F2# => romdata <= X"52818AB8";
    when 16#001F3# => romdata <= X"33709029";
    when 16#001F4# => romdata <= X"71317010";
    when 16#001F5# => romdata <= X"108181E8";
    when 16#001F6# => romdata <= X"05535555";
    when 16#001F7# => romdata <= X"B9C83F81";
    when 16#001F8# => romdata <= X"8AB83370";
    when 16#001F9# => romdata <= X"10108189";
    when 16#001FA# => romdata <= X"A8059CAE";
    when 16#001FB# => romdata <= X"710C5481";
    when 16#001FC# => romdata <= X"11515473";
    when 16#001FD# => romdata <= X"818AB834";
    when 16#001FE# => romdata <= X"80E5E852";
    when 16#001FF# => romdata <= X"7381FF06";
    when 16#00200# => romdata <= X"708A2981";
    when 16#00201# => romdata <= X"80C80552";
    when 16#00202# => romdata <= X"53B99B3F";
    when 16#00203# => romdata <= X"80E5F052";
    when 16#00204# => romdata <= X"818AB833";
    when 16#00205# => romdata <= X"70902971";
    when 16#00206# => romdata <= X"31701010";
    when 16#00207# => romdata <= X"8181E805";
    when 16#00208# => romdata <= X"535654B9";
    when 16#00209# => romdata <= X"813F818A";
    when 16#0020A# => romdata <= X"B8337010";
    when 16#0020B# => romdata <= X"108189A8";
    when 16#0020C# => romdata <= X"059E8971";
    when 16#0020D# => romdata <= X"0C548111";
    when 16#0020E# => romdata <= X"51557481";
    when 16#0020F# => romdata <= X"8AB83480";
    when 16#00210# => romdata <= X"E6885274";
    when 16#00211# => romdata <= X"81FF0670";
    when 16#00212# => romdata <= X"8A298180";
    when 16#00213# => romdata <= X"C8055253";
    when 16#00214# => romdata <= X"B8D43F80";
    when 16#00215# => romdata <= X"E6905281";
    when 16#00216# => romdata <= X"8AB83370";
    when 16#00217# => romdata <= X"90297131";
    when 16#00218# => romdata <= X"70101081";
    when 16#00219# => romdata <= X"81E80553";
    when 16#0021A# => romdata <= X"5555B8BA";
    when 16#0021B# => romdata <= X"3F818AB8";
    when 16#0021C# => romdata <= X"33701010";
    when 16#0021D# => romdata <= X"8189A805";
    when 16#0021E# => romdata <= X"A0BF710C";
    when 16#0021F# => romdata <= X"54811151";
    when 16#00220# => romdata <= X"5473818A";
    when 16#00221# => romdata <= X"B83480E6";
    when 16#00222# => romdata <= X"A8527381";
    when 16#00223# => romdata <= X"FF06708A";
    when 16#00224# => romdata <= X"298180C8";
    when 16#00225# => romdata <= X"055253B8";
    when 16#00226# => romdata <= X"8D3F80E6";
    when 16#00227# => romdata <= X"B052818A";
    when 16#00228# => romdata <= X"B8337090";
    when 16#00229# => romdata <= X"29713170";
    when 16#0022A# => romdata <= X"10108181";
    when 16#0022B# => romdata <= X"E8055356";
    when 16#0022C# => romdata <= X"54B7F33F";
    when 16#0022D# => romdata <= X"818AB833";
    when 16#0022E# => romdata <= X"70101081";
    when 16#0022F# => romdata <= X"89A805A6";
    when 16#00230# => romdata <= X"E8710C54";
    when 16#00231# => romdata <= X"81115155";
    when 16#00232# => romdata <= X"74818AB8";
    when 16#00233# => romdata <= X"3480E6C8";
    when 16#00234# => romdata <= X"527481FF";
    when 16#00235# => romdata <= X"06708A29";
    when 16#00236# => romdata <= X"8180C805";
    when 16#00237# => romdata <= X"5253B7C6";
    when 16#00238# => romdata <= X"3F80E6D0";
    when 16#00239# => romdata <= X"52818AB8";
    when 16#0023A# => romdata <= X"33709029";
    when 16#0023B# => romdata <= X"71317010";
    when 16#0023C# => romdata <= X"108181E8";
    when 16#0023D# => romdata <= X"05535555";
    when 16#0023E# => romdata <= X"B7AC3F81";
    when 16#0023F# => romdata <= X"8AB83370";
    when 16#00240# => romdata <= X"10108189";
    when 16#00241# => romdata <= X"A805A28F";
    when 16#00242# => romdata <= X"710C5481";
    when 16#00243# => romdata <= X"11515473";
    when 16#00244# => romdata <= X"818AB834";
    when 16#00245# => romdata <= X"80E6F852";
    when 16#00246# => romdata <= X"7381FF06";
    when 16#00247# => romdata <= X"708A2981";
    when 16#00248# => romdata <= X"80C80552";
    when 16#00249# => romdata <= X"53B6FF3F";
    when 16#0024A# => romdata <= X"80E6FC52";
    when 16#0024B# => romdata <= X"818AB833";
    when 16#0024C# => romdata <= X"70902971";
    when 16#0024D# => romdata <= X"31701010";
    when 16#0024E# => romdata <= X"8181E805";
    when 16#0024F# => romdata <= X"535654B6";
    when 16#00250# => romdata <= X"E53F818A";
    when 16#00251# => romdata <= X"B8337010";
    when 16#00252# => romdata <= X"108189A8";
    when 16#00253# => romdata <= X"05969071";
    when 16#00254# => romdata <= X"0C548111";
    when 16#00255# => romdata <= X"51557481";
    when 16#00256# => romdata <= X"8AB83480";
    when 16#00257# => romdata <= X"E7885274";
    when 16#00258# => romdata <= X"81FF0670";
    when 16#00259# => romdata <= X"8A298180";
    when 16#0025A# => romdata <= X"C8055253";
    when 16#0025B# => romdata <= X"B6B83F80";
    when 16#0025C# => romdata <= X"E7905281";
    when 16#0025D# => romdata <= X"8AB83370";
    when 16#0025E# => romdata <= X"90297131";
    when 16#0025F# => romdata <= X"70101081";
    when 16#00260# => romdata <= X"81E80553";
    when 16#00261# => romdata <= X"5555B69E";
    when 16#00262# => romdata <= X"3F818AB8";
    when 16#00263# => romdata <= X"33701010";
    when 16#00264# => romdata <= X"8189A805";
    when 16#00265# => romdata <= X"99D2710C";
    when 16#00266# => romdata <= X"54811151";
    when 16#00267# => romdata <= X"5473818A";
    when 16#00268# => romdata <= X"B83480E8";
    when 16#00269# => romdata <= X"EC527381";
    when 16#0026A# => romdata <= X"FF06708A";
    when 16#0026B# => romdata <= X"298180C8";
    when 16#0026C# => romdata <= X"055253B5";
    when 16#0026D# => romdata <= X"F13F80E7";
    when 16#0026E# => romdata <= X"9C52818A";
    when 16#0026F# => romdata <= X"B8337090";
    when 16#00270# => romdata <= X"29713170";
    when 16#00271# => romdata <= X"10108181";
    when 16#00272# => romdata <= X"E8055356";
    when 16#00273# => romdata <= X"54B5D73F";
    when 16#00274# => romdata <= X"818AB833";
    when 16#00275# => romdata <= X"70101081";
    when 16#00276# => romdata <= X"89A80596";
    when 16#00277# => romdata <= X"90710C54";
    when 16#00278# => romdata <= X"81115155";
    when 16#00279# => romdata <= X"74818AB8";
    when 16#0027A# => romdata <= X"3480E7AC";
    when 16#0027B# => romdata <= X"527481FF";
    when 16#0027C# => romdata <= X"06708A29";
    when 16#0027D# => romdata <= X"8180C805";
    when 16#0027E# => romdata <= X"5253B5AA";
    when 16#0027F# => romdata <= X"3F80E7B4";
    when 16#00280# => romdata <= X"52818AB8";
    when 16#00281# => romdata <= X"33709029";
    when 16#00282# => romdata <= X"71317010";
    when 16#00283# => romdata <= X"108181E8";
    when 16#00284# => romdata <= X"05535555";
    when 16#00285# => romdata <= X"B5903F81";
    when 16#00286# => romdata <= X"8AB83370";
    when 16#00287# => romdata <= X"10108189";
    when 16#00288# => romdata <= X"A8059CA2";
    when 16#00289# => romdata <= X"710C5481";
    when 16#0028A# => romdata <= X"11515473";
    when 16#0028B# => romdata <= X"818AB834";
    when 16#0028C# => romdata <= X"80E7C452";
    when 16#0028D# => romdata <= X"7381FF06";
    when 16#0028E# => romdata <= X"708A2981";
    when 16#0028F# => romdata <= X"80C80552";
    when 16#00290# => romdata <= X"53B4E33F";
    when 16#00291# => romdata <= X"80E7EC52";
    when 16#00292# => romdata <= X"818AB833";
    when 16#00293# => romdata <= X"70902971";
    when 16#00294# => romdata <= X"31701010";
    when 16#00295# => romdata <= X"8181E805";
    when 16#00296# => romdata <= X"535654B4";
    when 16#00297# => romdata <= X"C93F818A";
    when 16#00298# => romdata <= X"B8337010";
    when 16#00299# => romdata <= X"108189A8";
    when 16#0029A# => romdata <= X"058DB871";
    when 16#0029B# => romdata <= X"0C548111";
    when 16#0029C# => romdata <= X"51557481";
    when 16#0029D# => romdata <= X"8AB83480";
    when 16#0029E# => romdata <= X"E4F85274";
    when 16#0029F# => romdata <= X"81FF0670";
    when 16#002A0# => romdata <= X"8A298180";
    when 16#002A1# => romdata <= X"C8055253";
    when 16#002A2# => romdata <= X"B49C3F80";
    when 16#002A3# => romdata <= X"E7EC5281";
    when 16#002A4# => romdata <= X"8AB83370";
    when 16#002A5# => romdata <= X"90297131";
    when 16#002A6# => romdata <= X"70101081";
    when 16#002A7# => romdata <= X"81E80553";
    when 16#002A8# => romdata <= X"5555B482";
    when 16#002A9# => romdata <= X"3F818AB8";
    when 16#002AA# => romdata <= X"33701010";
    when 16#002AB# => romdata <= X"8189A805";
    when 16#002AC# => romdata <= X"8DBF710C";
    when 16#002AD# => romdata <= X"54810553";
    when 16#002AE# => romdata <= X"72818AB8";
    when 16#002AF# => romdata <= X"34F8803F";
    when 16#002B0# => romdata <= X"80E58051";
    when 16#002B1# => romdata <= X"A3E03F81";
    when 16#002B2# => romdata <= X"0B818AC4";
    when 16#002B3# => romdata <= X"34A7CA3F";
    when 16#002B4# => romdata <= X"8008AE38";
    when 16#002B5# => romdata <= X"818AC008";
    when 16#002B6# => romdata <= X"53728D38";
    when 16#002B7# => romdata <= X"818AC433";
    when 16#002B8# => romdata <= X"5372EA38";
    when 16#002B9# => romdata <= X"863D0D04";
    when 16#002BA# => romdata <= X"722D800B";
    when 16#002BB# => romdata <= X"818AC00C";
    when 16#002BC# => romdata <= X"80E58051";
    when 16#002BD# => romdata <= X"A3B03F81";
    when 16#002BE# => romdata <= X"8AC43353";
    when 16#002BF# => romdata <= X"72CF38E4";
    when 16#002C0# => romdata <= X"39A7A93F";
    when 16#002C1# => romdata <= X"800881FF";
    when 16#002C2# => romdata <= X"0651F582";
    when 16#002C3# => romdata <= X"3FFFBE39";
    when 16#002C4# => romdata <= X"F63D0D80";
    when 16#002C5# => romdata <= X"0B8189E8";
    when 16#002C6# => romdata <= X"338189E8";
    when 16#002C7# => romdata <= X"59555673";
    when 16#002C8# => romdata <= X"A02E0981";
    when 16#002C9# => romdata <= X"06963881";
    when 16#002CA# => romdata <= X"167081FF";
    when 16#002CB# => romdata <= X"068189E8";
    when 16#002CC# => romdata <= X"11703353";
    when 16#002CD# => romdata <= X"59575473";
    when 16#002CE# => romdata <= X"A02EEC38";
    when 16#002CF# => romdata <= X"80588077";
    when 16#002D0# => romdata <= X"33565474";
    when 16#002D1# => romdata <= X"742E8338";
    when 16#002D2# => romdata <= X"815474A0";
    when 16#002D3# => romdata <= X"2E81CE38";
    when 16#002D4# => romdata <= X"7381FB38";
    when 16#002D5# => romdata <= X"74A02E81";
    when 16#002D6# => romdata <= X"C4388118";
    when 16#002D7# => romdata <= X"7081FF06";
    when 16#002D8# => romdata <= X"59548178";
    when 16#002D9# => romdata <= X"26D83890";
    when 16#002DA# => romdata <= X"538C3DFC";
    when 16#002DB# => romdata <= X"05527651";
    when 16#002DC# => romdata <= X"B8CF3F80";
    when 16#002DD# => romdata <= X"0859800B";
    when 16#002DE# => romdata <= X"8189E833";
    when 16#002DF# => romdata <= X"8189E859";
    when 16#002E0# => romdata <= X"555673A0";
    when 16#002E1# => romdata <= X"2E098106";
    when 16#002E2# => romdata <= X"96388116";
    when 16#002E3# => romdata <= X"7081FF06";
    when 16#002E4# => romdata <= X"8189E811";
    when 16#002E5# => romdata <= X"70335759";
    when 16#002E6# => romdata <= X"575873A0";
    when 16#002E7# => romdata <= X"2EEC3880";
    when 16#002E8# => romdata <= X"58807733";
    when 16#002E9# => romdata <= X"56547474";
    when 16#002EA# => romdata <= X"2E833881";
    when 16#002EB# => romdata <= X"5474A02E";
    when 16#002EC# => romdata <= X"81AC3873";
    when 16#002ED# => romdata <= X"828C3874";
    when 16#002EE# => romdata <= X"A02E81A2";
    when 16#002EF# => romdata <= X"38811870";
    when 16#002F0# => romdata <= X"81FF0659";
    when 16#002F1# => romdata <= X"55827826";
    when 16#002F2# => romdata <= X"D8389053";
    when 16#002F3# => romdata <= X"8C3DF805";
    when 16#002F4# => romdata <= X"527651B7";
    when 16#002F5# => romdata <= X"EC3F8008";
    when 16#002F6# => romdata <= X"57800883";
    when 16#002F7# => romdata <= X"38905778";
    when 16#002F8# => romdata <= X"FC065580";
    when 16#002F9# => romdata <= X"56757727";
    when 16#002FA# => romdata <= X"AB387583";
    when 16#002FB# => romdata <= X"06597880";
    when 16#002FC# => romdata <= X"2E819C38";
    when 16#002FD# => romdata <= X"80E7CC51";
    when 16#002FE# => romdata <= X"A1AC3F74";
    when 16#002FF# => romdata <= X"70840556";
    when 16#00300# => romdata <= X"0852A051";
    when 16#00301# => romdata <= X"A1C33FA0";
    when 16#00302# => romdata <= X"51A1813F";
    when 16#00303# => romdata <= X"81165676";
    when 16#00304# => romdata <= X"7626D738";
    when 16#00305# => romdata <= X"8A51A0F4";
    when 16#00306# => romdata <= X"3F8C3D0D";
    when 16#00307# => romdata <= X"04811670";
    when 16#00308# => romdata <= X"81FF0681";
    when 16#00309# => romdata <= X"89E81170";
    when 16#0030A# => romdata <= X"335C5257";
    when 16#0030B# => romdata <= X"5778A02E";
    when 16#0030C# => romdata <= X"098106FE";
    when 16#0030D# => romdata <= X"A5388116";
    when 16#0030E# => romdata <= X"7081FF06";
    when 16#0030F# => romdata <= X"8189E811";
    when 16#00310# => romdata <= X"70335C52";
    when 16#00311# => romdata <= X"575778A0";
    when 16#00312# => romdata <= X"2ED338FE";
    when 16#00313# => romdata <= X"8D398116";
    when 16#00314# => romdata <= X"7081FF06";
    when 16#00315# => romdata <= X"8189E811";
    when 16#00316# => romdata <= X"595755FD";
    when 16#00317# => romdata <= X"E1398116";
    when 16#00318# => romdata <= X"7081FF06";
    when 16#00319# => romdata <= X"8189E811";
    when 16#0031A# => romdata <= X"70335752";
    when 16#0031B# => romdata <= X"575773A0";
    when 16#0031C# => romdata <= X"2E098106";
    when 16#0031D# => romdata <= X"FEC73881";
    when 16#0031E# => romdata <= X"167081FF";
    when 16#0031F# => romdata <= X"068189E8";
    when 16#00320# => romdata <= X"11703357";
    when 16#00321# => romdata <= X"52575773";
    when 16#00322# => romdata <= X"A02ED338";
    when 16#00323# => romdata <= X"FEAF3980";
    when 16#00324# => romdata <= X"E7D051A0";
    when 16#00325# => romdata <= X"913F7452";
    when 16#00326# => romdata <= X"A051A0AD";
    when 16#00327# => romdata <= X"3F80E7D4";
    when 16#00328# => romdata <= X"51A0833F";
    when 16#00329# => romdata <= X"80E7CC51";
    when 16#0032A# => romdata <= X"9FFC3F74";
    when 16#0032B# => romdata <= X"70840556";
    when 16#0032C# => romdata <= X"0852A051";
    when 16#0032D# => romdata <= X"A0933FA0";
    when 16#0032E# => romdata <= X"519FD13F";
    when 16#0032F# => romdata <= X"811656FE";
    when 16#00330# => romdata <= X"CE398116";
    when 16#00331# => romdata <= X"7081FF06";
    when 16#00332# => romdata <= X"8189E811";
    when 16#00333# => romdata <= X"595755FD";
    when 16#00334# => romdata <= X"D039F63D";
    when 16#00335# => romdata <= X"0D800B81";
    when 16#00336# => romdata <= X"89E83381";
    when 16#00337# => romdata <= X"89E85955";
    when 16#00338# => romdata <= X"5673A02E";
    when 16#00339# => romdata <= X"09810696";
    when 16#0033A# => romdata <= X"38811670";
    when 16#0033B# => romdata <= X"81FF0681";
    when 16#0033C# => romdata <= X"89E81170";
    when 16#0033D# => romdata <= X"33535957";
    when 16#0033E# => romdata <= X"5473A02E";
    when 16#0033F# => romdata <= X"EC388058";
    when 16#00340# => romdata <= X"80773356";
    when 16#00341# => romdata <= X"5474742E";
    when 16#00342# => romdata <= X"83388154";
    when 16#00343# => romdata <= X"74A02E81";
    when 16#00344# => romdata <= X"8F387381";
    when 16#00345# => romdata <= X"BC3874A0";
    when 16#00346# => romdata <= X"2E818538";
    when 16#00347# => romdata <= X"81187081";
    when 16#00348# => romdata <= X"FF065954";
    when 16#00349# => romdata <= X"817826D8";
    when 16#0034A# => romdata <= X"3890538C";
    when 16#0034B# => romdata <= X"3DFC0552";
    when 16#0034C# => romdata <= X"7651B58D";
    when 16#0034D# => romdata <= X"3F800859";
    when 16#0034E# => romdata <= X"800B8189";
    when 16#0034F# => romdata <= X"E8338189";
    when 16#00350# => romdata <= X"E8595556";
    when 16#00351# => romdata <= X"73A02E09";
    when 16#00352# => romdata <= X"81069638";
    when 16#00353# => romdata <= X"81167081";
    when 16#00354# => romdata <= X"FF068189";
    when 16#00355# => romdata <= X"E8117033";
    when 16#00356# => romdata <= X"57595758";
    when 16#00357# => romdata <= X"73A02EEC";
    when 16#00358# => romdata <= X"38805880";
    when 16#00359# => romdata <= X"77335654";
    when 16#0035A# => romdata <= X"74742E83";
    when 16#0035B# => romdata <= X"38815474";
    when 16#0035C# => romdata <= X"A02E80ED";
    when 16#0035D# => romdata <= X"3873819A";
    when 16#0035E# => romdata <= X"3874A02E";
    when 16#0035F# => romdata <= X"80E33881";
    when 16#00360# => romdata <= X"187081FF";
    when 16#00361# => romdata <= X"06595582";
    when 16#00362# => romdata <= X"7826D838";
    when 16#00363# => romdata <= X"90538C3D";
    when 16#00364# => romdata <= X"F8055276";
    when 16#00365# => romdata <= X"51B4AA3F";
    when 16#00366# => romdata <= X"8008790C";
    when 16#00367# => romdata <= X"8C3D0D04";
    when 16#00368# => romdata <= X"81167081";
    when 16#00369# => romdata <= X"FF068189";
    when 16#0036A# => romdata <= X"E8117033";
    when 16#0036B# => romdata <= X"5C525757";
    when 16#0036C# => romdata <= X"78A02E09";
    when 16#0036D# => romdata <= X"8106FEE4";
    when 16#0036E# => romdata <= X"38811670";
    when 16#0036F# => romdata <= X"81FF0681";
    when 16#00370# => romdata <= X"89E81170";
    when 16#00371# => romdata <= X"335C5257";
    when 16#00372# => romdata <= X"5778A02E";
    when 16#00373# => romdata <= X"D338FECC";
    when 16#00374# => romdata <= X"39811670";
    when 16#00375# => romdata <= X"81FF0681";
    when 16#00376# => romdata <= X"89E81159";
    when 16#00377# => romdata <= X"5755FEA0";
    when 16#00378# => romdata <= X"39811670";
    when 16#00379# => romdata <= X"81FF0681";
    when 16#0037A# => romdata <= X"89E81170";
    when 16#0037B# => romdata <= X"33575257";
    when 16#0037C# => romdata <= X"5773A02E";
    when 16#0037D# => romdata <= X"098106FF";
    when 16#0037E# => romdata <= X"86388116";
    when 16#0037F# => romdata <= X"7081FF06";
    when 16#00380# => romdata <= X"8189E811";
    when 16#00381# => romdata <= X"70335752";
    when 16#00382# => romdata <= X"575773A0";
    when 16#00383# => romdata <= X"2ED338FE";
    when 16#00384# => romdata <= X"EE398116";
    when 16#00385# => romdata <= X"7081FF06";
    when 16#00386# => romdata <= X"8189E811";
    when 16#00387# => romdata <= X"595755FE";
    when 16#00388# => romdata <= X"C239803D";
    when 16#00389# => romdata <= X"0D8C519C";
    when 16#0038A# => romdata <= X"E33F823D";
    when 16#0038B# => romdata <= X"0D04FB3D";
    when 16#0038C# => romdata <= X"0D80E7D8";
    when 16#0038D# => romdata <= X"519CEF3F";
    when 16#0038E# => romdata <= X"805680F0";
    when 16#0038F# => romdata <= X"BC087610";
    when 16#00390# => romdata <= X"81FE0688";
    when 16#00391# => romdata <= X"120C5481";
    when 16#00392# => romdata <= X"D00B8C15";
    when 16#00393# => romdata <= X"0C8C1408";
    when 16#00394# => romdata <= X"70812A81";
    when 16#00395# => romdata <= X"06515574";
    when 16#00396# => romdata <= X"F4388C14";
    when 16#00397# => romdata <= X"0870872A";
    when 16#00398# => romdata <= X"81065553";
    when 16#00399# => romdata <= X"73802E80";
    when 16#0039A# => romdata <= X"DE388116";
    when 16#0039B# => romdata <= X"7081FF06";
    when 16#0039C# => romdata <= X"70982B56";
    when 16#0039D# => romdata <= X"57537380";
    when 16#0039E# => romdata <= X"25C03880";
    when 16#0039F# => romdata <= X"E7E4519C";
    when 16#003A0# => romdata <= X"A53F80F0";
    when 16#003A1# => romdata <= X"B8087510";
    when 16#003A2# => romdata <= X"81FE0688";
    when 16#003A3# => romdata <= X"120C5481";
    when 16#003A4# => romdata <= X"D00B8C15";
    when 16#003A5# => romdata <= X"0C8C1408";
    when 16#003A6# => romdata <= X"70812A81";
    when 16#003A7# => romdata <= X"06515372";
    when 16#003A8# => romdata <= X"F4388C14";
    when 16#003A9# => romdata <= X"0870872A";
    when 16#003AA# => romdata <= X"81065553";
    when 16#003AB# => romdata <= X"73802E80";
    when 16#003AC# => romdata <= X"C0388115";
    when 16#003AD# => romdata <= X"7081FF06";
    when 16#003AE# => romdata <= X"70982B56";
    when 16#003AF# => romdata <= X"56567380";
    when 16#003B0# => romdata <= X"25C03887";
    when 16#003B1# => romdata <= X"3D0D0480";
    when 16#003B2# => romdata <= X"E7F0519B";
    when 16#003B3# => romdata <= X"D93F7552";
    when 16#003B4# => romdata <= X"88519BF5";
    when 16#003B5# => romdata <= X"3F80E880";
    when 16#003B6# => romdata <= X"519BCB3F";
    when 16#003B7# => romdata <= X"81167081";
    when 16#003B8# => romdata <= X"FF067098";
    when 16#003B9# => romdata <= X"2B565753";
    when 16#003BA# => romdata <= X"738025FE";
    when 16#003BB# => romdata <= X"CD38FF8B";
    when 16#003BC# => romdata <= X"3980E7F0";
    when 16#003BD# => romdata <= X"519BAF3F";
    when 16#003BE# => romdata <= X"74528851";
    when 16#003BF# => romdata <= X"9BCB3F80";
    when 16#003C0# => romdata <= X"E880519B";
    when 16#003C1# => romdata <= X"A13FFFAA";
    when 16#003C2# => romdata <= X"39F83D0D";
    when 16#003C3# => romdata <= X"80E89051";
    when 16#003C4# => romdata <= X"9B943F82";
    when 16#003C5# => romdata <= X"80519CD3";
    when 16#003C6# => romdata <= X"3F80E8A4";
    when 16#003C7# => romdata <= X"519B873F";
    when 16#003C8# => romdata <= X"80D05288";
    when 16#003C9# => romdata <= X"519BA23F";
    when 16#003CA# => romdata <= X"80E8C051";
    when 16#003CB# => romdata <= X"9AF83F80";
    when 16#003CC# => romdata <= X"5780F0BC";
    when 16#003CD# => romdata <= X"085581A1";
    when 16#003CE# => romdata <= X"0B88160C";
    when 16#003CF# => romdata <= X"81900B8C";
    when 16#003D0# => romdata <= X"160C8C15";
    when 16#003D1# => romdata <= X"0870812A";
    when 16#003D2# => romdata <= X"81065154";
    when 16#003D3# => romdata <= X"73F4388C";
    when 16#003D4# => romdata <= X"15087488";
    when 16#003D5# => romdata <= X"170C5380";
    when 16#003D6# => romdata <= X"E00B8C16";
    when 16#003D7# => romdata <= X"0C8C1508";
    when 16#003D8# => romdata <= X"70812A81";
    when 16#003D9# => romdata <= X"06575475";
    when 16#003DA# => romdata <= X"F4388C15";
    when 16#003DB# => romdata <= X"0870872A";
    when 16#003DC# => romdata <= X"81067887";
    when 16#003DD# => romdata <= X"06565156";
    when 16#003DE# => romdata <= X"75802EB3";
    when 16#003DF# => romdata <= X"3873872E";
    when 16#003E0# => romdata <= X"81803881";
    when 16#003E1# => romdata <= X"177083FF";
    when 16#003E2# => romdata <= X"FF065855";
    when 16#003E3# => romdata <= X"82807726";
    when 16#003E4# => romdata <= X"FF9F3880";
    when 16#003E5# => romdata <= X"F0BC0854";
    when 16#003E6# => romdata <= X"80E00B8C";
    when 16#003E7# => romdata <= X"150C8C14";
    when 16#003E8# => romdata <= X"0870812A";
    when 16#003E9# => romdata <= X"81065856";
    when 16#003EA# => romdata <= X"76F4388A";
    when 16#003EB# => romdata <= X"3D0D0488";
    when 16#003EC# => romdata <= X"15087081";
    when 16#003ED# => romdata <= X"FF0680E7";
    when 16#003EE# => romdata <= X"CC535654";
    when 16#003EF# => romdata <= X"99E83F74";
    when 16#003F0# => romdata <= X"5288519A";
    when 16#003F1# => romdata <= X"843F80EB";
    when 16#003F2# => romdata <= X"E45199DA";
    when 16#003F3# => romdata <= X"3F755474";
    when 16#003F4# => romdata <= X"80E62EBE";
    when 16#003F5# => romdata <= X"38748D32";
    when 16#003F6# => romdata <= X"70307080";
    when 16#003F7# => romdata <= X"25760752";
    when 16#003F8# => romdata <= X"57537280";
    when 16#003F9# => romdata <= X"C138748A";
    when 16#003FA# => romdata <= X"2EBC3876";
    when 16#003FB# => romdata <= X"87068B3D";
    when 16#003FC# => romdata <= X"7105F805";
    when 16#003FD# => romdata <= X"54547473";
    when 16#003FE# => romdata <= X"3473872E";
    when 16#003FF# => romdata <= X"098106FF";
    when 16#00400# => romdata <= X"82388A3D";
    when 16#00401# => romdata <= X"F8055199";
    when 16#00402# => romdata <= X"9D3F8A51";
    when 16#00403# => romdata <= X"98FE3FFE";
    when 16#00404# => romdata <= X"F2398175";
    when 16#00405# => romdata <= X"8D327030";
    when 16#00406# => romdata <= X"70802573";
    when 16#00407# => romdata <= X"07525854";
    when 16#00408# => romdata <= X"5472802E";
    when 16#00409# => romdata <= X"C1387687";
    when 16#0040A# => romdata <= X"068B3D71";
    when 16#0040B# => romdata <= X"05F80557";
    when 16#0040C# => romdata <= X"54A07634";
    when 16#0040D# => romdata <= X"73872E09";
    when 16#0040E# => romdata <= X"8106FEC7";
    when 16#0040F# => romdata <= X"38C439FB";
    when 16#00410# => romdata <= X"3D0D9C56";
    when 16#00411# => romdata <= X"80E8C451";
    when 16#00412# => romdata <= X"98DC3F75";
    when 16#00413# => romdata <= X"52885198";
    when 16#00414# => romdata <= X"F83F80F0";
    when 16#00415# => romdata <= X"BC085481";
    when 16#00416# => romdata <= X"EC0B8815";
    when 16#00417# => romdata <= X"0C81900B";
    when 16#00418# => romdata <= X"8C150C8C";
    when 16#00419# => romdata <= X"14087081";
    when 16#0041A# => romdata <= X"2A810651";
    when 16#0041B# => romdata <= X"5372F438";
    when 16#0041C# => romdata <= X"8C140876";
    when 16#0041D# => romdata <= X"88160C53";
    when 16#0041E# => romdata <= X"900B8C15";
    when 16#0041F# => romdata <= X"0C8C1408";
    when 16#00420# => romdata <= X"70812A81";
    when 16#00421# => romdata <= X"06515574";
    when 16#00422# => romdata <= X"F4388C14";
    when 16#00423# => romdata <= X"085381ED";
    when 16#00424# => romdata <= X"0B88150C";
    when 16#00425# => romdata <= X"81900B8C";
    when 16#00426# => romdata <= X"150C8C14";
    when 16#00427# => romdata <= X"0870812A";
    when 16#00428# => romdata <= X"81065155";
    when 16#00429# => romdata <= X"74F4388C";
    when 16#0042A# => romdata <= X"14087588";
    when 16#0042B# => romdata <= X"160C5380";
    when 16#0042C# => romdata <= X"E00B8C15";
    when 16#0042D# => romdata <= X"0C8C1408";
    when 16#0042E# => romdata <= X"70812A81";
    when 16#0042F# => romdata <= X"06515372";
    when 16#00430# => romdata <= X"F4388C14";
    when 16#00431# => romdata <= X"08881508";
    when 16#00432# => romdata <= X"7081FF06";
    when 16#00433# => romdata <= X"8C170870";
    when 16#00434# => romdata <= X"872A8132";
    when 16#00435# => romdata <= X"81065852";
    when 16#00436# => romdata <= X"57515373";
    when 16#00437# => romdata <= X"802EA738";
    when 16#00438# => romdata <= X"80E8D451";
    when 16#00439# => romdata <= X"97C03F74";
    when 16#0043A# => romdata <= X"52885197";
    when 16#0043B# => romdata <= X"DC3F8A51";
    when 16#0043C# => romdata <= X"979A3F81";
    when 16#0043D# => romdata <= X"167081FF";
    when 16#0043E# => romdata <= X"06575580";
    when 16#0043F# => romdata <= X"D57627FE";
    when 16#00440# => romdata <= X"C338873D";
    when 16#00441# => romdata <= X"0D0480E8";
    when 16#00442# => romdata <= X"DC51979A";
    when 16#00443# => romdata <= X"3FE039F6";
    when 16#00444# => romdata <= X"3D0D800B";
    when 16#00445# => romdata <= X"8189E833";
    when 16#00446# => romdata <= X"8189E859";
    when 16#00447# => romdata <= X"555673A0";
    when 16#00448# => romdata <= X"2E098106";
    when 16#00449# => romdata <= X"96388116";
    when 16#0044A# => romdata <= X"7081FF06";
    when 16#0044B# => romdata <= X"8189E811";
    when 16#0044C# => romdata <= X"70335359";
    when 16#0044D# => romdata <= X"575473A0";
    when 16#0044E# => romdata <= X"2EEC3880";
    when 16#0044F# => romdata <= X"58807733";
    when 16#00450# => romdata <= X"56547474";
    when 16#00451# => romdata <= X"2E833881";
    when 16#00452# => romdata <= X"5474A02E";
    when 16#00453# => romdata <= X"83883873";
    when 16#00454# => romdata <= X"83B53874";
    when 16#00455# => romdata <= X"A02E82FE";
    when 16#00456# => romdata <= X"38811870";
    when 16#00457# => romdata <= X"81FF0659";
    when 16#00458# => romdata <= X"54817826";
    when 16#00459# => romdata <= X"D8389053";
    when 16#0045A# => romdata <= X"8C3DFC05";
    when 16#0045B# => romdata <= X"527651AC";
    when 16#0045C# => romdata <= X"D03F8008";
    when 16#0045D# => romdata <= X"81FF0659";
    when 16#0045E# => romdata <= X"800B8189";
    when 16#0045F# => romdata <= X"E8338189";
    when 16#00460# => romdata <= X"E8595556";
    when 16#00461# => romdata <= X"73A02E09";
    when 16#00462# => romdata <= X"81069638";
    when 16#00463# => romdata <= X"81167081";
    when 16#00464# => romdata <= X"FF068189";
    when 16#00465# => romdata <= X"E8117033";
    when 16#00466# => romdata <= X"57595758";
    when 16#00467# => romdata <= X"73A02EEC";
    when 16#00468# => romdata <= X"38805880";
    when 16#00469# => romdata <= X"77335654";
    when 16#0046A# => romdata <= X"74742E83";
    when 16#0046B# => romdata <= X"38815474";
    when 16#0046C# => romdata <= X"A02E82E3";
    when 16#0046D# => romdata <= X"38738390";
    when 16#0046E# => romdata <= X"3874A02E";
    when 16#0046F# => romdata <= X"82D93881";
    when 16#00470# => romdata <= X"187081FF";
    when 16#00471# => romdata <= X"06595582";
    when 16#00472# => romdata <= X"7826D838";
    when 16#00473# => romdata <= X"90538C3D";
    when 16#00474# => romdata <= X"F8055276";
    when 16#00475# => romdata <= X"51ABEA3F";
    when 16#00476# => romdata <= X"800881FF";
    when 16#00477# => romdata <= X"0680F0BC";
    when 16#00478# => romdata <= X"08565681";
    when 16#00479# => romdata <= X"EC0B8816";
    when 16#0047A# => romdata <= X"0C81900B";
    when 16#0047B# => romdata <= X"8C160C8C";
    when 16#0047C# => romdata <= X"15087081";
    when 16#0047D# => romdata <= X"2A810659";
    when 16#0047E# => romdata <= X"5777F438";
    when 16#0047F# => romdata <= X"8C150879";
    when 16#00480# => romdata <= X"88170C54";
    when 16#00481# => romdata <= X"900B8C16";
    when 16#00482# => romdata <= X"0C8C1508";
    when 16#00483# => romdata <= X"70812A81";
    when 16#00484# => romdata <= X"06595777";
    when 16#00485# => romdata <= X"F4388C15";
    when 16#00486# => romdata <= X"08768817";
    when 16#00487# => romdata <= X"0C5480D0";
    when 16#00488# => romdata <= X"0B8C160C";
    when 16#00489# => romdata <= X"8C150870";
    when 16#0048A# => romdata <= X"812A8106";
    when 16#0048B# => romdata <= X"575475F4";
    when 16#0048C# => romdata <= X"388C1508";
    when 16#0048D# => romdata <= X"5481EC0B";
    when 16#0048E# => romdata <= X"88160C81";
    when 16#0048F# => romdata <= X"900B8C16";
    when 16#00490# => romdata <= X"0C8C1508";
    when 16#00491# => romdata <= X"70812A81";
    when 16#00492# => romdata <= X"06585876";
    when 16#00493# => romdata <= X"F4388C15";
    when 16#00494# => romdata <= X"08798817";
    when 16#00495# => romdata <= X"0C54900B";
    when 16#00496# => romdata <= X"8C160C8C";
    when 16#00497# => romdata <= X"15087081";
    when 16#00498# => romdata <= X"2A81065A";
    when 16#00499# => romdata <= X"5778F438";
    when 16#0049A# => romdata <= X"8C150854";
    when 16#0049B# => romdata <= X"81ED0B88";
    when 16#0049C# => romdata <= X"160C8190";
    when 16#0049D# => romdata <= X"0B8C160C";
    when 16#0049E# => romdata <= X"8C150870";
    when 16#0049F# => romdata <= X"812A8106";
    when 16#004A0# => romdata <= X"515675F4";
    when 16#004A1# => romdata <= X"388C1508";
    when 16#004A2# => romdata <= X"7688170C";
    when 16#004A3# => romdata <= X"5480E00B";
    when 16#004A4# => romdata <= X"8C160C8C";
    when 16#004A5# => romdata <= X"15087081";
    when 16#004A6# => romdata <= X"2A81065A";
    when 16#004A7# => romdata <= X"5778F438";
    when 16#004A8# => romdata <= X"8C150888";
    when 16#004A9# => romdata <= X"16087081";
    when 16#004AA# => romdata <= X"FF068C18";
    when 16#004AB# => romdata <= X"0870872A";
    when 16#004AC# => romdata <= X"81328106";
    when 16#004AD# => romdata <= X"595C5851";
    when 16#004AE# => romdata <= X"5474802E";
    when 16#004AF# => romdata <= X"819A3880";
    when 16#004B0# => romdata <= X"E8E45193";
    when 16#004B1# => romdata <= X"E13F7552";
    when 16#004B2# => romdata <= X"885193FD";
    when 16#004B3# => romdata <= X"3F8A5193";
    when 16#004B4# => romdata <= X"BB3F8C3D";
    when 16#004B5# => romdata <= X"0D048116";
    when 16#004B6# => romdata <= X"7081FF06";
    when 16#004B7# => romdata <= X"8189E811";
    when 16#004B8# => romdata <= X"70335C52";
    when 16#004B9# => romdata <= X"575778A0";
    when 16#004BA# => romdata <= X"2E098106";
    when 16#004BB# => romdata <= X"FCEB3881";
    when 16#004BC# => romdata <= X"167081FF";
    when 16#004BD# => romdata <= X"068189E8";
    when 16#004BE# => romdata <= X"1170335C";
    when 16#004BF# => romdata <= X"52575778";
    when 16#004C0# => romdata <= X"A02ED338";
    when 16#004C1# => romdata <= X"FCD33981";
    when 16#004C2# => romdata <= X"167081FF";
    when 16#004C3# => romdata <= X"068189E8";
    when 16#004C4# => romdata <= X"11595755";
    when 16#004C5# => romdata <= X"FCA73981";
    when 16#004C6# => romdata <= X"167081FF";
    when 16#004C7# => romdata <= X"068189E8";
    when 16#004C8# => romdata <= X"11703357";
    when 16#004C9# => romdata <= X"52575773";
    when 16#004CA# => romdata <= X"A02E0981";
    when 16#004CB# => romdata <= X"06FD9038";
    when 16#004CC# => romdata <= X"81167081";
    when 16#004CD# => romdata <= X"FF068189";
    when 16#004CE# => romdata <= X"E8117033";
    when 16#004CF# => romdata <= X"57525757";
    when 16#004D0# => romdata <= X"73A02ED3";
    when 16#004D1# => romdata <= X"38FCF839";
    when 16#004D2# => romdata <= X"81167081";
    when 16#004D3# => romdata <= X"FF068189";
    when 16#004D4# => romdata <= X"E8115957";
    when 16#004D5# => romdata <= X"55FCCC39";
    when 16#004D6# => romdata <= X"80E8F051";
    when 16#004D7# => romdata <= X"92C83F8A";
    when 16#004D8# => romdata <= X"5192A93F";
    when 16#004D9# => romdata <= X"8C3D0D04";
    when 16#004DA# => romdata <= X"FF3D0D80";
    when 16#004DB# => romdata <= X"F0BC0852";
    when 16#004DC# => romdata <= X"81EC0B88";
    when 16#004DD# => romdata <= X"130C8190";
    when 16#004DE# => romdata <= X"0B8C130C";
    when 16#004DF# => romdata <= X"8C120870";
    when 16#004E0# => romdata <= X"812A7081";
    when 16#004E1# => romdata <= X"06515151";
    when 16#004E2# => romdata <= X"70F2388C";
    when 16#004E3# => romdata <= X"1208519D";
    when 16#004E4# => romdata <= X"0B88130C";
    when 16#004E5# => romdata <= X"900B8C13";
    when 16#004E6# => romdata <= X"0C8C1208";
    when 16#004E7# => romdata <= X"70812A70";
    when 16#004E8# => romdata <= X"81065151";
    when 16#004E9# => romdata <= X"5170F238";
    when 16#004EA# => romdata <= X"8C120851";
    when 16#004EB# => romdata <= X"80C50B88";
    when 16#004EC# => romdata <= X"130C80D0";
    when 16#004ED# => romdata <= X"0B8C130C";
    when 16#004EE# => romdata <= X"8C120870";
    when 16#004EF# => romdata <= X"812A7081";
    when 16#004F0# => romdata <= X"06515151";
    when 16#004F1# => romdata <= X"70F2388C";
    when 16#004F2# => romdata <= X"12085181";
    when 16#004F3# => romdata <= X"EC0B8813";
    when 16#004F4# => romdata <= X"0C81900B";
    when 16#004F5# => romdata <= X"8C130C8C";
    when 16#004F6# => romdata <= X"12087081";
    when 16#004F7# => romdata <= X"2A708106";
    when 16#004F8# => romdata <= X"51515170";
    when 16#004F9# => romdata <= X"F2388C12";
    when 16#004FA# => romdata <= X"0851A10B";
    when 16#004FB# => romdata <= X"88130C90";
    when 16#004FC# => romdata <= X"0B8C130C";
    when 16#004FD# => romdata <= X"8C120870";
    when 16#004FE# => romdata <= X"812A7081";
    when 16#004FF# => romdata <= X"06515151";
    when 16#00500# => romdata <= X"70F2388C";
    when 16#00501# => romdata <= X"12085189";
    when 16#00502# => romdata <= X"0B88130C";
    when 16#00503# => romdata <= X"80D00B8C";
    when 16#00504# => romdata <= X"130C8C12";
    when 16#00505# => romdata <= X"0870812A";
    when 16#00506# => romdata <= X"70810651";
    when 16#00507# => romdata <= X"515170F2";
    when 16#00508# => romdata <= X"388C1208";
    when 16#00509# => romdata <= X"5181EC0B";
    when 16#0050A# => romdata <= X"88130C81";
    when 16#0050B# => romdata <= X"900B8C13";
    when 16#0050C# => romdata <= X"0C8C1208";
    when 16#0050D# => romdata <= X"70812A70";
    when 16#0050E# => romdata <= X"81065151";
    when 16#0050F# => romdata <= X"5170F238";
    when 16#00510# => romdata <= X"8C120851";
    when 16#00511# => romdata <= X"B30B8813";
    when 16#00512# => romdata <= X"0C900B8C";
    when 16#00513# => romdata <= X"130C8C12";
    when 16#00514# => romdata <= X"0870812A";
    when 16#00515# => romdata <= X"70810651";
    when 16#00516# => romdata <= X"515170F2";
    when 16#00517# => romdata <= X"388C1208";
    when 16#00518# => romdata <= X"51880B88";
    when 16#00519# => romdata <= X"130C80D0";
    when 16#0051A# => romdata <= X"0B8C130C";
    when 16#0051B# => romdata <= X"8C120870";
    when 16#0051C# => romdata <= X"812A7081";
    when 16#0051D# => romdata <= X"06515151";
    when 16#0051E# => romdata <= X"70F2388C";
    when 16#0051F# => romdata <= X"12085181";
    when 16#00520# => romdata <= X"EC0B8813";
    when 16#00521# => romdata <= X"0C81900B";
    when 16#00522# => romdata <= X"8C130C8C";
    when 16#00523# => romdata <= X"12087081";
    when 16#00524# => romdata <= X"2A708106";
    when 16#00525# => romdata <= X"51515170";
    when 16#00526# => romdata <= X"F2388C12";
    when 16#00527# => romdata <= X"0851B40B";
    when 16#00528# => romdata <= X"88130C90";
    when 16#00529# => romdata <= X"0B8C130C";
    when 16#0052A# => romdata <= X"8C120870";
    when 16#0052B# => romdata <= X"812A7081";
    when 16#0052C# => romdata <= X"06515151";
    when 16#0052D# => romdata <= X"70F2388C";
    when 16#0052E# => romdata <= X"12085196";
    when 16#0052F# => romdata <= X"0B88130C";
    when 16#00530# => romdata <= X"80D00B8C";
    when 16#00531# => romdata <= X"130C8C12";
    when 16#00532# => romdata <= X"0870812A";
    when 16#00533# => romdata <= X"70810651";
    when 16#00534# => romdata <= X"515170F2";
    when 16#00535# => romdata <= X"388C1208";
    when 16#00536# => romdata <= X"5181EC0B";
    when 16#00537# => romdata <= X"88130C81";
    when 16#00538# => romdata <= X"900B8C13";
    when 16#00539# => romdata <= X"0C8C1208";
    when 16#0053A# => romdata <= X"70812A70";
    when 16#0053B# => romdata <= X"81065151";
    when 16#0053C# => romdata <= X"5170F238";
    when 16#0053D# => romdata <= X"8C120851";
    when 16#0053E# => romdata <= X"B60B8813";
    when 16#0053F# => romdata <= X"0C900B8C";
    when 16#00540# => romdata <= X"130C8C12";
    when 16#00541# => romdata <= X"0870812A";
    when 16#00542# => romdata <= X"70810651";
    when 16#00543# => romdata <= X"515170F2";
    when 16#00544# => romdata <= X"388C1208";
    when 16#00545# => romdata <= X"5180E00B";
    when 16#00546# => romdata <= X"88130C80";
    when 16#00547# => romdata <= X"D00B8C13";
    when 16#00548# => romdata <= X"0C8C1208";
    when 16#00549# => romdata <= X"70812A70";
    when 16#0054A# => romdata <= X"81065151";
    when 16#0054B# => romdata <= X"5170F238";
    when 16#0054C# => romdata <= X"8C120851";
    when 16#0054D# => romdata <= X"81EC0B88";
    when 16#0054E# => romdata <= X"130C8190";
    when 16#0054F# => romdata <= X"0B8C130C";
    when 16#00550# => romdata <= X"8C120870";
    when 16#00551# => romdata <= X"812A7081";
    when 16#00552# => romdata <= X"06515151";
    when 16#00553# => romdata <= X"70F2388C";
    when 16#00554# => romdata <= X"12085180";
    when 16#00555# => romdata <= X"C90B8813";
    when 16#00556# => romdata <= X"0C900B8C";
    when 16#00557# => romdata <= X"130C8C12";
    when 16#00558# => romdata <= X"0870812A";
    when 16#00559# => romdata <= X"70810651";
    when 16#0055A# => romdata <= X"515170F2";
    when 16#0055B# => romdata <= X"388C1208";
    when 16#0055C# => romdata <= X"5181C00B";
    when 16#0055D# => romdata <= X"88130C80";
    when 16#0055E# => romdata <= X"D00B8C13";
    when 16#0055F# => romdata <= X"0C8C1208";
    when 16#00560# => romdata <= X"70812A70";
    when 16#00561# => romdata <= X"81065151";
    when 16#00562# => romdata <= X"5170F238";
    when 16#00563# => romdata <= X"8C120851";
    when 16#00564# => romdata <= X"833D0D04";
    when 16#00565# => romdata <= X"FE3D0D80";
    when 16#00566# => romdata <= X"E980518E";
    when 16#00567# => romdata <= X"893F80E9";
    when 16#00568# => romdata <= X"A0518E82";
    when 16#00569# => romdata <= X"3F80E9E8";
    when 16#0056A# => romdata <= X"518DFB3F";
    when 16#0056B# => romdata <= X"80EAB051";
    when 16#0056C# => romdata <= X"8DF43F80";
    when 16#0056D# => romdata <= X"F0C00870";
    when 16#0056E# => romdata <= X"0852528F";
    when 16#0056F# => romdata <= X"AE3F8008";
    when 16#00570# => romdata <= X"81FF0652";
    when 16#00571# => romdata <= X"718C2793";
    when 16#00572# => romdata <= X"38A0518D";
    when 16#00573# => romdata <= X"BF3F8112";
    when 16#00574# => romdata <= X"7081FF06";
    when 16#00575# => romdata <= X"53538C72";
    when 16#00576# => romdata <= X"26EF3880";
    when 16#00577# => romdata <= X"F0C00884";
    when 16#00578# => romdata <= X"11085252";
    when 16#00579# => romdata <= X"8F853F80";
    when 16#0057A# => romdata <= X"0881FF06";
    when 16#0057B# => romdata <= X"52718C27";
    when 16#0057C# => romdata <= X"9338A051";
    when 16#0057D# => romdata <= X"8D963F81";
    when 16#0057E# => romdata <= X"127081FF";
    when 16#0057F# => romdata <= X"0653538C";
    when 16#00580# => romdata <= X"7226EF38";
    when 16#00581# => romdata <= X"80F0C008";
    when 16#00582# => romdata <= X"88110852";
    when 16#00583# => romdata <= X"528EDC3F";
    when 16#00584# => romdata <= X"800881FF";
    when 16#00585# => romdata <= X"0652718C";
    when 16#00586# => romdata <= X"279338A0";
    when 16#00587# => romdata <= X"518CED3F";
    when 16#00588# => romdata <= X"81127081";
    when 16#00589# => romdata <= X"FF065353";
    when 16#0058A# => romdata <= X"8C7226EF";
    when 16#0058B# => romdata <= X"3880F0C0";
    when 16#0058C# => romdata <= X"088C1108";
    when 16#0058D# => romdata <= X"52528EB3";
    when 16#0058E# => romdata <= X"3F800881";
    when 16#0058F# => romdata <= X"FF065271";
    when 16#00590# => romdata <= X"8C279338";
    when 16#00591# => romdata <= X"A0518CC4";
    when 16#00592# => romdata <= X"3F811270";
    when 16#00593# => romdata <= X"81FF0653";
    when 16#00594# => romdata <= X"538C7226";
    when 16#00595# => romdata <= X"EF3880EA";
    when 16#00596# => romdata <= X"CC518CCA";
    when 16#00597# => romdata <= X"3F80F0C0";
    when 16#00598# => romdata <= X"08901108";
    when 16#00599# => romdata <= X"52528E83";
    when 16#0059A# => romdata <= X"3F800881";
    when 16#0059B# => romdata <= X"FF065271";
    when 16#0059C# => romdata <= X"8C279338";
    when 16#0059D# => romdata <= X"A0518C94";
    when 16#0059E# => romdata <= X"3F811270";
    when 16#0059F# => romdata <= X"81FF0653";
    when 16#005A0# => romdata <= X"538C7226";
    when 16#005A1# => romdata <= X"EF3880F0";
    when 16#005A2# => romdata <= X"C0089411";
    when 16#005A3# => romdata <= X"0852528D";
    when 16#005A4# => romdata <= X"DA3F8008";
    when 16#005A5# => romdata <= X"81FF0652";
    when 16#005A6# => romdata <= X"718C2793";
    when 16#005A7# => romdata <= X"38A0518B";
    when 16#005A8# => romdata <= X"EB3F8112";
    when 16#005A9# => romdata <= X"7081FF06";
    when 16#005AA# => romdata <= X"53538C72";
    when 16#005AB# => romdata <= X"26EF3880";
    when 16#005AC# => romdata <= X"F0C00898";
    when 16#005AD# => romdata <= X"11085252";
    when 16#005AE# => romdata <= X"8DB13F80";
    when 16#005AF# => romdata <= X"0881FF06";
    when 16#005B0# => romdata <= X"52718C27";
    when 16#005B1# => romdata <= X"9338A051";
    when 16#005B2# => romdata <= X"8BC23F81";
    when 16#005B3# => romdata <= X"127081FF";
    when 16#005B4# => romdata <= X"0653538C";
    when 16#005B5# => romdata <= X"7226EF38";
    when 16#005B6# => romdata <= X"80F0C008";
    when 16#005B7# => romdata <= X"9C110852";
    when 16#005B8# => romdata <= X"528D883F";
    when 16#005B9# => romdata <= X"800881FF";
    when 16#005BA# => romdata <= X"0652718C";
    when 16#005BB# => romdata <= X"279338A0";
    when 16#005BC# => romdata <= X"518B993F";
    when 16#005BD# => romdata <= X"81127081";
    when 16#005BE# => romdata <= X"FF065353";
    when 16#005BF# => romdata <= X"8C7226EF";
    when 16#005C0# => romdata <= X"3880EAE8";
    when 16#005C1# => romdata <= X"518B9F3F";
    when 16#005C2# => romdata <= X"80F0C008";
    when 16#005C3# => romdata <= X"53810BB0";
    when 16#005C4# => romdata <= X"140CB013";
    when 16#005C5# => romdata <= X"08527180";
    when 16#005C6# => romdata <= X"25F838A0";
    when 16#005C7# => romdata <= X"1308518C";
    when 16#005C8# => romdata <= X"CA3F8008";
    when 16#005C9# => romdata <= X"81FF0652";
    when 16#005CA# => romdata <= X"718C2793";
    when 16#005CB# => romdata <= X"38A0518A";
    when 16#005CC# => romdata <= X"DB3F8112";
    when 16#005CD# => romdata <= X"7081FF06";
    when 16#005CE# => romdata <= X"53538C72";
    when 16#005CF# => romdata <= X"26EF3880";
    when 16#005D0# => romdata <= X"F0C008A4";
    when 16#005D1# => romdata <= X"11085252";
    when 16#005D2# => romdata <= X"8CA13F80";
    when 16#005D3# => romdata <= X"0881FF06";
    when 16#005D4# => romdata <= X"52718C27";
    when 16#005D5# => romdata <= X"9338A051";
    when 16#005D6# => romdata <= X"8AB23F81";
    when 16#005D7# => romdata <= X"127081FF";
    when 16#005D8# => romdata <= X"0653538C";
    when 16#005D9# => romdata <= X"7226EF38";
    when 16#005DA# => romdata <= X"80F0C008";
    when 16#005DB# => romdata <= X"A8110852";
    when 16#005DC# => romdata <= X"528BF83F";
    when 16#005DD# => romdata <= X"800881FF";
    when 16#005DE# => romdata <= X"0652718C";
    when 16#005DF# => romdata <= X"279338A0";
    when 16#005E0# => romdata <= X"518A893F";
    when 16#005E1# => romdata <= X"81127081";
    when 16#005E2# => romdata <= X"FF065353";
    when 16#005E3# => romdata <= X"8C7226EF";
    when 16#005E4# => romdata <= X"3880F0C0";
    when 16#005E5# => romdata <= X"08AC1108";
    when 16#005E6# => romdata <= X"52528BCF";
    when 16#005E7# => romdata <= X"3F800881";
    when 16#005E8# => romdata <= X"FF065271";
    when 16#005E9# => romdata <= X"8C279338";
    when 16#005EA# => romdata <= X"A05189E0";
    when 16#005EB# => romdata <= X"3F811270";
    when 16#005EC# => romdata <= X"81FF0653";
    when 16#005ED# => romdata <= X"538C7226";
    when 16#005EE# => romdata <= X"EF3880EB";
    when 16#005EF# => romdata <= X"845189E6";
    when 16#005F0# => romdata <= X"3F80F0C0";
    when 16#005F1# => romdata <= X"08B01108";
    when 16#005F2# => romdata <= X"FE0A0652";
    when 16#005F3# => romdata <= X"538B9C3F";
    when 16#005F4# => romdata <= X"80F0C008";
    when 16#005F5# => romdata <= X"53800BB0";
    when 16#005F6# => romdata <= X"140C80EB";
    when 16#005F7# => romdata <= X"985189C6";
    when 16#005F8# => romdata <= X"3F80EBB0";
    when 16#005F9# => romdata <= X"5189BF3F";
    when 16#005FA# => romdata <= X"80F0C008";
    when 16#005FB# => romdata <= X"80C01108";
    when 16#005FC# => romdata <= X"52528AF7";
    when 16#005FD# => romdata <= X"3F800881";
    when 16#005FE# => romdata <= X"FF065271";
    when 16#005FF# => romdata <= X"98279338";
    when 16#00600# => romdata <= X"A0518988";
    when 16#00601# => romdata <= X"3F811270";
    when 16#00602# => romdata <= X"81FF0651";
    when 16#00603# => romdata <= X"52987226";
    when 16#00604# => romdata <= X"EF3880F0";
    when 16#00605# => romdata <= X"C00880C8";
    when 16#00606# => romdata <= X"11085253";
    when 16#00607# => romdata <= X"8ACD3F80";
    when 16#00608# => romdata <= X"0881FF06";
    when 16#00609# => romdata <= X"52719827";
    when 16#0060A# => romdata <= X"9338A051";
    when 16#0060B# => romdata <= X"88DE3F81";
    when 16#0060C# => romdata <= X"127081FF";
    when 16#0060D# => romdata <= X"06515298";
    when 16#0060E# => romdata <= X"7226EF38";
    when 16#0060F# => romdata <= X"80EBCC51";
    when 16#00610# => romdata <= X"88E43F80";
    when 16#00611# => romdata <= X"F0C00880";
    when 16#00612# => romdata <= X"C4110852";
    when 16#00613# => romdata <= X"538A9C3F";
    when 16#00614# => romdata <= X"800881FF";
    when 16#00615# => romdata <= X"06527198";
    when 16#00616# => romdata <= X"279338A0";
    when 16#00617# => romdata <= X"5188AD3F";
    when 16#00618# => romdata <= X"81127081";
    when 16#00619# => romdata <= X"FF065152";
    when 16#0061A# => romdata <= X"987226EF";
    when 16#0061B# => romdata <= X"3880F0C0";
    when 16#0061C# => romdata <= X"0880CC11";
    when 16#0061D# => romdata <= X"08525389";
    when 16#0061E# => romdata <= X"F23F8008";
    when 16#0061F# => romdata <= X"81FF0652";
    when 16#00620# => romdata <= X"71982793";
    when 16#00621# => romdata <= X"38A05188";
    when 16#00622# => romdata <= X"833F8112";
    when 16#00623# => romdata <= X"7081FF06";
    when 16#00624# => romdata <= X"51529872";
    when 16#00625# => romdata <= X"26EF388A";
    when 16#00626# => romdata <= X"5187F13F";
    when 16#00627# => romdata <= X"80F0C008";
    when 16#00628# => romdata <= X"B4110870";
    when 16#00629# => romdata <= X"81FF0680";
    when 16#0062A# => romdata <= X"EBE85452";
    when 16#0062B# => romdata <= X"545287F6";
    when 16#0062C# => romdata <= X"3F715189";
    when 16#0062D# => romdata <= X"B63FA051";
    when 16#0062E# => romdata <= X"87D23F71";
    when 16#0062F# => romdata <= X"86269338";
    when 16#00630# => romdata <= X"71101080";
    when 16#00631# => romdata <= X"EDB80553";
    when 16#00632# => romdata <= X"72080480";
    when 16#00633# => romdata <= X"EBFC5187";
    when 16#00634# => romdata <= X"D53F8A51";
    when 16#00635# => romdata <= X"87B63F84";
    when 16#00636# => romdata <= X"3D0D0480";
    when 16#00637# => romdata <= X"EC885187";
    when 16#00638# => romdata <= X"C53FEF39";
    when 16#00639# => romdata <= X"80EC9451";
    when 16#0063A# => romdata <= X"87BC3FE6";
    when 16#0063B# => romdata <= X"3980ECA0";
    when 16#0063C# => romdata <= X"5187B33F";
    when 16#0063D# => romdata <= X"DD3980EC";
    when 16#0063E# => romdata <= X"A45187AA";
    when 16#0063F# => romdata <= X"3FD43980";
    when 16#00640# => romdata <= X"ECB05187";
    when 16#00641# => romdata <= X"A13FCB39";
    when 16#00642# => romdata <= X"80ECBC51";
    when 16#00643# => romdata <= X"87983FC2";
    when 16#00644# => romdata <= X"39FC3D0D";
    when 16#00645# => romdata <= X"80F0C808";
    when 16#00646# => romdata <= X"7008810A";
    when 16#00647# => romdata <= X"068180C4";
    when 16#00648# => romdata <= X"0C538AAE";
    when 16#00649# => romdata <= X"3F8ADC3F";
    when 16#0064A# => romdata <= X"8180C408";
    when 16#0064B# => romdata <= X"B8F65452";
    when 16#0064C# => romdata <= X"7184388A";
    when 16#0064D# => romdata <= X"F5537281";
    when 16#0064E# => romdata <= X"8ACC0C71";
    when 16#0064F# => romdata <= X"802E8298";
    when 16#00650# => romdata <= X"3880E8C0";
    when 16#00651# => romdata <= X"5186DF3F";
    when 16#00652# => romdata <= X"8C5186C0";
    when 16#00653# => romdata <= X"3F80ECC8";
    when 16#00654# => romdata <= X"5186D33F";
    when 16#00655# => romdata <= X"8180C408";
    when 16#00656# => romdata <= X"802E80F2";
    when 16#00657# => romdata <= X"3880ECE0";
    when 16#00658# => romdata <= X"5186C33F";
    when 16#00659# => romdata <= X"8180C408";
    when 16#0065A# => romdata <= X"802E81C4";
    when 16#0065B# => romdata <= X"3880F0C0";
    when 16#0065C# => romdata <= X"0853800B";
    when 16#0065D# => romdata <= X"B4140CF8";
    when 16#0065E# => romdata <= X"9B3FF881";
    when 16#0065F# => romdata <= X"C08E8053";
    when 16#00660# => romdata <= X"9F0B80F0";
    when 16#00661# => romdata <= X"C8085555";
    when 16#00662# => romdata <= X"8180C408";
    when 16#00663# => romdata <= X"802E80FB";
    when 16#00664# => romdata <= X"387281FF";
    when 16#00665# => romdata <= X"0684150C";
    when 16#00666# => romdata <= X"818AC808";
    when 16#00667# => romdata <= X"5271802E";
    when 16#00668# => romdata <= X"9F38729F";
    when 16#00669# => romdata <= X"2A731007";
    when 16#0066A# => romdata <= X"5374802E";
    when 16#0066B# => romdata <= X"9E38FF15";
    when 16#0066C# => romdata <= X"7381FF06";
    when 16#0066D# => romdata <= X"84160C81";
    when 16#0066E# => romdata <= X"8AC80853";
    when 16#0066F# => romdata <= X"5571E338";
    when 16#00670# => romdata <= X"72812A73";
    when 16#00671# => romdata <= X"9F2B0753";
    when 16#00672# => romdata <= X"74E43890";
    when 16#00673# => romdata <= X"BE3F80EC";
    when 16#00674# => romdata <= X"EC5185D2";
    when 16#00675# => romdata <= X"3F80ED90";
    when 16#00676# => romdata <= X"5185CB3F";
    when 16#00677# => romdata <= X"B451878B";
    when 16#00678# => romdata <= X"3F80EDA0";
    when 16#00679# => romdata <= X"5185BF3F";
    when 16#0067A# => romdata <= X"80EDA851";
    when 16#0067B# => romdata <= X"85B83F81";
    when 16#0067C# => romdata <= X"80C408FE";
    when 16#0067D# => romdata <= X"F838B939";
    when 16#0067E# => romdata <= X"72812A73";
    when 16#0067F# => romdata <= X"9F2B0753";
    when 16#00680# => romdata <= X"80FD5188";
    when 16#00681# => romdata <= X"AA3F80F0";
    when 16#00682# => romdata <= X"C8085472";
    when 16#00683# => romdata <= X"81FF0684";
    when 16#00684# => romdata <= X"150C818A";
    when 16#00685# => romdata <= X"C8085574";
    when 16#00686# => romdata <= X"802EDD38";
    when 16#00687# => romdata <= X"729F2A73";
    when 16#00688# => romdata <= X"10075380";
    when 16#00689# => romdata <= X"FD518887";
    when 16#0068A# => romdata <= X"3F80F0C8";
    when 16#0068B# => romdata <= X"0854DC39";
    when 16#0068C# => romdata <= X"DAA73F80";
    when 16#0068D# => romdata <= X"F0C00853";
    when 16#0068E# => romdata <= X"800BB414";
    when 16#0068F# => romdata <= X"0CF6D53F";
    when 16#00690# => romdata <= X"F881C08E";
    when 16#00691# => romdata <= X"80539F0B";
    when 16#00692# => romdata <= X"80F0C808";
    when 16#00693# => romdata <= X"55558180";
    when 16#00694# => romdata <= X"C408FEBD";
    when 16#00695# => romdata <= X"38FFB439";
    when 16#00696# => romdata <= X"89C43F80";
    when 16#00697# => romdata <= X"F0BC0853";
    when 16#00698# => romdata <= X"99730C81";
    when 16#00699# => romdata <= X"800B8414";
    when 16#0069A# => romdata <= X"0C80F0B8";
    when 16#0069B# => romdata <= X"08549974";
    when 16#0069C# => romdata <= X"0C81800B";
    when 16#0069D# => romdata <= X"84150C81";
    when 16#0069E# => romdata <= X"EC0B8814";
    when 16#0069F# => romdata <= X"0C81900B";
    when 16#006A0# => romdata <= X"8C140C8C";
    when 16#006A1# => romdata <= X"13087081";
    when 16#006A2# => romdata <= X"2A810656";
    when 16#006A3# => romdata <= X"5474F438";
    when 16#006A4# => romdata <= X"8C130852";
    when 16#006A5# => romdata <= X"9D0B8814";
    when 16#006A6# => romdata <= X"0C900B8C";
    when 16#006A7# => romdata <= X"140C8C13";
    when 16#006A8# => romdata <= X"0870812A";
    when 16#006A9# => romdata <= X"81065654";
    when 16#006AA# => romdata <= X"74F4388C";
    when 16#006AB# => romdata <= X"13085280";
    when 16#006AC# => romdata <= X"C50B8814";
    when 16#006AD# => romdata <= X"0C80D00B";
    when 16#006AE# => romdata <= X"8C140C8C";
    when 16#006AF# => romdata <= X"13087081";
    when 16#006B0# => romdata <= X"2A810656";
    when 16#006B1# => romdata <= X"5474F438";
    when 16#006B2# => romdata <= X"8C130852";
    when 16#006B3# => romdata <= X"81EC0B88";
    when 16#006B4# => romdata <= X"140C8190";
    when 16#006B5# => romdata <= X"0B8C140C";
    when 16#006B6# => romdata <= X"8C130870";
    when 16#006B7# => romdata <= X"812A8106";
    when 16#006B8# => romdata <= X"565474F4";
    when 16#006B9# => romdata <= X"388C1308";
    when 16#006BA# => romdata <= X"52A10B88";
    when 16#006BB# => romdata <= X"140C900B";
    when 16#006BC# => romdata <= X"8C140C8C";
    when 16#006BD# => romdata <= X"13087081";
    when 16#006BE# => romdata <= X"2A810656";
    when 16#006BF# => romdata <= X"5474F438";
    when 16#006C0# => romdata <= X"8C130852";
    when 16#006C1# => romdata <= X"890B8814";
    when 16#006C2# => romdata <= X"0C80D00B";
    when 16#006C3# => romdata <= X"8C140C8C";
    when 16#006C4# => romdata <= X"13087081";
    when 16#006C5# => romdata <= X"2A810656";
    when 16#006C6# => romdata <= X"5474F438";
    when 16#006C7# => romdata <= X"8C130852";
    when 16#006C8# => romdata <= X"81EC0B88";
    when 16#006C9# => romdata <= X"140C8190";
    when 16#006CA# => romdata <= X"0B8C140C";
    when 16#006CB# => romdata <= X"8C130870";
    when 16#006CC# => romdata <= X"812A8106";
    when 16#006CD# => romdata <= X"565474F4";
    when 16#006CE# => romdata <= X"388C1308";
    when 16#006CF# => romdata <= X"52B30B88";
    when 16#006D0# => romdata <= X"140C900B";
    when 16#006D1# => romdata <= X"8C140C8C";
    when 16#006D2# => romdata <= X"13087081";
    when 16#006D3# => romdata <= X"2A810656";
    when 16#006D4# => romdata <= X"5474F438";
    when 16#006D5# => romdata <= X"8C130852";
    when 16#006D6# => romdata <= X"880B8814";
    when 16#006D7# => romdata <= X"0C80D00B";
    when 16#006D8# => romdata <= X"8C140C8C";
    when 16#006D9# => romdata <= X"13087081";
    when 16#006DA# => romdata <= X"2A810656";
    when 16#006DB# => romdata <= X"5474F438";
    when 16#006DC# => romdata <= X"8C130852";
    when 16#006DD# => romdata <= X"81EC0B88";
    when 16#006DE# => romdata <= X"140C8190";
    when 16#006DF# => romdata <= X"0B8C140C";
    when 16#006E0# => romdata <= X"8C130870";
    when 16#006E1# => romdata <= X"812A8106";
    when 16#006E2# => romdata <= X"565474F4";
    when 16#006E3# => romdata <= X"388C1308";
    when 16#006E4# => romdata <= X"52B40B88";
    when 16#006E5# => romdata <= X"140C900B";
    when 16#006E6# => romdata <= X"8C140C8C";
    when 16#006E7# => romdata <= X"13087081";
    when 16#006E8# => romdata <= X"2A810656";
    when 16#006E9# => romdata <= X"5474F438";
    when 16#006EA# => romdata <= X"8C130852";
    when 16#006EB# => romdata <= X"960B8814";
    when 16#006EC# => romdata <= X"0C80D00B";
    when 16#006ED# => romdata <= X"8C140C8C";
    when 16#006EE# => romdata <= X"13087081";
    when 16#006EF# => romdata <= X"2A810656";
    when 16#006F0# => romdata <= X"5474F438";
    when 16#006F1# => romdata <= X"8C130852";
    when 16#006F2# => romdata <= X"81EC0B88";
    when 16#006F3# => romdata <= X"140C8190";
    when 16#006F4# => romdata <= X"0B8C140C";
    when 16#006F5# => romdata <= X"8C130870";
    when 16#006F6# => romdata <= X"812A8106";
    when 16#006F7# => romdata <= X"565474F4";
    when 16#006F8# => romdata <= X"388C1308";
    when 16#006F9# => romdata <= X"52B60B88";
    when 16#006FA# => romdata <= X"140C900B";
    when 16#006FB# => romdata <= X"8C140C8C";
    when 16#006FC# => romdata <= X"13087081";
    when 16#006FD# => romdata <= X"2A810656";
    when 16#006FE# => romdata <= X"5474F438";
    when 16#006FF# => romdata <= X"8C130852";
    when 16#00700# => romdata <= X"80E00B88";
    when 16#00701# => romdata <= X"140C80D0";
    when 16#00702# => romdata <= X"0B8C140C";
    when 16#00703# => romdata <= X"8C130870";
    when 16#00704# => romdata <= X"812A8106";
    when 16#00705# => romdata <= X"565474F4";
    when 16#00706# => romdata <= X"388C1308";
    when 16#00707# => romdata <= X"5281EC0B";
    when 16#00708# => romdata <= X"88140C81";
    when 16#00709# => romdata <= X"900B8C14";
    when 16#0070A# => romdata <= X"0C8C1308";
    when 16#0070B# => romdata <= X"70812A81";
    when 16#0070C# => romdata <= X"06565474";
    when 16#0070D# => romdata <= X"F4388C13";
    when 16#0070E# => romdata <= X"085280C9";
    when 16#0070F# => romdata <= X"0B88140C";
    when 16#00710# => romdata <= X"900B8C14";
    when 16#00711# => romdata <= X"0C8C1308";
    when 16#00712# => romdata <= X"70812A81";
    when 16#00713# => romdata <= X"06565474";
    when 16#00714# => romdata <= X"F4388C13";
    when 16#00715# => romdata <= X"085281C0";
    when 16#00716# => romdata <= X"0B88140C";
    when 16#00717# => romdata <= X"80D00B8C";
    when 16#00718# => romdata <= X"140C8C13";
    when 16#00719# => romdata <= X"0870812A";
    when 16#0071A# => romdata <= X"81065654";
    when 16#0071B# => romdata <= X"74F4388C";
    when 16#0071C# => romdata <= X"130852F9";
    when 16#0071D# => romdata <= X"CC39FF3D";
    when 16#0071E# => romdata <= X"0D028F05";
    when 16#0071F# => romdata <= X"3380F0D4";
    when 16#00720# => romdata <= X"0852710C";
    when 16#00721# => romdata <= X"800B800C";
    when 16#00722# => romdata <= X"833D0D04";
    when 16#00723# => romdata <= X"FF3D0D02";
    when 16#00724# => romdata <= X"8F053351";
    when 16#00725# => romdata <= X"818ACC08";
    when 16#00726# => romdata <= X"52712D80";
    when 16#00727# => romdata <= X"0881FF06";
    when 16#00728# => romdata <= X"800C833D";
    when 16#00729# => romdata <= X"0D04FE3D";
    when 16#0072A# => romdata <= X"0D747033";
    when 16#0072B# => romdata <= X"53537180";
    when 16#0072C# => romdata <= X"2E933881";
    when 16#0072D# => romdata <= X"13725281";
    when 16#0072E# => romdata <= X"8ACC0853";
    when 16#0072F# => romdata <= X"53712D72";
    when 16#00730# => romdata <= X"335271EF";
    when 16#00731# => romdata <= X"38843D0D";
    when 16#00732# => romdata <= X"04F43D0D";
    when 16#00733# => romdata <= X"7F028405";
    when 16#00734# => romdata <= X"BB053355";
    when 16#00735# => romdata <= X"57880B8C";
    when 16#00736# => romdata <= X"3D5A5A89";
    when 16#00737# => romdata <= X"5380EDF8";
    when 16#00738# => romdata <= X"5278518A";
    when 16#00739# => romdata <= X"B33F737A";
    when 16#0073A# => romdata <= X"2E80FA38";
    when 16#0073B# => romdata <= X"79567390";
    when 16#0073C# => romdata <= X"2E80E738";
    when 16#0073D# => romdata <= X"02A70558";
    when 16#0073E# => romdata <= X"768F0654";
    when 16#0073F# => romdata <= X"738926BF";
    when 16#00740# => romdata <= X"387518B0";
    when 16#00741# => romdata <= X"15555573";
    when 16#00742# => romdata <= X"75347684";
    when 16#00743# => romdata <= X"2AFF1770";
    when 16#00744# => romdata <= X"81FF0658";
    when 16#00745# => romdata <= X"555775E0";
    when 16#00746# => romdata <= X"38791955";
    when 16#00747# => romdata <= X"75753478";
    when 16#00748# => romdata <= X"70335555";
    when 16#00749# => romdata <= X"73802E93";
    when 16#0074A# => romdata <= X"38811574";
    when 16#0074B# => romdata <= X"52818ACC";
    when 16#0074C# => romdata <= X"08575575";
    when 16#0074D# => romdata <= X"2D743354";
    when 16#0074E# => romdata <= X"73EF388E";
    when 16#0074F# => romdata <= X"3D0D0475";
    when 16#00750# => romdata <= X"18B71555";
    when 16#00751# => romdata <= X"55737534";
    when 16#00752# => romdata <= X"76842AFF";
    when 16#00753# => romdata <= X"177081FF";
    when 16#00754# => romdata <= X"06585557";
    when 16#00755# => romdata <= X"75FFA138";
    when 16#00756# => romdata <= X"C0398470";
    when 16#00757# => romdata <= X"575A02A7";
    when 16#00758# => romdata <= X"0558FF94";
    when 16#00759# => romdata <= X"39827057";
    when 16#0075A# => romdata <= X"5AF439F2";
    when 16#0075B# => romdata <= X"3D0D608C";
    when 16#0075C# => romdata <= X"3D705B5B";
    when 16#0075D# => romdata <= X"53807356";
    when 16#0075E# => romdata <= X"57767324";
    when 16#0075F# => romdata <= X"81803878";
    when 16#00760# => romdata <= X"17548A52";
    when 16#00761# => romdata <= X"745184E2";
    when 16#00762# => romdata <= X"3F8008B0";
    when 16#00763# => romdata <= X"05537274";
    when 16#00764# => romdata <= X"34811757";
    when 16#00765# => romdata <= X"8A527451";
    when 16#00766# => romdata <= X"84AB3F80";
    when 16#00767# => romdata <= X"08558008";
    when 16#00768# => romdata <= X"DE388008";
    when 16#00769# => romdata <= X"779F2A18";
    when 16#0076A# => romdata <= X"70812C5A";
    when 16#0076B# => romdata <= X"56568078";
    when 16#0076C# => romdata <= X"259E3878";
    when 16#0076D# => romdata <= X"17FF0555";
    when 16#0076E# => romdata <= X"75197033";
    when 16#0076F# => romdata <= X"55537433";
    when 16#00770# => romdata <= X"73347375";
    when 16#00771# => romdata <= X"348116FF";
    when 16#00772# => romdata <= X"16565677";
    when 16#00773# => romdata <= X"7624E938";
    when 16#00774# => romdata <= X"76195680";
    when 16#00775# => romdata <= X"76347681";
    when 16#00776# => romdata <= X"FF067A70";
    when 16#00777# => romdata <= X"33555654";
    when 16#00778# => romdata <= X"72802E93";
    when 16#00779# => romdata <= X"38811573";
    when 16#0077A# => romdata <= X"52818ACC";
    when 16#0077B# => romdata <= X"08585576";
    when 16#0077C# => romdata <= X"2D743353";
    when 16#0077D# => romdata <= X"72EF3873";
    when 16#0077E# => romdata <= X"800C903D";
    when 16#0077F# => romdata <= X"0D04AD7A";
    when 16#00780# => romdata <= X"3402A905";
    when 16#00781# => romdata <= X"73307119";
    when 16#00782# => romdata <= X"5656598A";
    when 16#00783# => romdata <= X"52745183";
    when 16#00784# => romdata <= X"D93F8008";
    when 16#00785# => romdata <= X"B0055372";
    when 16#00786# => romdata <= X"74348117";
    when 16#00787# => romdata <= X"578A5274";
    when 16#00788# => romdata <= X"5183A23F";
    when 16#00789# => romdata <= X"80085580";
    when 16#0078A# => romdata <= X"08FED438";
    when 16#0078B# => romdata <= X"FEF439FD";
    when 16#0078C# => romdata <= X"3D0D80F0";
    when 16#0078D# => romdata <= X"CC0876B2";
    when 16#0078E# => romdata <= X"E4299412";
    when 16#0078F# => romdata <= X"0C54850B";
    when 16#00790# => romdata <= X"98150C98";
    when 16#00791# => romdata <= X"14087081";
    when 16#00792# => romdata <= X"06515372";
    when 16#00793# => romdata <= X"F638853D";
    when 16#00794# => romdata <= X"0D04803D";
    when 16#00795# => romdata <= X"0D80F0CC";
    when 16#00796# => romdata <= X"0851870B";
    when 16#00797# => romdata <= X"84120CFF";
    when 16#00798# => romdata <= X"0BB4120C";
    when 16#00799# => romdata <= X"A70BB812";
    when 16#0079A# => romdata <= X"0C87E80B";
    when 16#0079B# => romdata <= X"A4120CA7";
    when 16#0079C# => romdata <= X"0BA8120C";
    when 16#0079D# => romdata <= X"B2E40B94";
    when 16#0079E# => romdata <= X"120C870B";
    when 16#0079F# => romdata <= X"98120C82";
    when 16#007A0# => romdata <= X"3D0D0480";
    when 16#007A1# => romdata <= X"3D0D80F0";
    when 16#007A2# => romdata <= X"D00851B8";
    when 16#007A3# => romdata <= X"0B8C120C";
    when 16#007A4# => romdata <= X"830B8812";
    when 16#007A5# => romdata <= X"0C823D0D";
    when 16#007A6# => romdata <= X"04803D0D";
    when 16#007A7# => romdata <= X"80F0D008";
    when 16#007A8# => romdata <= X"84110881";
    when 16#007A9# => romdata <= X"06800C51";
    when 16#007AA# => romdata <= X"823D0D04";
    when 16#007AB# => romdata <= X"FF3D0D80";
    when 16#007AC# => romdata <= X"F0D00852";
    when 16#007AD# => romdata <= X"84120870";
    when 16#007AE# => romdata <= X"81065151";
    when 16#007AF# => romdata <= X"70802EF4";
    when 16#007B0# => romdata <= X"38710870";
    when 16#007B1# => romdata <= X"81FF0680";
    when 16#007B2# => romdata <= X"0C51833D";
    when 16#007B3# => romdata <= X"0D04FE3D";
    when 16#007B4# => romdata <= X"0D029305";
    when 16#007B5# => romdata <= X"3353728A";
    when 16#007B6# => romdata <= X"2E9C3880";
    when 16#007B7# => romdata <= X"F0D00852";
    when 16#007B8# => romdata <= X"84120870";
    when 16#007B9# => romdata <= X"892A7081";
    when 16#007BA# => romdata <= X"06515151";
    when 16#007BB# => romdata <= X"70F23872";
    when 16#007BC# => romdata <= X"720C843D";
    when 16#007BD# => romdata <= X"0D0480F0";
    when 16#007BE# => romdata <= X"D0085284";
    when 16#007BF# => romdata <= X"12087089";
    when 16#007C0# => romdata <= X"2A708106";
    when 16#007C1# => romdata <= X"51515170";
    when 16#007C2# => romdata <= X"F2388D72";
    when 16#007C3# => romdata <= X"0C841208";
    when 16#007C4# => romdata <= X"70892A70";
    when 16#007C5# => romdata <= X"81065151";
    when 16#007C6# => romdata <= X"5170C538";
    when 16#007C7# => romdata <= X"D239803D";
    when 16#007C8# => romdata <= X"0D80F0C4";
    when 16#007C9# => romdata <= X"0851800B";
    when 16#007CA# => romdata <= X"84120C83";
    when 16#007CB# => romdata <= X"FE800B88";
    when 16#007CC# => romdata <= X"120C800B";
    when 16#007CD# => romdata <= X"818AD034";
    when 16#007CE# => romdata <= X"800B818A";
    when 16#007CF# => romdata <= X"D434823D";
    when 16#007D0# => romdata <= X"0D04FA3D";
    when 16#007D1# => romdata <= X"0D02A305";
    when 16#007D2# => romdata <= X"3380F0C4";
    when 16#007D3# => romdata <= X"08818AD0";
    when 16#007D4# => romdata <= X"337081FF";
    when 16#007D5# => romdata <= X"06701010";
    when 16#007D6# => romdata <= X"11818AD4";
    when 16#007D7# => romdata <= X"337081FF";
    when 16#007D8# => romdata <= X"06729029";
    when 16#007D9# => romdata <= X"1170882B";
    when 16#007DA# => romdata <= X"7807770C";
    when 16#007DB# => romdata <= X"535B5B55";
    when 16#007DC# => romdata <= X"55595454";
    when 16#007DD# => romdata <= X"738A2E98";
    when 16#007DE# => romdata <= X"387480CF";
    when 16#007DF# => romdata <= X"2E923873";
    when 16#007E0# => romdata <= X"8C2EA438";
    when 16#007E1# => romdata <= X"81165372";
    when 16#007E2# => romdata <= X"818AD434";
    when 16#007E3# => romdata <= X"883D0D04";
    when 16#007E4# => romdata <= X"71A326A3";
    when 16#007E5# => romdata <= X"38811752";
    when 16#007E6# => romdata <= X"71818AD0";
    when 16#007E7# => romdata <= X"34800B81";
    when 16#007E8# => romdata <= X"8AD43488";
    when 16#007E9# => romdata <= X"3D0D0480";
    when 16#007EA# => romdata <= X"5271882B";
    when 16#007EB# => romdata <= X"730C8112";
    when 16#007EC# => romdata <= X"52979072";
    when 16#007ED# => romdata <= X"26F33880";
    when 16#007EE# => romdata <= X"0B818AD0";
    when 16#007EF# => romdata <= X"34800B81";
    when 16#007F0# => romdata <= X"8AD434DF";
    when 16#007F1# => romdata <= X"398C0802";
    when 16#007F2# => romdata <= X"8C0CFD3D";
    when 16#007F3# => romdata <= X"0D80538C";
    when 16#007F4# => romdata <= X"088C0508";
    when 16#007F5# => romdata <= X"528C0888";
    when 16#007F6# => romdata <= X"05085182";
    when 16#007F7# => romdata <= X"DE3F8008";
    when 16#007F8# => romdata <= X"70800C54";
    when 16#007F9# => romdata <= X"853D0D8C";
    when 16#007FA# => romdata <= X"0C048C08";
    when 16#007FB# => romdata <= X"028C0CFD";
    when 16#007FC# => romdata <= X"3D0D8153";
    when 16#007FD# => romdata <= X"8C088C05";
    when 16#007FE# => romdata <= X"08528C08";
    when 16#007FF# => romdata <= X"88050851";
    when 16#00800# => romdata <= X"82B93F80";
    when 16#00801# => romdata <= X"0870800C";
    when 16#00802# => romdata <= X"54853D0D";
    when 16#00803# => romdata <= X"8C0C048C";
    when 16#00804# => romdata <= X"08028C0C";
    when 16#00805# => romdata <= X"F93D0D80";
    when 16#00806# => romdata <= X"0B8C08FC";
    when 16#00807# => romdata <= X"050C8C08";
    when 16#00808# => romdata <= X"88050880";
    when 16#00809# => romdata <= X"25AB388C";
    when 16#0080A# => romdata <= X"08880508";
    when 16#0080B# => romdata <= X"308C0888";
    when 16#0080C# => romdata <= X"050C800B";
    when 16#0080D# => romdata <= X"8C08F405";
    when 16#0080E# => romdata <= X"0C8C08FC";
    when 16#0080F# => romdata <= X"05088838";
    when 16#00810# => romdata <= X"810B8C08";
    when 16#00811# => romdata <= X"F4050C8C";
    when 16#00812# => romdata <= X"08F40508";
    when 16#00813# => romdata <= X"8C08FC05";
    when 16#00814# => romdata <= X"0C8C088C";
    when 16#00815# => romdata <= X"05088025";
    when 16#00816# => romdata <= X"AB388C08";
    when 16#00817# => romdata <= X"8C050830";
    when 16#00818# => romdata <= X"8C088C05";
    when 16#00819# => romdata <= X"0C800B8C";
    when 16#0081A# => romdata <= X"08F0050C";
    when 16#0081B# => romdata <= X"8C08FC05";
    when 16#0081C# => romdata <= X"08883881";
    when 16#0081D# => romdata <= X"0B8C08F0";
    when 16#0081E# => romdata <= X"050C8C08";
    when 16#0081F# => romdata <= X"F005088C";
    when 16#00820# => romdata <= X"08FC050C";
    when 16#00821# => romdata <= X"80538C08";
    when 16#00822# => romdata <= X"8C050852";
    when 16#00823# => romdata <= X"8C088805";
    when 16#00824# => romdata <= X"085181A7";
    when 16#00825# => romdata <= X"3F800870";
    when 16#00826# => romdata <= X"8C08F805";
    when 16#00827# => romdata <= X"0C548C08";
    when 16#00828# => romdata <= X"FC050880";
    when 16#00829# => romdata <= X"2E8C388C";
    when 16#0082A# => romdata <= X"08F80508";
    when 16#0082B# => romdata <= X"308C08F8";
    when 16#0082C# => romdata <= X"050C8C08";
    when 16#0082D# => romdata <= X"F8050870";
    when 16#0082E# => romdata <= X"800C5489";
    when 16#0082F# => romdata <= X"3D0D8C0C";
    when 16#00830# => romdata <= X"048C0802";
    when 16#00831# => romdata <= X"8C0CFB3D";
    when 16#00832# => romdata <= X"0D800B8C";
    when 16#00833# => romdata <= X"08FC050C";
    when 16#00834# => romdata <= X"8C088805";
    when 16#00835# => romdata <= X"08802593";
    when 16#00836# => romdata <= X"388C0888";
    when 16#00837# => romdata <= X"0508308C";
    when 16#00838# => romdata <= X"0888050C";
    when 16#00839# => romdata <= X"810B8C08";
    when 16#0083A# => romdata <= X"FC050C8C";
    when 16#0083B# => romdata <= X"088C0508";
    when 16#0083C# => romdata <= X"80258C38";
    when 16#0083D# => romdata <= X"8C088C05";
    when 16#0083E# => romdata <= X"08308C08";
    when 16#0083F# => romdata <= X"8C050C81";
    when 16#00840# => romdata <= X"538C088C";
    when 16#00841# => romdata <= X"0508528C";
    when 16#00842# => romdata <= X"08880508";
    when 16#00843# => romdata <= X"51AD3F80";
    when 16#00844# => romdata <= X"08708C08";
    when 16#00845# => romdata <= X"F8050C54";
    when 16#00846# => romdata <= X"8C08FC05";
    when 16#00847# => romdata <= X"08802E8C";
    when 16#00848# => romdata <= X"388C08F8";
    when 16#00849# => romdata <= X"0508308C";
    when 16#0084A# => romdata <= X"08F8050C";
    when 16#0084B# => romdata <= X"8C08F805";
    when 16#0084C# => romdata <= X"0870800C";
    when 16#0084D# => romdata <= X"54873D0D";
    when 16#0084E# => romdata <= X"8C0C048C";
    when 16#0084F# => romdata <= X"08028C0C";
    when 16#00850# => romdata <= X"FD3D0D81";
    when 16#00851# => romdata <= X"0B8C08FC";
    when 16#00852# => romdata <= X"050C800B";
    when 16#00853# => romdata <= X"8C08F805";
    when 16#00854# => romdata <= X"0C8C088C";
    when 16#00855# => romdata <= X"05088C08";
    when 16#00856# => romdata <= X"88050827";
    when 16#00857# => romdata <= X"AC388C08";
    when 16#00858# => romdata <= X"FC050880";
    when 16#00859# => romdata <= X"2EA33880";
    when 16#0085A# => romdata <= X"0B8C088C";
    when 16#0085B# => romdata <= X"05082499";
    when 16#0085C# => romdata <= X"388C088C";
    when 16#0085D# => romdata <= X"0508108C";
    when 16#0085E# => romdata <= X"088C050C";
    when 16#0085F# => romdata <= X"8C08FC05";
    when 16#00860# => romdata <= X"08108C08";
    when 16#00861# => romdata <= X"FC050CC9";
    when 16#00862# => romdata <= X"398C08FC";
    when 16#00863# => romdata <= X"0508802E";
    when 16#00864# => romdata <= X"80C9388C";
    when 16#00865# => romdata <= X"088C0508";
    when 16#00866# => romdata <= X"8C088805";
    when 16#00867# => romdata <= X"0826A138";
    when 16#00868# => romdata <= X"8C088805";
    when 16#00869# => romdata <= X"088C088C";
    when 16#0086A# => romdata <= X"0508318C";
    when 16#0086B# => romdata <= X"0888050C";
    when 16#0086C# => romdata <= X"8C08F805";
    when 16#0086D# => romdata <= X"088C08FC";
    when 16#0086E# => romdata <= X"0508078C";
    when 16#0086F# => romdata <= X"08F8050C";
    when 16#00870# => romdata <= X"8C08FC05";
    when 16#00871# => romdata <= X"08812A8C";
    when 16#00872# => romdata <= X"08FC050C";
    when 16#00873# => romdata <= X"8C088C05";
    when 16#00874# => romdata <= X"08812A8C";
    when 16#00875# => romdata <= X"088C050C";
    when 16#00876# => romdata <= X"FFAF398C";
    when 16#00877# => romdata <= X"08900508";
    when 16#00878# => romdata <= X"802E8F38";
    when 16#00879# => romdata <= X"8C088805";
    when 16#0087A# => romdata <= X"08708C08";
    when 16#0087B# => romdata <= X"F4050C51";
    when 16#0087C# => romdata <= X"8D398C08";
    when 16#0087D# => romdata <= X"F8050870";
    when 16#0087E# => romdata <= X"8C08F405";
    when 16#0087F# => romdata <= X"0C518C08";
    when 16#00880# => romdata <= X"F4050880";
    when 16#00881# => romdata <= X"0C853D0D";
    when 16#00882# => romdata <= X"8C0C0480";
    when 16#00883# => romdata <= X"3D0D8651";
    when 16#00884# => romdata <= X"84963F81";
    when 16#00885# => romdata <= X"519F873F";
    when 16#00886# => romdata <= X"FC3D0D76";
    when 16#00887# => romdata <= X"70797B55";
    when 16#00888# => romdata <= X"5555558F";
    when 16#00889# => romdata <= X"72278C38";
    when 16#0088A# => romdata <= X"72750783";
    when 16#0088B# => romdata <= X"06517080";
    when 16#0088C# => romdata <= X"2EA738FF";
    when 16#0088D# => romdata <= X"125271FF";
    when 16#0088E# => romdata <= X"2E983872";
    when 16#0088F# => romdata <= X"70810554";
    when 16#00890# => romdata <= X"33747081";
    when 16#00891# => romdata <= X"055634FF";
    when 16#00892# => romdata <= X"125271FF";
    when 16#00893# => romdata <= X"2E098106";
    when 16#00894# => romdata <= X"EA387480";
    when 16#00895# => romdata <= X"0C863D0D";
    when 16#00896# => romdata <= X"04745172";
    when 16#00897# => romdata <= X"70840554";
    when 16#00898# => romdata <= X"08717084";
    when 16#00899# => romdata <= X"05530C72";
    when 16#0089A# => romdata <= X"70840554";
    when 16#0089B# => romdata <= X"08717084";
    when 16#0089C# => romdata <= X"05530C72";
    when 16#0089D# => romdata <= X"70840554";
    when 16#0089E# => romdata <= X"08717084";
    when 16#0089F# => romdata <= X"05530C72";
    when 16#008A0# => romdata <= X"70840554";
    when 16#008A1# => romdata <= X"08717084";
    when 16#008A2# => romdata <= X"05530CF0";
    when 16#008A3# => romdata <= X"1252718F";
    when 16#008A4# => romdata <= X"26C93883";
    when 16#008A5# => romdata <= X"72279538";
    when 16#008A6# => romdata <= X"72708405";
    when 16#008A7# => romdata <= X"54087170";
    when 16#008A8# => romdata <= X"8405530C";
    when 16#008A9# => romdata <= X"FC125271";
    when 16#008AA# => romdata <= X"8326ED38";
    when 16#008AB# => romdata <= X"7054FF83";
    when 16#008AC# => romdata <= X"39FD3D0D";
    when 16#008AD# => romdata <= X"755384D8";
    when 16#008AE# => romdata <= X"1308802E";
    when 16#008AF# => romdata <= X"8A388053";
    when 16#008B0# => romdata <= X"72800C85";
    when 16#008B1# => romdata <= X"3D0D0481";
    when 16#008B2# => romdata <= X"80527251";
    when 16#008B3# => romdata <= X"8A883F80";
    when 16#008B4# => romdata <= X"0884D814";
    when 16#008B5# => romdata <= X"0CFF5380";
    when 16#008B6# => romdata <= X"08802EE4";
    when 16#008B7# => romdata <= X"38800854";
    when 16#008B8# => romdata <= X"9F538074";
    when 16#008B9# => romdata <= X"70840556";
    when 16#008BA# => romdata <= X"0CFF1353";
    when 16#008BB# => romdata <= X"807324CE";
    when 16#008BC# => romdata <= X"38807470";
    when 16#008BD# => romdata <= X"8405560C";
    when 16#008BE# => romdata <= X"FF135372";
    when 16#008BF# => romdata <= X"8025E338";
    when 16#008C0# => romdata <= X"FFBC39FD";
    when 16#008C1# => romdata <= X"3D0D7577";
    when 16#008C2# => romdata <= X"55539F74";
    when 16#008C3# => romdata <= X"278D3896";
    when 16#008C4# => romdata <= X"730CFF52";
    when 16#008C5# => romdata <= X"71800C85";
    when 16#008C6# => romdata <= X"3D0D0484";
    when 16#008C7# => romdata <= X"D8130852";
    when 16#008C8# => romdata <= X"71802E93";
    when 16#008C9# => romdata <= X"38731010";
    when 16#008CA# => romdata <= X"12700879";
    when 16#008CB# => romdata <= X"720C5152";
    when 16#008CC# => romdata <= X"71800C85";
    when 16#008CD# => romdata <= X"3D0D0472";
    when 16#008CE# => romdata <= X"51FEF63F";
    when 16#008CF# => romdata <= X"FF528008";
    when 16#008D0# => romdata <= X"D33884D8";
    when 16#008D1# => romdata <= X"13087410";
    when 16#008D2# => romdata <= X"10117008";
    when 16#008D3# => romdata <= X"7A720C51";
    when 16#008D4# => romdata <= X"5152DD39";
    when 16#008D5# => romdata <= X"F93D0D79";
    when 16#008D6# => romdata <= X"7B585676";
    when 16#008D7# => romdata <= X"9F2680E8";
    when 16#008D8# => romdata <= X"3884D816";
    when 16#008D9# => romdata <= X"08547380";
    when 16#008DA# => romdata <= X"2EAA3876";
    when 16#008DB# => romdata <= X"10101470";
    when 16#008DC# => romdata <= X"08555573";
    when 16#008DD# => romdata <= X"802EBA38";
    when 16#008DE# => romdata <= X"80587381";
    when 16#008DF# => romdata <= X"2E8F3873";
    when 16#008E0# => romdata <= X"FF2EA338";
    when 16#008E1# => romdata <= X"80750C76";
    when 16#008E2# => romdata <= X"51732D80";
    when 16#008E3# => romdata <= X"5877800C";
    when 16#008E4# => romdata <= X"893D0D04";
    when 16#008E5# => romdata <= X"7551FE99";
    when 16#008E6# => romdata <= X"3FFF5880";
    when 16#008E7# => romdata <= X"08EF3884";
    when 16#008E8# => romdata <= X"D8160854";
    when 16#008E9# => romdata <= X"C6399676";
    when 16#008EA# => romdata <= X"0C810B80";
    when 16#008EB# => romdata <= X"0C893D0D";
    when 16#008EC# => romdata <= X"04755181";
    when 16#008ED# => romdata <= X"ED3F7653";
    when 16#008EE# => romdata <= X"80085275";
    when 16#008EF# => romdata <= X"5181AD3F";
    when 16#008F0# => romdata <= X"8008800C";
    when 16#008F1# => romdata <= X"893D0D04";
    when 16#008F2# => romdata <= X"96760CFF";
    when 16#008F3# => romdata <= X"0B800C89";
    when 16#008F4# => romdata <= X"3D0D04FC";
    when 16#008F5# => romdata <= X"3D0D7678";
    when 16#008F6# => romdata <= X"5653FF54";
    when 16#008F7# => romdata <= X"749F26B1";
    when 16#008F8# => romdata <= X"3884D813";
    when 16#008F9# => romdata <= X"08527180";
    when 16#008FA# => romdata <= X"2EAE3874";
    when 16#008FB# => romdata <= X"10101270";
    when 16#008FC# => romdata <= X"08535381";
    when 16#008FD# => romdata <= X"5471802E";
    when 16#008FE# => romdata <= X"98388254";
    when 16#008FF# => romdata <= X"71FF2E91";
    when 16#00900# => romdata <= X"38835471";
    when 16#00901# => romdata <= X"812E8A38";
    when 16#00902# => romdata <= X"80730C74";
    when 16#00903# => romdata <= X"51712D80";
    when 16#00904# => romdata <= X"5473800C";
    when 16#00905# => romdata <= X"863D0D04";
    when 16#00906# => romdata <= X"7251FD95";
    when 16#00907# => romdata <= X"3F8008F1";
    when 16#00908# => romdata <= X"3884D813";
    when 16#00909# => romdata <= X"0852C439";
    when 16#0090A# => romdata <= X"FF3D0D73";
    when 16#0090B# => romdata <= X"5280F0D8";
    when 16#0090C# => romdata <= X"0851FEA0";
    when 16#0090D# => romdata <= X"3F833D0D";
    when 16#0090E# => romdata <= X"04FE3D0D";
    when 16#0090F# => romdata <= X"75537452";
    when 16#00910# => romdata <= X"80F0D808";
    when 16#00911# => romdata <= X"51FDBC3F";
    when 16#00912# => romdata <= X"843D0D04";
    when 16#00913# => romdata <= X"803D0D80";
    when 16#00914# => romdata <= X"F0D80851";
    when 16#00915# => romdata <= X"FCDB3F82";
    when 16#00916# => romdata <= X"3D0D04FF";
    when 16#00917# => romdata <= X"3D0D7352";
    when 16#00918# => romdata <= X"80F0D808";
    when 16#00919# => romdata <= X"51FEEC3F";
    when 16#0091A# => romdata <= X"833D0D04";
    when 16#0091B# => romdata <= X"FC3D0D80";
    when 16#0091C# => romdata <= X"0B818AE0";
    when 16#0091D# => romdata <= X"0C785277";
    when 16#0091E# => romdata <= X"5199973F";
    when 16#0091F# => romdata <= X"80085480";
    when 16#00920# => romdata <= X"08FF2E88";
    when 16#00921# => romdata <= X"3873800C";
    when 16#00922# => romdata <= X"863D0D04";
    when 16#00923# => romdata <= X"818AE008";
    when 16#00924# => romdata <= X"5574802E";
    when 16#00925# => romdata <= X"F0387675";
    when 16#00926# => romdata <= X"710C5373";
    when 16#00927# => romdata <= X"800C863D";
    when 16#00928# => romdata <= X"0D0498E9";
    when 16#00929# => romdata <= X"3F04FC3D";
    when 16#0092A# => romdata <= X"0D767079";
    when 16#0092B# => romdata <= X"70730783";
    when 16#0092C# => romdata <= X"06545454";
    when 16#0092D# => romdata <= X"557080C3";
    when 16#0092E# => romdata <= X"38717008";
    when 16#0092F# => romdata <= X"700970F7";
    when 16#00930# => romdata <= X"FBFDFF13";
    when 16#00931# => romdata <= X"0670F884";
    when 16#00932# => romdata <= X"82818006";
    when 16#00933# => romdata <= X"51515353";
    when 16#00934# => romdata <= X"5470A638";
    when 16#00935# => romdata <= X"84147274";
    when 16#00936# => romdata <= X"70840556";
    when 16#00937# => romdata <= X"0C700870";
    when 16#00938# => romdata <= X"0970F7FB";
    when 16#00939# => romdata <= X"FDFF1306";
    when 16#0093A# => romdata <= X"70F88482";
    when 16#0093B# => romdata <= X"81800651";
    when 16#0093C# => romdata <= X"51535354";
    when 16#0093D# => romdata <= X"70802EDC";
    when 16#0093E# => romdata <= X"38735271";
    when 16#0093F# => romdata <= X"70810553";
    when 16#00940# => romdata <= X"33517073";
    when 16#00941# => romdata <= X"70810555";
    when 16#00942# => romdata <= X"3470F038";
    when 16#00943# => romdata <= X"74800C86";
    when 16#00944# => romdata <= X"3D0D04FD";
    when 16#00945# => romdata <= X"3D0D7570";
    when 16#00946# => romdata <= X"71830653";
    when 16#00947# => romdata <= X"555270B8";
    when 16#00948# => romdata <= X"38717008";
    when 16#00949# => romdata <= X"7009F7FB";
    when 16#0094A# => romdata <= X"FDFF1206";
    when 16#0094B# => romdata <= X"70F88482";
    when 16#0094C# => romdata <= X"81800651";
    when 16#0094D# => romdata <= X"51525370";
    when 16#0094E# => romdata <= X"9D388413";
    when 16#0094F# => romdata <= X"70087009";
    when 16#00950# => romdata <= X"F7FBFDFF";
    when 16#00951# => romdata <= X"120670F8";
    when 16#00952# => romdata <= X"84828180";
    when 16#00953# => romdata <= X"06515152";
    when 16#00954# => romdata <= X"5370802E";
    when 16#00955# => romdata <= X"E5387252";
    when 16#00956# => romdata <= X"71335170";
    when 16#00957# => romdata <= X"802E8A38";
    when 16#00958# => romdata <= X"81127033";
    when 16#00959# => romdata <= X"525270F8";
    when 16#0095A# => romdata <= X"38717431";
    when 16#0095B# => romdata <= X"800C853D";
    when 16#0095C# => romdata <= X"0D04FA3D";
    when 16#0095D# => romdata <= X"0D787A7C";
    when 16#0095E# => romdata <= X"70545555";
    when 16#0095F# => romdata <= X"5272802E";
    when 16#00960# => romdata <= X"80D93871";
    when 16#00961# => romdata <= X"74078306";
    when 16#00962# => romdata <= X"5170802E";
    when 16#00963# => romdata <= X"80D438FF";
    when 16#00964# => romdata <= X"135372FF";
    when 16#00965# => romdata <= X"2EB13871";
    when 16#00966# => romdata <= X"33743356";
    when 16#00967# => romdata <= X"5174712E";
    when 16#00968# => romdata <= X"098106A9";
    when 16#00969# => romdata <= X"3872802E";
    when 16#0096A# => romdata <= X"81873870";
    when 16#0096B# => romdata <= X"81FF0651";
    when 16#0096C# => romdata <= X"70802E80";
    when 16#0096D# => romdata <= X"FC388112";
    when 16#0096E# => romdata <= X"8115FF15";
    when 16#0096F# => romdata <= X"55555272";
    when 16#00970# => romdata <= X"FF2E0981";
    when 16#00971# => romdata <= X"06D13871";
    when 16#00972# => romdata <= X"33743356";
    when 16#00973# => romdata <= X"517081FF";
    when 16#00974# => romdata <= X"067581FF";
    when 16#00975# => romdata <= X"06717131";
    when 16#00976# => romdata <= X"51525270";
    when 16#00977# => romdata <= X"800C883D";
    when 16#00978# => romdata <= X"0D047174";
    when 16#00979# => romdata <= X"57558373";
    when 16#0097A# => romdata <= X"27883871";
    when 16#0097B# => romdata <= X"0874082E";
    when 16#0097C# => romdata <= X"88387476";
    when 16#0097D# => romdata <= X"5552FF97";
    when 16#0097E# => romdata <= X"39FC1353";
    when 16#0097F# => romdata <= X"72802EB1";
    when 16#00980# => romdata <= X"38740870";
    when 16#00981# => romdata <= X"09F7FBFD";
    when 16#00982# => romdata <= X"FF120670";
    when 16#00983# => romdata <= X"F8848281";
    when 16#00984# => romdata <= X"80065151";
    when 16#00985# => romdata <= X"51709A38";
    when 16#00986# => romdata <= X"84158417";
    when 16#00987# => romdata <= X"57558373";
    when 16#00988# => romdata <= X"27D03874";
    when 16#00989# => romdata <= X"0876082E";
    when 16#0098A# => romdata <= X"D0387476";
    when 16#0098B# => romdata <= X"5552FEDF";
    when 16#0098C# => romdata <= X"39800B80";
    when 16#0098D# => romdata <= X"0C883D0D";
    when 16#0098E# => romdata <= X"04F33D0D";
    when 16#0098F# => romdata <= X"60626472";
    when 16#00990# => romdata <= X"5A5A5D5D";
    when 16#00991# => romdata <= X"805E7670";
    when 16#00992# => romdata <= X"81055833";
    when 16#00993# => romdata <= X"80EE8511";
    when 16#00994# => romdata <= X"3370832A";
    when 16#00995# => romdata <= X"70810651";
    when 16#00996# => romdata <= X"55555672";
    when 16#00997# => romdata <= X"E93875AD";
    when 16#00998# => romdata <= X"2E81FF38";
    when 16#00999# => romdata <= X"75AB2E81";
    when 16#0099A# => romdata <= X"FB387730";
    when 16#0099B# => romdata <= X"70790780";
    when 16#0099C# => romdata <= X"25799032";
    when 16#0099D# => romdata <= X"70307072";
    when 16#0099E# => romdata <= X"07802573";
    when 16#0099F# => romdata <= X"07535757";
    when 16#009A0# => romdata <= X"51537280";
    when 16#009A1# => romdata <= X"2E873875";
    when 16#009A2# => romdata <= X"B02E81E2";
    when 16#009A3# => romdata <= X"38778A38";
    when 16#009A4# => romdata <= X"885875B0";
    when 16#009A5# => romdata <= X"2E83388A";
    when 16#009A6# => romdata <= X"587752FF";
    when 16#009A7# => romdata <= X"51F2A63F";
    when 16#009A8# => romdata <= X"80087853";
    when 16#009A9# => romdata <= X"5AFF51F2";
    when 16#009AA# => romdata <= X"C13F8008";
    when 16#009AB# => romdata <= X"5B80705A";
    when 16#009AC# => romdata <= X"5580EE85";
    when 16#009AD# => romdata <= X"16337082";
    when 16#009AE# => romdata <= X"2A708106";
    when 16#009AF# => romdata <= X"51545472";
    when 16#009B0# => romdata <= X"802E80C1";
    when 16#009B1# => romdata <= X"38D01656";
    when 16#009B2# => romdata <= X"75782580";
    when 16#009B3# => romdata <= X"D7388079";
    when 16#009B4# => romdata <= X"24757B26";
    when 16#009B5# => romdata <= X"07537293";
    when 16#009B6# => romdata <= X"38747A2E";
    when 16#009B7# => romdata <= X"80EB387A";
    when 16#009B8# => romdata <= X"762580ED";
    when 16#009B9# => romdata <= X"3872802E";
    when 16#009BA# => romdata <= X"80E738FF";
    when 16#009BB# => romdata <= X"77708105";
    when 16#009BC# => romdata <= X"59335759";
    when 16#009BD# => romdata <= X"80EE8516";
    when 16#009BE# => romdata <= X"3370822A";
    when 16#009BF# => romdata <= X"70810651";
    when 16#009C0# => romdata <= X"545472C1";
    when 16#009C1# => romdata <= X"38738306";
    when 16#009C2# => romdata <= X"5372802E";
    when 16#009C3# => romdata <= X"97387381";
    when 16#009C4# => romdata <= X"06C91755";
    when 16#009C5# => romdata <= X"53728538";
    when 16#009C6# => romdata <= X"FFA91654";
    when 16#009C7# => romdata <= X"73567776";
    when 16#009C8# => romdata <= X"24FFAB38";
    when 16#009C9# => romdata <= X"80792481";
    when 16#009CA# => romdata <= X"89387D80";
    when 16#009CB# => romdata <= X"2E843874";
    when 16#009CC# => romdata <= X"30557B80";
    when 16#009CD# => romdata <= X"2E8C38FF";
    when 16#009CE# => romdata <= X"17537883";
    when 16#009CF# => romdata <= X"387C5372";
    when 16#009D0# => romdata <= X"7C0C7480";
    when 16#009D1# => romdata <= X"0C8F3D0D";
    when 16#009D2# => romdata <= X"04815375";
    when 16#009D3# => romdata <= X"7B24FF95";
    when 16#009D4# => romdata <= X"38817579";
    when 16#009D5# => romdata <= X"29177870";
    when 16#009D6# => romdata <= X"81055A33";
    when 16#009D7# => romdata <= X"585659FF";
    when 16#009D8# => romdata <= X"9339815E";
    when 16#009D9# => romdata <= X"76708105";
    when 16#009DA# => romdata <= X"583356FD";
    when 16#009DB# => romdata <= X"FD398077";
    when 16#009DC# => romdata <= X"33545472";
    when 16#009DD# => romdata <= X"80F82E80";
    when 16#009DE# => romdata <= X"C3387280";
    when 16#009DF# => romdata <= X"D8327030";
    when 16#009E0# => romdata <= X"70802576";
    when 16#009E1# => romdata <= X"07515153";
    when 16#009E2# => romdata <= X"72802EFE";
    when 16#009E3# => romdata <= X"80388117";
    when 16#009E4# => romdata <= X"33821858";
    when 16#009E5# => romdata <= X"56907053";
    when 16#009E6# => romdata <= X"58FF51F0";
    when 16#009E7# => romdata <= X"A83F8008";
    when 16#009E8# => romdata <= X"78535AFF";
    when 16#009E9# => romdata <= X"51F0C33F";
    when 16#009EA# => romdata <= X"80085B80";
    when 16#009EB# => romdata <= X"705A55FE";
    when 16#009EC# => romdata <= X"8039FF60";
    when 16#009ED# => romdata <= X"5455A273";
    when 16#009EE# => romdata <= X"0CFEF739";
    when 16#009EF# => romdata <= X"8154FFBA";
    when 16#009F0# => romdata <= X"39FD3D0D";
    when 16#009F1# => romdata <= X"77547653";
    when 16#009F2# => romdata <= X"755280F0";
    when 16#009F3# => romdata <= X"D80851FC";
    when 16#009F4# => romdata <= X"E83F853D";
    when 16#009F5# => romdata <= X"0D04F33D";
    when 16#009F6# => romdata <= X"0D7F618B";
    when 16#009F7# => romdata <= X"1170F806";
    when 16#009F8# => romdata <= X"5C55555E";
    when 16#009F9# => romdata <= X"72962683";
    when 16#009FA# => romdata <= X"38905980";
    when 16#009FB# => romdata <= X"7924747A";
    when 16#009FC# => romdata <= X"26075380";
    when 16#009FD# => romdata <= X"5472742E";
    when 16#009FE# => romdata <= X"09810680";
    when 16#009FF# => romdata <= X"CB387D51";
    when 16#00A00# => romdata <= X"8BCA3F78";
    when 16#00A01# => romdata <= X"83F72680";
    when 16#00A02# => romdata <= X"C6387883";
    when 16#00A03# => romdata <= X"2A701010";
    when 16#00A04# => romdata <= X"1080F894";
    when 16#00A05# => romdata <= X"058C1108";
    when 16#00A06# => romdata <= X"59595A76";
    when 16#00A07# => romdata <= X"782E83B0";
    when 16#00A08# => romdata <= X"38841708";
    when 16#00A09# => romdata <= X"FC06568C";
    when 16#00A0A# => romdata <= X"17088818";
    when 16#00A0B# => romdata <= X"08718C12";
    when 16#00A0C# => romdata <= X"0C88120C";
    when 16#00A0D# => romdata <= X"58751784";
    when 16#00A0E# => romdata <= X"11088107";
    when 16#00A0F# => romdata <= X"84120C53";
    when 16#00A10# => romdata <= X"7D518B89";
    when 16#00A11# => romdata <= X"3F881754";
    when 16#00A12# => romdata <= X"73800C8F";
    when 16#00A13# => romdata <= X"3D0D0478";
    when 16#00A14# => romdata <= X"892A7983";
    when 16#00A15# => romdata <= X"2A5B5372";
    when 16#00A16# => romdata <= X"802EBF38";
    when 16#00A17# => romdata <= X"78862AB8";
    when 16#00A18# => romdata <= X"055A8473";
    when 16#00A19# => romdata <= X"27B43880";
    when 16#00A1A# => romdata <= X"DB135A94";
    when 16#00A1B# => romdata <= X"7327AB38";
    when 16#00A1C# => romdata <= X"788C2A80";
    when 16#00A1D# => romdata <= X"EE055A80";
    when 16#00A1E# => romdata <= X"D473279E";
    when 16#00A1F# => romdata <= X"38788F2A";
    when 16#00A20# => romdata <= X"80F7055A";
    when 16#00A21# => romdata <= X"82D47327";
    when 16#00A22# => romdata <= X"91387892";
    when 16#00A23# => romdata <= X"2A80FC05";
    when 16#00A24# => romdata <= X"5A8AD473";
    when 16#00A25# => romdata <= X"27843880";
    when 16#00A26# => romdata <= X"FE5A7910";
    when 16#00A27# => romdata <= X"101080F8";
    when 16#00A28# => romdata <= X"94058C11";
    when 16#00A29# => romdata <= X"08585576";
    when 16#00A2A# => romdata <= X"752EA338";
    when 16#00A2B# => romdata <= X"841708FC";
    when 16#00A2C# => romdata <= X"06707A31";
    when 16#00A2D# => romdata <= X"5556738F";
    when 16#00A2E# => romdata <= X"2488D538";
    when 16#00A2F# => romdata <= X"738025FE";
    when 16#00A30# => romdata <= X"E6388C17";
    when 16#00A31# => romdata <= X"08577675";
    when 16#00A32# => romdata <= X"2E098106";
    when 16#00A33# => romdata <= X"DF38811A";
    when 16#00A34# => romdata <= X"5A80F8A4";
    when 16#00A35# => romdata <= X"08577680";
    when 16#00A36# => romdata <= X"F89C2E82";
    when 16#00A37# => romdata <= X"C0388417";
    when 16#00A38# => romdata <= X"08FC0670";
    when 16#00A39# => romdata <= X"7A315556";
    when 16#00A3A# => romdata <= X"738F2481";
    when 16#00A3B# => romdata <= X"F93880F8";
    when 16#00A3C# => romdata <= X"9C0B80F8";
    when 16#00A3D# => romdata <= X"A80C80F8";
    when 16#00A3E# => romdata <= X"9C0B80F8";
    when 16#00A3F# => romdata <= X"A40C7380";
    when 16#00A40# => romdata <= X"25FEB238";
    when 16#00A41# => romdata <= X"83FF7627";
    when 16#00A42# => romdata <= X"83DF3875";
    when 16#00A43# => romdata <= X"892A7683";
    when 16#00A44# => romdata <= X"2A555372";
    when 16#00A45# => romdata <= X"802EBF38";
    when 16#00A46# => romdata <= X"75862AB8";
    when 16#00A47# => romdata <= X"05548473";
    when 16#00A48# => romdata <= X"27B43880";
    when 16#00A49# => romdata <= X"DB135494";
    when 16#00A4A# => romdata <= X"7327AB38";
    when 16#00A4B# => romdata <= X"758C2A80";
    when 16#00A4C# => romdata <= X"EE055480";
    when 16#00A4D# => romdata <= X"D473279E";
    when 16#00A4E# => romdata <= X"38758F2A";
    when 16#00A4F# => romdata <= X"80F70554";
    when 16#00A50# => romdata <= X"82D47327";
    when 16#00A51# => romdata <= X"91387592";
    when 16#00A52# => romdata <= X"2A80FC05";
    when 16#00A53# => romdata <= X"548AD473";
    when 16#00A54# => romdata <= X"27843880";
    when 16#00A55# => romdata <= X"FE547310";
    when 16#00A56# => romdata <= X"101080F8";
    when 16#00A57# => romdata <= X"94058811";
    when 16#00A58# => romdata <= X"08565874";
    when 16#00A59# => romdata <= X"782E86CF";
    when 16#00A5A# => romdata <= X"38841508";
    when 16#00A5B# => romdata <= X"FC065375";
    when 16#00A5C# => romdata <= X"73278D38";
    when 16#00A5D# => romdata <= X"88150855";
    when 16#00A5E# => romdata <= X"74782E09";
    when 16#00A5F# => romdata <= X"8106EA38";
    when 16#00A60# => romdata <= X"8C150880";
    when 16#00A61# => romdata <= X"F8940B84";
    when 16#00A62# => romdata <= X"0508718C";
    when 16#00A63# => romdata <= X"1A0C7688";
    when 16#00A64# => romdata <= X"1A0C7888";
    when 16#00A65# => romdata <= X"130C788C";
    when 16#00A66# => romdata <= X"180C5D58";
    when 16#00A67# => romdata <= X"7953807A";
    when 16#00A68# => romdata <= X"2483E638";
    when 16#00A69# => romdata <= X"72822C81";
    when 16#00A6A# => romdata <= X"712B5C53";
    when 16#00A6B# => romdata <= X"7A7C2681";
    when 16#00A6C# => romdata <= X"98387B7B";
    when 16#00A6D# => romdata <= X"06537282";
    when 16#00A6E# => romdata <= X"F13879FC";
    when 16#00A6F# => romdata <= X"0684055A";
    when 16#00A70# => romdata <= X"7A10707D";
    when 16#00A71# => romdata <= X"06545B72";
    when 16#00A72# => romdata <= X"82E03884";
    when 16#00A73# => romdata <= X"1A5AF139";
    when 16#00A74# => romdata <= X"88178C11";
    when 16#00A75# => romdata <= X"08585876";
    when 16#00A76# => romdata <= X"782E0981";
    when 16#00A77# => romdata <= X"06FCC238";
    when 16#00A78# => romdata <= X"821A5AFD";
    when 16#00A79# => romdata <= X"EC397817";
    when 16#00A7A# => romdata <= X"79810784";
    when 16#00A7B# => romdata <= X"190C7080";
    when 16#00A7C# => romdata <= X"F8A80C70";
    when 16#00A7D# => romdata <= X"80F8A40C";
    when 16#00A7E# => romdata <= X"80F89C0B";
    when 16#00A7F# => romdata <= X"8C120C8C";
    when 16#00A80# => romdata <= X"11088812";
    when 16#00A81# => romdata <= X"0C748107";
    when 16#00A82# => romdata <= X"84120C74";
    when 16#00A83# => romdata <= X"1175710C";
    when 16#00A84# => romdata <= X"51537D51";
    when 16#00A85# => romdata <= X"87B73F88";
    when 16#00A86# => romdata <= X"1754FCAC";
    when 16#00A87# => romdata <= X"3980F894";
    when 16#00A88# => romdata <= X"0B840508";
    when 16#00A89# => romdata <= X"7A545C79";
    when 16#00A8A# => romdata <= X"8025FEF8";
    when 16#00A8B# => romdata <= X"3882DA39";
    when 16#00A8C# => romdata <= X"7A097C06";
    when 16#00A8D# => romdata <= X"7080F894";
    when 16#00A8E# => romdata <= X"0B84050C";
    when 16#00A8F# => romdata <= X"5C7A105B";
    when 16#00A90# => romdata <= X"7A7C2685";
    when 16#00A91# => romdata <= X"387A85B8";
    when 16#00A92# => romdata <= X"3880F894";
    when 16#00A93# => romdata <= X"0B880508";
    when 16#00A94# => romdata <= X"70841208";
    when 16#00A95# => romdata <= X"FC06707C";
    when 16#00A96# => romdata <= X"317C7226";
    when 16#00A97# => romdata <= X"8F722507";
    when 16#00A98# => romdata <= X"57575C5D";
    when 16#00A99# => romdata <= X"5572802E";
    when 16#00A9A# => romdata <= X"80DB3879";
    when 16#00A9B# => romdata <= X"7A1680F8";
    when 16#00A9C# => romdata <= X"8C081B90";
    when 16#00A9D# => romdata <= X"115A5557";
    when 16#00A9E# => romdata <= X"5B80F888";
    when 16#00A9F# => romdata <= X"08FF2E88";
    when 16#00AA0# => romdata <= X"38A08F13";
    when 16#00AA1# => romdata <= X"E0800657";
    when 16#00AA2# => romdata <= X"76527D51";
    when 16#00AA3# => romdata <= X"86C03F80";
    when 16#00AA4# => romdata <= X"08548008";
    when 16#00AA5# => romdata <= X"FF2E9038";
    when 16#00AA6# => romdata <= X"80087627";
    when 16#00AA7# => romdata <= X"82993874";
    when 16#00AA8# => romdata <= X"80F8942E";
    when 16#00AA9# => romdata <= X"82913880";
    when 16#00AAA# => romdata <= X"F8940B88";
    when 16#00AAB# => romdata <= X"05085584";
    when 16#00AAC# => romdata <= X"1508FC06";
    when 16#00AAD# => romdata <= X"707A317A";
    when 16#00AAE# => romdata <= X"72268F72";
    when 16#00AAF# => romdata <= X"25075255";
    when 16#00AB0# => romdata <= X"537283E6";
    when 16#00AB1# => romdata <= X"38747981";
    when 16#00AB2# => romdata <= X"0784170C";
    when 16#00AB3# => romdata <= X"79167080";
    when 16#00AB4# => romdata <= X"F8940B88";
    when 16#00AB5# => romdata <= X"050C7581";
    when 16#00AB6# => romdata <= X"0784120C";
    when 16#00AB7# => romdata <= X"547E5257";
    when 16#00AB8# => romdata <= X"85EB3F88";
    when 16#00AB9# => romdata <= X"1754FAE0";
    when 16#00ABA# => romdata <= X"3975832A";
    when 16#00ABB# => romdata <= X"70545480";
    when 16#00ABC# => romdata <= X"7424819B";
    when 16#00ABD# => romdata <= X"3872822C";
    when 16#00ABE# => romdata <= X"81712B80";
    when 16#00ABF# => romdata <= X"F8980807";
    when 16#00AC0# => romdata <= X"7080F894";
    when 16#00AC1# => romdata <= X"0B84050C";
    when 16#00AC2# => romdata <= X"75101010";
    when 16#00AC3# => romdata <= X"80F89405";
    when 16#00AC4# => romdata <= X"88110858";
    when 16#00AC5# => romdata <= X"5A5D5377";
    when 16#00AC6# => romdata <= X"8C180C74";
    when 16#00AC7# => romdata <= X"88180C76";
    when 16#00AC8# => romdata <= X"88190C76";
    when 16#00AC9# => romdata <= X"8C160CFC";
    when 16#00ACA# => romdata <= X"F339797A";
    when 16#00ACB# => romdata <= X"10101080";
    when 16#00ACC# => romdata <= X"F8940570";
    when 16#00ACD# => romdata <= X"57595D8C";
    when 16#00ACE# => romdata <= X"15085776";
    when 16#00ACF# => romdata <= X"752EA338";
    when 16#00AD0# => romdata <= X"841708FC";
    when 16#00AD1# => romdata <= X"06707A31";
    when 16#00AD2# => romdata <= X"5556738F";
    when 16#00AD3# => romdata <= X"2483CA38";
    when 16#00AD4# => romdata <= X"73802584";
    when 16#00AD5# => romdata <= X"81388C17";
    when 16#00AD6# => romdata <= X"08577675";
    when 16#00AD7# => romdata <= X"2E098106";
    when 16#00AD8# => romdata <= X"DF388815";
    when 16#00AD9# => romdata <= X"811B7083";
    when 16#00ADA# => romdata <= X"06555B55";
    when 16#00ADB# => romdata <= X"72C9387C";
    when 16#00ADC# => romdata <= X"83065372";
    when 16#00ADD# => romdata <= X"802EFDB8";
    when 16#00ADE# => romdata <= X"38FF1DF8";
    when 16#00ADF# => romdata <= X"19595D88";
    when 16#00AE0# => romdata <= X"1808782E";
    when 16#00AE1# => romdata <= X"EA38FDB5";
    when 16#00AE2# => romdata <= X"39831A53";
    when 16#00AE3# => romdata <= X"FC963983";
    when 16#00AE4# => romdata <= X"1470822C";
    when 16#00AE5# => romdata <= X"81712B80";
    when 16#00AE6# => romdata <= X"F8980807";
    when 16#00AE7# => romdata <= X"7080F894";
    when 16#00AE8# => romdata <= X"0B84050C";
    when 16#00AE9# => romdata <= X"76101010";
    when 16#00AEA# => romdata <= X"80F89405";
    when 16#00AEB# => romdata <= X"88110859";
    when 16#00AEC# => romdata <= X"5B5E5153";
    when 16#00AED# => romdata <= X"FEE13980";
    when 16#00AEE# => romdata <= X"F7D80817";
    when 16#00AEF# => romdata <= X"58800876";
    when 16#00AF0# => romdata <= X"2E818D38";
    when 16#00AF1# => romdata <= X"80F88808";
    when 16#00AF2# => romdata <= X"FF2E83EC";
    when 16#00AF3# => romdata <= X"38737631";
    when 16#00AF4# => romdata <= X"1880F7D8";
    when 16#00AF5# => romdata <= X"0C738706";
    when 16#00AF6# => romdata <= X"70575372";
    when 16#00AF7# => romdata <= X"802E8838";
    when 16#00AF8# => romdata <= X"88733170";
    when 16#00AF9# => romdata <= X"15555676";
    when 16#00AFA# => romdata <= X"149FFF06";
    when 16#00AFB# => romdata <= X"A0807131";
    when 16#00AFC# => romdata <= X"1770547F";
    when 16#00AFD# => romdata <= X"53575383";
    when 16#00AFE# => romdata <= X"D53F8008";
    when 16#00AFF# => romdata <= X"538008FF";
    when 16#00B00# => romdata <= X"2E81A038";
    when 16#00B01# => romdata <= X"80F7D808";
    when 16#00B02# => romdata <= X"167080F7";
    when 16#00B03# => romdata <= X"D80C7475";
    when 16#00B04# => romdata <= X"80F8940B";
    when 16#00B05# => romdata <= X"88050C74";
    when 16#00B06# => romdata <= X"76311870";
    when 16#00B07# => romdata <= X"81075155";
    when 16#00B08# => romdata <= X"56587B80";
    when 16#00B09# => romdata <= X"F8942E83";
    when 16#00B0A# => romdata <= X"9C38798F";
    when 16#00B0B# => romdata <= X"2682CB38";
    when 16#00B0C# => romdata <= X"810B8415";
    when 16#00B0D# => romdata <= X"0C841508";
    when 16#00B0E# => romdata <= X"FC06707A";
    when 16#00B0F# => romdata <= X"317A7226";
    when 16#00B10# => romdata <= X"8F722507";
    when 16#00B11# => romdata <= X"52555372";
    when 16#00B12# => romdata <= X"802EFCF9";
    when 16#00B13# => romdata <= X"3880DB39";
    when 16#00B14# => romdata <= X"80089FFF";
    when 16#00B15# => romdata <= X"065372FE";
    when 16#00B16# => romdata <= X"EB387780";
    when 16#00B17# => romdata <= X"F7D80C80";
    when 16#00B18# => romdata <= X"F8940B88";
    when 16#00B19# => romdata <= X"05087B18";
    when 16#00B1A# => romdata <= X"81078412";
    when 16#00B1B# => romdata <= X"0C5580F8";
    when 16#00B1C# => romdata <= X"84087827";
    when 16#00B1D# => romdata <= X"86387780";
    when 16#00B1E# => romdata <= X"F8840C80";
    when 16#00B1F# => romdata <= X"F8800878";
    when 16#00B20# => romdata <= X"27FCAC38";
    when 16#00B21# => romdata <= X"7780F880";
    when 16#00B22# => romdata <= X"0C841508";
    when 16#00B23# => romdata <= X"FC06707A";
    when 16#00B24# => romdata <= X"317A7226";
    when 16#00B25# => romdata <= X"8F722507";
    when 16#00B26# => romdata <= X"52555372";
    when 16#00B27# => romdata <= X"802EFCA5";
    when 16#00B28# => romdata <= X"38883980";
    when 16#00B29# => romdata <= X"745456FE";
    when 16#00B2A# => romdata <= X"DB397D51";
    when 16#00B2B# => romdata <= X"829F3F80";
    when 16#00B2C# => romdata <= X"0B800C8F";
    when 16#00B2D# => romdata <= X"3D0D0473";
    when 16#00B2E# => romdata <= X"53807424";
    when 16#00B2F# => romdata <= X"A9387282";
    when 16#00B30# => romdata <= X"2C81712B";
    when 16#00B31# => romdata <= X"80F89808";
    when 16#00B32# => romdata <= X"077080F8";
    when 16#00B33# => romdata <= X"940B8405";
    when 16#00B34# => romdata <= X"0C5D5377";
    when 16#00B35# => romdata <= X"8C180C74";
    when 16#00B36# => romdata <= X"88180C76";
    when 16#00B37# => romdata <= X"88190C76";
    when 16#00B38# => romdata <= X"8C160CF9";
    when 16#00B39# => romdata <= X"B7398314";
    when 16#00B3A# => romdata <= X"70822C81";
    when 16#00B3B# => romdata <= X"712B80F8";
    when 16#00B3C# => romdata <= X"98080770";
    when 16#00B3D# => romdata <= X"80F8940B";
    when 16#00B3E# => romdata <= X"84050C5E";
    when 16#00B3F# => romdata <= X"5153D439";
    when 16#00B40# => romdata <= X"7B7B0653";
    when 16#00B41# => romdata <= X"72FCA338";
    when 16#00B42# => romdata <= X"841A7B10";
    when 16#00B43# => romdata <= X"5C5AF139";
    when 16#00B44# => romdata <= X"FF1A8111";
    when 16#00B45# => romdata <= X"515AF7B9";
    when 16#00B46# => romdata <= X"39781779";
    when 16#00B47# => romdata <= X"81078419";
    when 16#00B48# => romdata <= X"0C8C1808";
    when 16#00B49# => romdata <= X"88190871";
    when 16#00B4A# => romdata <= X"8C120C88";
    when 16#00B4B# => romdata <= X"120C5970";
    when 16#00B4C# => romdata <= X"80F8A80C";
    when 16#00B4D# => romdata <= X"7080F8A4";
    when 16#00B4E# => romdata <= X"0C80F89C";
    when 16#00B4F# => romdata <= X"0B8C120C";
    when 16#00B50# => romdata <= X"8C110888";
    when 16#00B51# => romdata <= X"120C7481";
    when 16#00B52# => romdata <= X"0784120C";
    when 16#00B53# => romdata <= X"74117571";
    when 16#00B54# => romdata <= X"0C5153F9";
    when 16#00B55# => romdata <= X"BD397517";
    when 16#00B56# => romdata <= X"84110881";
    when 16#00B57# => romdata <= X"0784120C";
    when 16#00B58# => romdata <= X"538C1708";
    when 16#00B59# => romdata <= X"88180871";
    when 16#00B5A# => romdata <= X"8C120C88";
    when 16#00B5B# => romdata <= X"120C587D";
    when 16#00B5C# => romdata <= X"5180DA3F";
    when 16#00B5D# => romdata <= X"881754F5";
    when 16#00B5E# => romdata <= X"CF397284";
    when 16#00B5F# => romdata <= X"150CF41A";
    when 16#00B60# => romdata <= X"F8067084";
    when 16#00B61# => romdata <= X"1E088106";
    when 16#00B62# => romdata <= X"07841E0C";
    when 16#00B63# => romdata <= X"701D545B";
    when 16#00B64# => romdata <= X"850B8414";
    when 16#00B65# => romdata <= X"0C850B88";
    when 16#00B66# => romdata <= X"140C8F7B";
    when 16#00B67# => romdata <= X"27FDCF38";
    when 16#00B68# => romdata <= X"881C527D";
    when 16#00B69# => romdata <= X"5182903F";
    when 16#00B6A# => romdata <= X"80F8940B";
    when 16#00B6B# => romdata <= X"88050880";
    when 16#00B6C# => romdata <= X"F7D80859";
    when 16#00B6D# => romdata <= X"55FDB739";
    when 16#00B6E# => romdata <= X"7780F7D8";
    when 16#00B6F# => romdata <= X"0C7380F8";
    when 16#00B70# => romdata <= X"880CFC91";
    when 16#00B71# => romdata <= X"39728415";
    when 16#00B72# => romdata <= X"0CFDA339";
    when 16#00B73# => romdata <= X"0404FD3D";
    when 16#00B74# => romdata <= X"0D800B81";
    when 16#00B75# => romdata <= X"8AE00C76";
    when 16#00B76# => romdata <= X"5186CC3F";
    when 16#00B77# => romdata <= X"80085380";
    when 16#00B78# => romdata <= X"08FF2E88";
    when 16#00B79# => romdata <= X"3872800C";
    when 16#00B7A# => romdata <= X"853D0D04";
    when 16#00B7B# => romdata <= X"818AE008";
    when 16#00B7C# => romdata <= X"5473802E";
    when 16#00B7D# => romdata <= X"F0387574";
    when 16#00B7E# => romdata <= X"710C5272";
    when 16#00B7F# => romdata <= X"800C853D";
    when 16#00B80# => romdata <= X"0D04FB3D";
    when 16#00B81# => romdata <= X"0D777052";
    when 16#00B82# => romdata <= X"56C23F80";
    when 16#00B83# => romdata <= X"F8940B88";
    when 16#00B84# => romdata <= X"05088411";
    when 16#00B85# => romdata <= X"08FC0670";
    when 16#00B86# => romdata <= X"7B319FEF";
    when 16#00B87# => romdata <= X"05E08006";
    when 16#00B88# => romdata <= X"E0800556";
    when 16#00B89# => romdata <= X"5653A080";
    when 16#00B8A# => romdata <= X"74249438";
    when 16#00B8B# => romdata <= X"80527551";
    when 16#00B8C# => romdata <= X"FF9C3F80";
    when 16#00B8D# => romdata <= X"F89C0815";
    when 16#00B8E# => romdata <= X"53728008";
    when 16#00B8F# => romdata <= X"2E8F3875";
    when 16#00B90# => romdata <= X"51FF8A3F";
    when 16#00B91# => romdata <= X"80537280";
    when 16#00B92# => romdata <= X"0C873D0D";
    when 16#00B93# => romdata <= X"04733052";
    when 16#00B94# => romdata <= X"7551FEFA";
    when 16#00B95# => romdata <= X"3F8008FF";
    when 16#00B96# => romdata <= X"2EA83880";
    when 16#00B97# => romdata <= X"F8940B88";
    when 16#00B98# => romdata <= X"05087575";
    when 16#00B99# => romdata <= X"31810784";
    when 16#00B9A# => romdata <= X"120C5380";
    when 16#00B9B# => romdata <= X"F7D80874";
    when 16#00B9C# => romdata <= X"3180F7D8";
    when 16#00B9D# => romdata <= X"0C7551FE";
    when 16#00B9E# => romdata <= X"D43F810B";
    when 16#00B9F# => romdata <= X"800C873D";
    when 16#00BA0# => romdata <= X"0D048052";
    when 16#00BA1# => romdata <= X"7551FEC6";
    when 16#00BA2# => romdata <= X"3F80F894";
    when 16#00BA3# => romdata <= X"0B880508";
    when 16#00BA4# => romdata <= X"80087131";
    when 16#00BA5# => romdata <= X"56538F75";
    when 16#00BA6# => romdata <= X"25FFA438";
    when 16#00BA7# => romdata <= X"800880F8";
    when 16#00BA8# => romdata <= X"88083180";
    when 16#00BA9# => romdata <= X"F7D80C74";
    when 16#00BAA# => romdata <= X"81078414";
    when 16#00BAB# => romdata <= X"0C7551FE";
    when 16#00BAC# => romdata <= X"9C3F8053";
    when 16#00BAD# => romdata <= X"FF9039F6";
    when 16#00BAE# => romdata <= X"3D0D7C7E";
    when 16#00BAF# => romdata <= X"545B7280";
    when 16#00BB0# => romdata <= X"2E828338";
    when 16#00BB1# => romdata <= X"7A51FE84";
    when 16#00BB2# => romdata <= X"3FF81384";
    when 16#00BB3# => romdata <= X"110870FE";
    when 16#00BB4# => romdata <= X"06701384";
    when 16#00BB5# => romdata <= X"1108FC06";
    when 16#00BB6# => romdata <= X"5D585954";
    when 16#00BB7# => romdata <= X"5880F89C";
    when 16#00BB8# => romdata <= X"08752E82";
    when 16#00BB9# => romdata <= X"DE387884";
    when 16#00BBA# => romdata <= X"160C8073";
    when 16#00BBB# => romdata <= X"8106545A";
    when 16#00BBC# => romdata <= X"727A2E81";
    when 16#00BBD# => romdata <= X"D5387815";
    when 16#00BBE# => romdata <= X"84110881";
    when 16#00BBF# => romdata <= X"06515372";
    when 16#00BC0# => romdata <= X"A0387817";
    when 16#00BC1# => romdata <= X"577981E6";
    when 16#00BC2# => romdata <= X"38881508";
    when 16#00BC3# => romdata <= X"537280F8";
    when 16#00BC4# => romdata <= X"9C2E82F9";
    when 16#00BC5# => romdata <= X"388C1508";
    when 16#00BC6# => romdata <= X"708C150C";
    when 16#00BC7# => romdata <= X"7388120C";
    when 16#00BC8# => romdata <= X"56768107";
    when 16#00BC9# => romdata <= X"84190C76";
    when 16#00BCA# => romdata <= X"1877710C";
    when 16#00BCB# => romdata <= X"53798191";
    when 16#00BCC# => romdata <= X"3883FF77";
    when 16#00BCD# => romdata <= X"2781C838";
    when 16#00BCE# => romdata <= X"76892A77";
    when 16#00BCF# => romdata <= X"832A5653";
    when 16#00BD0# => romdata <= X"72802EBF";
    when 16#00BD1# => romdata <= X"3876862A";
    when 16#00BD2# => romdata <= X"B8055584";
    when 16#00BD3# => romdata <= X"7327B438";
    when 16#00BD4# => romdata <= X"80DB1355";
    when 16#00BD5# => romdata <= X"947327AB";
    when 16#00BD6# => romdata <= X"38768C2A";
    when 16#00BD7# => romdata <= X"80EE0555";
    when 16#00BD8# => romdata <= X"80D47327";
    when 16#00BD9# => romdata <= X"9E38768F";
    when 16#00BDA# => romdata <= X"2A80F705";
    when 16#00BDB# => romdata <= X"5582D473";
    when 16#00BDC# => romdata <= X"27913876";
    when 16#00BDD# => romdata <= X"922A80FC";
    when 16#00BDE# => romdata <= X"05558AD4";
    when 16#00BDF# => romdata <= X"73278438";
    when 16#00BE0# => romdata <= X"80FE5574";
    when 16#00BE1# => romdata <= X"10101080";
    when 16#00BE2# => romdata <= X"F8940588";
    when 16#00BE3# => romdata <= X"11085556";
    when 16#00BE4# => romdata <= X"73762E82";
    when 16#00BE5# => romdata <= X"B3388414";
    when 16#00BE6# => romdata <= X"08FC0653";
    when 16#00BE7# => romdata <= X"7673278D";
    when 16#00BE8# => romdata <= X"38881408";
    when 16#00BE9# => romdata <= X"5473762E";
    when 16#00BEA# => romdata <= X"098106EA";
    when 16#00BEB# => romdata <= X"388C1408";
    when 16#00BEC# => romdata <= X"708C1A0C";
    when 16#00BED# => romdata <= X"74881A0C";
    when 16#00BEE# => romdata <= X"7888120C";
    when 16#00BEF# => romdata <= X"56778C15";
    when 16#00BF0# => romdata <= X"0C7A51FC";
    when 16#00BF1# => romdata <= X"883F8C3D";
    when 16#00BF2# => romdata <= X"0D047708";
    when 16#00BF3# => romdata <= X"78713159";
    when 16#00BF4# => romdata <= X"77058819";
    when 16#00BF5# => romdata <= X"08545772";
    when 16#00BF6# => romdata <= X"80F89C2E";
    when 16#00BF7# => romdata <= X"80E0388C";
    when 16#00BF8# => romdata <= X"1808708C";
    when 16#00BF9# => romdata <= X"150C7388";
    when 16#00BFA# => romdata <= X"120C56FE";
    when 16#00BFB# => romdata <= X"89398815";
    when 16#00BFC# => romdata <= X"088C1608";
    when 16#00BFD# => romdata <= X"708C130C";
    when 16#00BFE# => romdata <= X"5788170C";
    when 16#00BFF# => romdata <= X"FEA33976";
    when 16#00C00# => romdata <= X"832A7054";
    when 16#00C01# => romdata <= X"55807524";
    when 16#00C02# => romdata <= X"81983872";
    when 16#00C03# => romdata <= X"822C8171";
    when 16#00C04# => romdata <= X"2B80F898";
    when 16#00C05# => romdata <= X"080780F8";
    when 16#00C06# => romdata <= X"940B8405";
    when 16#00C07# => romdata <= X"0C537410";
    when 16#00C08# => romdata <= X"101080F8";
    when 16#00C09# => romdata <= X"94058811";
    when 16#00C0A# => romdata <= X"08555675";
    when 16#00C0B# => romdata <= X"8C190C73";
    when 16#00C0C# => romdata <= X"88190C77";
    when 16#00C0D# => romdata <= X"88170C77";
    when 16#00C0E# => romdata <= X"8C150CFF";
    when 16#00C0F# => romdata <= X"8439815A";
    when 16#00C10# => romdata <= X"FDB43978";
    when 16#00C11# => romdata <= X"17738106";
    when 16#00C12# => romdata <= X"54577298";
    when 16#00C13# => romdata <= X"38770878";
    when 16#00C14# => romdata <= X"71315977";
    when 16#00C15# => romdata <= X"058C1908";
    when 16#00C16# => romdata <= X"881A0871";
    when 16#00C17# => romdata <= X"8C120C88";
    when 16#00C18# => romdata <= X"120C5757";
    when 16#00C19# => romdata <= X"76810784";
    when 16#00C1A# => romdata <= X"190C7780";
    when 16#00C1B# => romdata <= X"F8940B88";
    when 16#00C1C# => romdata <= X"050C80F8";
    when 16#00C1D# => romdata <= X"90087726";
    when 16#00C1E# => romdata <= X"FEC73880";
    when 16#00C1F# => romdata <= X"F88C0852";
    when 16#00C20# => romdata <= X"7A51FAFE";
    when 16#00C21# => romdata <= X"3F7A51FA";
    when 16#00C22# => romdata <= X"C43FFEBA";
    when 16#00C23# => romdata <= X"3981788C";
    when 16#00C24# => romdata <= X"150C7888";
    when 16#00C25# => romdata <= X"150C738C";
    when 16#00C26# => romdata <= X"1A0C7388";
    when 16#00C27# => romdata <= X"1A0C5AFD";
    when 16#00C28# => romdata <= X"80398315";
    when 16#00C29# => romdata <= X"70822C81";
    when 16#00C2A# => romdata <= X"712B80F8";
    when 16#00C2B# => romdata <= X"98080780";
    when 16#00C2C# => romdata <= X"F8940B84";
    when 16#00C2D# => romdata <= X"050C5153";
    when 16#00C2E# => romdata <= X"74101010";
    when 16#00C2F# => romdata <= X"80F89405";
    when 16#00C30# => romdata <= X"88110855";
    when 16#00C31# => romdata <= X"56FEE439";
    when 16#00C32# => romdata <= X"74538075";
    when 16#00C33# => romdata <= X"24A73872";
    when 16#00C34# => romdata <= X"822C8171";
    when 16#00C35# => romdata <= X"2B80F898";
    when 16#00C36# => romdata <= X"080780F8";
    when 16#00C37# => romdata <= X"940B8405";
    when 16#00C38# => romdata <= X"0C53758C";
    when 16#00C39# => romdata <= X"190C7388";
    when 16#00C3A# => romdata <= X"190C7788";
    when 16#00C3B# => romdata <= X"170C778C";
    when 16#00C3C# => romdata <= X"150CFDCD";
    when 16#00C3D# => romdata <= X"39831570";
    when 16#00C3E# => romdata <= X"822C8171";
    when 16#00C3F# => romdata <= X"2B80F898";
    when 16#00C40# => romdata <= X"080780F8";
    when 16#00C41# => romdata <= X"940B8405";
    when 16#00C42# => romdata <= X"0C5153D6";
    when 16#00C43# => romdata <= X"39810B80";
    when 16#00C44# => romdata <= X"0C04803D";
    when 16#00C45# => romdata <= X"0D72812E";
    when 16#00C46# => romdata <= X"8938800B";
    when 16#00C47# => romdata <= X"800C823D";
    when 16#00C48# => romdata <= X"0D047351";
    when 16#00C49# => romdata <= X"80F83FFE";
    when 16#00C4A# => romdata <= X"3D0D818A";
    when 16#00C4B# => romdata <= X"D8085170";
    when 16#00C4C# => romdata <= X"8A38818A";
    when 16#00C4D# => romdata <= X"E470818A";
    when 16#00C4E# => romdata <= X"D80C5170";
    when 16#00C4F# => romdata <= X"75125252";
    when 16#00C50# => romdata <= X"FF537087";
    when 16#00C51# => romdata <= X"FB808026";
    when 16#00C52# => romdata <= X"88387081";
    when 16#00C53# => romdata <= X"8AD80C71";
    when 16#00C54# => romdata <= X"5372800C";
    when 16#00C55# => romdata <= X"843D0D04";
    when 16#00C56# => romdata <= X"FD3D0D80";
    when 16#00C57# => romdata <= X"0B80F0AC";
    when 16#00C58# => romdata <= X"08545472";
    when 16#00C59# => romdata <= X"812E9C38";
    when 16#00C5A# => romdata <= X"73818ADC";
    when 16#00C5B# => romdata <= X"0CFFA6B3";
    when 16#00C5C# => romdata <= X"3FFFA58C";
    when 16#00C5D# => romdata <= X"3F81809C";
    when 16#00C5E# => romdata <= X"528151CF";
    when 16#00C5F# => romdata <= X"943F8008";
    when 16#00C60# => romdata <= X"51A23F72";
    when 16#00C61# => romdata <= X"818ADC0C";
    when 16#00C62# => romdata <= X"FFA6983F";
    when 16#00C63# => romdata <= X"FFA4F13F";
    when 16#00C64# => romdata <= X"81809C52";
    when 16#00C65# => romdata <= X"8151CEF9";
    when 16#00C66# => romdata <= X"3F800851";
    when 16#00C67# => romdata <= X"873F00FF";
    when 16#00C68# => romdata <= X"3900FF39";
    when 16#00C69# => romdata <= X"F73D0D7B";
    when 16#00C6A# => romdata <= X"80F0D808";
    when 16#00C6B# => romdata <= X"82C81108";
    when 16#00C6C# => romdata <= X"5A545A77";
    when 16#00C6D# => romdata <= X"802E80DA";
    when 16#00C6E# => romdata <= X"38818818";
    when 16#00C6F# => romdata <= X"841908FF";
    when 16#00C70# => romdata <= X"0581712B";
    when 16#00C71# => romdata <= X"59555980";
    when 16#00C72# => romdata <= X"742480EA";
    when 16#00C73# => romdata <= X"38807424";
    when 16#00C74# => romdata <= X"B5387382";
    when 16#00C75# => romdata <= X"2B781188";
    when 16#00C76# => romdata <= X"05565681";
    when 16#00C77# => romdata <= X"80190877";
    when 16#00C78# => romdata <= X"06537280";
    when 16#00C79# => romdata <= X"2EB63878";
    when 16#00C7A# => romdata <= X"16700853";
    when 16#00C7B# => romdata <= X"53795174";
    when 16#00C7C# => romdata <= X"0853722D";
    when 16#00C7D# => romdata <= X"FF14FC17";
    when 16#00C7E# => romdata <= X"FC177981";
    when 16#00C7F# => romdata <= X"2C5A5757";
    when 16#00C80# => romdata <= X"54738025";
    when 16#00C81# => romdata <= X"D6387708";
    when 16#00C82# => romdata <= X"5877FFAD";
    when 16#00C83# => romdata <= X"3880F0D8";
    when 16#00C84# => romdata <= X"0853BC13";
    when 16#00C85# => romdata <= X"08A53879";
    when 16#00C86# => romdata <= X"51FF833F";
    when 16#00C87# => romdata <= X"74085372";
    when 16#00C88# => romdata <= X"2DFF14FC";
    when 16#00C89# => romdata <= X"17FC1779";
    when 16#00C8A# => romdata <= X"812C5A57";
    when 16#00C8B# => romdata <= X"57547380";
    when 16#00C8C# => romdata <= X"25FFA838";
    when 16#00C8D# => romdata <= X"D1398057";
    when 16#00C8E# => romdata <= X"FF933972";
    when 16#00C8F# => romdata <= X"51BC1308";
    when 16#00C90# => romdata <= X"53722D79";
    when 16#00C91# => romdata <= X"51FED73F";
    when 16#00C92# => romdata <= X"FF3D0D81";
    when 16#00C93# => romdata <= X"80A40BFC";
    when 16#00C94# => romdata <= X"05700852";
    when 16#00C95# => romdata <= X"5270FF2E";
    when 16#00C96# => romdata <= X"9138702D";
    when 16#00C97# => romdata <= X"FC127008";
    when 16#00C98# => romdata <= X"525270FF";
    when 16#00C99# => romdata <= X"2E098106";
    when 16#00C9A# => romdata <= X"F138833D";
    when 16#00C9B# => romdata <= X"0D0404FF";
    when 16#00C9C# => romdata <= X"A59E3F04";
    when 16#00C9D# => romdata <= X"00000040";
    when 16#00C9E# => romdata <= X"68656C70";
    when 16#00C9F# => romdata <= X"00000000";
    when 16#00CA0# => romdata <= X"3E200000";
    when 16#00CA1# => romdata <= X"636F6D6D";
    when 16#00CA2# => romdata <= X"616E6420";
    when 16#00CA3# => romdata <= X"6E6F7420";
    when 16#00CA4# => romdata <= X"666F756E";
    when 16#00CA5# => romdata <= X"642E0A00";
    when 16#00CA6# => romdata <= X"73757070";
    when 16#00CA7# => romdata <= X"6F727465";
    when 16#00CA8# => romdata <= X"6420636F";
    when 16#00CA9# => romdata <= X"6D6D616E";
    when 16#00CAA# => romdata <= X"64733A0A";
    when 16#00CAB# => romdata <= X"0A000000";
    when 16#00CAC# => romdata <= X"202D2000";
    when 16#00CAD# => romdata <= X"62706D00";
    when 16#00CAE# => romdata <= X"73686F77";
    when 16#00CAF# => romdata <= X"2042504D";
    when 16#00CB0# => romdata <= X"20726567";
    when 16#00CB1# => romdata <= X"69737465";
    when 16#00CB2# => romdata <= X"72730000";
    when 16#00CB3# => romdata <= X"63686563";
    when 16#00CB4# => romdata <= X"6B000000";
    when 16#00CB5# => romdata <= X"63686563";
    when 16#00CB6# => romdata <= X"6B204932";
    when 16#00CB7# => romdata <= X"43206164";
    when 16#00CB8# => romdata <= X"64726573";
    when 16#00CB9# => romdata <= X"73000000";
    when 16#00CBA# => romdata <= X"65646964";
    when 16#00CBB# => romdata <= X"00000000";
    when 16#00CBC# => romdata <= X"72656164";
    when 16#00CBD# => romdata <= X"20454449";
    when 16#00CBE# => romdata <= X"44206469";
    when 16#00CBF# => romdata <= X"73706C61";
    when 16#00CC0# => romdata <= X"79206461";
    when 16#00CC1# => romdata <= X"74610000";
    when 16#00CC2# => romdata <= X"63726561";
    when 16#00CC3# => romdata <= X"64000000";
    when 16#00CC4# => romdata <= X"72656164";
    when 16#00CC5# => romdata <= X"20636872";
    when 16#00CC6# => romdata <= X"6F6E7465";
    when 16#00CC7# => romdata <= X"6C207265";
    when 16#00CC8# => romdata <= X"67697374";
    when 16#00CC9# => romdata <= X"65727300";
    when 16#00CCA# => romdata <= X"63696E69";
    when 16#00CCB# => romdata <= X"74000000";
    when 16#00CCC# => romdata <= X"696E6974";
    when 16#00CCD# => romdata <= X"20636872";
    when 16#00CCE# => romdata <= X"6F6E7465";
    when 16#00CCF# => romdata <= X"6C207265";
    when 16#00CD0# => romdata <= X"67697374";
    when 16#00CD1# => romdata <= X"65727300";
    when 16#00CD2# => romdata <= X"63777269";
    when 16#00CD3# => romdata <= X"74650000";
    when 16#00CD4# => romdata <= X"77726974";
    when 16#00CD5# => romdata <= X"65206368";
    when 16#00CD6# => romdata <= X"726F6E74";
    when 16#00CD7# => romdata <= X"656C2072";
    when 16#00CD8# => romdata <= X"65676973";
    when 16#00CD9# => romdata <= X"74657220";
    when 16#00CDA# => romdata <= X"3C726567";
    when 16#00CDB# => romdata <= X"3E203C76";
    when 16#00CDC# => romdata <= X"616C7565";
    when 16#00CDD# => romdata <= X"3E000000";
    when 16#00CDE# => romdata <= X"6D656D00";
    when 16#00CDF# => romdata <= X"616C6961";
    when 16#00CE0# => romdata <= X"7320666F";
    when 16#00CE1# => romdata <= X"72207800";
    when 16#00CE2# => romdata <= X"776D656D";
    when 16#00CE3# => romdata <= X"00000000";
    when 16#00CE4# => romdata <= X"77726974";
    when 16#00CE5# => romdata <= X"6520776F";
    when 16#00CE6# => romdata <= X"72640000";
    when 16#00CE7# => romdata <= X"6558616D";
    when 16#00CE8# => romdata <= X"696E6520";
    when 16#00CE9# => romdata <= X"6D656D6F";
    when 16#00CEA# => romdata <= X"72790000";
    when 16#00CEB# => romdata <= X"636C6561";
    when 16#00CEC# => romdata <= X"72000000";
    when 16#00CED# => romdata <= X"636C6561";
    when 16#00CEE# => romdata <= X"72207363";
    when 16#00CEF# => romdata <= X"7265656E";
    when 16#00CF0# => romdata <= X"00000000";
    when 16#00CF1# => romdata <= X"71756974";
    when 16#00CF2# => romdata <= X"00000000";
    when 16#00CF3# => romdata <= X"30780000";
    when 16#00CF4# => romdata <= X"0A307800";
    when 16#00CF5# => romdata <= X"203A2000";
    when 16#00CF6# => romdata <= X"69326320";
    when 16#00CF7# => romdata <= X"4456490A";
    when 16#00CF8# => romdata <= X"00000000";
    when 16#00CF9# => romdata <= X"69326320";
    when 16#00CFA# => romdata <= X"464D430A";
    when 16#00CFB# => romdata <= X"00000000";
    when 16#00CFC# => romdata <= X"69326320";
    when 16#00CFD# => romdata <= X"61646472";
    when 16#00CFE# => romdata <= X"6573733A";
    when 16#00CFF# => romdata <= X"20307800";
    when 16#00D00# => romdata <= X"2020202D";
    when 16#00D01# => romdata <= X"2D3E2020";
    when 16#00D02# => romdata <= X"2041434B";
    when 16#00D03# => romdata <= X"0A000000";
    when 16#00D04# => romdata <= X"72656164";
    when 16#00D05# => romdata <= X"20454449";
    when 16#00D06# => romdata <= X"44206461";
    when 16#00D07# => romdata <= X"74612028";
    when 16#00D08# => romdata <= X"00000000";
    when 16#00D09# => romdata <= X"20627974";
    when 16#00D0A# => romdata <= X"65732920";
    when 16#00D0B# => romdata <= X"66726F6D";
    when 16#00D0C# => romdata <= X"20493243";
    when 16#00D0D# => romdata <= X"2D616464";
    when 16#00D0E# => romdata <= X"72657373";
    when 16#00D0F# => romdata <= X"20307800";
    when 16#00D10# => romdata <= X"0A0A0000";
    when 16#00D11# => romdata <= X"6368726F";
    when 16#00D12# => romdata <= X"6E74656C";
    when 16#00D13# => romdata <= X"20726567";
    when 16#00D14# => romdata <= X"20307800";
    when 16#00D15# => romdata <= X"3A203078";
    when 16#00D16# => romdata <= X"00000000";
    when 16#00D17# => romdata <= X"206E6163";
    when 16#00D18# => romdata <= X"6B000000";
    when 16#00D19# => romdata <= X"76616C75";
    when 16#00D1A# => romdata <= X"653A2030";
    when 16#00D1B# => romdata <= X"78000000";
    when 16#00D1C# => romdata <= X"6572726F";
    when 16#00D1D# => romdata <= X"7220286E";
    when 16#00D1E# => romdata <= X"61636B29";
    when 16#00D1F# => romdata <= X"00000000";
    when 16#00D20# => romdata <= X"6265616D";
    when 16#00D21# => romdata <= X"20706F73";
    when 16#00D22# => romdata <= X"6974696F";
    when 16#00D23# => romdata <= X"6E206D6F";
    when 16#00D24# => romdata <= X"6E69746F";
    when 16#00D25# => romdata <= X"72207265";
    when 16#00D26# => romdata <= X"67697374";
    when 16#00D27# => romdata <= X"65727300";
    when 16#00D28# => romdata <= X"0A202020";
    when 16#00D29# => romdata <= X"20202020";
    when 16#00D2A# => romdata <= X"20202020";
    when 16#00D2B# => romdata <= X"20202020";
    when 16#00D2C# => romdata <= X"20202020";
    when 16#00D2D# => romdata <= X"20202020";
    when 16#00D2E# => romdata <= X"20636861";
    when 16#00D2F# => romdata <= X"6E6E656C";
    when 16#00D30# => romdata <= X"20302020";
    when 16#00D31# => romdata <= X"20636861";
    when 16#00D32# => romdata <= X"6E6E656C";
    when 16#00D33# => romdata <= X"20312020";
    when 16#00D34# => romdata <= X"20636861";
    when 16#00D35# => romdata <= X"6E6E656C";
    when 16#00D36# => romdata <= X"20322020";
    when 16#00D37# => romdata <= X"20636861";
    when 16#00D38# => romdata <= X"6E6E656C";
    when 16#00D39# => romdata <= X"20330000";
    when 16#00D3A# => romdata <= X"0A202020";
    when 16#00D3B# => romdata <= X"20202020";
    when 16#00D3C# => romdata <= X"20202020";
    when 16#00D3D# => romdata <= X"20202020";
    when 16#00D3E# => romdata <= X"20202020";
    when 16#00D3F# => romdata <= X"20202020";
    when 16#00D40# => romdata <= X"202D2D2D";
    when 16#00D41# => romdata <= X"2D20686F";
    when 16#00D42# => romdata <= X"72697A6F";
    when 16#00D43# => romdata <= X"6E74616C";
    when 16#00D44# => romdata <= X"202D2D2D";
    when 16#00D45# => romdata <= X"2D2D2020";
    when 16#00D46# => romdata <= X"202D2D2D";
    when 16#00D47# => romdata <= X"2D2D2D20";
    when 16#00D48# => romdata <= X"76657274";
    when 16#00D49# => romdata <= X"6963616C";
    when 16#00D4A# => romdata <= X"202D2D2D";
    when 16#00D4B# => romdata <= X"2D2D0000";
    when 16#00D4C# => romdata <= X"0A736361";
    when 16#00D4D# => romdata <= X"6C657220";
    when 16#00D4E# => romdata <= X"76616C75";
    when 16#00D4F# => romdata <= X"65732020";
    when 16#00D50# => romdata <= X"20202020";
    when 16#00D51# => romdata <= X"20202020";
    when 16#00D52# => romdata <= X"20000000";
    when 16#00D53# => romdata <= X"0A6E6F69";
    when 16#00D54# => romdata <= X"73652063";
    when 16#00D55# => romdata <= X"6F6D7065";
    when 16#00D56# => romdata <= X"6E736174";
    when 16#00D57# => romdata <= X"696F6E20";
    when 16#00D58# => romdata <= X"20202020";
    when 16#00D59# => romdata <= X"20000000";
    when 16#00D5A# => romdata <= X"0A6D6561";
    when 16#00D5B# => romdata <= X"73757265";
    when 16#00D5C# => romdata <= X"6D656E74";
    when 16#00D5D# => romdata <= X"20202020";
    when 16#00D5E# => romdata <= X"20202020";
    when 16#00D5F# => romdata <= X"20202020";
    when 16#00D60# => romdata <= X"20000000";
    when 16#00D61# => romdata <= X"0A73756D";
    when 16#00D62# => romdata <= X"20636861";
    when 16#00D63# => romdata <= X"6E6E656C";
    when 16#00D64# => romdata <= X"2020203A";
    when 16#00D65# => romdata <= X"20000000";
    when 16#00D66# => romdata <= X"0A706F73";
    when 16#00D67# => romdata <= X"6974696F";
    when 16#00D68# => romdata <= X"6E20636F";
    when 16#00D69# => romdata <= X"6D707574";
    when 16#00D6A# => romdata <= X"6174696F";
    when 16#00D6B# => romdata <= X"6E000000";
    when 16#00D6C# => romdata <= X"0A202073";
    when 16#00D6D# => romdata <= X"63616C65";
    when 16#00D6E# => romdata <= X"72207661";
    when 16#00D6F# => romdata <= X"6C756573";
    when 16#00D70# => romdata <= X"20202020";
    when 16#00D71# => romdata <= X"20202020";
    when 16#00D72# => romdata <= X"20000000";
    when 16#00D73# => romdata <= X"0A20206F";
    when 16#00D74# => romdata <= X"66667365";
    when 16#00D75# => romdata <= X"74202020";
    when 16#00D76# => romdata <= X"20202020";
    when 16#00D77# => romdata <= X"20202020";
    when 16#00D78# => romdata <= X"20202020";
    when 16#00D79# => romdata <= X"20000000";
    when 16#00D7A# => romdata <= X"0A6F7574";
    when 16#00D7B# => romdata <= X"70757420";
    when 16#00D7C# => romdata <= X"73656C65";
    when 16#00D7D# => romdata <= X"6374203A";
    when 16#00D7E# => romdata <= X"20000000";
    when 16#00D7F# => romdata <= X"6368616E";
    when 16#00D80# => romdata <= X"6E656C20";
    when 16#00D81# => romdata <= X"30000000";
    when 16#00D82# => romdata <= X"76657274";
    when 16#00D83# => romdata <= X"6963616C";
    when 16#00D84# => romdata <= X"00000000";
    when 16#00D85# => romdata <= X"686F7269";
    when 16#00D86# => romdata <= X"7A6F6E74";
    when 16#00D87# => romdata <= X"616C0000";
    when 16#00D88# => romdata <= X"73756D00";
    when 16#00D89# => romdata <= X"6368616E";
    when 16#00D8A# => romdata <= X"6E656C20";
    when 16#00D8B# => romdata <= X"33000000";
    when 16#00D8C# => romdata <= X"6368616E";
    when 16#00D8D# => romdata <= X"6E656C20";
    when 16#00D8E# => romdata <= X"32000000";
    when 16#00D8F# => romdata <= X"6368616E";
    when 16#00D90# => romdata <= X"6E656C20";
    when 16#00D91# => romdata <= X"31000000";
    when 16#00D92# => romdata <= X"6265616D";
    when 16#00D93# => romdata <= X"20706F73";
    when 16#00D94# => romdata <= X"6974696F";
    when 16#00D95# => romdata <= X"6E206D6F";
    when 16#00D96# => romdata <= X"6E69746F";
    when 16#00D97# => romdata <= X"72000000";
    when 16#00D98# => romdata <= X"20286F6E";
    when 16#00D99# => romdata <= X"2073696D";
    when 16#00D9A# => romdata <= X"290A0000";
    when 16#00D9B# => romdata <= X"0A636F6D";
    when 16#00D9C# => romdata <= X"70696C65";
    when 16#00D9D# => romdata <= X"643A204D";
    when 16#00D9E# => romdata <= X"61792020";
    when 16#00D9F# => romdata <= X"32203230";
    when 16#00DA0# => romdata <= X"31312020";
    when 16#00DA1# => romdata <= X"31313A34";
    when 16#00DA2# => romdata <= X"303A3339";
    when 16#00DA3# => romdata <= X"00000000";
    when 16#00DA4# => romdata <= X"0A737973";
    when 16#00DA5# => romdata <= X"74656D20";
    when 16#00DA6# => romdata <= X"636C6F63";
    when 16#00DA7# => romdata <= X"6B3A2000";
    when 16#00DA8# => romdata <= X"204D487A";
    when 16#00DA9# => romdata <= X"0A000000";
    when 16#00DAA# => romdata <= X"44454255";
    when 16#00DAB# => romdata <= X"47204D4F";
    when 16#00DAC# => romdata <= X"4445204F";
    when 16#00DAD# => romdata <= X"4E0A0000";
    when 16#00DAE# => romdata <= X"000018CB";
    when 16#00DAF# => romdata <= X"00001908";
    when 16#00DB0# => romdata <= X"000018FF";
    when 16#00DB1# => romdata <= X"000018F6";
    when 16#00DB2# => romdata <= X"000018ED";
    when 16#00DB3# => romdata <= X"000018E4";
    when 16#00DB4# => romdata <= X"000018DB";
    when 16#00DB5# => romdata <= X"30622020";
    when 16#00DB6# => romdata <= X"20202020";
    when 16#00DB7# => romdata <= X"20202020";
    when 16#00DB8# => romdata <= X"20202020";
    when 16#00DB9# => romdata <= X"20202020";
    when 16#00DBA# => romdata <= X"20202020";
    when 16#00DBB# => romdata <= X"20202020";
    when 16#00DBC# => romdata <= X"20202020";
    when 16#00DBD# => romdata <= X"20200000";
    when 16#00DBE# => romdata <= X"20202020";
    when 16#00DBF# => romdata <= X"20202020";
    when 16#00DC0# => romdata <= X"00000000";
    when 16#00DC1# => romdata <= X"00202020";
    when 16#00DC2# => romdata <= X"20202020";
    when 16#00DC3# => romdata <= X"20202828";
    when 16#00DC4# => romdata <= X"28282820";
    when 16#00DC5# => romdata <= X"20202020";
    when 16#00DC6# => romdata <= X"20202020";
    when 16#00DC7# => romdata <= X"20202020";
    when 16#00DC8# => romdata <= X"20202020";
    when 16#00DC9# => romdata <= X"20881010";
    when 16#00DCA# => romdata <= X"10101010";
    when 16#00DCB# => romdata <= X"10101010";
    when 16#00DCC# => romdata <= X"10101010";
    when 16#00DCD# => romdata <= X"10040404";
    when 16#00DCE# => romdata <= X"04040404";
    when 16#00DCF# => romdata <= X"04040410";
    when 16#00DD0# => romdata <= X"10101010";
    when 16#00DD1# => romdata <= X"10104141";
    when 16#00DD2# => romdata <= X"41414141";
    when 16#00DD3# => romdata <= X"01010101";
    when 16#00DD4# => romdata <= X"01010101";
    when 16#00DD5# => romdata <= X"01010101";
    when 16#00DD6# => romdata <= X"01010101";
    when 16#00DD7# => romdata <= X"01010101";
    when 16#00DD8# => romdata <= X"10101010";
    when 16#00DD9# => romdata <= X"10104242";
    when 16#00DDA# => romdata <= X"42424242";
    when 16#00DDB# => romdata <= X"02020202";
    when 16#00DDC# => romdata <= X"02020202";
    when 16#00DDD# => romdata <= X"02020202";
    when 16#00DDE# => romdata <= X"02020202";
    when 16#00DDF# => romdata <= X"02020202";
    when 16#00DE0# => romdata <= X"10101010";
    when 16#00DE1# => romdata <= X"20000000";
    when 16#00DE2# => romdata <= X"00000000";
    when 16#00DE3# => romdata <= X"00000000";
    when 16#00DE4# => romdata <= X"00000000";
    when 16#00DE5# => romdata <= X"00000000";
    when 16#00DE6# => romdata <= X"00000000";
    when 16#00DE7# => romdata <= X"00000000";
    when 16#00DE8# => romdata <= X"00000000";
    when 16#00DE9# => romdata <= X"00000000";
    when 16#00DEA# => romdata <= X"00000000";
    when 16#00DEB# => romdata <= X"00000000";
    when 16#00DEC# => romdata <= X"00000000";
    when 16#00DED# => romdata <= X"00000000";
    when 16#00DEE# => romdata <= X"00000000";
    when 16#00DEF# => romdata <= X"00000000";
    when 16#00DF0# => romdata <= X"00000000";
    when 16#00DF1# => romdata <= X"00000000";
    when 16#00DF2# => romdata <= X"00000000";
    when 16#00DF3# => romdata <= X"00000000";
    when 16#00DF4# => romdata <= X"00000000";
    when 16#00DF5# => romdata <= X"00000000";
    when 16#00DF6# => romdata <= X"00000000";
    when 16#00DF7# => romdata <= X"00000000";
    when 16#00DF8# => romdata <= X"00000000";
    when 16#00DF9# => romdata <= X"00000000";
    when 16#00DFA# => romdata <= X"00000000";
    when 16#00DFB# => romdata <= X"00000000";
    when 16#00DFC# => romdata <= X"00000000";
    when 16#00DFD# => romdata <= X"00000000";
    when 16#00DFE# => romdata <= X"00000000";
    when 16#00DFF# => romdata <= X"00000000";
    when 16#00E00# => romdata <= X"00000000";
    when 16#00E01# => romdata <= X"00000000";
    when 16#00E02# => romdata <= X"43000000";
    when 16#00E03# => romdata <= X"64756D6D";
    when 16#00E04# => romdata <= X"792E6578";
    when 16#00E05# => romdata <= X"65000000";
    when 16#00E06# => romdata <= X"00FFFFFF";
    when 16#00E07# => romdata <= X"FF00FFFF";
    when 16#00E08# => romdata <= X"FFFF00FF";
    when 16#00E09# => romdata <= X"FFFFFF00";
    when 16#00E0A# => romdata <= X"00000000";
    when 16#00E0B# => romdata <= X"00000000";
    when 16#00E0C# => romdata <= X"00000000";
    when 16#00E0D# => romdata <= X"0000402C";
    when 16#00E0E# => romdata <= X"80000A00";
    when 16#00E0F# => romdata <= X"80000700";
    when 16#00E10# => romdata <= X"80000800";
    when 16#00E11# => romdata <= X"80000600";
    when 16#00E12# => romdata <= X"80000400";
    when 16#00E13# => romdata <= X"80000200";
    when 16#00E14# => romdata <= X"80000100";
    when 16#00E15# => romdata <= X"80000000";
    when 16#00E16# => romdata <= X"0000385C";
    when 16#00E17# => romdata <= X"00000000";
    when 16#00E18# => romdata <= X"00003AC4";
    when 16#00E19# => romdata <= X"00003B20";
    when 16#00E1A# => romdata <= X"00003B7C";
    when 16#00E1B# => romdata <= X"00000000";
    when 16#00E1C# => romdata <= X"00000000";
    when 16#00E1D# => romdata <= X"00000000";
    when 16#00E1E# => romdata <= X"00000000";
    when 16#00E1F# => romdata <= X"00000000";
    when 16#00E20# => romdata <= X"00000000";
    when 16#00E21# => romdata <= X"00000000";
    when 16#00E22# => romdata <= X"00000000";
    when 16#00E23# => romdata <= X"00000000";
    when 16#00E24# => romdata <= X"00003808";
    when 16#00E25# => romdata <= X"00000000";
    when 16#00E26# => romdata <= X"00000000";
    when 16#00E27# => romdata <= X"00000000";
    when 16#00E28# => romdata <= X"00000000";
    when 16#00E29# => romdata <= X"00000000";
    when 16#00E2A# => romdata <= X"00000000";
    when 16#00E2B# => romdata <= X"00000000";
    when 16#00E2C# => romdata <= X"00000000";
    when 16#00E2D# => romdata <= X"00000000";
    when 16#00E2E# => romdata <= X"00000000";
    when 16#00E2F# => romdata <= X"00000000";
    when 16#00E30# => romdata <= X"00000000";
    when 16#00E31# => romdata <= X"00000000";
    when 16#00E32# => romdata <= X"00000000";
    when 16#00E33# => romdata <= X"00000000";
    when 16#00E34# => romdata <= X"00000000";
    when 16#00E35# => romdata <= X"00000000";
    when 16#00E36# => romdata <= X"00000000";
    when 16#00E37# => romdata <= X"00000000";
    when 16#00E38# => romdata <= X"00000000";
    when 16#00E39# => romdata <= X"00000000";
    when 16#00E3A# => romdata <= X"00000000";
    when 16#00E3B# => romdata <= X"00000000";
    when 16#00E3C# => romdata <= X"00000000";
    when 16#00E3D# => romdata <= X"00000000";
    when 16#00E3E# => romdata <= X"00000000";
    when 16#00E3F# => romdata <= X"00000000";
    when 16#00E40# => romdata <= X"00000000";
    when 16#00E41# => romdata <= X"00000001";
    when 16#00E42# => romdata <= X"330EABCD";
    when 16#00E43# => romdata <= X"1234E66D";
    when 16#00E44# => romdata <= X"DEEC0005";
    when 16#00E45# => romdata <= X"000B0000";
    when 16#00E46# => romdata <= X"00000000";
    when 16#00E47# => romdata <= X"00000000";
    when 16#00E48# => romdata <= X"00000000";
    when 16#00E49# => romdata <= X"00000000";
    when 16#00E4A# => romdata <= X"00000000";
    when 16#00E4B# => romdata <= X"00000000";
    when 16#00E4C# => romdata <= X"00000000";
    when 16#00E4D# => romdata <= X"00000000";
    when 16#00E4E# => romdata <= X"00000000";
    when 16#00E4F# => romdata <= X"00000000";
    when 16#00E50# => romdata <= X"00000000";
    when 16#00E51# => romdata <= X"00000000";
    when 16#00E52# => romdata <= X"00000000";
    when 16#00E53# => romdata <= X"00000000";
    when 16#00E54# => romdata <= X"00000000";
    when 16#00E55# => romdata <= X"00000000";
    when 16#00E56# => romdata <= X"00000000";
    when 16#00E57# => romdata <= X"00000000";
    when 16#00E58# => romdata <= X"00000000";
    when 16#00E59# => romdata <= X"00000000";
    when 16#00E5A# => romdata <= X"00000000";
    when 16#00E5B# => romdata <= X"00000000";
    when 16#00E5C# => romdata <= X"00000000";
    when 16#00E5D# => romdata <= X"00000000";
    when 16#00E5E# => romdata <= X"00000000";
    when 16#00E5F# => romdata <= X"00000000";
    when 16#00E60# => romdata <= X"00000000";
    when 16#00E61# => romdata <= X"00000000";
    when 16#00E62# => romdata <= X"00000000";
    when 16#00E63# => romdata <= X"00000000";
    when 16#00E64# => romdata <= X"00000000";
    when 16#00E65# => romdata <= X"00000000";
    when 16#00E66# => romdata <= X"00000000";
    when 16#00E67# => romdata <= X"00000000";
    when 16#00E68# => romdata <= X"00000000";
    when 16#00E69# => romdata <= X"00000000";
    when 16#00E6A# => romdata <= X"00000000";
    when 16#00E6B# => romdata <= X"00000000";
    when 16#00E6C# => romdata <= X"00000000";
    when 16#00E6D# => romdata <= X"00000000";
    when 16#00E6E# => romdata <= X"00000000";
    when 16#00E6F# => romdata <= X"00000000";
    when 16#00E70# => romdata <= X"00000000";
    when 16#00E71# => romdata <= X"00000000";
    when 16#00E72# => romdata <= X"00000000";
    when 16#00E73# => romdata <= X"00000000";
    when 16#00E74# => romdata <= X"00000000";
    when 16#00E75# => romdata <= X"00000000";
    when 16#00E76# => romdata <= X"00000000";
    when 16#00E77# => romdata <= X"00000000";
    when 16#00E78# => romdata <= X"00000000";
    when 16#00E79# => romdata <= X"00000000";
    when 16#00E7A# => romdata <= X"00000000";
    when 16#00E7B# => romdata <= X"00000000";
    when 16#00E7C# => romdata <= X"00000000";
    when 16#00E7D# => romdata <= X"00000000";
    when 16#00E7E# => romdata <= X"00000000";
    when 16#00E7F# => romdata <= X"00000000";
    when 16#00E80# => romdata <= X"00000000";
    when 16#00E81# => romdata <= X"00000000";
    when 16#00E82# => romdata <= X"00000000";
    when 16#00E83# => romdata <= X"00000000";
    when 16#00E84# => romdata <= X"00000000";
    when 16#00E85# => romdata <= X"00000000";
    when 16#00E86# => romdata <= X"00000000";
    when 16#00E87# => romdata <= X"00000000";
    when 16#00E88# => romdata <= X"00000000";
    when 16#00E89# => romdata <= X"00000000";
    when 16#00E8A# => romdata <= X"00000000";
    when 16#00E8B# => romdata <= X"00000000";
    when 16#00E8C# => romdata <= X"00000000";
    when 16#00E8D# => romdata <= X"00000000";
    when 16#00E8E# => romdata <= X"00000000";
    when 16#00E8F# => romdata <= X"00000000";
    when 16#00E90# => romdata <= X"00000000";
    when 16#00E91# => romdata <= X"00000000";
    when 16#00E92# => romdata <= X"00000000";
    when 16#00E93# => romdata <= X"00000000";
    when 16#00E94# => romdata <= X"00000000";
    when 16#00E95# => romdata <= X"00000000";
    when 16#00E96# => romdata <= X"00000000";
    when 16#00E97# => romdata <= X"00000000";
    when 16#00E98# => romdata <= X"00000000";
    when 16#00E99# => romdata <= X"00000000";
    when 16#00E9A# => romdata <= X"00000000";
    when 16#00E9B# => romdata <= X"00000000";
    when 16#00E9C# => romdata <= X"00000000";
    when 16#00E9D# => romdata <= X"00000000";
    when 16#00E9E# => romdata <= X"00000000";
    when 16#00E9F# => romdata <= X"00000000";
    when 16#00EA0# => romdata <= X"00000000";
    when 16#00EA1# => romdata <= X"00000000";
    when 16#00EA2# => romdata <= X"00000000";
    when 16#00EA3# => romdata <= X"00000000";
    when 16#00EA4# => romdata <= X"00000000";
    when 16#00EA5# => romdata <= X"00000000";
    when 16#00EA6# => romdata <= X"00000000";
    when 16#00EA7# => romdata <= X"00000000";
    when 16#00EA8# => romdata <= X"00000000";
    when 16#00EA9# => romdata <= X"00000000";
    when 16#00EAA# => romdata <= X"00000000";
    when 16#00EAB# => romdata <= X"00000000";
    when 16#00EAC# => romdata <= X"00000000";
    when 16#00EAD# => romdata <= X"00000000";
    when 16#00EAE# => romdata <= X"00000000";
    when 16#00EAF# => romdata <= X"00000000";
    when 16#00EB0# => romdata <= X"00000000";
    when 16#00EB1# => romdata <= X"00000000";
    when 16#00EB2# => romdata <= X"00000000";
    when 16#00EB3# => romdata <= X"00000000";
    when 16#00EB4# => romdata <= X"00000000";
    when 16#00EB5# => romdata <= X"00000000";
    when 16#00EB6# => romdata <= X"00000000";
    when 16#00EB7# => romdata <= X"00000000";
    when 16#00EB8# => romdata <= X"00000000";
    when 16#00EB9# => romdata <= X"00000000";
    when 16#00EBA# => romdata <= X"00000000";
    when 16#00EBB# => romdata <= X"00000000";
    when 16#00EBC# => romdata <= X"00000000";
    when 16#00EBD# => romdata <= X"00000000";
    when 16#00EBE# => romdata <= X"00000000";
    when 16#00EBF# => romdata <= X"00000000";
    when 16#00EC0# => romdata <= X"00000000";
    when 16#00EC1# => romdata <= X"00000000";
    when 16#00EC2# => romdata <= X"00000000";
    when 16#00EC3# => romdata <= X"00000000";
    when 16#00EC4# => romdata <= X"00000000";
    when 16#00EC5# => romdata <= X"00000000";
    when 16#00EC6# => romdata <= X"00000000";
    when 16#00EC7# => romdata <= X"00000000";
    when 16#00EC8# => romdata <= X"00000000";
    when 16#00EC9# => romdata <= X"00000000";
    when 16#00ECA# => romdata <= X"00000000";
    when 16#00ECB# => romdata <= X"00000000";
    when 16#00ECC# => romdata <= X"00000000";
    when 16#00ECD# => romdata <= X"00000000";
    when 16#00ECE# => romdata <= X"00000000";
    when 16#00ECF# => romdata <= X"00000000";
    when 16#00ED0# => romdata <= X"00000000";
    when 16#00ED1# => romdata <= X"00000000";
    when 16#00ED2# => romdata <= X"00000000";
    when 16#00ED3# => romdata <= X"00000000";
    when 16#00ED4# => romdata <= X"00000000";
    when 16#00ED5# => romdata <= X"00000000";
    when 16#00ED6# => romdata <= X"00000000";
    when 16#00ED7# => romdata <= X"00000000";
    when 16#00ED8# => romdata <= X"00000000";
    when 16#00ED9# => romdata <= X"00000000";
    when 16#00EDA# => romdata <= X"00000000";
    when 16#00EDB# => romdata <= X"00000000";
    when 16#00EDC# => romdata <= X"00000000";
    when 16#00EDD# => romdata <= X"00000000";
    when 16#00EDE# => romdata <= X"00000000";
    when 16#00EDF# => romdata <= X"00000000";
    when 16#00EE0# => romdata <= X"00000000";
    when 16#00EE1# => romdata <= X"00000000";
    when 16#00EE2# => romdata <= X"00000000";
    when 16#00EE3# => romdata <= X"00000000";
    when 16#00EE4# => romdata <= X"00000000";
    when 16#00EE5# => romdata <= X"00000000";
    when 16#00EE6# => romdata <= X"00000000";
    when 16#00EE7# => romdata <= X"00000000";
    when 16#00EE8# => romdata <= X"00000000";
    when 16#00EE9# => romdata <= X"00000000";
    when 16#00EEA# => romdata <= X"00000000";
    when 16#00EEB# => romdata <= X"00000000";
    when 16#00EEC# => romdata <= X"00000000";
    when 16#00EED# => romdata <= X"00000000";
    when 16#00EEE# => romdata <= X"00000000";
    when 16#00EEF# => romdata <= X"00000000";
    when 16#00EF0# => romdata <= X"00000000";
    when 16#00EF1# => romdata <= X"00000000";
    when 16#00EF2# => romdata <= X"00000000";
    when 16#00EF3# => romdata <= X"00000000";
    when 16#00EF4# => romdata <= X"00000000";
    when 16#00EF5# => romdata <= X"00000000";
    when 16#00EF6# => romdata <= X"00000000";
    when 16#00EF7# => romdata <= X"00000000";
    when 16#00EF8# => romdata <= X"00000000";
    when 16#00EF9# => romdata <= X"00000000";
    when 16#00EFA# => romdata <= X"00000000";
    when 16#00EFB# => romdata <= X"00000000";
    when 16#00EFC# => romdata <= X"00000000";
    when 16#00EFD# => romdata <= X"00000000";
    when 16#00EFE# => romdata <= X"00000000";
    when 16#00EFF# => romdata <= X"00000000";
    when 16#00F00# => romdata <= X"00000000";
    when 16#00F01# => romdata <= X"00000000";
    when 16#00F02# => romdata <= X"FFFFFFFF";
    when 16#00F03# => romdata <= X"00000000";
    when 16#00F04# => romdata <= X"00020000";
    when 16#00F05# => romdata <= X"00000000";
    when 16#00F06# => romdata <= X"00000000";
    when 16#00F07# => romdata <= X"00003C14";
    when 16#00F08# => romdata <= X"00003C14";
    when 16#00F09# => romdata <= X"00003C1C";
    when 16#00F0A# => romdata <= X"00003C1C";
    when 16#00F0B# => romdata <= X"00003C24";
    when 16#00F0C# => romdata <= X"00003C24";
    when 16#00F0D# => romdata <= X"00003C2C";
    when 16#00F0E# => romdata <= X"00003C2C";
    when 16#00F0F# => romdata <= X"00003C34";
    when 16#00F10# => romdata <= X"00003C34";
    when 16#00F11# => romdata <= X"00003C3C";
    when 16#00F12# => romdata <= X"00003C3C";
    when 16#00F13# => romdata <= X"00003C44";
    when 16#00F14# => romdata <= X"00003C44";
    when 16#00F15# => romdata <= X"00003C4C";
    when 16#00F16# => romdata <= X"00003C4C";
    when 16#00F17# => romdata <= X"00003C54";
    when 16#00F18# => romdata <= X"00003C54";
    when 16#00F19# => romdata <= X"00003C5C";
    when 16#00F1A# => romdata <= X"00003C5C";
    when 16#00F1B# => romdata <= X"00003C64";
    when 16#00F1C# => romdata <= X"00003C64";
    when 16#00F1D# => romdata <= X"00003C6C";
    when 16#00F1E# => romdata <= X"00003C6C";
    when 16#00F1F# => romdata <= X"00003C74";
    when 16#00F20# => romdata <= X"00003C74";
    when 16#00F21# => romdata <= X"00003C7C";
    when 16#00F22# => romdata <= X"00003C7C";
    when 16#00F23# => romdata <= X"00003C84";
    when 16#00F24# => romdata <= X"00003C84";
    when 16#00F25# => romdata <= X"00003C8C";
    when 16#00F26# => romdata <= X"00003C8C";
    when 16#00F27# => romdata <= X"00003C94";
    when 16#00F28# => romdata <= X"00003C94";
    when 16#00F29# => romdata <= X"00003C9C";
    when 16#00F2A# => romdata <= X"00003C9C";
    when 16#00F2B# => romdata <= X"00003CA4";
    when 16#00F2C# => romdata <= X"00003CA4";
    when 16#00F2D# => romdata <= X"00003CAC";
    when 16#00F2E# => romdata <= X"00003CAC";
    when 16#00F2F# => romdata <= X"00003CB4";
    when 16#00F30# => romdata <= X"00003CB4";
    when 16#00F31# => romdata <= X"00003CBC";
    when 16#00F32# => romdata <= X"00003CBC";
    when 16#00F33# => romdata <= X"00003CC4";
    when 16#00F34# => romdata <= X"00003CC4";
    when 16#00F35# => romdata <= X"00003CCC";
    when 16#00F36# => romdata <= X"00003CCC";
    when 16#00F37# => romdata <= X"00003CD4";
    when 16#00F38# => romdata <= X"00003CD4";
    when 16#00F39# => romdata <= X"00003CDC";
    when 16#00F3A# => romdata <= X"00003CDC";
    when 16#00F3B# => romdata <= X"00003CE4";
    when 16#00F3C# => romdata <= X"00003CE4";
    when 16#00F3D# => romdata <= X"00003CEC";
    when 16#00F3E# => romdata <= X"00003CEC";
    when 16#00F3F# => romdata <= X"00003CF4";
    when 16#00F40# => romdata <= X"00003CF4";
    when 16#00F41# => romdata <= X"00003CFC";
    when 16#00F42# => romdata <= X"00003CFC";
    when 16#00F43# => romdata <= X"00003D04";
    when 16#00F44# => romdata <= X"00003D04";
    when 16#00F45# => romdata <= X"00003D0C";
    when 16#00F46# => romdata <= X"00003D0C";
    when 16#00F47# => romdata <= X"00003D14";
    when 16#00F48# => romdata <= X"00003D14";
    when 16#00F49# => romdata <= X"00003D1C";
    when 16#00F4A# => romdata <= X"00003D1C";
    when 16#00F4B# => romdata <= X"00003D24";
    when 16#00F4C# => romdata <= X"00003D24";
    when 16#00F4D# => romdata <= X"00003D2C";
    when 16#00F4E# => romdata <= X"00003D2C";
    when 16#00F4F# => romdata <= X"00003D34";
    when 16#00F50# => romdata <= X"00003D34";
    when 16#00F51# => romdata <= X"00003D3C";
    when 16#00F52# => romdata <= X"00003D3C";
    when 16#00F53# => romdata <= X"00003D44";
    when 16#00F54# => romdata <= X"00003D44";
    when 16#00F55# => romdata <= X"00003D4C";
    when 16#00F56# => romdata <= X"00003D4C";
    when 16#00F57# => romdata <= X"00003D54";
    when 16#00F58# => romdata <= X"00003D54";
    when 16#00F59# => romdata <= X"00003D5C";
    when 16#00F5A# => romdata <= X"00003D5C";
    when 16#00F5B# => romdata <= X"00003D64";
    when 16#00F5C# => romdata <= X"00003D64";
    when 16#00F5D# => romdata <= X"00003D6C";
    when 16#00F5E# => romdata <= X"00003D6C";
    when 16#00F5F# => romdata <= X"00003D74";
    when 16#00F60# => romdata <= X"00003D74";
    when 16#00F61# => romdata <= X"00003D7C";
    when 16#00F62# => romdata <= X"00003D7C";
    when 16#00F63# => romdata <= X"00003D84";
    when 16#00F64# => romdata <= X"00003D84";
    when 16#00F65# => romdata <= X"00003D8C";
    when 16#00F66# => romdata <= X"00003D8C";
    when 16#00F67# => romdata <= X"00003D94";
    when 16#00F68# => romdata <= X"00003D94";
    when 16#00F69# => romdata <= X"00003D9C";
    when 16#00F6A# => romdata <= X"00003D9C";
    when 16#00F6B# => romdata <= X"00003DA4";
    when 16#00F6C# => romdata <= X"00003DA4";
    when 16#00F6D# => romdata <= X"00003DAC";
    when 16#00F6E# => romdata <= X"00003DAC";
    when 16#00F6F# => romdata <= X"00003DB4";
    when 16#00F70# => romdata <= X"00003DB4";
    when 16#00F71# => romdata <= X"00003DBC";
    when 16#00F72# => romdata <= X"00003DBC";
    when 16#00F73# => romdata <= X"00003DC4";
    when 16#00F74# => romdata <= X"00003DC4";
    when 16#00F75# => romdata <= X"00003DCC";
    when 16#00F76# => romdata <= X"00003DCC";
    when 16#00F77# => romdata <= X"00003DD4";
    when 16#00F78# => romdata <= X"00003DD4";
    when 16#00F79# => romdata <= X"00003DDC";
    when 16#00F7A# => romdata <= X"00003DDC";
    when 16#00F7B# => romdata <= X"00003DE4";
    when 16#00F7C# => romdata <= X"00003DE4";
    when 16#00F7D# => romdata <= X"00003DEC";
    when 16#00F7E# => romdata <= X"00003DEC";
    when 16#00F7F# => romdata <= X"00003DF4";
    when 16#00F80# => romdata <= X"00003DF4";
    when 16#00F81# => romdata <= X"00003DFC";
    when 16#00F82# => romdata <= X"00003DFC";
    when 16#00F83# => romdata <= X"00003E04";
    when 16#00F84# => romdata <= X"00003E04";
    when 16#00F85# => romdata <= X"00003E0C";
    when 16#00F86# => romdata <= X"00003E0C";
    when 16#00F87# => romdata <= X"00003E14";
    when 16#00F88# => romdata <= X"00003E14";
    when 16#00F89# => romdata <= X"00003E1C";
    when 16#00F8A# => romdata <= X"00003E1C";
    when 16#00F8B# => romdata <= X"00003E24";
    when 16#00F8C# => romdata <= X"00003E24";
    when 16#00F8D# => romdata <= X"00003E2C";
    when 16#00F8E# => romdata <= X"00003E2C";
    when 16#00F8F# => romdata <= X"00003E34";
    when 16#00F90# => romdata <= X"00003E34";
    when 16#00F91# => romdata <= X"00003E3C";
    when 16#00F92# => romdata <= X"00003E3C";
    when 16#00F93# => romdata <= X"00003E44";
    when 16#00F94# => romdata <= X"00003E44";
    when 16#00F95# => romdata <= X"00003E4C";
    when 16#00F96# => romdata <= X"00003E4C";
    when 16#00F97# => romdata <= X"00003E54";
    when 16#00F98# => romdata <= X"00003E54";
    when 16#00F99# => romdata <= X"00003E5C";
    when 16#00F9A# => romdata <= X"00003E5C";
    when 16#00F9B# => romdata <= X"00003E64";
    when 16#00F9C# => romdata <= X"00003E64";
    when 16#00F9D# => romdata <= X"00003E6C";
    when 16#00F9E# => romdata <= X"00003E6C";
    when 16#00F9F# => romdata <= X"00003E74";
    when 16#00FA0# => romdata <= X"00003E74";
    when 16#00FA1# => romdata <= X"00003E7C";
    when 16#00FA2# => romdata <= X"00003E7C";
    when 16#00FA3# => romdata <= X"00003E84";
    when 16#00FA4# => romdata <= X"00003E84";
    when 16#00FA5# => romdata <= X"00003E8C";
    when 16#00FA6# => romdata <= X"00003E8C";
    when 16#00FA7# => romdata <= X"00003E94";
    when 16#00FA8# => romdata <= X"00003E94";
    when 16#00FA9# => romdata <= X"00003E9C";
    when 16#00FAA# => romdata <= X"00003E9C";
    when 16#00FAB# => romdata <= X"00003EA4";
    when 16#00FAC# => romdata <= X"00003EA4";
    when 16#00FAD# => romdata <= X"00003EAC";
    when 16#00FAE# => romdata <= X"00003EAC";
    when 16#00FAF# => romdata <= X"00003EB4";
    when 16#00FB0# => romdata <= X"00003EB4";
    when 16#00FB1# => romdata <= X"00003EBC";
    when 16#00FB2# => romdata <= X"00003EBC";
    when 16#00FB3# => romdata <= X"00003EC4";
    when 16#00FB4# => romdata <= X"00003EC4";
    when 16#00FB5# => romdata <= X"00003ECC";
    when 16#00FB6# => romdata <= X"00003ECC";
    when 16#00FB7# => romdata <= X"00003ED4";
    when 16#00FB8# => romdata <= X"00003ED4";
    when 16#00FB9# => romdata <= X"00003EDC";
    when 16#00FBA# => romdata <= X"00003EDC";
    when 16#00FBB# => romdata <= X"00003EE4";
    when 16#00FBC# => romdata <= X"00003EE4";
    when 16#00FBD# => romdata <= X"00003EEC";
    when 16#00FBE# => romdata <= X"00003EEC";
    when 16#00FBF# => romdata <= X"00003EF4";
    when 16#00FC0# => romdata <= X"00003EF4";
    when 16#00FC1# => romdata <= X"00003EFC";
    when 16#00FC2# => romdata <= X"00003EFC";
    when 16#00FC3# => romdata <= X"00003F04";
    when 16#00FC4# => romdata <= X"00003F04";
    when 16#00FC5# => romdata <= X"00003F0C";
    when 16#00FC6# => romdata <= X"00003F0C";
    when 16#00FC7# => romdata <= X"00003F14";
    when 16#00FC8# => romdata <= X"00003F14";
    when 16#00FC9# => romdata <= X"00003F1C";
    when 16#00FCA# => romdata <= X"00003F1C";
    when 16#00FCB# => romdata <= X"00003F24";
    when 16#00FCC# => romdata <= X"00003F24";
    when 16#00FCD# => romdata <= X"00003F2C";
    when 16#00FCE# => romdata <= X"00003F2C";
    when 16#00FCF# => romdata <= X"00003F34";
    when 16#00FD0# => romdata <= X"00003F34";
    when 16#00FD1# => romdata <= X"00003F3C";
    when 16#00FD2# => romdata <= X"00003F3C";
    when 16#00FD3# => romdata <= X"00003F44";
    when 16#00FD4# => romdata <= X"00003F44";
    when 16#00FD5# => romdata <= X"00003F4C";
    when 16#00FD6# => romdata <= X"00003F4C";
    when 16#00FD7# => romdata <= X"00003F54";
    when 16#00FD8# => romdata <= X"00003F54";
    when 16#00FD9# => romdata <= X"00003F5C";
    when 16#00FDA# => romdata <= X"00003F5C";
    when 16#00FDB# => romdata <= X"00003F64";
    when 16#00FDC# => romdata <= X"00003F64";
    when 16#00FDD# => romdata <= X"00003F6C";
    when 16#00FDE# => romdata <= X"00003F6C";
    when 16#00FDF# => romdata <= X"00003F74";
    when 16#00FE0# => romdata <= X"00003F74";
    when 16#00FE1# => romdata <= X"00003F7C";
    when 16#00FE2# => romdata <= X"00003F7C";
    when 16#00FE3# => romdata <= X"00003F84";
    when 16#00FE4# => romdata <= X"00003F84";
    when 16#00FE5# => romdata <= X"00003F8C";
    when 16#00FE6# => romdata <= X"00003F8C";
    when 16#00FE7# => romdata <= X"00003F94";
    when 16#00FE8# => romdata <= X"00003F94";
    when 16#00FE9# => romdata <= X"00003F9C";
    when 16#00FEA# => romdata <= X"00003F9C";
    when 16#00FEB# => romdata <= X"00003FA4";
    when 16#00FEC# => romdata <= X"00003FA4";
    when 16#00FED# => romdata <= X"00003FAC";
    when 16#00FEE# => romdata <= X"00003FAC";
    when 16#00FEF# => romdata <= X"00003FB4";
    when 16#00FF0# => romdata <= X"00003FB4";
    when 16#00FF1# => romdata <= X"00003FBC";
    when 16#00FF2# => romdata <= X"00003FBC";
    when 16#00FF3# => romdata <= X"00003FC4";
    when 16#00FF4# => romdata <= X"00003FC4";
    when 16#00FF5# => romdata <= X"00003FCC";
    when 16#00FF6# => romdata <= X"00003FCC";
    when 16#00FF7# => romdata <= X"00003FD4";
    when 16#00FF8# => romdata <= X"00003FD4";
    when 16#00FF9# => romdata <= X"00003FDC";
    when 16#00FFA# => romdata <= X"00003FDC";
    when 16#00FFB# => romdata <= X"00003FE4";
    when 16#00FFC# => romdata <= X"00003FE4";
    when 16#00FFD# => romdata <= X"00003FEC";
    when 16#00FFE# => romdata <= X"00003FEC";
    when 16#00FFF# => romdata <= X"00003FF4";
    when 16#01000# => romdata <= X"00003FF4";
    when 16#01001# => romdata <= X"00003FFC";
    when 16#01002# => romdata <= X"00003FFC";
    when 16#01003# => romdata <= X"00004004";
    when 16#01004# => romdata <= X"00004004";
    when 16#01005# => romdata <= X"0000400C";
    when 16#01006# => romdata <= X"0000400C";
    when 16#01007# => romdata <= X"0000380C";
    when 16#01008# => romdata <= X"FFFFFFFF";
    when 16#01009# => romdata <= X"00000000";
    when 16#0100A# => romdata <= X"FFFFFFFF";
    when 16#0100B# => romdata <= X"00000000";
    when 16#0100C# => romdata <= X"00000000";
    when 16#0100D# => romdata <= X"00000000";
    when others => romdata <= (others => '-');
    end case;
  end process;
  -- pragma translate_off
  bootmsg : report_version 
  generic map ("ahbrom" & tost(hindex) &
  ": 32-bit AHB ROM Module,  " & tost(bytes/4) & " words, " & tost(abits-2) & " address bits" );
  -- pragma translate_on
  end;
