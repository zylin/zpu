-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"0bbaa40c",
     3 => x"3a0b0b0b",
     4 => x"b2de0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"0bb3a02d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b0bba",
   162 => x"90738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0bad",
   171 => x"c92d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bae",
   179 => x"fb2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"0bbaa00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"81fb3fac",
   257 => x"c03f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104ba",
   280 => x"a008802e",
   281 => x"a338baa4",
   282 => x"08822ebd",
   283 => x"38838080",
   284 => x"0b0b0b80",
   285 => x"c1d80c82",
   286 => x"a0800b80",
   287 => x"c1dc0c82",
   288 => x"90800b80",
   289 => x"c1e00c04",
   290 => x"f8808080",
   291 => x"a40b0b0b",
   292 => x"80c1d80c",
   293 => x"f8808082",
   294 => x"800b80c1",
   295 => x"dc0cf880",
   296 => x"8084800b",
   297 => x"80c1e00c",
   298 => x"0480c0a8",
   299 => x"808c0b0b",
   300 => x"0b80c1d8",
   301 => x"0c80c0a8",
   302 => x"80940b80",
   303 => x"c1dc0c0b",
   304 => x"0b0bb4f0",
   305 => x"0b80c1e0",
   306 => x"0c04ff3d",
   307 => x"0d80c1e4",
   308 => x"335170a4",
   309 => x"38baac08",
   310 => x"70085252",
   311 => x"70802e92",
   312 => x"388412ba",
   313 => x"ac0c702d",
   314 => x"baac0870",
   315 => x"08525270",
   316 => x"f038810b",
   317 => x"80c1e434",
   318 => x"833d0d04",
   319 => x"04803d0d",
   320 => x"0b0b80c1",
   321 => x"d408802e",
   322 => x"8e380b0b",
   323 => x"0b0b800b",
   324 => x"802e0981",
   325 => x"06853882",
   326 => x"3d0d040b",
   327 => x"0b80c1d4",
   328 => x"510b0b0b",
   329 => x"f5da3f82",
   330 => x"3d0d0404",
   331 => x"fd3d0dba",
   332 => x"b80876b0",
   333 => x"ea299412",
   334 => x"0c54850b",
   335 => x"98150c98",
   336 => x"14087081",
   337 => x"06515372",
   338 => x"f638853d",
   339 => x"0d04ff3d",
   340 => x"0dbab808",
   341 => x"74101075",
   342 => x"10059412",
   343 => x"0c52850b",
   344 => x"98130c98",
   345 => x"12087081",
   346 => x"06515170",
   347 => x"f638833d",
   348 => x"0d04803d",
   349 => x"0d725180",
   350 => x"71278738",
   351 => x"ff115170",
   352 => x"fb38823d",
   353 => x"0d04803d",
   354 => x"0dbab808",
   355 => x"51870b84",
   356 => x"120c823d",
   357 => x"0d04803d",
   358 => x"0dbabc08",
   359 => x"51b60b8c",
   360 => x"120c830b",
   361 => x"88120c82",
   362 => x"3d0d04ff",
   363 => x"3d0dbabc",
   364 => x"08528412",
   365 => x"08708106",
   366 => x"51517080",
   367 => x"2ef43871",
   368 => x"087081ff",
   369 => x"06800c51",
   370 => x"833d0d04",
   371 => x"fe3d0d02",
   372 => x"930533ba",
   373 => x"bc085353",
   374 => x"84120870",
   375 => x"892a7081",
   376 => x"06515151",
   377 => x"70f23872",
   378 => x"720c843d",
   379 => x"0d04fe3d",
   380 => x"0d029305",
   381 => x"3353728a",
   382 => x"2e9b38ba",
   383 => x"bc085284",
   384 => x"12087089",
   385 => x"2a708106",
   386 => x"51515170",
   387 => x"f2387272",
   388 => x"0c843d0d",
   389 => x"04babc08",
   390 => x"52841208",
   391 => x"70892a70",
   392 => x"81065151",
   393 => x"5170f238",
   394 => x"8d720c84",
   395 => x"12087089",
   396 => x"2a708106",
   397 => x"51515170",
   398 => x"c638d339",
   399 => x"fd3d0d75",
   400 => x"70335254",
   401 => x"70802ea7",
   402 => x"3870babc",
   403 => x"08535381",
   404 => x"1454728a",
   405 => x"2e9d3884",
   406 => x"12087089",
   407 => x"2a708106",
   408 => x"51515170",
   409 => x"f2387272",
   410 => x"0c733353",
   411 => x"72e13885",
   412 => x"3d0d0484",
   413 => x"12087089",
   414 => x"2a708106",
   415 => x"51515170",
   416 => x"f2388d72",
   417 => x"0c841208",
   418 => x"70892a70",
   419 => x"81065151",
   420 => x"5170c438",
   421 => x"d139f53d",
   422 => x"0d7e0284",
   423 => x"05b70533",
   424 => x"8c3d5b55",
   425 => x"578b53b4",
   426 => x"f4527851",
   427 => x"a4973f82",
   428 => x"5673882e",
   429 => x"96388456",
   430 => x"73902e8f",
   431 => x"38885673",
   432 => x"a02e8838",
   433 => x"74567480",
   434 => x"2ea73802",
   435 => x"a5055876",
   436 => x"8f065473",
   437 => x"892680cb",
   438 => x"387518b0",
   439 => x"15555573",
   440 => x"75347684",
   441 => x"2aff1770",
   442 => x"81ff0658",
   443 => x"555775df",
   444 => x"38787933",
   445 => x"55577380",
   446 => x"2ea53873",
   447 => x"babc0856",
   448 => x"56811757",
   449 => x"758a2eb7",
   450 => x"38841508",
   451 => x"70892a81",
   452 => x"06595477",
   453 => x"f4387575",
   454 => x"0c763356",
   455 => x"75e3388d",
   456 => x"3d0d0475",
   457 => x"18b71555",
   458 => x"55737534",
   459 => x"76842aff",
   460 => x"177081ff",
   461 => x"06585557",
   462 => x"75ff9438",
   463 => x"ffb33984",
   464 => x"15087089",
   465 => x"2a810659",
   466 => x"5477f438",
   467 => x"8d750c84",
   468 => x"15087089",
   469 => x"2a810659",
   470 => x"5477ffad",
   471 => x"38ffb739",
   472 => x"f83d0d7a",
   473 => x"7c595380",
   474 => x"73565776",
   475 => x"732480dc",
   476 => x"38771754",
   477 => x"8a527451",
   478 => x"9eaa3f80",
   479 => x"08b00553",
   480 => x"72743481",
   481 => x"17578a52",
   482 => x"74519df3",
   483 => x"3f800855",
   484 => x"8008de38",
   485 => x"8008779f",
   486 => x"2a187081",
   487 => x"2c5b5656",
   488 => x"8079259e",
   489 => x"387717ff",
   490 => x"05557518",
   491 => x"70335553",
   492 => x"74337334",
   493 => x"73753481",
   494 => x"16ff1656",
   495 => x"56787624",
   496 => x"e9387618",
   497 => x"56807634",
   498 => x"8a3d0d04",
   499 => x"ad787081",
   500 => x"055a3472",
   501 => x"30781855",
   502 => x"558a5274",
   503 => x"519dc53f",
   504 => x"8008b005",
   505 => x"53727434",
   506 => x"8117578a",
   507 => x"5274519d",
   508 => x"8e3f8008",
   509 => x"558008fe",
   510 => x"f838ff98",
   511 => x"39803d0d",
   512 => x"bab40851",
   513 => x"81ff0b88",
   514 => x"120c823d",
   515 => x"0d04fb3d",
   516 => x"0d8880e0",
   517 => x"870bbab4",
   518 => x"08bab808",
   519 => x"7284130c",
   520 => x"565755af",
   521 => x"d7c20b94",
   522 => x"150c850b",
   523 => x"98150c98",
   524 => x"14087081",
   525 => x"06515372",
   526 => x"f638749f",
   527 => x"2a751007",
   528 => x"7084180c",
   529 => x"55afd7c2",
   530 => x"0b94150c",
   531 => x"850b9815",
   532 => x"0cdd39fd",
   533 => x"3d0dbab4",
   534 => x"085480d5",
   535 => x"0b84150c",
   536 => x"babc0852",
   537 => x"84120881",
   538 => x"06517080",
   539 => x"2ef63871",
   540 => x"087081ff",
   541 => x"06f61152",
   542 => x"545170ae",
   543 => x"268b3870",
   544 => x"1010b788",
   545 => x"05517008",
   546 => x"04841208",
   547 => x"70892a70",
   548 => x"81065151",
   549 => x"5170f238",
   550 => x"ab720c72",
   551 => x"8a2ea638",
   552 => x"84120870",
   553 => x"892a7081",
   554 => x"06515151",
   555 => x"70f23872",
   556 => x"720c8412",
   557 => x"0870892a",
   558 => x"81065153",
   559 => x"72f438ad",
   560 => x"720cffa0",
   561 => x"39841208",
   562 => x"70892a70",
   563 => x"81065151",
   564 => x"5170f238",
   565 => x"8d720c84",
   566 => x"12087089",
   567 => x"2a708106",
   568 => x"51515170",
   569 => x"ffba38c7",
   570 => x"3981ff0b",
   571 => x"84150cfe",
   572 => x"f33980ff",
   573 => x"0b84150c",
   574 => x"feea39bf",
   575 => x"0b84150c",
   576 => x"fee2399f",
   577 => x"0b84150c",
   578 => x"feda398f",
   579 => x"0b84150c",
   580 => x"fed23987",
   581 => x"0b84150c",
   582 => x"feca3983",
   583 => x"0b84150c",
   584 => x"fec23981",
   585 => x"0b84150c",
   586 => x"feba3980",
   587 => x"0b84150c",
   588 => x"feb239ff",
   589 => x"3d0dbab4",
   590 => x"08527108",
   591 => x"708f0670",
   592 => x"71842b07",
   593 => x"84150c51",
   594 => x"51710870",
   595 => x"8f067071",
   596 => x"842b0784",
   597 => x"150c5151",
   598 => x"e139d53d",
   599 => x"0dbab008",
   600 => x"58ff0b84",
   601 => x"190cfdaa",
   602 => x"d50b8819",
   603 => x"0c85adaa",
   604 => x"d5aa0b8c",
   605 => x"190ca4b4",
   606 => x"0b94190c",
   607 => x"8186a10b",
   608 => x"98190cb5",
   609 => x"800bb580",
   610 => x"33555773",
   611 => x"802ea638",
   612 => x"73babc08",
   613 => x"56568117",
   614 => x"57758a2e",
   615 => x"8cfe3884",
   616 => x"15087089",
   617 => x"2a810651",
   618 => x"5978f438",
   619 => x"75750c76",
   620 => x"335675e2",
   621 => x"38b5940b",
   622 => x"b5943355",
   623 => x"5773802e",
   624 => x"a638babc",
   625 => x"08745755",
   626 => x"81175775",
   627 => x"8a2e8ced",
   628 => x"38841508",
   629 => x"70892a81",
   630 => x"06515978",
   631 => x"f4387575",
   632 => x"0c763356",
   633 => x"75e23877",
   634 => x"08a63d5a",
   635 => x"568b53b4",
   636 => x"f4527851",
   637 => x"9dcf3f88",
   638 => x"02840581",
   639 => x"91055957",
   640 => x"758f0654",
   641 => x"7389268c",
   642 => x"d5387618",
   643 => x"b0155555",
   644 => x"73753475",
   645 => x"842aff18",
   646 => x"7081ff06",
   647 => x"59565676",
   648 => x"df387879",
   649 => x"33555773",
   650 => x"802ea638",
   651 => x"babc0874",
   652 => x"57558117",
   653 => x"57758a2e",
   654 => x"8cc03884",
   655 => x"15087089",
   656 => x"2a810659",
   657 => x"5977f438",
   658 => x"75750c76",
   659 => x"335675e2",
   660 => x"38b5a40b",
   661 => x"b5a43355",
   662 => x"5773802e",
   663 => x"a638babc",
   664 => x"08745755",
   665 => x"81175775",
   666 => x"8a2e8caf",
   667 => x"38841508",
   668 => x"70892a81",
   669 => x"06595977",
   670 => x"f4387575",
   671 => x"0c763356",
   672 => x"75e238ba",
   673 => x"b0088411",
   674 => x"08a43d5b",
   675 => x"57578b53",
   676 => x"b4f45278",
   677 => x"519cae3f",
   678 => x"88028405",
   679 => x"81850559",
   680 => x"57758f06",
   681 => x"54738926",
   682 => x"918b3876",
   683 => x"18b01555",
   684 => x"55737534",
   685 => x"75842aff",
   686 => x"187081ff",
   687 => x"06595656",
   688 => x"76df3878",
   689 => x"79335557",
   690 => x"73802ea6",
   691 => x"38babc08",
   692 => x"74575581",
   693 => x"1757758a",
   694 => x"2e8be138",
   695 => x"84150870",
   696 => x"892a8106",
   697 => x"595977f4",
   698 => x"3875750c",
   699 => x"76335675",
   700 => x"e238b5b4",
   701 => x"0bb5b433",
   702 => x"55577380",
   703 => x"2ea638ba",
   704 => x"bc087457",
   705 => x"55811757",
   706 => x"758a2e8b",
   707 => x"d0388415",
   708 => x"0870892a",
   709 => x"81065959",
   710 => x"77f43875",
   711 => x"750c7633",
   712 => x"5675e238",
   713 => x"bab00888",
   714 => x"1108a13d",
   715 => x"5b57578b",
   716 => x"53b4f452",
   717 => x"78519b8d",
   718 => x"3f880284",
   719 => x"0580f905",
   720 => x"5957758f",
   721 => x"06547389",
   722 => x"268fe138",
   723 => x"7618b015",
   724 => x"55557375",
   725 => x"3475842a",
   726 => x"ff187081",
   727 => x"ff065956",
   728 => x"5676df38",
   729 => x"78793355",
   730 => x"5773802e",
   731 => x"a638babc",
   732 => x"08745755",
   733 => x"81175775",
   734 => x"8a2e8b82",
   735 => x"38841508",
   736 => x"70892a81",
   737 => x"06595977",
   738 => x"f4387575",
   739 => x"0c763356",
   740 => x"75e238b5",
   741 => x"c40bb5c4",
   742 => x"33555773",
   743 => x"802ea638",
   744 => x"babc0874",
   745 => x"57558117",
   746 => x"57758a2e",
   747 => x"8af13884",
   748 => x"15087089",
   749 => x"2a810659",
   750 => x"5977f438",
   751 => x"75750c76",
   752 => x"335675e2",
   753 => x"38bab008",
   754 => x"8c11089e",
   755 => x"3d5b5757",
   756 => x"8b53b4f4",
   757 => x"52785199",
   758 => x"ec3f8802",
   759 => x"840580ed",
   760 => x"05595775",
   761 => x"8f065473",
   762 => x"89268eb7",
   763 => x"387618b0",
   764 => x"15555573",
   765 => x"75347584",
   766 => x"2aff1870",
   767 => x"81ff0659",
   768 => x"565676df",
   769 => x"38787933",
   770 => x"55577380",
   771 => x"2ea638ba",
   772 => x"bc087457",
   773 => x"55811757",
   774 => x"758a2e8a",
   775 => x"a3388415",
   776 => x"0870892a",
   777 => x"81065959",
   778 => x"77f43875",
   779 => x"750c7633",
   780 => x"5675e238",
   781 => x"b5d40bb5",
   782 => x"d4335557",
   783 => x"73802ea6",
   784 => x"38babc08",
   785 => x"74575581",
   786 => x"1757758a",
   787 => x"2e8a9238",
   788 => x"84150870",
   789 => x"892a8106",
   790 => x"595977f4",
   791 => x"3875750c",
   792 => x"76335675",
   793 => x"e238bab0",
   794 => x"08901108",
   795 => x"9b3d5b57",
   796 => x"578b53b4",
   797 => x"f4527851",
   798 => x"98cb3f88",
   799 => x"02840580",
   800 => x"e1055957",
   801 => x"758f0654",
   802 => x"7389268d",
   803 => x"8d387618",
   804 => x"b0155555",
   805 => x"73753475",
   806 => x"842aff18",
   807 => x"7081ff06",
   808 => x"59565676",
   809 => x"df387879",
   810 => x"33555773",
   811 => x"802ea638",
   812 => x"babc0874",
   813 => x"57558117",
   814 => x"57758a2e",
   815 => x"89c43884",
   816 => x"15087089",
   817 => x"2a810659",
   818 => x"5977f438",
   819 => x"75750c76",
   820 => x"335675e2",
   821 => x"38b5e40b",
   822 => x"b5e43355",
   823 => x"5773802e",
   824 => x"a638babc",
   825 => x"08745755",
   826 => x"81175775",
   827 => x"8a2e89b3",
   828 => x"38841508",
   829 => x"70892a81",
   830 => x"06595977",
   831 => x"f4387575",
   832 => x"0c763356",
   833 => x"75e238ba",
   834 => x"b0089411",
   835 => x"08983d5b",
   836 => x"57578b53",
   837 => x"b4f45278",
   838 => x"5197aa3f",
   839 => x"88028405",
   840 => x"80d50559",
   841 => x"57758f06",
   842 => x"54738926",
   843 => x"8be33876",
   844 => x"18b01555",
   845 => x"55737534",
   846 => x"75842aff",
   847 => x"187081ff",
   848 => x"06595656",
   849 => x"76df3878",
   850 => x"79335557",
   851 => x"73802ea6",
   852 => x"38babc08",
   853 => x"74575581",
   854 => x"1757758a",
   855 => x"2e88e538",
   856 => x"84150870",
   857 => x"892a8106",
   858 => x"595977f4",
   859 => x"3875750c",
   860 => x"76335675",
   861 => x"e238b5f4",
   862 => x"0bb5f433",
   863 => x"55577380",
   864 => x"2ea638ba",
   865 => x"bc087457",
   866 => x"55811757",
   867 => x"758a2e88",
   868 => x"d4388415",
   869 => x"0870892a",
   870 => x"81065959",
   871 => x"77f43875",
   872 => x"750c7633",
   873 => x"5675e238",
   874 => x"bab00898",
   875 => x"1108953d",
   876 => x"5b57578b",
   877 => x"53b4f452",
   878 => x"78519689",
   879 => x"3f880284",
   880 => x"0580c905",
   881 => x"5957758f",
   882 => x"06547389",
   883 => x"268ab938",
   884 => x"7618b015",
   885 => x"55557375",
   886 => x"3475842a",
   887 => x"ff187081",
   888 => x"ff065956",
   889 => x"5676df38",
   890 => x"78793355",
   891 => x"5773802e",
   892 => x"a638babc",
   893 => x"08745755",
   894 => x"81175775",
   895 => x"8a2e8886",
   896 => x"38841508",
   897 => x"70892a81",
   898 => x"06595977",
   899 => x"f4387575",
   900 => x"0c763356",
   901 => x"75e238b6",
   902 => x"840bb684",
   903 => x"33555773",
   904 => x"802ea638",
   905 => x"babc0874",
   906 => x"57558117",
   907 => x"57758a2e",
   908 => x"87f53884",
   909 => x"15087089",
   910 => x"2a810659",
   911 => x"5977f438",
   912 => x"75750c76",
   913 => x"335675e2",
   914 => x"38bab008",
   915 => x"9c110892",
   916 => x"3d5b5757",
   917 => x"8b53b4f4",
   918 => x"52785194",
   919 => x"e83f8802",
   920 => x"8405bd05",
   921 => x"5957758f",
   922 => x"06547389",
   923 => x"26899038",
   924 => x"7618b015",
   925 => x"55557375",
   926 => x"3475842a",
   927 => x"ff187081",
   928 => x"ff065956",
   929 => x"5676df38",
   930 => x"78793355",
   931 => x"5773802e",
   932 => x"a638babc",
   933 => x"08745755",
   934 => x"81175775",
   935 => x"8a2e87a8",
   936 => x"38841508",
   937 => x"70892a81",
   938 => x"06595977",
   939 => x"f4387575",
   940 => x"0c763356",
   941 => x"75e238b6",
   942 => x"940bb694",
   943 => x"33555773",
   944 => x"802ea638",
   945 => x"babc0874",
   946 => x"57558117",
   947 => x"57758a2e",
   948 => x"87973884",
   949 => x"15087089",
   950 => x"2a810659",
   951 => x"5977f438",
   952 => x"75750c76",
   953 => x"335675e2",
   954 => x"38bab008",
   955 => x"a011088f",
   956 => x"3d5b5757",
   957 => x"8b53b4f4",
   958 => x"52785193",
   959 => x"c83f8802",
   960 => x"8405b105",
   961 => x"5957758f",
   962 => x"06547389",
   963 => x"2687e738",
   964 => x"7618b015",
   965 => x"55557375",
   966 => x"3475842a",
   967 => x"ff187081",
   968 => x"ff065956",
   969 => x"5676df38",
   970 => x"78793355",
   971 => x"5773802e",
   972 => x"a638babc",
   973 => x"08745755",
   974 => x"81175775",
   975 => x"8a2e86ca",
   976 => x"38841508",
   977 => x"70892a81",
   978 => x"06595977",
   979 => x"f4387575",
   980 => x"0c763356",
   981 => x"75e238b6",
   982 => x"a40bb6a4",
   983 => x"33555773",
   984 => x"802ea638",
   985 => x"babc0874",
   986 => x"57558117",
   987 => x"57758a2e",
   988 => x"86b93884",
   989 => x"15087089",
   990 => x"2a810659",
   991 => x"5977f438",
   992 => x"75750c76",
   993 => x"335675e2",
   994 => x"38bab008",
   995 => x"a411088c",
   996 => x"3d5b5757",
   997 => x"8b53b4f4",
   998 => x"52785192",
   999 => x"a83f8802",
  1000 => x"8405a505",
  1001 => x"5957758f",
  1002 => x"06547389",
  1003 => x"2686be38",
  1004 => x"7618b015",
  1005 => x"55557375",
  1006 => x"3475842a",
  1007 => x"ff187081",
  1008 => x"ff065956",
  1009 => x"5676df38",
  1010 => x"78793355",
  1011 => x"5773802e",
  1012 => x"86ec38ba",
  1013 => x"bc087457",
  1014 => x"55811757",
  1015 => x"758a2e85",
  1016 => x"eb388415",
  1017 => x"0870892a",
  1018 => x"81065959",
  1019 => x"77f43875",
  1020 => x"750c7633",
  1021 => x"5675e238",
  1022 => x"84150870",
  1023 => x"892a8106",
  1024 => x"575875f4",
  1025 => x"388d750c",
  1026 => x"84150870",
  1027 => x"892a8106",
  1028 => x"555673f4",
  1029 => x"388a750c",
  1030 => x"ad3d0d04",
  1031 => x"84150870",
  1032 => x"892a8106",
  1033 => x"515473f4",
  1034 => x"388d750c",
  1035 => x"84150870",
  1036 => x"892a8106",
  1037 => x"515978f2",
  1038 => x"e638f2f0",
  1039 => x"39841508",
  1040 => x"70892a81",
  1041 => x"06515473",
  1042 => x"f4388d75",
  1043 => x"0c841508",
  1044 => x"70892a81",
  1045 => x"06515978",
  1046 => x"f2f738f3",
  1047 => x"81397618",
  1048 => x"b7155555",
  1049 => x"73753475",
  1050 => x"842aff18",
  1051 => x"7081ff06",
  1052 => x"59565676",
  1053 => x"f38a38f3",
  1054 => x"a9398415",
  1055 => x"0870892a",
  1056 => x"81065959",
  1057 => x"77f4388d",
  1058 => x"750c8415",
  1059 => x"0870892a",
  1060 => x"81065959",
  1061 => x"77f3a438",
  1062 => x"f3ae3984",
  1063 => x"15087089",
  1064 => x"2a810659",
  1065 => x"5977f438",
  1066 => x"8d750c84",
  1067 => x"15087089",
  1068 => x"2a810659",
  1069 => x"5977f3b5",
  1070 => x"38f3bf39",
  1071 => x"84150870",
  1072 => x"892a8106",
  1073 => x"595977f4",
  1074 => x"388d750c",
  1075 => x"84150870",
  1076 => x"892a8106",
  1077 => x"595977f4",
  1078 => x"8338f48d",
  1079 => x"39841508",
  1080 => x"70892a81",
  1081 => x"06595977",
  1082 => x"f4388d75",
  1083 => x"0c841508",
  1084 => x"70892a81",
  1085 => x"06595977",
  1086 => x"f49438f4",
  1087 => x"9e398415",
  1088 => x"0870892a",
  1089 => x"81065959",
  1090 => x"77f4388d",
  1091 => x"750c8415",
  1092 => x"0870892a",
  1093 => x"81065959",
  1094 => x"77f4e238",
  1095 => x"f4ec3984",
  1096 => x"15087089",
  1097 => x"2a810659",
  1098 => x"5977f438",
  1099 => x"8d750c84",
  1100 => x"15087089",
  1101 => x"2a810659",
  1102 => x"5977f4f3",
  1103 => x"38f4fd39",
  1104 => x"84150870",
  1105 => x"892a8106",
  1106 => x"595977f4",
  1107 => x"388d750c",
  1108 => x"84150870",
  1109 => x"892a8106",
  1110 => x"595977f5",
  1111 => x"c138f5cb",
  1112 => x"39841508",
  1113 => x"70892a81",
  1114 => x"06595977",
  1115 => x"f4388d75",
  1116 => x"0c841508",
  1117 => x"70892a81",
  1118 => x"06595977",
  1119 => x"f5d238f5",
  1120 => x"dc398415",
  1121 => x"0870892a",
  1122 => x"81065959",
  1123 => x"77f4388d",
  1124 => x"750c8415",
  1125 => x"0870892a",
  1126 => x"81065959",
  1127 => x"77f6a038",
  1128 => x"f6aa3984",
  1129 => x"15087089",
  1130 => x"2a810659",
  1131 => x"5977f438",
  1132 => x"8d750c84",
  1133 => x"15087089",
  1134 => x"2a810659",
  1135 => x"5977f6b1",
  1136 => x"38f6bb39",
  1137 => x"84150870",
  1138 => x"892a8106",
  1139 => x"595977f4",
  1140 => x"388d750c",
  1141 => x"84150870",
  1142 => x"892a8106",
  1143 => x"595977f6",
  1144 => x"ff38f789",
  1145 => x"39841508",
  1146 => x"70892a81",
  1147 => x"06595977",
  1148 => x"f4388d75",
  1149 => x"0c841508",
  1150 => x"70892a81",
  1151 => x"06595977",
  1152 => x"f79038f7",
  1153 => x"9a398415",
  1154 => x"0870892a",
  1155 => x"81065959",
  1156 => x"77f4388d",
  1157 => x"750c8415",
  1158 => x"0870892a",
  1159 => x"81065959",
  1160 => x"77f7de38",
  1161 => x"f7e83984",
  1162 => x"15087089",
  1163 => x"2a810659",
  1164 => x"5977f438",
  1165 => x"8d750c84",
  1166 => x"15087089",
  1167 => x"2a810659",
  1168 => x"5977f7ef",
  1169 => x"38f7f939",
  1170 => x"84150870",
  1171 => x"892a8106",
  1172 => x"595977f4",
  1173 => x"388d750c",
  1174 => x"84150870",
  1175 => x"892a8106",
  1176 => x"595977f8",
  1177 => x"bc38f8c6",
  1178 => x"39841508",
  1179 => x"70892a81",
  1180 => x"06595977",
  1181 => x"f4388d75",
  1182 => x"0c841508",
  1183 => x"70892a81",
  1184 => x"06595977",
  1185 => x"f8cd38f8",
  1186 => x"d7398415",
  1187 => x"0870892a",
  1188 => x"81065959",
  1189 => x"77f4388d",
  1190 => x"750c8415",
  1191 => x"0870892a",
  1192 => x"81065959",
  1193 => x"77f99a38",
  1194 => x"f9a43984",
  1195 => x"15087089",
  1196 => x"2a810659",
  1197 => x"5977f438",
  1198 => x"8d750c84",
  1199 => x"15087089",
  1200 => x"2a810659",
  1201 => x"5977f9ab",
  1202 => x"38f9b539",
  1203 => x"84150870",
  1204 => x"892a8106",
  1205 => x"595977f4",
  1206 => x"388d750c",
  1207 => x"84150870",
  1208 => x"892a8106",
  1209 => x"595977f9",
  1210 => x"f938fa83",
  1211 => x"397618b7",
  1212 => x"155555f9",
  1213 => x"c1397618",
  1214 => x"b7155555",
  1215 => x"f8983976",
  1216 => x"18b71555",
  1217 => x"55f6ef39",
  1218 => x"7618b715",
  1219 => x"5555f5c6",
  1220 => x"397618b7",
  1221 => x"155555f4",
  1222 => x"9c397618",
  1223 => x"b7155555",
  1224 => x"f2f23976",
  1225 => x"18b71555",
  1226 => x"55f1c839",
  1227 => x"7618b715",
  1228 => x"5555f09e",
  1229 => x"397618b7",
  1230 => x"155555ee",
  1231 => x"f439babc",
  1232 => x"08841108",
  1233 => x"70892a81",
  1234 => x"06585955",
  1235 => x"75f9a938",
  1236 => x"f9b33980",
  1237 => x"3d0dbab0",
  1238 => x"08519171",
  1239 => x"0cff39fc",
  1240 => x"3d0d029a",
  1241 => x"05220284",
  1242 => x"059e0522",
  1243 => x"028805a2",
  1244 => x"0522bab0",
  1245 => x"08555654",
  1246 => x"55901208",
  1247 => x"70832a70",
  1248 => x"81065151",
  1249 => x"5170f238",
  1250 => x"74902b73",
  1251 => x"8b2b0774",
  1252 => x"862b0781",
  1253 => x"0790130c",
  1254 => x"863d0d04",
  1255 => x"fd3d0d02",
  1256 => x"96052202",
  1257 => x"84059a05",
  1258 => x"22bab008",
  1259 => x"54545490",
  1260 => x"12087083",
  1261 => x"2a708106",
  1262 => x"51515170",
  1263 => x"f238738b",
  1264 => x"2b73862b",
  1265 => x"07820790",
  1266 => x"130c9012",
  1267 => x"0870902a",
  1268 => x"800c5385",
  1269 => x"3d0d04fa",
  1270 => x"3d0dbab4",
  1271 => x"08700881",
  1272 => x"0a06bab8",
  1273 => x"08555855",
  1274 => x"870b8414",
  1275 => x"0cbabc08",
  1276 => x"54b60b8c",
  1277 => x"150c830b",
  1278 => x"88150cb6",
  1279 => x"b40bb6b4",
  1280 => x"33545672",
  1281 => x"802ea438",
  1282 => x"72558116",
  1283 => x"56748a2e",
  1284 => x"81e23884",
  1285 => x"14087089",
  1286 => x"2a708106",
  1287 => x"51515372",
  1288 => x"f2387474",
  1289 => x"0c753355",
  1290 => x"74e038b6",
  1291 => x"b80bb6b8",
  1292 => x"33545672",
  1293 => x"802ea438",
  1294 => x"72558116",
  1295 => x"56748a2e",
  1296 => x"81d73884",
  1297 => x"14087089",
  1298 => x"2a708106",
  1299 => x"51515372",
  1300 => x"f2387474",
  1301 => x"0c753355",
  1302 => x"74e03876",
  1303 => x"802e82d9",
  1304 => x"38b6c40b",
  1305 => x"b6c43354",
  1306 => x"5672802e",
  1307 => x"a2387255",
  1308 => x"81165674",
  1309 => x"8a2e81c6",
  1310 => x"38841408",
  1311 => x"70892a81",
  1312 => x"06515372",
  1313 => x"f4387474",
  1314 => x"0c753355",
  1315 => x"74e238b6",
  1316 => x"d40bb6d4",
  1317 => x"33545672",
  1318 => x"802ea238",
  1319 => x"72558116",
  1320 => x"56748a2e",
  1321 => x"81b93884",
  1322 => x"14087089",
  1323 => x"2a810651",
  1324 => x"5372f438",
  1325 => x"74740c75",
  1326 => x"335574e2",
  1327 => x"38e99b3f",
  1328 => x"bab40856",
  1329 => x"80d50b84",
  1330 => x"170cbabc",
  1331 => x"08548414",
  1332 => x"08810655",
  1333 => x"74802ef6",
  1334 => x"38730870",
  1335 => x"81ff06f6",
  1336 => x"11525653",
  1337 => x"72ae2681",
  1338 => x"97387210",
  1339 => x"10b8c405",
  1340 => x"57760804",
  1341 => x"84140870",
  1342 => x"892a7081",
  1343 => x"06515153",
  1344 => x"72f2388d",
  1345 => x"740c8414",
  1346 => x"0870892a",
  1347 => x"70810651",
  1348 => x"515372fd",
  1349 => x"fe38fe8a",
  1350 => x"39841408",
  1351 => x"70892a70",
  1352 => x"81065151",
  1353 => x"5372f238",
  1354 => x"8d740c84",
  1355 => x"14087089",
  1356 => x"2a708106",
  1357 => x"51515372",
  1358 => x"fe8938fe",
  1359 => x"95398414",
  1360 => x"0870892a",
  1361 => x"81065157",
  1362 => x"76f4388d",
  1363 => x"740c8414",
  1364 => x"0870892a",
  1365 => x"81065153",
  1366 => x"72fe9e38",
  1367 => x"fea83984",
  1368 => x"14087089",
  1369 => x"2a810651",
  1370 => x"5776f438",
  1371 => x"8d740c84",
  1372 => x"14087089",
  1373 => x"2a810651",
  1374 => x"5372feab",
  1375 => x"38feb539",
  1376 => x"84140870",
  1377 => x"892a8106",
  1378 => x"515372f4",
  1379 => x"38ab740c",
  1380 => x"748a2e80",
  1381 => x"ff388414",
  1382 => x"0870892a",
  1383 => x"81065153",
  1384 => x"72f43874",
  1385 => x"740c8414",
  1386 => x"0870892a",
  1387 => x"81065653",
  1388 => x"74f438ad",
  1389 => x"740cfe96",
  1390 => x"39b6f80b",
  1391 => x"b6f83354",
  1392 => x"5672802e",
  1393 => x"fdc93872",
  1394 => x"81175755",
  1395 => x"748a2ea5",
  1396 => x"38841408",
  1397 => x"70892a81",
  1398 => x"06515372",
  1399 => x"f4387474",
  1400 => x"0c753355",
  1401 => x"74802efd",
  1402 => x"a6388116",
  1403 => x"56748a2e",
  1404 => x"098106dd",
  1405 => x"38841408",
  1406 => x"70892a81",
  1407 => x"06515776",
  1408 => x"f4388d74",
  1409 => x"0c841408",
  1410 => x"70892a81",
  1411 => x"06515372",
  1412 => x"c038cb39",
  1413 => x"84140870",
  1414 => x"892a8106",
  1415 => x"515776f4",
  1416 => x"388d740c",
  1417 => x"84140870",
  1418 => x"892a8106",
  1419 => x"515372fe",
  1420 => x"e538feef",
  1421 => x"3981ff0b",
  1422 => x"84170cfd",
  1423 => x"913980ff",
  1424 => x"0b84170c",
  1425 => x"fd8839bf",
  1426 => x"0b84170c",
  1427 => x"fd80399f",
  1428 => x"0b84170c",
  1429 => x"fcf8398f",
  1430 => x"0b84170c",
  1431 => x"fcf03987",
  1432 => x"0b84170c",
  1433 => x"fce83983",
  1434 => x"0b84170c",
  1435 => x"fce03981",
  1436 => x"0b84170c",
  1437 => x"fcd83980",
  1438 => x"0b84170c",
  1439 => x"fcd0398c",
  1440 => x"08028c0c",
  1441 => x"fd3d0d80",
  1442 => x"538c088c",
  1443 => x"0508528c",
  1444 => x"08880508",
  1445 => x"5182de3f",
  1446 => x"80087080",
  1447 => x"0c54853d",
  1448 => x"0d8c0c04",
  1449 => x"8c08028c",
  1450 => x"0cfd3d0d",
  1451 => x"81538c08",
  1452 => x"8c050852",
  1453 => x"8c088805",
  1454 => x"085182b9",
  1455 => x"3f800870",
  1456 => x"800c5485",
  1457 => x"3d0d8c0c",
  1458 => x"048c0802",
  1459 => x"8c0cf93d",
  1460 => x"0d800b8c",
  1461 => x"08fc050c",
  1462 => x"8c088805",
  1463 => x"088025ab",
  1464 => x"388c0888",
  1465 => x"0508308c",
  1466 => x"0888050c",
  1467 => x"800b8c08",
  1468 => x"f4050c8c",
  1469 => x"08fc0508",
  1470 => x"8838810b",
  1471 => x"8c08f405",
  1472 => x"0c8c08f4",
  1473 => x"05088c08",
  1474 => x"fc050c8c",
  1475 => x"088c0508",
  1476 => x"8025ab38",
  1477 => x"8c088c05",
  1478 => x"08308c08",
  1479 => x"8c050c80",
  1480 => x"0b8c08f0",
  1481 => x"050c8c08",
  1482 => x"fc050888",
  1483 => x"38810b8c",
  1484 => x"08f0050c",
  1485 => x"8c08f005",
  1486 => x"088c08fc",
  1487 => x"050c8053",
  1488 => x"8c088c05",
  1489 => x"08528c08",
  1490 => x"88050851",
  1491 => x"81a73f80",
  1492 => x"08708c08",
  1493 => x"f8050c54",
  1494 => x"8c08fc05",
  1495 => x"08802e8c",
  1496 => x"388c08f8",
  1497 => x"0508308c",
  1498 => x"08f8050c",
  1499 => x"8c08f805",
  1500 => x"0870800c",
  1501 => x"54893d0d",
  1502 => x"8c0c048c",
  1503 => x"08028c0c",
  1504 => x"fb3d0d80",
  1505 => x"0b8c08fc",
  1506 => x"050c8c08",
  1507 => x"88050880",
  1508 => x"2593388c",
  1509 => x"08880508",
  1510 => x"308c0888",
  1511 => x"050c810b",
  1512 => x"8c08fc05",
  1513 => x"0c8c088c",
  1514 => x"05088025",
  1515 => x"8c388c08",
  1516 => x"8c050830",
  1517 => x"8c088c05",
  1518 => x"0c81538c",
  1519 => x"088c0508",
  1520 => x"528c0888",
  1521 => x"050851ad",
  1522 => x"3f800870",
  1523 => x"8c08f805",
  1524 => x"0c548c08",
  1525 => x"fc050880",
  1526 => x"2e8c388c",
  1527 => x"08f80508",
  1528 => x"308c08f8",
  1529 => x"050c8c08",
  1530 => x"f8050870",
  1531 => x"800c5487",
  1532 => x"3d0d8c0c",
  1533 => x"048c0802",
  1534 => x"8c0cfd3d",
  1535 => x"0d810b8c",
  1536 => x"08fc050c",
  1537 => x"800b8c08",
  1538 => x"f8050c8c",
  1539 => x"088c0508",
  1540 => x"8c088805",
  1541 => x"0827ac38",
  1542 => x"8c08fc05",
  1543 => x"08802ea3",
  1544 => x"38800b8c",
  1545 => x"088c0508",
  1546 => x"2499388c",
  1547 => x"088c0508",
  1548 => x"108c088c",
  1549 => x"050c8c08",
  1550 => x"fc050810",
  1551 => x"8c08fc05",
  1552 => x"0cc9398c",
  1553 => x"08fc0508",
  1554 => x"802e80c9",
  1555 => x"388c088c",
  1556 => x"05088c08",
  1557 => x"88050826",
  1558 => x"a1388c08",
  1559 => x"8805088c",
  1560 => x"088c0508",
  1561 => x"318c0888",
  1562 => x"050c8c08",
  1563 => x"f805088c",
  1564 => x"08fc0508",
  1565 => x"078c08f8",
  1566 => x"050c8c08",
  1567 => x"fc050881",
  1568 => x"2a8c08fc",
  1569 => x"050c8c08",
  1570 => x"8c050881",
  1571 => x"2a8c088c",
  1572 => x"050cffaf",
  1573 => x"398c0890",
  1574 => x"0508802e",
  1575 => x"8f388c08",
  1576 => x"88050870",
  1577 => x"8c08f405",
  1578 => x"0c518d39",
  1579 => x"8c08f805",
  1580 => x"08708c08",
  1581 => x"f4050c51",
  1582 => x"8c08f405",
  1583 => x"08800c85",
  1584 => x"3d0d8c0c",
  1585 => x"04fc3d0d",
  1586 => x"7670797b",
  1587 => x"55555555",
  1588 => x"8f72278c",
  1589 => x"38727507",
  1590 => x"83065170",
  1591 => x"802ea738",
  1592 => x"ff125271",
  1593 => x"ff2e9838",
  1594 => x"72708105",
  1595 => x"54337470",
  1596 => x"81055634",
  1597 => x"ff125271",
  1598 => x"ff2e0981",
  1599 => x"06ea3874",
  1600 => x"800c863d",
  1601 => x"0d047451",
  1602 => x"72708405",
  1603 => x"54087170",
  1604 => x"8405530c",
  1605 => x"72708405",
  1606 => x"54087170",
  1607 => x"8405530c",
  1608 => x"72708405",
  1609 => x"54087170",
  1610 => x"8405530c",
  1611 => x"72708405",
  1612 => x"54087170",
  1613 => x"8405530c",
  1614 => x"f0125271",
  1615 => x"8f26c938",
  1616 => x"83722795",
  1617 => x"38727084",
  1618 => x"05540871",
  1619 => x"70840553",
  1620 => x"0cfc1252",
  1621 => x"718326ed",
  1622 => x"387054ff",
  1623 => x"8339fd3d",
  1624 => x"0d800bba",
  1625 => x"a4085454",
  1626 => x"72812e99",
  1627 => x"387380c1",
  1628 => x"e80cd5eb",
  1629 => x"3fd5893f",
  1630 => x"bac05281",
  1631 => x"51f4d83f",
  1632 => x"8008519f",
  1633 => x"3f7280c1",
  1634 => x"e80cd5d3",
  1635 => x"3fd4f13f",
  1636 => x"bac05281",
  1637 => x"51f4c03f",
  1638 => x"80085187",
  1639 => x"3f00ff39",
  1640 => x"00ff39f7",
  1641 => x"3d0d7bba",
  1642 => x"c40882c8",
  1643 => x"11085a54",
  1644 => x"5a77802e",
  1645 => x"80d93881",
  1646 => x"88188419",
  1647 => x"08ff0581",
  1648 => x"712b5955",
  1649 => x"59807424",
  1650 => x"80e93880",
  1651 => x"7424b538",
  1652 => x"73822b78",
  1653 => x"11880556",
  1654 => x"56818019",
  1655 => x"08770653",
  1656 => x"72802eb5",
  1657 => x"38781670",
  1658 => x"08535379",
  1659 => x"51740853",
  1660 => x"722dff14",
  1661 => x"fc17fc17",
  1662 => x"79812c5a",
  1663 => x"57575473",
  1664 => x"8025d638",
  1665 => x"77085877",
  1666 => x"ffad38ba",
  1667 => x"c40853bc",
  1668 => x"1308a538",
  1669 => x"7951ff85",
  1670 => x"3f740853",
  1671 => x"722dff14",
  1672 => x"fc17fc17",
  1673 => x"79812c5a",
  1674 => x"57575473",
  1675 => x"8025ffa9",
  1676 => x"38d23980",
  1677 => x"57ff9439",
  1678 => x"7251bc13",
  1679 => x"0853722d",
  1680 => x"7951fed9",
  1681 => x"3fff3d0d",
  1682 => x"80c1c80b",
  1683 => x"fc057008",
  1684 => x"525270ff",
  1685 => x"2e913870",
  1686 => x"2dfc1270",
  1687 => x"08525270",
  1688 => x"ff2e0981",
  1689 => x"06f13883",
  1690 => x"3d0d0404",
  1691 => x"d4dc3f04",
  1692 => x"00000040",
  1693 => x"30782020",
  1694 => x"20202020",
  1695 => x"20200000",
  1696 => x"0a677265",
  1697 => x"74682072",
  1698 => x"65676973",
  1699 => x"74657273",
  1700 => x"3a000000",
  1701 => x"0a636f6e",
  1702 => x"74726f6c",
  1703 => x"3a202020",
  1704 => x"20202000",
  1705 => x"0a737461",
  1706 => x"7475733a",
  1707 => x"20202020",
  1708 => x"20202000",
  1709 => x"0a6d6163",
  1710 => x"5f6d7362",
  1711 => x"3a202020",
  1712 => x"20202000",
  1713 => x"0a6d6163",
  1714 => x"5f6c7362",
  1715 => x"3a202020",
  1716 => x"20202000",
  1717 => x"0a6d6469",
  1718 => x"6f5f636f",
  1719 => x"6e74726f",
  1720 => x"6c3a2000",
  1721 => x"0a74785f",
  1722 => x"706f696e",
  1723 => x"7465723a",
  1724 => x"20202000",
  1725 => x"0a72785f",
  1726 => x"706f696e",
  1727 => x"7465723a",
  1728 => x"20202000",
  1729 => x"0a656463",
  1730 => x"6c5f6970",
  1731 => x"3a202020",
  1732 => x"20202000",
  1733 => x"0a686173",
  1734 => x"685f6d73",
  1735 => x"623a2020",
  1736 => x"20202000",
  1737 => x"0a686173",
  1738 => x"685f6c73",
  1739 => x"623a2020",
  1740 => x"20202000",
  1741 => x"0a0a0000",
  1742 => x"5a505520",
  1743 => x"74657374",
  1744 => x"20000000",
  1745 => x"286f6e20",
  1746 => x"73696d75",
  1747 => x"6c61746f",
  1748 => x"72290a00",
  1749 => x"636f6d70",
  1750 => x"696c6564",
  1751 => x"3a204175",
  1752 => x"67202036",
  1753 => x"20323031",
  1754 => x"30202031",
  1755 => x"363a3036",
  1756 => x"3a30320a",
  1757 => x"00000000",
  1758 => x"286f6e20",
  1759 => x"68617264",
  1760 => x"77617265",
  1761 => x"290a0000",
  1762 => x"00000864",
  1763 => x"00000889",
  1764 => x"00000889",
  1765 => x"00000864",
  1766 => x"00000889",
  1767 => x"00000889",
  1768 => x"00000889",
  1769 => x"00000889",
  1770 => x"00000889",
  1771 => x"00000889",
  1772 => x"00000889",
  1773 => x"00000889",
  1774 => x"00000889",
  1775 => x"00000889",
  1776 => x"00000889",
  1777 => x"00000889",
  1778 => x"00000889",
  1779 => x"00000889",
  1780 => x"00000889",
  1781 => x"00000889",
  1782 => x"00000889",
  1783 => x"00000889",
  1784 => x"00000889",
  1785 => x"00000889",
  1786 => x"00000889",
  1787 => x"00000889",
  1788 => x"00000889",
  1789 => x"00000889",
  1790 => x"00000889",
  1791 => x"00000889",
  1792 => x"00000889",
  1793 => x"00000889",
  1794 => x"00000889",
  1795 => x"00000889",
  1796 => x"00000889",
  1797 => x"00000889",
  1798 => x"00000889",
  1799 => x"00000889",
  1800 => x"0000092b",
  1801 => x"00000923",
  1802 => x"0000091b",
  1803 => x"00000913",
  1804 => x"0000090b",
  1805 => x"00000903",
  1806 => x"000008fb",
  1807 => x"000008f2",
  1808 => x"000008e9",
  1809 => x"000014ce",
  1810 => x"00001580",
  1811 => x"00001580",
  1812 => x"000014ce",
  1813 => x"00001580",
  1814 => x"00001580",
  1815 => x"00001580",
  1816 => x"00001580",
  1817 => x"00001580",
  1818 => x"00001580",
  1819 => x"00001580",
  1820 => x"00001580",
  1821 => x"00001580",
  1822 => x"00001580",
  1823 => x"00001580",
  1824 => x"00001580",
  1825 => x"00001580",
  1826 => x"00001580",
  1827 => x"00001580",
  1828 => x"00001580",
  1829 => x"00001580",
  1830 => x"00001580",
  1831 => x"00001580",
  1832 => x"00001580",
  1833 => x"00001580",
  1834 => x"00001580",
  1835 => x"00001580",
  1836 => x"00001580",
  1837 => x"00001580",
  1838 => x"00001580",
  1839 => x"00001580",
  1840 => x"00001580",
  1841 => x"00001580",
  1842 => x"00001580",
  1843 => x"00001580",
  1844 => x"00001580",
  1845 => x"00001580",
  1846 => x"00001580",
  1847 => x"00001677",
  1848 => x"0000166f",
  1849 => x"00001667",
  1850 => x"0000165f",
  1851 => x"00001657",
  1852 => x"0000164f",
  1853 => x"00001647",
  1854 => x"0000163e",
  1855 => x"00001635",
  1856 => x"64756d6d",
  1857 => x"792e6578",
  1858 => x"65000000",
  1859 => x"43000000",
  1860 => x"00ffffff",
  1861 => x"ff00ffff",
  1862 => x"ffff00ff",
  1863 => x"ffffff00",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"00000000",
  1867 => x"000020d0",
  1868 => x"80000c00",
  1869 => x"80000800",
  1870 => x"80000200",
  1871 => x"80000100",
  1872 => x"00001d00",
  1873 => x"00001d48",
  1874 => x"00000000",
  1875 => x"00001fb0",
  1876 => x"0000200c",
  1877 => x"00002068",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00000000",
  1887 => x"00001d0c",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000001",
  1917 => x"330eabcd",
  1918 => x"1234e66d",
  1919 => x"deec0005",
  1920 => x"000b0000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000000",
  1928 => x"00000000",
  1929 => x"00000000",
  1930 => x"00000000",
  1931 => x"00000000",
  1932 => x"00000000",
  1933 => x"00000000",
  1934 => x"00000000",
  1935 => x"00000000",
  1936 => x"00000000",
  1937 => x"00000000",
  1938 => x"00000000",
  1939 => x"00000000",
  1940 => x"00000000",
  1941 => x"00000000",
  1942 => x"00000000",
  1943 => x"00000000",
  1944 => x"00000000",
  1945 => x"00000000",
  1946 => x"00000000",
  1947 => x"00000000",
  1948 => x"00000000",
  1949 => x"00000000",
  1950 => x"00000000",
  1951 => x"00000000",
  1952 => x"00000000",
  1953 => x"00000000",
  1954 => x"00000000",
  1955 => x"00000000",
  1956 => x"00000000",
  1957 => x"00000000",
  1958 => x"00000000",
  1959 => x"00000000",
  1960 => x"00000000",
  1961 => x"00000000",
  1962 => x"00000000",
  1963 => x"00000000",
  1964 => x"00000000",
  1965 => x"00000000",
  1966 => x"00000000",
  1967 => x"00000000",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00000000",
  1972 => x"00000000",
  1973 => x"00000000",
  1974 => x"00000000",
  1975 => x"00000000",
  1976 => x"00000000",
  1977 => x"00000000",
  1978 => x"00000000",
  1979 => x"00000000",
  1980 => x"00000000",
  1981 => x"00000000",
  1982 => x"00000000",
  1983 => x"00000000",
  1984 => x"00000000",
  1985 => x"00000000",
  1986 => x"00000000",
  1987 => x"00000000",
  1988 => x"00000000",
  1989 => x"00000000",
  1990 => x"00000000",
  1991 => x"00000000",
  1992 => x"00000000",
  1993 => x"00000000",
  1994 => x"00000000",
  1995 => x"00000000",
  1996 => x"00000000",
  1997 => x"00000000",
  1998 => x"00000000",
  1999 => x"00000000",
  2000 => x"00000000",
  2001 => x"00000000",
  2002 => x"00000000",
  2003 => x"00000000",
  2004 => x"00000000",
  2005 => x"00000000",
  2006 => x"00000000",
  2007 => x"00000000",
  2008 => x"00000000",
  2009 => x"00000000",
  2010 => x"00000000",
  2011 => x"00000000",
  2012 => x"00000000",
  2013 => x"00000000",
  2014 => x"00000000",
  2015 => x"00000000",
  2016 => x"00000000",
  2017 => x"00000000",
  2018 => x"00000000",
  2019 => x"00000000",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"00000000",
  2023 => x"00000000",
  2024 => x"00000000",
  2025 => x"00000000",
  2026 => x"00000000",
  2027 => x"00000000",
  2028 => x"00000000",
  2029 => x"00000000",
  2030 => x"00000000",
  2031 => x"00000000",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"00000000",
  2035 => x"00000000",
  2036 => x"00000000",
  2037 => x"00000000",
  2038 => x"00000000",
  2039 => x"00000000",
  2040 => x"00000000",
  2041 => x"00000000",
  2042 => x"00000000",
  2043 => x"00000000",
  2044 => x"00000000",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"00000000",
  2048 => x"00000000",
  2049 => x"00000000",
  2050 => x"00000000",
  2051 => x"00000000",
  2052 => x"00000000",
  2053 => x"00000000",
  2054 => x"00000000",
  2055 => x"00000000",
  2056 => x"00000000",
  2057 => x"00000000",
  2058 => x"00000000",
  2059 => x"00000000",
  2060 => x"00000000",
  2061 => x"00000000",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"00000000",
  2065 => x"00000000",
  2066 => x"00000000",
  2067 => x"00000000",
  2068 => x"00000000",
  2069 => x"00000000",
  2070 => x"00000000",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"ffffffff",
  2098 => x"00000000",
  2099 => x"ffffffff",
  2100 => x"00000000",
  2101 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
