-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpu_config.all;
use work.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80d5f40c",
     3 => x"3a0b0b80",
     4 => x"c4fb0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80c5c22d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c3040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a6",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80d5",
   162 => x"e0738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88a90400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b0bad",
   171 => x"aa2d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b0bad",
   179 => x"ee2d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80d5f00c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82fd3fbf",
   257 => x"a03f0410",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10105351",
   266 => x"047381ff",
   267 => x"06738306",
   268 => x"09810583",
   269 => x"05101010",
   270 => x"2b0772fc",
   271 => x"060c5151",
   272 => x"043c0472",
   273 => x"72807281",
   274 => x"06ff0509",
   275 => x"72060571",
   276 => x"1052720a",
   277 => x"100a5372",
   278 => x"ed385151",
   279 => x"535104ff",
   280 => x"3d0d0b0b",
   281 => x"80e5e408",
   282 => x"52710870",
   283 => x"882a8132",
   284 => x"70810651",
   285 => x"515170f1",
   286 => x"3873720c",
   287 => x"833d0d04",
   288 => x"80d5f008",
   289 => x"802ea438",
   290 => x"80d5f408",
   291 => x"822ebd38",
   292 => x"8380800b",
   293 => x"0b0b80e5",
   294 => x"e40c82a0",
   295 => x"800b80e5",
   296 => x"e80c8290",
   297 => x"800b80e5",
   298 => x"ec0c04f8",
   299 => x"808080a4",
   300 => x"0b0b0b80",
   301 => x"e5e40cf8",
   302 => x"80808280",
   303 => x"0b80e5e8",
   304 => x"0cf88080",
   305 => x"84800b80",
   306 => x"e5ec0c04",
   307 => x"80c0a880",
   308 => x"8c0b0b0b",
   309 => x"80e5e40c",
   310 => x"80c0a880",
   311 => x"940b80e5",
   312 => x"e80c0b0b",
   313 => x"80c7d00b",
   314 => x"80e5ec0c",
   315 => x"04f23d0d",
   316 => x"6080e5e8",
   317 => x"08565d82",
   318 => x"750c8059",
   319 => x"805a800b",
   320 => x"8f3d5d5b",
   321 => x"7a101015",
   322 => x"70087108",
   323 => x"719f2c7e",
   324 => x"852b5855",
   325 => x"557d5359",
   326 => x"5799993f",
   327 => x"7d7f7a72",
   328 => x"077c7207",
   329 => x"71716081",
   330 => x"05415f5d",
   331 => x"5b595755",
   332 => x"817b278f",
   333 => x"38767d0c",
   334 => x"77841e0c",
   335 => x"7c800c90",
   336 => x"3d0d0480",
   337 => x"e5e80855",
   338 => x"ffba3970",
   339 => x"7080e5f0",
   340 => x"335170a7",
   341 => x"3880d5fc",
   342 => x"08700852",
   343 => x"5270802e",
   344 => x"94388412",
   345 => x"80d5fc0c",
   346 => x"702d80d5",
   347 => x"fc087008",
   348 => x"525270ee",
   349 => x"38810b80",
   350 => x"e5f03450",
   351 => x"50040470",
   352 => x"0b0b80e5",
   353 => x"e008802e",
   354 => x"8e380b0b",
   355 => x"0b0b800b",
   356 => x"802e0981",
   357 => x"06833850",
   358 => x"040b0b80",
   359 => x"e5e0510b",
   360 => x"0b0bf4dc",
   361 => x"3f500404",
   362 => x"ff3d0d02",
   363 => x"8f053352",
   364 => x"718a2e8a",
   365 => x"387151fd",
   366 => x"a63f833d",
   367 => x"0d048d51",
   368 => x"fd9d3f71",
   369 => x"51fd983f",
   370 => x"833d0d04",
   371 => x"ce3d0db5",
   372 => x"3d707084",
   373 => x"0552088b",
   374 => x"a85c56a5",
   375 => x"3d5e5c80",
   376 => x"75708105",
   377 => x"5733765b",
   378 => x"55587378",
   379 => x"2e80c138",
   380 => x"8e3d5b73",
   381 => x"a52e0981",
   382 => x"0680c538",
   383 => x"78708105",
   384 => x"5a335473",
   385 => x"80e42e81",
   386 => x"b6387380",
   387 => x"e42480c6",
   388 => x"387380e3",
   389 => x"2ea13880",
   390 => x"52a55179",
   391 => x"2d805273",
   392 => x"51792d82",
   393 => x"18587870",
   394 => x"81055a33",
   395 => x"5473c438",
   396 => x"77800cb4",
   397 => x"3d0d047b",
   398 => x"841d8312",
   399 => x"33565d57",
   400 => x"80527351",
   401 => x"792d8118",
   402 => x"79708105",
   403 => x"5b335558",
   404 => x"73ffa038",
   405 => x"db397380",
   406 => x"f32e0981",
   407 => x"06ffb838",
   408 => x"7b841d71",
   409 => x"08595d56",
   410 => x"80773355",
   411 => x"5673762e",
   412 => x"8d388116",
   413 => x"70187033",
   414 => x"57555674",
   415 => x"f538ff16",
   416 => x"55807625",
   417 => x"ffa03876",
   418 => x"70810558",
   419 => x"33548052",
   420 => x"7351792d",
   421 => x"811875ff",
   422 => x"17575758",
   423 => x"807625ff",
   424 => x"85387670",
   425 => x"81055833",
   426 => x"54805273",
   427 => x"51792d81",
   428 => x"1875ff17",
   429 => x"57575875",
   430 => x"8024cc38",
   431 => x"fee8397b",
   432 => x"841d7108",
   433 => x"70719f2c",
   434 => x"5953595d",
   435 => x"56807524",
   436 => x"81913875",
   437 => x"7d7c5856",
   438 => x"54805773",
   439 => x"772e0981",
   440 => x"06b638b0",
   441 => x"7b3402b5",
   442 => x"05567a76",
   443 => x"2e9738ff",
   444 => x"16567533",
   445 => x"75708105",
   446 => x"57348117",
   447 => x"577a762e",
   448 => x"098106eb",
   449 => x"38807534",
   450 => x"767dff12",
   451 => x"57585675",
   452 => x"8024fef3",
   453 => x"38fe8f39",
   454 => x"8a527351",
   455 => x"9fd03f80",
   456 => x"0880c7d4",
   457 => x"05337670",
   458 => x"81055834",
   459 => x"8a527351",
   460 => x"9ef83f80",
   461 => x"08548008",
   462 => x"802effae",
   463 => x"388a5273",
   464 => x"519fab3f",
   465 => x"800880c7",
   466 => x"d4053376",
   467 => x"70810558",
   468 => x"348a5273",
   469 => x"519ed33f",
   470 => x"80085480",
   471 => x"08ffb938",
   472 => x"ff883974",
   473 => x"527653b4",
   474 => x"3dffb805",
   475 => x"51949a3f",
   476 => x"a33d0856",
   477 => x"fedd3980",
   478 => x"3d0d80c1",
   479 => x"0b81b4bc",
   480 => x"34800b81",
   481 => x"b6980c70",
   482 => x"800c823d",
   483 => x"0d04ff3d",
   484 => x"0d800b81",
   485 => x"b4bc3352",
   486 => x"527080c1",
   487 => x"2e993871",
   488 => x"81b69808",
   489 => x"0781b698",
   490 => x"0c80c20b",
   491 => x"81b4c034",
   492 => x"70800c83",
   493 => x"3d0d0481",
   494 => x"0b81b698",
   495 => x"080781b6",
   496 => x"980c80c2",
   497 => x"0b81b4c0",
   498 => x"3470800c",
   499 => x"833d0d04",
   500 => x"fd3d0d75",
   501 => x"70088a05",
   502 => x"535381b4",
   503 => x"bc335170",
   504 => x"80c12e8b",
   505 => x"3873f338",
   506 => x"70800c85",
   507 => x"3d0d04ff",
   508 => x"127081b4",
   509 => x"b8083174",
   510 => x"0c800c85",
   511 => x"3d0d04fc",
   512 => x"3d0d81b4",
   513 => x"c4085574",
   514 => x"802e8c38",
   515 => x"76750871",
   516 => x"0c81b4c4",
   517 => x"0856548c",
   518 => x"155381b4",
   519 => x"b808528a",
   520 => x"518fd43f",
   521 => x"73800c86",
   522 => x"3d0d04fb",
   523 => x"3d0d7770",
   524 => x"085656b0",
   525 => x"5381b4c4",
   526 => x"08527451",
   527 => x"ab943f85",
   528 => x"0b8c170c",
   529 => x"850b8c16",
   530 => x"0c750875",
   531 => x"0c81b4c4",
   532 => x"08547380",
   533 => x"2e8a3873",
   534 => x"08750c81",
   535 => x"b4c40854",
   536 => x"8c145381",
   537 => x"b4b80852",
   538 => x"8a518f8b",
   539 => x"3f841508",
   540 => x"ad38860b",
   541 => x"8c160c88",
   542 => x"15528816",
   543 => x"08518e97",
   544 => x"3f81b4c4",
   545 => x"08700876",
   546 => x"0c548c15",
   547 => x"7054548a",
   548 => x"52730851",
   549 => x"8ee13f73",
   550 => x"800c873d",
   551 => x"0d047508",
   552 => x"54b05373",
   553 => x"527551aa",
   554 => x"a93f7380",
   555 => x"0c873d0d",
   556 => x"04d93d0d",
   557 => x"b0519dcf",
   558 => x"3f800881",
   559 => x"b4b40cb0",
   560 => x"519dc43f",
   561 => x"800881b4",
   562 => x"c40c81b4",
   563 => x"b4088008",
   564 => x"0c800b80",
   565 => x"0884050c",
   566 => x"820b8008",
   567 => x"88050ca8",
   568 => x"0b80088c",
   569 => x"050c9f53",
   570 => x"80c7e052",
   571 => x"80089005",
   572 => x"51a9df3f",
   573 => x"a13d5e9f",
   574 => x"5380c880",
   575 => x"527d51a9",
   576 => x"d13f8a0b",
   577 => x"80f2f80c",
   578 => x"80d2a451",
   579 => x"f9be3f80",
   580 => x"c8a051f9",
   581 => x"b73f80d2",
   582 => x"a451f9b0",
   583 => x"3f80d684",
   584 => x"08802e89",
   585 => x"d33880c8",
   586 => x"d051f9a0",
   587 => x"3f80d2a4",
   588 => x"51f9993f",
   589 => x"80d68008",
   590 => x"5280c8fc",
   591 => x"51f98d3f",
   592 => x"80e69451",
   593 => x"b2ff3f81",
   594 => x"0b9a3d5e",
   595 => x"5b800b80",
   596 => x"d6800825",
   597 => x"82d43890",
   598 => x"3d5f80c1",
   599 => x"0b81b4bc",
   600 => x"34810b81",
   601 => x"b6980c80",
   602 => x"c20b81b4",
   603 => x"c0348240",
   604 => x"835a9f53",
   605 => x"80c9ac52",
   606 => x"7c51a8d6",
   607 => x"3f814180",
   608 => x"7d537e52",
   609 => x"568e943f",
   610 => x"8008762e",
   611 => x"09810683",
   612 => x"38815675",
   613 => x"81b6980c",
   614 => x"7f705856",
   615 => x"758325a2",
   616 => x"38751010",
   617 => x"16fd0542",
   618 => x"a93dffa4",
   619 => x"05538352",
   620 => x"76518cc3",
   621 => x"3f7f8105",
   622 => x"70417058",
   623 => x"56837624",
   624 => x"e0386154",
   625 => x"755380e6",
   626 => x"9c5281b4",
   627 => x"d0518cb7",
   628 => x"3f81b4c4",
   629 => x"08700858",
   630 => x"58b05377",
   631 => x"527651a7",
   632 => x"f13f850b",
   633 => x"8c190c85",
   634 => x"0b8c180c",
   635 => x"7708770c",
   636 => x"81b4c408",
   637 => x"5675802e",
   638 => x"8a387508",
   639 => x"770c81b4",
   640 => x"c408568c",
   641 => x"165381b4",
   642 => x"b808528a",
   643 => x"518be83f",
   644 => x"84170887",
   645 => x"ea38860b",
   646 => x"8c180c88",
   647 => x"17528818",
   648 => x"08518af3",
   649 => x"3f81b4c4",
   650 => x"08700878",
   651 => x"0c568c17",
   652 => x"7054598a",
   653 => x"52780851",
   654 => x"8bbd3f80",
   655 => x"c10b81b4",
   656 => x"c0335757",
   657 => x"767626a2",
   658 => x"3880c352",
   659 => x"76518ca1",
   660 => x"3f800861",
   661 => x"2e89e438",
   662 => x"81177081",
   663 => x"ff0681b4",
   664 => x"c0335858",
   665 => x"58757727",
   666 => x"e0387960",
   667 => x"29627054",
   668 => x"71535b59",
   669 => x"98b43f80",
   670 => x"0840787a",
   671 => x"31708729",
   672 => x"80083180",
   673 => x"088a0581",
   674 => x"b4bc3381",
   675 => x"b4b8085e",
   676 => x"5b525a56",
   677 => x"7780c12e",
   678 => x"89ce387b",
   679 => x"f738811b",
   680 => x"5b80d680",
   681 => x"087b25fd",
   682 => x"b13881b4",
   683 => x"ac51b095",
   684 => x"3f80c9cc",
   685 => x"51f6953f",
   686 => x"80d2a451",
   687 => x"f68e3f80",
   688 => x"c9dc51f6",
   689 => x"873f80d2",
   690 => x"a451f680",
   691 => x"3f81b4b8",
   692 => x"085280ca",
   693 => x"9451f5f4",
   694 => x"3f855280",
   695 => x"cab051f5",
   696 => x"eb3f81b6",
   697 => x"98085280",
   698 => x"cacc51f5",
   699 => x"df3f8152",
   700 => x"80cab051",
   701 => x"f5d63f81",
   702 => x"b4bc3352",
   703 => x"80cae851",
   704 => x"f5ca3f80",
   705 => x"c15280cb",
   706 => x"8451f5c0",
   707 => x"3f81b4c0",
   708 => x"335280cb",
   709 => x"a051f5b4",
   710 => x"3f80c252",
   711 => x"80cb8451",
   712 => x"f5aa3f81",
   713 => x"b4f00852",
   714 => x"80cbbc51",
   715 => x"f59e3f87",
   716 => x"5280cab0",
   717 => x"51f5953f",
   718 => x"80f2f808",
   719 => x"5280cbd8",
   720 => x"51f5893f",
   721 => x"80cbf451",
   722 => x"f5823f80",
   723 => x"cca051f4",
   724 => x"fb3f81b4",
   725 => x"c4087008",
   726 => x"535a80cc",
   727 => x"ac51f4ec",
   728 => x"3f80ccc8",
   729 => x"51f4e53f",
   730 => x"81b4c408",
   731 => x"84110853",
   732 => x"5680ccfc",
   733 => x"51f4d53f",
   734 => x"805280ca",
   735 => x"b051f4cc",
   736 => x"3f81b4c4",
   737 => x"08881108",
   738 => x"535880cd",
   739 => x"9851f4bc",
   740 => x"3f825280",
   741 => x"cab051f4",
   742 => x"b33f81b4",
   743 => x"c4088c11",
   744 => x"08535780",
   745 => x"cdb451f4",
   746 => x"a33f9152",
   747 => x"80cab051",
   748 => x"f49a3f81",
   749 => x"b4c40890",
   750 => x"055280cd",
   751 => x"d051f48c",
   752 => x"3f80cdec",
   753 => x"51f4853f",
   754 => x"80cea451",
   755 => x"f3fe3f81",
   756 => x"b4b40870",
   757 => x"08535f80",
   758 => x"ccac51f3",
   759 => x"ef3f80ce",
   760 => x"b851f3e8",
   761 => x"3f81b4b4",
   762 => x"08841108",
   763 => x"535b80cc",
   764 => x"fc51f3d8",
   765 => x"3f805280",
   766 => x"cab051f3",
   767 => x"cf3f81b4",
   768 => x"b4088811",
   769 => x"08535c80",
   770 => x"cd9851f3",
   771 => x"bf3f8152",
   772 => x"80cab051",
   773 => x"f3b63f81",
   774 => x"b4b4088c",
   775 => x"1108535a",
   776 => x"80cdb451",
   777 => x"f3a63f92",
   778 => x"5280cab0",
   779 => x"51f39d3f",
   780 => x"81b4b408",
   781 => x"90055280",
   782 => x"cdd051f3",
   783 => x"8f3f80cd",
   784 => x"ec51f388",
   785 => x"3f7f5280",
   786 => x"cef851f2",
   787 => x"ff3f8552",
   788 => x"80cab051",
   789 => x"f2f63f78",
   790 => x"5280cf94",
   791 => x"51f2ed3f",
   792 => x"8d5280ca",
   793 => x"b051f2e4",
   794 => x"3f615280",
   795 => x"cfb051f2",
   796 => x"db3f8752",
   797 => x"80cab051",
   798 => x"f2d23f60",
   799 => x"5280cfcc",
   800 => x"51f2c93f",
   801 => x"815280ca",
   802 => x"b051f2c0",
   803 => x"3f7d5280",
   804 => x"cfe851f2",
   805 => x"b73f80d0",
   806 => x"8451f2b0",
   807 => x"3f7c5280",
   808 => x"d0bc51f2",
   809 => x"a73f80d0",
   810 => x"d851f2a0",
   811 => x"3f80d2a4",
   812 => x"51f2993f",
   813 => x"81b4ac08",
   814 => x"81b4b008",
   815 => x"80e69408",
   816 => x"80e69808",
   817 => x"72713170",
   818 => x"74267574",
   819 => x"31707231",
   820 => x"80e68c0c",
   821 => x"444480e6",
   822 => x"900c80e6",
   823 => x"90085680",
   824 => x"d190555c",
   825 => x"595758f1",
   826 => x"e33f80e6",
   827 => x"8c085680",
   828 => x"762582a3",
   829 => x"3880d680",
   830 => x"0870719f",
   831 => x"2c9a3d53",
   832 => x"565680e6",
   833 => x"8c0880e6",
   834 => x"90084153",
   835 => x"7f547052",
   836 => x"5a89eb3f",
   837 => x"66685f80",
   838 => x"e5fc0c7d",
   839 => x"80e6800c",
   840 => x"80d68008",
   841 => x"709f2c58",
   842 => x"568058bd",
   843 => x"84c07855",
   844 => x"55765275",
   845 => x"53795187",
   846 => x"d13f953d",
   847 => x"80e68c08",
   848 => x"80e69008",
   849 => x"41557f56",
   850 => x"67694053",
   851 => x"7e547052",
   852 => x"5c89ab3f",
   853 => x"64665e80",
   854 => x"e6840c7c",
   855 => x"80e6880c",
   856 => x"80d68008",
   857 => x"709f2c40",
   858 => x"58805783",
   859 => x"dceb9480",
   860 => x"7755557e",
   861 => x"5277537b",
   862 => x"51878f3f",
   863 => x"64665d5b",
   864 => x"805e8ddd",
   865 => x"7e555580",
   866 => x"e68c0880",
   867 => x"e6900859",
   868 => x"52775379",
   869 => x"5186f33f",
   870 => x"66684054",
   871 => x"7e557a52",
   872 => x"7b53a93d",
   873 => x"ffa80551",
   874 => x"88d43f62",
   875 => x"645e81b4",
   876 => x"c80c7c81",
   877 => x"b4cc0c80",
   878 => x"d1a051f0",
   879 => x"8f3f80e6",
   880 => x"80085280",
   881 => x"d1d051f0",
   882 => x"833f80d1",
   883 => x"d851effc",
   884 => x"3f80e688",
   885 => x"085280d1",
   886 => x"d051eff0",
   887 => x"3f81b4cc",
   888 => x"085280d2",
   889 => x"8851efe4",
   890 => x"3f80d2a4",
   891 => x"51efdd3f",
   892 => x"800b800c",
   893 => x"a93d0d04",
   894 => x"80d2a851",
   895 => x"f6ac3977",
   896 => x"0857b053",
   897 => x"76527751",
   898 => x"9fc83f80",
   899 => x"c10b81b4",
   900 => x"c0335757",
   901 => x"f8ae3975",
   902 => x"8a3880e6",
   903 => x"90088126",
   904 => x"fdd33880",
   905 => x"d2d851ef",
   906 => x"a33f80d3",
   907 => x"9051ef9c",
   908 => x"3f80d2a4",
   909 => x"51ef953f",
   910 => x"80d68008",
   911 => x"70719f2c",
   912 => x"9a3d5356",
   913 => x"5680e68c",
   914 => x"0880e690",
   915 => x"0841537f",
   916 => x"5470525a",
   917 => x"87a83f66",
   918 => x"685f80e5",
   919 => x"fc0c7d80",
   920 => x"e6800c80",
   921 => x"d6800870",
   922 => x"9f2c5856",
   923 => x"8058bd84",
   924 => x"c0785555",
   925 => x"76527553",
   926 => x"7951858e",
   927 => x"3f953d80",
   928 => x"e68c0880",
   929 => x"e6900841",
   930 => x"557f5667",
   931 => x"6940537e",
   932 => x"5470525c",
   933 => x"86e83f64",
   934 => x"665e80e6",
   935 => x"840c7c80",
   936 => x"e6880c80",
   937 => x"d6800870",
   938 => x"9f2c4058",
   939 => x"805783dc",
   940 => x"eb948077",
   941 => x"55557e52",
   942 => x"77537b51",
   943 => x"84cc3f64",
   944 => x"665d5b80",
   945 => x"5e8ddd7e",
   946 => x"555580e6",
   947 => x"8c0880e6",
   948 => x"90085952",
   949 => x"77537951",
   950 => x"84b03f66",
   951 => x"6840547e",
   952 => x"557a527b",
   953 => x"53a93dff",
   954 => x"a8055186",
   955 => x"913f6264",
   956 => x"5e81b4c8",
   957 => x"0c7c81b4",
   958 => x"cc0c80d1",
   959 => x"a051edcc",
   960 => x"3f80e680",
   961 => x"085280d1",
   962 => x"d051edc0",
   963 => x"3f80d1d8",
   964 => x"51edb93f",
   965 => x"80e68808",
   966 => x"5280d1d0",
   967 => x"51edad3f",
   968 => x"81b4cc08",
   969 => x"5280d288",
   970 => x"51eda13f",
   971 => x"80d2a451",
   972 => x"ed9a3f80",
   973 => x"0b800ca9",
   974 => x"3d0d04a9",
   975 => x"3dffa005",
   976 => x"52805180",
   977 => x"d23f9f53",
   978 => x"80d3b052",
   979 => x"7c519d82",
   980 => x"3f7a7b81",
   981 => x"b4b80c81",
   982 => x"187081ff",
   983 => x"0681b4c0",
   984 => x"33595959",
   985 => x"5af5fe39",
   986 => x"ff16707b",
   987 => x"31600c5c",
   988 => x"800b811c",
   989 => x"5c5c80d6",
   990 => x"80087b25",
   991 => x"f3dc38f6",
   992 => x"a939ff3d",
   993 => x"0d738232",
   994 => x"70307072",
   995 => x"07802580",
   996 => x"0c525283",
   997 => x"3d0d04fe",
   998 => x"3d0d7476",
   999 => x"71535452",
  1000 => x"71822e83",
  1001 => x"38835171",
  1002 => x"812e9a38",
  1003 => x"8172269f",
  1004 => x"3871822e",
  1005 => x"b8387184",
  1006 => x"2ea93870",
  1007 => x"730c7080",
  1008 => x"0c843d0d",
  1009 => x"0480e40b",
  1010 => x"81b4b808",
  1011 => x"258b3880",
  1012 => x"730c7080",
  1013 => x"0c843d0d",
  1014 => x"0483730c",
  1015 => x"70800c84",
  1016 => x"3d0d0482",
  1017 => x"730c7080",
  1018 => x"0c843d0d",
  1019 => x"0481730c",
  1020 => x"70800c84",
  1021 => x"3d0d0480",
  1022 => x"3d0d7474",
  1023 => x"14820571",
  1024 => x"0c800c82",
  1025 => x"3d0d04f7",
  1026 => x"3d0d7b7d",
  1027 => x"7f618512",
  1028 => x"70822b75",
  1029 => x"11707471",
  1030 => x"70840553",
  1031 => x"0c5a5a5d",
  1032 => x"5b760c79",
  1033 => x"80f8180c",
  1034 => x"79861252",
  1035 => x"57585a5a",
  1036 => x"76762499",
  1037 => x"3876b329",
  1038 => x"822b7911",
  1039 => x"51537673",
  1040 => x"70840555",
  1041 => x"0c811454",
  1042 => x"757425f2",
  1043 => x"387681cc",
  1044 => x"2919fc11",
  1045 => x"088105fc",
  1046 => x"120c7a19",
  1047 => x"70089fa0",
  1048 => x"130c5856",
  1049 => x"850b81b4",
  1050 => x"b80c7580",
  1051 => x"0c8b3d0d",
  1052 => x"04fe3d0d",
  1053 => x"02930533",
  1054 => x"51800284",
  1055 => x"05970533",
  1056 => x"54527073",
  1057 => x"2e883871",
  1058 => x"800c843d",
  1059 => x"0d047081",
  1060 => x"b4bc3481",
  1061 => x"0b800c84",
  1062 => x"3d0d04f8",
  1063 => x"3d0d7a7c",
  1064 => x"5956820b",
  1065 => x"83195555",
  1066 => x"74167033",
  1067 => x"75335b51",
  1068 => x"5372792e",
  1069 => x"80c63880",
  1070 => x"c10b8116",
  1071 => x"81165656",
  1072 => x"57827525",
  1073 => x"e338ffa9",
  1074 => x"177081ff",
  1075 => x"06555973",
  1076 => x"82268338",
  1077 => x"87558153",
  1078 => x"7680d22e",
  1079 => x"98387752",
  1080 => x"75519bc3",
  1081 => x"3f805372",
  1082 => x"80082589",
  1083 => x"38871581",
  1084 => x"b4b80c81",
  1085 => x"5372800c",
  1086 => x"8a3d0d04",
  1087 => x"7281b4bc",
  1088 => x"34827525",
  1089 => x"ffa238ff",
  1090 => x"bd39ef3d",
  1091 => x"0d636567",
  1092 => x"5b427943",
  1093 => x"67695940",
  1094 => x"77415a80",
  1095 => x"5d805e61",
  1096 => x"7083ffff",
  1097 => x"0671902a",
  1098 => x"627083ff",
  1099 => x"ff067190",
  1100 => x"2a747229",
  1101 => x"74732975",
  1102 => x"73297774",
  1103 => x"2973902a",
  1104 => x"05721151",
  1105 => x"5856535f",
  1106 => x"5a575a58",
  1107 => x"55587373",
  1108 => x"27863884",
  1109 => x"80801656",
  1110 => x"73902a16",
  1111 => x"5b7883ff",
  1112 => x"ff067484",
  1113 => x"80802905",
  1114 => x"5c7a7c5a",
  1115 => x"5d785e77",
  1116 => x"7f296178",
  1117 => x"29057d05",
  1118 => x"5d7c7e56",
  1119 => x"7a0c7484",
  1120 => x"1b0c7980",
  1121 => x"0c933d0d",
  1122 => x"04f93d0d",
  1123 => x"797b7d54",
  1124 => x"58725977",
  1125 => x"30797030",
  1126 => x"7072079f",
  1127 => x"2a737131",
  1128 => x"5a525977",
  1129 => x"7956730c",
  1130 => x"53738413",
  1131 => x"0c54800c",
  1132 => x"893d0d04",
  1133 => x"f93d0d79",
  1134 => x"7b7d7f56",
  1135 => x"54525472",
  1136 => x"802ea038",
  1137 => x"70577158",
  1138 => x"a0733152",
  1139 => x"807225a1",
  1140 => x"38777074",
  1141 => x"2b577073",
  1142 => x"2a78752b",
  1143 => x"07565174",
  1144 => x"76535170",
  1145 => x"740c7184",
  1146 => x"150c7380",
  1147 => x"0c893d0d",
  1148 => x"04805677",
  1149 => x"72302b55",
  1150 => x"74765351",
  1151 => x"e639e43d",
  1152 => x"0d6ea13d",
  1153 => x"08a33d08",
  1154 => x"59575f80",
  1155 => x"764d774e",
  1156 => x"a33d08a5",
  1157 => x"3d08574b",
  1158 => x"754c5e7d",
  1159 => x"6c2486fb",
  1160 => x"38806a24",
  1161 => x"878f3869",
  1162 => x"6b58566b",
  1163 => x"6d5d467b",
  1164 => x"47754476",
  1165 => x"45646468",
  1166 => x"685c5c56",
  1167 => x"567481e7",
  1168 => x"38787627",
  1169 => x"82c73875",
  1170 => x"81ff2683",
  1171 => x"2b5583ff",
  1172 => x"ff76278c",
  1173 => x"389055fe",
  1174 => x"800a7627",
  1175 => x"83389855",
  1176 => x"75752a80",
  1177 => x"d3d00570",
  1178 => x"33a07731",
  1179 => x"71315755",
  1180 => x"5774802e",
  1181 => x"95387575",
  1182 => x"2ba07631",
  1183 => x"7a772b7c",
  1184 => x"722a077c",
  1185 => x"782b5d5b",
  1186 => x"59567590",
  1187 => x"2a7683ff",
  1188 => x"ff067154",
  1189 => x"7a535957",
  1190 => x"88803f80",
  1191 => x"085b87ea",
  1192 => x"3f800880",
  1193 => x"0879297c",
  1194 => x"902b7c90",
  1195 => x"2a075656",
  1196 => x"59737527",
  1197 => x"94388008",
  1198 => x"ff057615",
  1199 => x"55597574",
  1200 => x"26873874",
  1201 => x"742687b9",
  1202 => x"38765273",
  1203 => x"75315187",
  1204 => x"c93f8008",
  1205 => x"5587b33f",
  1206 => x"80088008",
  1207 => x"79297b83",
  1208 => x"ffff0677",
  1209 => x"902b0756",
  1210 => x"59577378",
  1211 => x"27963880",
  1212 => x"08ff0576",
  1213 => x"15555775",
  1214 => x"74268938",
  1215 => x"77742677",
  1216 => x"71315856",
  1217 => x"78902b77",
  1218 => x"0758805b",
  1219 => x"7a407741",
  1220 => x"7f615654",
  1221 => x"7d80d938",
  1222 => x"737f0c74",
  1223 => x"7f84050c",
  1224 => x"7e800c9e",
  1225 => x"3d0d0480",
  1226 => x"705c5874",
  1227 => x"7926dd38",
  1228 => x"7481ff26",
  1229 => x"832b5774",
  1230 => x"83ffff26",
  1231 => x"82a53874",
  1232 => x"772a80d3",
  1233 => x"d0057033",
  1234 => x"a0793171",
  1235 => x"31595c5d",
  1236 => x"7682b338",
  1237 => x"76547479",
  1238 => x"27833881",
  1239 => x"54797627",
  1240 => x"74075981",
  1241 => x"5878ffa2",
  1242 => x"38765880",
  1243 => x"5bff9d39",
  1244 => x"73527453",
  1245 => x"9e3de805",
  1246 => x"51fc8e3f",
  1247 => x"6769567f",
  1248 => x"0c747f84",
  1249 => x"050c7e80",
  1250 => x"0c9e3d0d",
  1251 => x"0475802e",
  1252 => x"81c43875",
  1253 => x"81ff2683",
  1254 => x"2b5583ff",
  1255 => x"ff76278c",
  1256 => x"389055fe",
  1257 => x"800a7627",
  1258 => x"83389855",
  1259 => x"75752a80",
  1260 => x"d3d00570",
  1261 => x"33a07731",
  1262 => x"7131575e",
  1263 => x"54748491",
  1264 => x"38787631",
  1265 => x"54817690",
  1266 => x"2a7783ff",
  1267 => x"ff065f5d",
  1268 => x"5b7b5273",
  1269 => x"5185c33f",
  1270 => x"80085785",
  1271 => x"ad3f8008",
  1272 => x"80087e29",
  1273 => x"78902b7c",
  1274 => x"902a0756",
  1275 => x"56597375",
  1276 => x"27943880",
  1277 => x"08ff0576",
  1278 => x"15555975",
  1279 => x"74268738",
  1280 => x"74742684",
  1281 => x"f3387b52",
  1282 => x"73753151",
  1283 => x"858c3f80",
  1284 => x"085584f6",
  1285 => x"3f800880",
  1286 => x"087e297b",
  1287 => x"83ffff06",
  1288 => x"77902b07",
  1289 => x"56595773",
  1290 => x"78279638",
  1291 => x"8008ff05",
  1292 => x"76155557",
  1293 => x"75742689",
  1294 => x"38777426",
  1295 => x"77713158",
  1296 => x"5a78902b",
  1297 => x"77077b41",
  1298 => x"417f6156",
  1299 => x"547d802e",
  1300 => x"fdc638fe",
  1301 => x"9b397552",
  1302 => x"815184ae",
  1303 => x"3f800856",
  1304 => x"feb13990",
  1305 => x"57fe800a",
  1306 => x"7527fdd3",
  1307 => x"38987571",
  1308 => x"2a80d3d0",
  1309 => x"057033a0",
  1310 => x"73317131",
  1311 => x"535d5e57",
  1312 => x"76802efd",
  1313 => x"cf38a077",
  1314 => x"3175782b",
  1315 => x"77722a07",
  1316 => x"77792b7b",
  1317 => x"7a2b7d74",
  1318 => x"2a077d7b",
  1319 => x"2b73902a",
  1320 => x"7483ffff",
  1321 => x"0671597f",
  1322 => x"772a585e",
  1323 => x"5c415f58",
  1324 => x"5c5483e6",
  1325 => x"3f800854",
  1326 => x"83d03f80",
  1327 => x"08800879",
  1328 => x"2975902b",
  1329 => x"7e902a07",
  1330 => x"56565973",
  1331 => x"75279938",
  1332 => x"8008ff05",
  1333 => x"7b155559",
  1334 => x"7a74268c",
  1335 => x"38737527",
  1336 => x"8738ff19",
  1337 => x"7b155559",
  1338 => x"76527375",
  1339 => x"315183aa",
  1340 => x"3f800855",
  1341 => x"83943f80",
  1342 => x"08800879",
  1343 => x"297d83ff",
  1344 => x"ff067790",
  1345 => x"2b075659",
  1346 => x"57737827",
  1347 => x"99388008",
  1348 => x"ff057b15",
  1349 => x"55577a74",
  1350 => x"268c3873",
  1351 => x"78278738",
  1352 => x"ff177b15",
  1353 => x"55577378",
  1354 => x"3179902b",
  1355 => x"78077083",
  1356 => x"ffff0671",
  1357 => x"902a7983",
  1358 => x"ffff067a",
  1359 => x"902a7372",
  1360 => x"29737329",
  1361 => x"74732976",
  1362 => x"74297390",
  1363 => x"2a057205",
  1364 => x"5755435f",
  1365 => x"5b585a57",
  1366 => x"595a747c",
  1367 => x"27863884",
  1368 => x"80801757",
  1369 => x"74902a17",
  1370 => x"7983ffff",
  1371 => x"06768480",
  1372 => x"80290557",
  1373 => x"57767a26",
  1374 => x"9a38767a",
  1375 => x"32703070",
  1376 => x"72078025",
  1377 => x"565a5b7c",
  1378 => x"7627fafe",
  1379 => x"3873802e",
  1380 => x"faf838ff",
  1381 => x"1858805b",
  1382 => x"faf239ff",
  1383 => x"76537754",
  1384 => x"9f3de805",
  1385 => x"525ef7e1",
  1386 => x"3f676957",
  1387 => x"4c754d69",
  1388 => x"8025f8f3",
  1389 => x"387d096a",
  1390 => x"6c5c537a",
  1391 => x"549f3de8",
  1392 => x"05525ef7",
  1393 => x"c43f6769",
  1394 => x"714c704d",
  1395 => x"5856f8db",
  1396 => x"39a07531",
  1397 => x"76762b7a",
  1398 => x"772b7c73",
  1399 => x"2a077c78",
  1400 => x"2b72902a",
  1401 => x"7383ffff",
  1402 => x"0671587e",
  1403 => x"762a5742",
  1404 => x"405d5d57",
  1405 => x"5881a33f",
  1406 => x"80085781",
  1407 => x"8d3f8008",
  1408 => x"80087e29",
  1409 => x"78902b7d",
  1410 => x"902a0756",
  1411 => x"56597375",
  1412 => x"27993880",
  1413 => x"08ff0576",
  1414 => x"15555975",
  1415 => x"74268c38",
  1416 => x"73752787",
  1417 => x"38ff1976",
  1418 => x"1555597b",
  1419 => x"52737531",
  1420 => x"5180e73f",
  1421 => x"80085580",
  1422 => x"d13f8008",
  1423 => x"80087e29",
  1424 => x"7c83ffff",
  1425 => x"06707890",
  1426 => x"2b075156",
  1427 => x"58587377",
  1428 => x"27993880",
  1429 => x"08ff0576",
  1430 => x"15555875",
  1431 => x"74268c38",
  1432 => x"73772787",
  1433 => x"38ff1876",
  1434 => x"15555878",
  1435 => x"902b7807",
  1436 => x"74783155",
  1437 => x"5bfada39",
  1438 => x"ff197615",
  1439 => x"5559fb86",
  1440 => x"39ff1976",
  1441 => x"155559f8",
  1442 => x"c0397070",
  1443 => x"70805375",
  1444 => x"52745181",
  1445 => x"913f5050",
  1446 => x"50047070",
  1447 => x"70815375",
  1448 => x"52745181",
  1449 => x"813f5050",
  1450 => x"5004fb3d",
  1451 => x"0d777955",
  1452 => x"55805675",
  1453 => x"7524ab38",
  1454 => x"8074249d",
  1455 => x"38805373",
  1456 => x"52745180",
  1457 => x"e13f8008",
  1458 => x"5475802e",
  1459 => x"85388008",
  1460 => x"30547380",
  1461 => x"0c873d0d",
  1462 => x"04733076",
  1463 => x"81325754",
  1464 => x"dc397430",
  1465 => x"55815673",
  1466 => x"8025d238",
  1467 => x"ec39fa3d",
  1468 => x"0d787a57",
  1469 => x"55805776",
  1470 => x"7524a438",
  1471 => x"759f2c54",
  1472 => x"81537574",
  1473 => x"32743152",
  1474 => x"74519b3f",
  1475 => x"80085476",
  1476 => x"802e8538",
  1477 => x"80083054",
  1478 => x"73800c88",
  1479 => x"3d0d0474",
  1480 => x"30558157",
  1481 => x"d739fc3d",
  1482 => x"0d767853",
  1483 => x"54815380",
  1484 => x"74732652",
  1485 => x"5572802e",
  1486 => x"98387080",
  1487 => x"2eab3880",
  1488 => x"7224a638",
  1489 => x"71107310",
  1490 => x"75722653",
  1491 => x"545272ea",
  1492 => x"38735178",
  1493 => x"83387451",
  1494 => x"70800c86",
  1495 => x"3d0d0472",
  1496 => x"0a100a72",
  1497 => x"0a100a53",
  1498 => x"5372802e",
  1499 => x"e4387174",
  1500 => x"26ed3873",
  1501 => x"72317574",
  1502 => x"07740a10",
  1503 => x"0a740a10",
  1504 => x"0a555556",
  1505 => x"54e33970",
  1506 => x"70735280",
  1507 => x"decc0851",
  1508 => x"933f5050",
  1509 => x"04707073",
  1510 => x"5280decc",
  1511 => x"085190ce",
  1512 => x"3f505004",
  1513 => x"f43d0d7e",
  1514 => x"608b1170",
  1515 => x"f8065b55",
  1516 => x"555d7296",
  1517 => x"26833890",
  1518 => x"58807824",
  1519 => x"74792607",
  1520 => x"55805474",
  1521 => x"742e0981",
  1522 => x"0680ca38",
  1523 => x"7c518d9e",
  1524 => x"3f7783f7",
  1525 => x"2680c538",
  1526 => x"77832a70",
  1527 => x"10101080",
  1528 => x"d6c4058c",
  1529 => x"11085858",
  1530 => x"5475772e",
  1531 => x"81f03884",
  1532 => x"1608fc06",
  1533 => x"8c170888",
  1534 => x"1808718c",
  1535 => x"120c8812",
  1536 => x"0c5b7605",
  1537 => x"84110881",
  1538 => x"0784120c",
  1539 => x"537c518c",
  1540 => x"de3f8816",
  1541 => x"5473800c",
  1542 => x"8e3d0d04",
  1543 => x"77892a78",
  1544 => x"832a5854",
  1545 => x"73802ebf",
  1546 => x"3877862a",
  1547 => x"b8055784",
  1548 => x"7427b438",
  1549 => x"80db1457",
  1550 => x"947427ab",
  1551 => x"38778c2a",
  1552 => x"80ee0557",
  1553 => x"80d47427",
  1554 => x"9e38778f",
  1555 => x"2a80f705",
  1556 => x"5782d474",
  1557 => x"27913877",
  1558 => x"922a80fc",
  1559 => x"05578ad4",
  1560 => x"74278438",
  1561 => x"80fe5776",
  1562 => x"10101080",
  1563 => x"d6c4058c",
  1564 => x"11085653",
  1565 => x"74732ea3",
  1566 => x"38841508",
  1567 => x"fc067079",
  1568 => x"31555673",
  1569 => x"8f2488e4",
  1570 => x"38738025",
  1571 => x"88e6388c",
  1572 => x"15085574",
  1573 => x"732e0981",
  1574 => x"06df3881",
  1575 => x"175980d6",
  1576 => x"d4085675",
  1577 => x"80d6cc2e",
  1578 => x"82cc3884",
  1579 => x"1608fc06",
  1580 => x"70793155",
  1581 => x"55738f24",
  1582 => x"bb3880d6",
  1583 => x"cc0b80d6",
  1584 => x"d80c80d6",
  1585 => x"cc0b80d6",
  1586 => x"d40c8074",
  1587 => x"2480db38",
  1588 => x"74168411",
  1589 => x"08810784",
  1590 => x"120c53fe",
  1591 => x"b0398816",
  1592 => x"8c110857",
  1593 => x"5975792e",
  1594 => x"098106fe",
  1595 => x"82388214",
  1596 => x"59ffab39",
  1597 => x"77167881",
  1598 => x"0784180c",
  1599 => x"7080d6d8",
  1600 => x"0c7080d6",
  1601 => x"d40c80d6",
  1602 => x"cc0b8c12",
  1603 => x"0c8c1108",
  1604 => x"88120c74",
  1605 => x"81078412",
  1606 => x"0c740574",
  1607 => x"710c5b7c",
  1608 => x"518acc3f",
  1609 => x"881654fd",
  1610 => x"ec3983ff",
  1611 => x"75278391",
  1612 => x"3874892a",
  1613 => x"75832a54",
  1614 => x"5473802e",
  1615 => x"bf387486",
  1616 => x"2ab80553",
  1617 => x"847427b4",
  1618 => x"3880db14",
  1619 => x"53947427",
  1620 => x"ab38748c",
  1621 => x"2a80ee05",
  1622 => x"5380d474",
  1623 => x"279e3874",
  1624 => x"8f2a80f7",
  1625 => x"055382d4",
  1626 => x"74279138",
  1627 => x"74922a80",
  1628 => x"fc05538a",
  1629 => x"d4742784",
  1630 => x"3880fe53",
  1631 => x"72101010",
  1632 => x"80d6c405",
  1633 => x"88110855",
  1634 => x"5773772e",
  1635 => x"868b3884",
  1636 => x"1408fc06",
  1637 => x"5b747b27",
  1638 => x"8d388814",
  1639 => x"08547377",
  1640 => x"2e098106",
  1641 => x"ea388c14",
  1642 => x"0880d6c4",
  1643 => x"0b840508",
  1644 => x"718c190c",
  1645 => x"7588190c",
  1646 => x"7788130c",
  1647 => x"5c57758c",
  1648 => x"150c7853",
  1649 => x"80792483",
  1650 => x"98387282",
  1651 => x"2c81712b",
  1652 => x"5656747b",
  1653 => x"2680ca38",
  1654 => x"7a750657",
  1655 => x"7682a338",
  1656 => x"78fc0684",
  1657 => x"05597410",
  1658 => x"707c0655",
  1659 => x"55738292",
  1660 => x"38841959",
  1661 => x"f13980d6",
  1662 => x"c40b8405",
  1663 => x"0879545b",
  1664 => x"788025c6",
  1665 => x"3882da39",
  1666 => x"74097b06",
  1667 => x"7080d6c4",
  1668 => x"0b84050c",
  1669 => x"5b741055",
  1670 => x"747b2685",
  1671 => x"387485bc",
  1672 => x"3880d6c4",
  1673 => x"0b880508",
  1674 => x"70841208",
  1675 => x"fc06707b",
  1676 => x"317b7226",
  1677 => x"8f722507",
  1678 => x"5d575c5c",
  1679 => x"5578802e",
  1680 => x"80d93879",
  1681 => x"1580d6bc",
  1682 => x"08199011",
  1683 => x"59545680",
  1684 => x"d6b808ff",
  1685 => x"2e8838a0",
  1686 => x"8f13e080",
  1687 => x"06577652",
  1688 => x"7c51888c",
  1689 => x"3f800854",
  1690 => x"8008ff2e",
  1691 => x"90388008",
  1692 => x"762782a7",
  1693 => x"387480d6",
  1694 => x"c42e829f",
  1695 => x"3880d6c4",
  1696 => x"0b880508",
  1697 => x"55841508",
  1698 => x"fc067079",
  1699 => x"31797226",
  1700 => x"8f722507",
  1701 => x"5d555a7a",
  1702 => x"83f23877",
  1703 => x"81078416",
  1704 => x"0c771570",
  1705 => x"80d6c40b",
  1706 => x"88050c74",
  1707 => x"81078412",
  1708 => x"0c567c51",
  1709 => x"87b93f88",
  1710 => x"15547380",
  1711 => x"0c8e3d0d",
  1712 => x"0474832a",
  1713 => x"70545480",
  1714 => x"7424819b",
  1715 => x"3872822c",
  1716 => x"81712b80",
  1717 => x"d6c80807",
  1718 => x"7080d6c4",
  1719 => x"0b84050c",
  1720 => x"75101010",
  1721 => x"80d6c405",
  1722 => x"88110871",
  1723 => x"8c1b0c70",
  1724 => x"881b0c79",
  1725 => x"88130c57",
  1726 => x"555c5575",
  1727 => x"8c150cfd",
  1728 => x"c1397879",
  1729 => x"10101080",
  1730 => x"d6c40570",
  1731 => x"565b5c8c",
  1732 => x"14085675",
  1733 => x"742ea338",
  1734 => x"841608fc",
  1735 => x"06707931",
  1736 => x"5853768f",
  1737 => x"2483f138",
  1738 => x"76802584",
  1739 => x"af388c16",
  1740 => x"08567574",
  1741 => x"2e098106",
  1742 => x"df388814",
  1743 => x"811a7083",
  1744 => x"06555a54",
  1745 => x"72c9387b",
  1746 => x"83065675",
  1747 => x"802efdb8",
  1748 => x"38ff1cf8",
  1749 => x"1b5b5c88",
  1750 => x"1a087a2e",
  1751 => x"ea38fdb5",
  1752 => x"39831953",
  1753 => x"fce43983",
  1754 => x"1470822c",
  1755 => x"81712b80",
  1756 => x"d6c80807",
  1757 => x"7080d6c4",
  1758 => x"0b84050c",
  1759 => x"76101010",
  1760 => x"80d6c405",
  1761 => x"88110871",
  1762 => x"8c1c0c70",
  1763 => x"881c0c7a",
  1764 => x"88130c58",
  1765 => x"535d5653",
  1766 => x"fee13980",
  1767 => x"d6880817",
  1768 => x"59800876",
  1769 => x"2e818b38",
  1770 => x"80d6b808",
  1771 => x"ff2e848e",
  1772 => x"38737631",
  1773 => x"1980d688",
  1774 => x"0c738706",
  1775 => x"70565372",
  1776 => x"802e8838",
  1777 => x"88733170",
  1778 => x"15555576",
  1779 => x"149fff06",
  1780 => x"a0807131",
  1781 => x"1670547e",
  1782 => x"53515385",
  1783 => x"933f8008",
  1784 => x"568008ff",
  1785 => x"2e819e38",
  1786 => x"80d68808",
  1787 => x"137080d6",
  1788 => x"880c7475",
  1789 => x"80d6c40b",
  1790 => x"88050c77",
  1791 => x"76311581",
  1792 => x"07555659",
  1793 => x"7a80d6c4",
  1794 => x"2e83c038",
  1795 => x"798f2682",
  1796 => x"ef38810b",
  1797 => x"84150c84",
  1798 => x"1508fc06",
  1799 => x"70793179",
  1800 => x"72268f72",
  1801 => x"25075d55",
  1802 => x"5a7a802e",
  1803 => x"fced3880",
  1804 => x"db398008",
  1805 => x"9fff0655",
  1806 => x"74feed38",
  1807 => x"7880d688",
  1808 => x"0c80d6c4",
  1809 => x"0b880508",
  1810 => x"7a188107",
  1811 => x"84120c55",
  1812 => x"80d6b408",
  1813 => x"79278638",
  1814 => x"7880d6b4",
  1815 => x"0c80d6b0",
  1816 => x"087927fc",
  1817 => x"a0387880",
  1818 => x"d6b00c84",
  1819 => x"1508fc06",
  1820 => x"70793179",
  1821 => x"72268f72",
  1822 => x"25075d55",
  1823 => x"5a7a802e",
  1824 => x"fc993888",
  1825 => x"39807457",
  1826 => x"53fedd39",
  1827 => x"7c5183df",
  1828 => x"3f800b80",
  1829 => x"0c8e3d0d",
  1830 => x"04807324",
  1831 => x"a5387282",
  1832 => x"2c81712b",
  1833 => x"80d6c808",
  1834 => x"077080d6",
  1835 => x"c40b8405",
  1836 => x"0c5c5a76",
  1837 => x"8c170c73",
  1838 => x"88170c75",
  1839 => x"88180cf9",
  1840 => x"fd398313",
  1841 => x"70822c81",
  1842 => x"712b80d6",
  1843 => x"c8080770",
  1844 => x"80d6c40b",
  1845 => x"84050c5d",
  1846 => x"5b53d839",
  1847 => x"7a75065c",
  1848 => x"7bfc9f38",
  1849 => x"84197510",
  1850 => x"5659f139",
  1851 => x"ff178105",
  1852 => x"59f7ab39",
  1853 => x"8c150888",
  1854 => x"1608718c",
  1855 => x"120c8812",
  1856 => x"0c597515",
  1857 => x"84110881",
  1858 => x"0784120c",
  1859 => x"587c5182",
  1860 => x"de3f8815",
  1861 => x"54fba339",
  1862 => x"77167881",
  1863 => x"0784180c",
  1864 => x"8c170888",
  1865 => x"1808718c",
  1866 => x"120c8812",
  1867 => x"0c5c7080",
  1868 => x"d6d80c70",
  1869 => x"80d6d40c",
  1870 => x"80d6cc0b",
  1871 => x"8c120c8c",
  1872 => x"11088812",
  1873 => x"0c778107",
  1874 => x"84120c77",
  1875 => x"0577710c",
  1876 => x"557c5182",
  1877 => x"9a3f8816",
  1878 => x"54f5ba39",
  1879 => x"72168411",
  1880 => x"08810784",
  1881 => x"120c588c",
  1882 => x"16088817",
  1883 => x"08718c12",
  1884 => x"0c88120c",
  1885 => x"577c5181",
  1886 => x"f63f8816",
  1887 => x"54f59639",
  1888 => x"7284150c",
  1889 => x"f41af806",
  1890 => x"70841d08",
  1891 => x"81060784",
  1892 => x"1d0c701c",
  1893 => x"5556850b",
  1894 => x"84150c85",
  1895 => x"0b88150c",
  1896 => x"8f7627fd",
  1897 => x"ab38881b",
  1898 => x"527c5184",
  1899 => x"c13f80d6",
  1900 => x"c40b8805",
  1901 => x"0880d688",
  1902 => x"085a55fd",
  1903 => x"93397880",
  1904 => x"d6880c73",
  1905 => x"80d6b80c",
  1906 => x"fbef3972",
  1907 => x"84150cfc",
  1908 => x"ff39fb3d",
  1909 => x"0d77707a",
  1910 => x"7c585553",
  1911 => x"568f7527",
  1912 => x"80e63872",
  1913 => x"76078306",
  1914 => x"517080dc",
  1915 => x"38757352",
  1916 => x"54707084",
  1917 => x"05520874",
  1918 => x"70840556",
  1919 => x"0c737170",
  1920 => x"84055308",
  1921 => x"71708405",
  1922 => x"530c7170",
  1923 => x"84055308",
  1924 => x"71708405",
  1925 => x"530c7170",
  1926 => x"84055308",
  1927 => x"71708405",
  1928 => x"530cf016",
  1929 => x"5654748f",
  1930 => x"26c73883",
  1931 => x"75279538",
  1932 => x"70708405",
  1933 => x"52087470",
  1934 => x"8405560c",
  1935 => x"fc155574",
  1936 => x"8326ed38",
  1937 => x"73715452",
  1938 => x"ff155170",
  1939 => x"ff2e9838",
  1940 => x"72708105",
  1941 => x"54337270",
  1942 => x"81055434",
  1943 => x"ff115170",
  1944 => x"ff2e0981",
  1945 => x"06ea3875",
  1946 => x"800c873d",
  1947 => x"0d040404",
  1948 => x"70707070",
  1949 => x"800b81b6",
  1950 => x"9c0c7651",
  1951 => x"87cc3f80",
  1952 => x"08538008",
  1953 => x"ff2e8938",
  1954 => x"72800c50",
  1955 => x"50505004",
  1956 => x"81b69c08",
  1957 => x"5473802e",
  1958 => x"ef387574",
  1959 => x"710c5272",
  1960 => x"800c5050",
  1961 => x"505004fb",
  1962 => x"3d0d7779",
  1963 => x"70720783",
  1964 => x"06535452",
  1965 => x"70933871",
  1966 => x"73730854",
  1967 => x"56547173",
  1968 => x"082e80c4",
  1969 => x"38737554",
  1970 => x"52713370",
  1971 => x"81ff0652",
  1972 => x"5470802e",
  1973 => x"9d387233",
  1974 => x"5570752e",
  1975 => x"09810695",
  1976 => x"38811281",
  1977 => x"14713370",
  1978 => x"81ff0654",
  1979 => x"56545270",
  1980 => x"e5387233",
  1981 => x"557381ff",
  1982 => x"067581ff",
  1983 => x"06717131",
  1984 => x"800c5552",
  1985 => x"873d0d04",
  1986 => x"7109f7fb",
  1987 => x"fdff1306",
  1988 => x"f8848281",
  1989 => x"80065271",
  1990 => x"97388414",
  1991 => x"84167108",
  1992 => x"54565471",
  1993 => x"75082ee0",
  1994 => x"38737554",
  1995 => x"52ff9a39",
  1996 => x"800b800c",
  1997 => x"873d0d04",
  1998 => x"fb3d0d77",
  1999 => x"705256fe",
  2000 => x"ad3f80d6",
  2001 => x"c40b8805",
  2002 => x"08841108",
  2003 => x"fc06707b",
  2004 => x"319fef05",
  2005 => x"e08006e0",
  2006 => x"80055255",
  2007 => x"55a08075",
  2008 => x"24943880",
  2009 => x"527551fe",
  2010 => x"873f80d6",
  2011 => x"cc081453",
  2012 => x"7280082e",
  2013 => x"8f387551",
  2014 => x"fdf53f80",
  2015 => x"5372800c",
  2016 => x"873d0d04",
  2017 => x"74305275",
  2018 => x"51fde53f",
  2019 => x"8008ff2e",
  2020 => x"a83880d6",
  2021 => x"c40b8805",
  2022 => x"08747631",
  2023 => x"81078412",
  2024 => x"0c5380d6",
  2025 => x"88087531",
  2026 => x"80d6880c",
  2027 => x"7551fdbf",
  2028 => x"3f810b80",
  2029 => x"0c873d0d",
  2030 => x"04805275",
  2031 => x"51fdb13f",
  2032 => x"80d6c40b",
  2033 => x"88050880",
  2034 => x"08713154",
  2035 => x"548f7325",
  2036 => x"ffa43880",
  2037 => x"0880d6b8",
  2038 => x"083180d6",
  2039 => x"880c7281",
  2040 => x"0784150c",
  2041 => x"7551fd87",
  2042 => x"3f8053ff",
  2043 => x"9039f73d",
  2044 => x"0d7b7d54",
  2045 => x"5a72802e",
  2046 => x"82833879",
  2047 => x"51fcef3f",
  2048 => x"f8138411",
  2049 => x"0870fe06",
  2050 => x"70138411",
  2051 => x"08fc065c",
  2052 => x"57585457",
  2053 => x"80d6cc08",
  2054 => x"742e82de",
  2055 => x"38778415",
  2056 => x"0c807381",
  2057 => x"06565974",
  2058 => x"792e81d5",
  2059 => x"38771484",
  2060 => x"11088106",
  2061 => x"565374a0",
  2062 => x"38771656",
  2063 => x"7881e638",
  2064 => x"88140855",
  2065 => x"7480d6cc",
  2066 => x"2e82f938",
  2067 => x"8c140870",
  2068 => x"8c170c75",
  2069 => x"88120c58",
  2070 => x"75810784",
  2071 => x"180c7517",
  2072 => x"76710c54",
  2073 => x"78819138",
  2074 => x"83ff7627",
  2075 => x"81c83875",
  2076 => x"892a7683",
  2077 => x"2a545473",
  2078 => x"802ebf38",
  2079 => x"75862ab8",
  2080 => x"05538474",
  2081 => x"27b43880",
  2082 => x"db145394",
  2083 => x"7427ab38",
  2084 => x"758c2a80",
  2085 => x"ee055380",
  2086 => x"d474279e",
  2087 => x"38758f2a",
  2088 => x"80f70553",
  2089 => x"82d47427",
  2090 => x"91387592",
  2091 => x"2a80fc05",
  2092 => x"538ad474",
  2093 => x"27843880",
  2094 => x"fe537210",
  2095 => x"101080d6",
  2096 => x"c4058811",
  2097 => x"08555573",
  2098 => x"752e82bf",
  2099 => x"38841408",
  2100 => x"fc065975",
  2101 => x"79278d38",
  2102 => x"88140854",
  2103 => x"73752e09",
  2104 => x"8106ea38",
  2105 => x"8c140870",
  2106 => x"8c190c74",
  2107 => x"88190c77",
  2108 => x"88120c55",
  2109 => x"768c150c",
  2110 => x"7951faf3",
  2111 => x"3f8b3d0d",
  2112 => x"04760877",
  2113 => x"71315876",
  2114 => x"05881808",
  2115 => x"56567480",
  2116 => x"d6cc2e80",
  2117 => x"e0388c17",
  2118 => x"08708c17",
  2119 => x"0c758812",
  2120 => x"0c53fe89",
  2121 => x"39881408",
  2122 => x"8c150870",
  2123 => x"8c130c59",
  2124 => x"88190cfe",
  2125 => x"a3397583",
  2126 => x"2a705454",
  2127 => x"80742481",
  2128 => x"98387282",
  2129 => x"2c81712b",
  2130 => x"80d6c808",
  2131 => x"0780d6c4",
  2132 => x"0b84050c",
  2133 => x"74101010",
  2134 => x"80d6c405",
  2135 => x"88110871",
  2136 => x"8c1b0c70",
  2137 => x"881b0c79",
  2138 => x"88130c56",
  2139 => x"5a55768c",
  2140 => x"150cff84",
  2141 => x"398159fd",
  2142 => x"b4397716",
  2143 => x"73810654",
  2144 => x"55729838",
  2145 => x"76087771",
  2146 => x"31587505",
  2147 => x"8c180888",
  2148 => x"1908718c",
  2149 => x"120c8812",
  2150 => x"0c555574",
  2151 => x"81078418",
  2152 => x"0c7680d6",
  2153 => x"c40b8805",
  2154 => x"0c80d6c0",
  2155 => x"087526fe",
  2156 => x"c73880d6",
  2157 => x"bc085279",
  2158 => x"51fafd3f",
  2159 => x"7951f9af",
  2160 => x"3ffeba39",
  2161 => x"81778c17",
  2162 => x"0c778817",
  2163 => x"0c758c19",
  2164 => x"0c758819",
  2165 => x"0c59fd80",
  2166 => x"39831470",
  2167 => x"822c8171",
  2168 => x"2b80d6c8",
  2169 => x"080780d6",
  2170 => x"c40b8405",
  2171 => x"0c751010",
  2172 => x"1080d6c4",
  2173 => x"05881108",
  2174 => x"718c1c0c",
  2175 => x"70881c0c",
  2176 => x"7a88130c",
  2177 => x"575b5653",
  2178 => x"fee43980",
  2179 => x"7324a338",
  2180 => x"72822c81",
  2181 => x"712b80d6",
  2182 => x"c8080780",
  2183 => x"d6c40b84",
  2184 => x"050c5874",
  2185 => x"8c180c73",
  2186 => x"88180c76",
  2187 => x"88160cfd",
  2188 => x"c3398313",
  2189 => x"70822c81",
  2190 => x"712b80d6",
  2191 => x"c8080780",
  2192 => x"d6c40b84",
  2193 => x"050c5953",
  2194 => x"da397070",
  2195 => x"7080e5f4",
  2196 => x"08893881",
  2197 => x"b6a00b80",
  2198 => x"e5f40c80",
  2199 => x"e5f40875",
  2200 => x"115252ff",
  2201 => x"537087fb",
  2202 => x"80802688",
  2203 => x"387080e5",
  2204 => x"f40c7153",
  2205 => x"72800c50",
  2206 => x"505004fd",
  2207 => x"3d0d800b",
  2208 => x"80d5f408",
  2209 => x"54547281",
  2210 => x"2e9b3873",
  2211 => x"80e5f80c",
  2212 => x"c3ee3fc2",
  2213 => x"eb3f80e5",
  2214 => x"cc528151",
  2215 => x"cc933f80",
  2216 => x"085180dd",
  2217 => x"3f7280e5",
  2218 => x"f80cc3d4",
  2219 => x"3fc2d13f",
  2220 => x"80e5cc52",
  2221 => x"8151cbf9",
  2222 => x"3f800851",
  2223 => x"80c33f00",
  2224 => x"ff3900ff",
  2225 => x"39f43d0d",
  2226 => x"7e80e5ec",
  2227 => x"08700870",
  2228 => x"81ff0692",
  2229 => x"3df80555",
  2230 => x"515a5759",
  2231 => x"c48f3f80",
  2232 => x"5477557b",
  2233 => x"7d585276",
  2234 => x"538e3df0",
  2235 => x"0551de8e",
  2236 => x"3f797b58",
  2237 => x"790c7684",
  2238 => x"1a0c7880",
  2239 => x"0c8e3d0d",
  2240 => x"04f73d0d",
  2241 => x"7b80decc",
  2242 => x"0882c811",
  2243 => x"085a545a",
  2244 => x"77802e80",
  2245 => x"da388188",
  2246 => x"18841908",
  2247 => x"ff058171",
  2248 => x"2b595559",
  2249 => x"80742480",
  2250 => x"ea388074",
  2251 => x"24b53873",
  2252 => x"822b7811",
  2253 => x"88055656",
  2254 => x"81801908",
  2255 => x"77065372",
  2256 => x"802eb638",
  2257 => x"78167008",
  2258 => x"53537951",
  2259 => x"74085372",
  2260 => x"2dff14fc",
  2261 => x"17fc1779",
  2262 => x"812c5a57",
  2263 => x"57547380",
  2264 => x"25d63877",
  2265 => x"085877ff",
  2266 => x"ad3880de",
  2267 => x"cc0853bc",
  2268 => x"1308a538",
  2269 => x"7951fec7",
  2270 => x"3f740853",
  2271 => x"722dff14",
  2272 => x"fc17fc17",
  2273 => x"79812c5a",
  2274 => x"57575473",
  2275 => x"8025ffa8",
  2276 => x"38d13980",
  2277 => x"57ff9339",
  2278 => x"7251bc13",
  2279 => x"0854732d",
  2280 => x"7951fe9b",
  2281 => x"3f707080",
  2282 => x"e5d40bfc",
  2283 => x"05700852",
  2284 => x"5270ff2e",
  2285 => x"9138702d",
  2286 => x"fc127008",
  2287 => x"525270ff",
  2288 => x"2e098106",
  2289 => x"f1385050",
  2290 => x"0404c2ff",
  2291 => x"3f040000",
  2292 => x"00000040",
  2293 => x"30313233",
  2294 => x"34353637",
  2295 => x"38390000",
  2296 => x"44485259",
  2297 => x"53544f4e",
  2298 => x"45205052",
  2299 => x"4f475241",
  2300 => x"4d2c2053",
  2301 => x"4f4d4520",
  2302 => x"53545249",
  2303 => x"4e470000",
  2304 => x"44485259",
  2305 => x"53544f4e",
  2306 => x"45205052",
  2307 => x"4f475241",
  2308 => x"4d2c2031",
  2309 => x"27535420",
  2310 => x"53545249",
  2311 => x"4e470000",
  2312 => x"44687279",
  2313 => x"73746f6e",
  2314 => x"65204265",
  2315 => x"6e63686d",
  2316 => x"61726b2c",
  2317 => x"20566572",
  2318 => x"73696f6e",
  2319 => x"20322e31",
  2320 => x"20284c61",
  2321 => x"6e677561",
  2322 => x"67653a20",
  2323 => x"43290a00",
  2324 => x"50726f67",
  2325 => x"72616d20",
  2326 => x"636f6d70",
  2327 => x"696c6564",
  2328 => x"20776974",
  2329 => x"68202772",
  2330 => x"65676973",
  2331 => x"74657227",
  2332 => x"20617474",
  2333 => x"72696275",
  2334 => x"74650a00",
  2335 => x"45786563",
  2336 => x"7574696f",
  2337 => x"6e207374",
  2338 => x"61727473",
  2339 => x"2c202564",
  2340 => x"2072756e",
  2341 => x"73207468",
  2342 => x"726f7567",
  2343 => x"68204468",
  2344 => x"72797374",
  2345 => x"6f6e650a",
  2346 => x"00000000",
  2347 => x"44485259",
  2348 => x"53544f4e",
  2349 => x"45205052",
  2350 => x"4f475241",
  2351 => x"4d2c2032",
  2352 => x"274e4420",
  2353 => x"53545249",
  2354 => x"4e470000",
  2355 => x"45786563",
  2356 => x"7574696f",
  2357 => x"6e20656e",
  2358 => x"64730a00",
  2359 => x"46696e61",
  2360 => x"6c207661",
  2361 => x"6c756573",
  2362 => x"206f6620",
  2363 => x"74686520",
  2364 => x"76617269",
  2365 => x"61626c65",
  2366 => x"73207573",
  2367 => x"65642069",
  2368 => x"6e207468",
  2369 => x"65206265",
  2370 => x"6e63686d",
  2371 => x"61726b3a",
  2372 => x"0a000000",
  2373 => x"496e745f",
  2374 => x"476c6f62",
  2375 => x"3a202020",
  2376 => x"20202020",
  2377 => x"20202020",
  2378 => x"2025640a",
  2379 => x"00000000",
  2380 => x"20202020",
  2381 => x"20202020",
  2382 => x"73686f75",
  2383 => x"6c642062",
  2384 => x"653a2020",
  2385 => x"2025640a",
  2386 => x"00000000",
  2387 => x"426f6f6c",
  2388 => x"5f476c6f",
  2389 => x"623a2020",
  2390 => x"20202020",
  2391 => x"20202020",
  2392 => x"2025640a",
  2393 => x"00000000",
  2394 => x"43685f31",
  2395 => x"5f476c6f",
  2396 => x"623a2020",
  2397 => x"20202020",
  2398 => x"20202020",
  2399 => x"2025630a",
  2400 => x"00000000",
  2401 => x"20202020",
  2402 => x"20202020",
  2403 => x"73686f75",
  2404 => x"6c642062",
  2405 => x"653a2020",
  2406 => x"2025630a",
  2407 => x"00000000",
  2408 => x"43685f32",
  2409 => x"5f476c6f",
  2410 => x"623a2020",
  2411 => x"20202020",
  2412 => x"20202020",
  2413 => x"2025630a",
  2414 => x"00000000",
  2415 => x"4172725f",
  2416 => x"315f476c",
  2417 => x"6f625b38",
  2418 => x"5d3a2020",
  2419 => x"20202020",
  2420 => x"2025640a",
  2421 => x"00000000",
  2422 => x"4172725f",
  2423 => x"325f476c",
  2424 => x"6f625b38",
  2425 => x"5d5b375d",
  2426 => x"3a202020",
  2427 => x"2025640a",
  2428 => x"00000000",
  2429 => x"20202020",
  2430 => x"20202020",
  2431 => x"73686f75",
  2432 => x"6c642062",
  2433 => x"653a2020",
  2434 => x"204e756d",
  2435 => x"6265725f",
  2436 => x"4f665f52",
  2437 => x"756e7320",
  2438 => x"2b203130",
  2439 => x"0a000000",
  2440 => x"5074725f",
  2441 => x"476c6f62",
  2442 => x"2d3e0a00",
  2443 => x"20205074",
  2444 => x"725f436f",
  2445 => x"6d703a20",
  2446 => x"20202020",
  2447 => x"20202020",
  2448 => x"2025640a",
  2449 => x"00000000",
  2450 => x"20202020",
  2451 => x"20202020",
  2452 => x"73686f75",
  2453 => x"6c642062",
  2454 => x"653a2020",
  2455 => x"2028696d",
  2456 => x"706c656d",
  2457 => x"656e7461",
  2458 => x"74696f6e",
  2459 => x"2d646570",
  2460 => x"656e6465",
  2461 => x"6e74290a",
  2462 => x"00000000",
  2463 => x"20204469",
  2464 => x"7363723a",
  2465 => x"20202020",
  2466 => x"20202020",
  2467 => x"20202020",
  2468 => x"2025640a",
  2469 => x"00000000",
  2470 => x"2020456e",
  2471 => x"756d5f43",
  2472 => x"6f6d703a",
  2473 => x"20202020",
  2474 => x"20202020",
  2475 => x"2025640a",
  2476 => x"00000000",
  2477 => x"2020496e",
  2478 => x"745f436f",
  2479 => x"6d703a20",
  2480 => x"20202020",
  2481 => x"20202020",
  2482 => x"2025640a",
  2483 => x"00000000",
  2484 => x"20205374",
  2485 => x"725f436f",
  2486 => x"6d703a20",
  2487 => x"20202020",
  2488 => x"20202020",
  2489 => x"2025730a",
  2490 => x"00000000",
  2491 => x"20202020",
  2492 => x"20202020",
  2493 => x"73686f75",
  2494 => x"6c642062",
  2495 => x"653a2020",
  2496 => x"20444852",
  2497 => x"5953544f",
  2498 => x"4e452050",
  2499 => x"524f4752",
  2500 => x"414d2c20",
  2501 => x"534f4d45",
  2502 => x"20535452",
  2503 => x"494e470a",
  2504 => x"00000000",
  2505 => x"4e657874",
  2506 => x"5f507472",
  2507 => x"5f476c6f",
  2508 => x"622d3e0a",
  2509 => x"00000000",
  2510 => x"20202020",
  2511 => x"20202020",
  2512 => x"73686f75",
  2513 => x"6c642062",
  2514 => x"653a2020",
  2515 => x"2028696d",
  2516 => x"706c656d",
  2517 => x"656e7461",
  2518 => x"74696f6e",
  2519 => x"2d646570",
  2520 => x"656e6465",
  2521 => x"6e74292c",
  2522 => x"2073616d",
  2523 => x"65206173",
  2524 => x"2061626f",
  2525 => x"76650a00",
  2526 => x"496e745f",
  2527 => x"315f4c6f",
  2528 => x"633a2020",
  2529 => x"20202020",
  2530 => x"20202020",
  2531 => x"2025640a",
  2532 => x"00000000",
  2533 => x"496e745f",
  2534 => x"325f4c6f",
  2535 => x"633a2020",
  2536 => x"20202020",
  2537 => x"20202020",
  2538 => x"2025640a",
  2539 => x"00000000",
  2540 => x"496e745f",
  2541 => x"335f4c6f",
  2542 => x"633a2020",
  2543 => x"20202020",
  2544 => x"20202020",
  2545 => x"2025640a",
  2546 => x"00000000",
  2547 => x"456e756d",
  2548 => x"5f4c6f63",
  2549 => x"3a202020",
  2550 => x"20202020",
  2551 => x"20202020",
  2552 => x"2025640a",
  2553 => x"00000000",
  2554 => x"5374725f",
  2555 => x"315f4c6f",
  2556 => x"633a2020",
  2557 => x"20202020",
  2558 => x"20202020",
  2559 => x"2025730a",
  2560 => x"00000000",
  2561 => x"20202020",
  2562 => x"20202020",
  2563 => x"73686f75",
  2564 => x"6c642062",
  2565 => x"653a2020",
  2566 => x"20444852",
  2567 => x"5953544f",
  2568 => x"4e452050",
  2569 => x"524f4752",
  2570 => x"414d2c20",
  2571 => x"31275354",
  2572 => x"20535452",
  2573 => x"494e470a",
  2574 => x"00000000",
  2575 => x"5374725f",
  2576 => x"325f4c6f",
  2577 => x"633a2020",
  2578 => x"20202020",
  2579 => x"20202020",
  2580 => x"2025730a",
  2581 => x"00000000",
  2582 => x"20202020",
  2583 => x"20202020",
  2584 => x"73686f75",
  2585 => x"6c642062",
  2586 => x"653a2020",
  2587 => x"20444852",
  2588 => x"5953544f",
  2589 => x"4e452050",
  2590 => x"524f4752",
  2591 => x"414d2c20",
  2592 => x"32274e44",
  2593 => x"20535452",
  2594 => x"494e470a",
  2595 => x"00000000",
  2596 => x"55736572",
  2597 => x"2074696d",
  2598 => x"653a2025",
  2599 => x"640a0000",
  2600 => x"4d696372",
  2601 => x"6f736563",
  2602 => x"6f6e6473",
  2603 => x"20666f72",
  2604 => x"206f6e65",
  2605 => x"2072756e",
  2606 => x"20746872",
  2607 => x"6f756768",
  2608 => x"20446872",
  2609 => x"7973746f",
  2610 => x"6e653a20",
  2611 => x"00000000",
  2612 => x"2564200a",
  2613 => x"00000000",
  2614 => x"44687279",
  2615 => x"73746f6e",
  2616 => x"65732070",
  2617 => x"65722053",
  2618 => x"65636f6e",
  2619 => x"643a2020",
  2620 => x"20202020",
  2621 => x"20202020",
  2622 => x"20202020",
  2623 => x"20202020",
  2624 => x"20202020",
  2625 => x"00000000",
  2626 => x"56415820",
  2627 => x"4d495053",
  2628 => x"20726174",
  2629 => x"696e6720",
  2630 => x"2a203130",
  2631 => x"3030203d",
  2632 => x"20256420",
  2633 => x"0a000000",
  2634 => x"50726f67",
  2635 => x"72616d20",
  2636 => x"636f6d70",
  2637 => x"696c6564",
  2638 => x"20776974",
  2639 => x"686f7574",
  2640 => x"20277265",
  2641 => x"67697374",
  2642 => x"65722720",
  2643 => x"61747472",
  2644 => x"69627574",
  2645 => x"650a0000",
  2646 => x"4d656173",
  2647 => x"75726564",
  2648 => x"2074696d",
  2649 => x"6520746f",
  2650 => x"6f20736d",
  2651 => x"616c6c20",
  2652 => x"746f206f",
  2653 => x"62746169",
  2654 => x"6e206d65",
  2655 => x"616e696e",
  2656 => x"6766756c",
  2657 => x"20726573",
  2658 => x"756c7473",
  2659 => x"0a000000",
  2660 => x"506c6561",
  2661 => x"73652069",
  2662 => x"6e637265",
  2663 => x"61736520",
  2664 => x"6e756d62",
  2665 => x"6572206f",
  2666 => x"66207275",
  2667 => x"6e730a00",
  2668 => x"44485259",
  2669 => x"53544f4e",
  2670 => x"45205052",
  2671 => x"4f475241",
  2672 => x"4d2c2033",
  2673 => x"27524420",
  2674 => x"53545249",
  2675 => x"4e470000",
  2676 => x"00010202",
  2677 => x"03030303",
  2678 => x"04040404",
  2679 => x"04040404",
  2680 => x"05050505",
  2681 => x"05050505",
  2682 => x"05050505",
  2683 => x"05050505",
  2684 => x"06060606",
  2685 => x"06060606",
  2686 => x"06060606",
  2687 => x"06060606",
  2688 => x"06060606",
  2689 => x"06060606",
  2690 => x"06060606",
  2691 => x"06060606",
  2692 => x"07070707",
  2693 => x"07070707",
  2694 => x"07070707",
  2695 => x"07070707",
  2696 => x"07070707",
  2697 => x"07070707",
  2698 => x"07070707",
  2699 => x"07070707",
  2700 => x"07070707",
  2701 => x"07070707",
  2702 => x"07070707",
  2703 => x"07070707",
  2704 => x"07070707",
  2705 => x"07070707",
  2706 => x"07070707",
  2707 => x"07070707",
  2708 => x"08080808",
  2709 => x"08080808",
  2710 => x"08080808",
  2711 => x"08080808",
  2712 => x"08080808",
  2713 => x"08080808",
  2714 => x"08080808",
  2715 => x"08080808",
  2716 => x"08080808",
  2717 => x"08080808",
  2718 => x"08080808",
  2719 => x"08080808",
  2720 => x"08080808",
  2721 => x"08080808",
  2722 => x"08080808",
  2723 => x"08080808",
  2724 => x"08080808",
  2725 => x"08080808",
  2726 => x"08080808",
  2727 => x"08080808",
  2728 => x"08080808",
  2729 => x"08080808",
  2730 => x"08080808",
  2731 => x"08080808",
  2732 => x"08080808",
  2733 => x"08080808",
  2734 => x"08080808",
  2735 => x"08080808",
  2736 => x"08080808",
  2737 => x"08080808",
  2738 => x"08080808",
  2739 => x"08080808",
  2740 => x"43000000",
  2741 => x"64756d6d",
  2742 => x"792e6578",
  2743 => x"65000000",
  2744 => x"00ffffff",
  2745 => x"ff00ffff",
  2746 => x"ffff00ff",
  2747 => x"ffffff00",
  2748 => x"00000000",
  2749 => x"00000000",
  2750 => x"00000000",
  2751 => x"000032dc",
  2752 => x"0000c350",
  2753 => x"00000000",
  2754 => x"00000000",
  2755 => x"00000000",
  2756 => x"00000000",
  2757 => x"00000000",
  2758 => x"00000000",
  2759 => x"00000000",
  2760 => x"00000000",
  2761 => x"00000000",
  2762 => x"00000000",
  2763 => x"00000000",
  2764 => x"00000000",
  2765 => x"00000000",
  2766 => x"ffffffff",
  2767 => x"00000000",
  2768 => x"00020000",
  2769 => x"00000000",
  2770 => x"00000000",
  2771 => x"00002b44",
  2772 => x"00002b44",
  2773 => x"00002b4c",
  2774 => x"00002b4c",
  2775 => x"00002b54",
  2776 => x"00002b54",
  2777 => x"00002b5c",
  2778 => x"00002b5c",
  2779 => x"00002b64",
  2780 => x"00002b64",
  2781 => x"00002b6c",
  2782 => x"00002b6c",
  2783 => x"00002b74",
  2784 => x"00002b74",
  2785 => x"00002b7c",
  2786 => x"00002b7c",
  2787 => x"00002b84",
  2788 => x"00002b84",
  2789 => x"00002b8c",
  2790 => x"00002b8c",
  2791 => x"00002b94",
  2792 => x"00002b94",
  2793 => x"00002b9c",
  2794 => x"00002b9c",
  2795 => x"00002ba4",
  2796 => x"00002ba4",
  2797 => x"00002bac",
  2798 => x"00002bac",
  2799 => x"00002bb4",
  2800 => x"00002bb4",
  2801 => x"00002bbc",
  2802 => x"00002bbc",
  2803 => x"00002bc4",
  2804 => x"00002bc4",
  2805 => x"00002bcc",
  2806 => x"00002bcc",
  2807 => x"00002bd4",
  2808 => x"00002bd4",
  2809 => x"00002bdc",
  2810 => x"00002bdc",
  2811 => x"00002be4",
  2812 => x"00002be4",
  2813 => x"00002bec",
  2814 => x"00002bec",
  2815 => x"00002bf4",
  2816 => x"00002bf4",
  2817 => x"00002bfc",
  2818 => x"00002bfc",
  2819 => x"00002c04",
  2820 => x"00002c04",
  2821 => x"00002c0c",
  2822 => x"00002c0c",
  2823 => x"00002c14",
  2824 => x"00002c14",
  2825 => x"00002c1c",
  2826 => x"00002c1c",
  2827 => x"00002c24",
  2828 => x"00002c24",
  2829 => x"00002c2c",
  2830 => x"00002c2c",
  2831 => x"00002c34",
  2832 => x"00002c34",
  2833 => x"00002c3c",
  2834 => x"00002c3c",
  2835 => x"00002c44",
  2836 => x"00002c44",
  2837 => x"00002c4c",
  2838 => x"00002c4c",
  2839 => x"00002c54",
  2840 => x"00002c54",
  2841 => x"00002c5c",
  2842 => x"00002c5c",
  2843 => x"00002c64",
  2844 => x"00002c64",
  2845 => x"00002c6c",
  2846 => x"00002c6c",
  2847 => x"00002c74",
  2848 => x"00002c74",
  2849 => x"00002c7c",
  2850 => x"00002c7c",
  2851 => x"00002c84",
  2852 => x"00002c84",
  2853 => x"00002c8c",
  2854 => x"00002c8c",
  2855 => x"00002c94",
  2856 => x"00002c94",
  2857 => x"00002c9c",
  2858 => x"00002c9c",
  2859 => x"00002ca4",
  2860 => x"00002ca4",
  2861 => x"00002cac",
  2862 => x"00002cac",
  2863 => x"00002cb4",
  2864 => x"00002cb4",
  2865 => x"00002cbc",
  2866 => x"00002cbc",
  2867 => x"00002cc4",
  2868 => x"00002cc4",
  2869 => x"00002ccc",
  2870 => x"00002ccc",
  2871 => x"00002cd4",
  2872 => x"00002cd4",
  2873 => x"00002cdc",
  2874 => x"00002cdc",
  2875 => x"00002ce4",
  2876 => x"00002ce4",
  2877 => x"00002cec",
  2878 => x"00002cec",
  2879 => x"00002cf4",
  2880 => x"00002cf4",
  2881 => x"00002cfc",
  2882 => x"00002cfc",
  2883 => x"00002d04",
  2884 => x"00002d04",
  2885 => x"00002d0c",
  2886 => x"00002d0c",
  2887 => x"00002d14",
  2888 => x"00002d14",
  2889 => x"00002d1c",
  2890 => x"00002d1c",
  2891 => x"00002d24",
  2892 => x"00002d24",
  2893 => x"00002d2c",
  2894 => x"00002d2c",
  2895 => x"00002d34",
  2896 => x"00002d34",
  2897 => x"00002d3c",
  2898 => x"00002d3c",
  2899 => x"00002d44",
  2900 => x"00002d44",
  2901 => x"00002d4c",
  2902 => x"00002d4c",
  2903 => x"00002d54",
  2904 => x"00002d54",
  2905 => x"00002d5c",
  2906 => x"00002d5c",
  2907 => x"00002d64",
  2908 => x"00002d64",
  2909 => x"00002d6c",
  2910 => x"00002d6c",
  2911 => x"00002d74",
  2912 => x"00002d74",
  2913 => x"00002d7c",
  2914 => x"00002d7c",
  2915 => x"00002d84",
  2916 => x"00002d84",
  2917 => x"00002d8c",
  2918 => x"00002d8c",
  2919 => x"00002d94",
  2920 => x"00002d94",
  2921 => x"00002d9c",
  2922 => x"00002d9c",
  2923 => x"00002da4",
  2924 => x"00002da4",
  2925 => x"00002dac",
  2926 => x"00002dac",
  2927 => x"00002db4",
  2928 => x"00002db4",
  2929 => x"00002dbc",
  2930 => x"00002dbc",
  2931 => x"00002dc4",
  2932 => x"00002dc4",
  2933 => x"00002dcc",
  2934 => x"00002dcc",
  2935 => x"00002dd4",
  2936 => x"00002dd4",
  2937 => x"00002ddc",
  2938 => x"00002ddc",
  2939 => x"00002de4",
  2940 => x"00002de4",
  2941 => x"00002dec",
  2942 => x"00002dec",
  2943 => x"00002df4",
  2944 => x"00002df4",
  2945 => x"00002dfc",
  2946 => x"00002dfc",
  2947 => x"00002e04",
  2948 => x"00002e04",
  2949 => x"00002e0c",
  2950 => x"00002e0c",
  2951 => x"00002e14",
  2952 => x"00002e14",
  2953 => x"00002e1c",
  2954 => x"00002e1c",
  2955 => x"00002e24",
  2956 => x"00002e24",
  2957 => x"00002e2c",
  2958 => x"00002e2c",
  2959 => x"00002e34",
  2960 => x"00002e34",
  2961 => x"00002e3c",
  2962 => x"00002e3c",
  2963 => x"00002e44",
  2964 => x"00002e44",
  2965 => x"00002e4c",
  2966 => x"00002e4c",
  2967 => x"00002e54",
  2968 => x"00002e54",
  2969 => x"00002e5c",
  2970 => x"00002e5c",
  2971 => x"00002e64",
  2972 => x"00002e64",
  2973 => x"00002e6c",
  2974 => x"00002e6c",
  2975 => x"00002e74",
  2976 => x"00002e74",
  2977 => x"00002e7c",
  2978 => x"00002e7c",
  2979 => x"00002e84",
  2980 => x"00002e84",
  2981 => x"00002e8c",
  2982 => x"00002e8c",
  2983 => x"00002e94",
  2984 => x"00002e94",
  2985 => x"00002e9c",
  2986 => x"00002e9c",
  2987 => x"00002ea4",
  2988 => x"00002ea4",
  2989 => x"00002eac",
  2990 => x"00002eac",
  2991 => x"00002eb4",
  2992 => x"00002eb4",
  2993 => x"00002ebc",
  2994 => x"00002ebc",
  2995 => x"00002ec4",
  2996 => x"00002ec4",
  2997 => x"00002ecc",
  2998 => x"00002ecc",
  2999 => x"00002ed4",
  3000 => x"00002ed4",
  3001 => x"00002edc",
  3002 => x"00002edc",
  3003 => x"00002ee4",
  3004 => x"00002ee4",
  3005 => x"00002eec",
  3006 => x"00002eec",
  3007 => x"00002ef4",
  3008 => x"00002ef4",
  3009 => x"00002efc",
  3010 => x"00002efc",
  3011 => x"00002f04",
  3012 => x"00002f04",
  3013 => x"00002f0c",
  3014 => x"00002f0c",
  3015 => x"00002f14",
  3016 => x"00002f14",
  3017 => x"00002f1c",
  3018 => x"00002f1c",
  3019 => x"00002f24",
  3020 => x"00002f24",
  3021 => x"00002f2c",
  3022 => x"00002f2c",
  3023 => x"00002f34",
  3024 => x"00002f34",
  3025 => x"00002f3c",
  3026 => x"00002f3c",
  3027 => x"00002f50",
  3028 => x"00000000",
  3029 => x"000031b8",
  3030 => x"00003214",
  3031 => x"00003270",
  3032 => x"00000000",
  3033 => x"00000000",
  3034 => x"00000000",
  3035 => x"00000000",
  3036 => x"00000000",
  3037 => x"00000000",
  3038 => x"00000000",
  3039 => x"00000000",
  3040 => x"00000000",
  3041 => x"00002ad0",
  3042 => x"00000000",
  3043 => x"00000000",
  3044 => x"00000000",
  3045 => x"00000000",
  3046 => x"00000000",
  3047 => x"00000000",
  3048 => x"00000000",
  3049 => x"00000000",
  3050 => x"00000000",
  3051 => x"00000000",
  3052 => x"00000000",
  3053 => x"00000000",
  3054 => x"00000000",
  3055 => x"00000000",
  3056 => x"00000000",
  3057 => x"00000000",
  3058 => x"00000000",
  3059 => x"00000000",
  3060 => x"00000000",
  3061 => x"00000000",
  3062 => x"00000000",
  3063 => x"00000000",
  3064 => x"00000000",
  3065 => x"00000000",
  3066 => x"00000000",
  3067 => x"00000000",
  3068 => x"00000000",
  3069 => x"00000000",
  3070 => x"00000001",
  3071 => x"330eabcd",
  3072 => x"1234e66d",
  3073 => x"deec0005",
  3074 => x"000b0000",
  3075 => x"00000000",
  3076 => x"00000000",
  3077 => x"00000000",
  3078 => x"00000000",
  3079 => x"00000000",
  3080 => x"00000000",
  3081 => x"00000000",
  3082 => x"00000000",
  3083 => x"00000000",
  3084 => x"00000000",
  3085 => x"00000000",
  3086 => x"00000000",
  3087 => x"00000000",
  3088 => x"00000000",
  3089 => x"00000000",
  3090 => x"00000000",
  3091 => x"00000000",
  3092 => x"00000000",
  3093 => x"00000000",
  3094 => x"00000000",
  3095 => x"00000000",
  3096 => x"00000000",
  3097 => x"00000000",
  3098 => x"00000000",
  3099 => x"00000000",
  3100 => x"00000000",
  3101 => x"00000000",
  3102 => x"00000000",
  3103 => x"00000000",
  3104 => x"00000000",
  3105 => x"00000000",
  3106 => x"00000000",
  3107 => x"00000000",
  3108 => x"00000000",
  3109 => x"00000000",
  3110 => x"00000000",
  3111 => x"00000000",
  3112 => x"00000000",
  3113 => x"00000000",
  3114 => x"00000000",
  3115 => x"00000000",
  3116 => x"00000000",
  3117 => x"00000000",
  3118 => x"00000000",
  3119 => x"00000000",
  3120 => x"00000000",
  3121 => x"00000000",
  3122 => x"00000000",
  3123 => x"00000000",
  3124 => x"00000000",
  3125 => x"00000000",
  3126 => x"00000000",
  3127 => x"00000000",
  3128 => x"00000000",
  3129 => x"00000000",
  3130 => x"00000000",
  3131 => x"00000000",
  3132 => x"00000000",
  3133 => x"00000000",
  3134 => x"00000000",
  3135 => x"00000000",
  3136 => x"00000000",
  3137 => x"00000000",
  3138 => x"00000000",
  3139 => x"00000000",
  3140 => x"00000000",
  3141 => x"00000000",
  3142 => x"00000000",
  3143 => x"00000000",
  3144 => x"00000000",
  3145 => x"00000000",
  3146 => x"00000000",
  3147 => x"00000000",
  3148 => x"00000000",
  3149 => x"00000000",
  3150 => x"00000000",
  3151 => x"00000000",
  3152 => x"00000000",
  3153 => x"00000000",
  3154 => x"00000000",
  3155 => x"00000000",
  3156 => x"00000000",
  3157 => x"00000000",
  3158 => x"00000000",
  3159 => x"00000000",
  3160 => x"00000000",
  3161 => x"00000000",
  3162 => x"00000000",
  3163 => x"00000000",
  3164 => x"00000000",
  3165 => x"00000000",
  3166 => x"00000000",
  3167 => x"00000000",
  3168 => x"00000000",
  3169 => x"00000000",
  3170 => x"00000000",
  3171 => x"00000000",
  3172 => x"00000000",
  3173 => x"00000000",
  3174 => x"00000000",
  3175 => x"00000000",
  3176 => x"00000000",
  3177 => x"00000000",
  3178 => x"00000000",
  3179 => x"00000000",
  3180 => x"00000000",
  3181 => x"00000000",
  3182 => x"00000000",
  3183 => x"00000000",
  3184 => x"00000000",
  3185 => x"00000000",
  3186 => x"00000000",
  3187 => x"00000000",
  3188 => x"00000000",
  3189 => x"00000000",
  3190 => x"00000000",
  3191 => x"00000000",
  3192 => x"00000000",
  3193 => x"00000000",
  3194 => x"00000000",
  3195 => x"00000000",
  3196 => x"00000000",
  3197 => x"00000000",
  3198 => x"00000000",
  3199 => x"00000000",
  3200 => x"00000000",
  3201 => x"00000000",
  3202 => x"00000000",
  3203 => x"00000000",
  3204 => x"00000000",
  3205 => x"00000000",
  3206 => x"00000000",
  3207 => x"00000000",
  3208 => x"00000000",
  3209 => x"00000000",
  3210 => x"00000000",
  3211 => x"00000000",
  3212 => x"00000000",
  3213 => x"00000000",
  3214 => x"00000000",
  3215 => x"00000000",
  3216 => x"00000000",
  3217 => x"00000000",
  3218 => x"00000000",
  3219 => x"00000000",
  3220 => x"00000000",
  3221 => x"00000000",
  3222 => x"00000000",
  3223 => x"00000000",
  3224 => x"00000000",
  3225 => x"00000000",
  3226 => x"00000000",
  3227 => x"00000000",
  3228 => x"00000000",
  3229 => x"00000000",
  3230 => x"00000000",
  3231 => x"00000000",
  3232 => x"00000000",
  3233 => x"00000000",
  3234 => x"00000000",
  3235 => x"00000000",
  3236 => x"00000000",
  3237 => x"00000000",
  3238 => x"00000000",
  3239 => x"00000000",
  3240 => x"00000000",
  3241 => x"00000000",
  3242 => x"00000000",
  3243 => x"00000000",
  3244 => x"00000000",
  3245 => x"00000000",
  3246 => x"00000000",
  3247 => x"00000000",
  3248 => x"00000000",
  3249 => x"00000000",
  3250 => x"00000000",
  3251 => x"00002ad4",
  3252 => x"ffffffff",
  3253 => x"00000000",
  3254 => x"ffffffff",
  3255 => x"00000000",
  3256 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
