-- ZPU
--
-- Copyright 2004-2009 oharboe - Oyvind Harboe - oyvind.harboe@zylin.com
-- 
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library zpu;
use zpu.zpu_config.all;
use zpu.zpupkg.all;

entity dualport_ram is
port (clk : in std_logic;
	memAWriteEnable : in std_logic;
	memAAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memAWrite : in std_logic_vector(wordSize-1 downto 0);
	memARead : out std_logic_vector(wordSize-1 downto 0);
	memBWriteEnable : in std_logic;
	memBAddr : in std_logic_vector(maxAddrBitBRAM downto minAddrBit);
	memBWrite : in std_logic_vector(wordSize-1 downto 0);
	memBRead : out std_logic_vector(wordSize-1 downto 0));
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"82700b0b",
     2 => x"80f0d80c",
     3 => x"3a0b0b80",
     4 => x"e18b0400",
     5 => x"00000000",
     6 => x"00000000",
     7 => x"00000000",
     8 => x"80088408",
     9 => x"88080b0b",
    10 => x"80e1d42d",
    11 => x"880c840c",
    12 => x"800c0400",
    13 => x"00000000",
    14 => x"00000000",
    15 => x"00000000",
    16 => x"71fd0608",
    17 => x"72830609",
    18 => x"81058205",
    19 => x"832b2a83",
    20 => x"ffff0652",
    21 => x"04000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"83ffff73",
    26 => x"83060981",
    27 => x"05820583",
    28 => x"2b2b0906",
    29 => x"7383ffff",
    30 => x"0b0b0b0b",
    31 => x"83a70400",
    32 => x"72098105",
    33 => x"72057373",
    34 => x"09060906",
    35 => x"73097306",
    36 => x"070a8106",
    37 => x"53510400",
    38 => x"00000000",
    39 => x"00000000",
    40 => x"72722473",
    41 => x"732e0753",
    42 => x"51040000",
    43 => x"00000000",
    44 => x"00000000",
    45 => x"00000000",
    46 => x"00000000",
    47 => x"00000000",
    48 => x"71737109",
    49 => x"71068106",
    50 => x"30720a10",
    51 => x"0a720a10",
    52 => x"0a31050a",
    53 => x"81065151",
    54 => x"53510400",
    55 => x"00000000",
    56 => x"72722673",
    57 => x"732e0753",
    58 => x"51040000",
    59 => x"00000000",
    60 => x"00000000",
    61 => x"00000000",
    62 => x"00000000",
    63 => x"00000000",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"00000000",
    67 => x"00000000",
    68 => x"00000000",
    69 => x"00000000",
    70 => x"00000000",
    71 => x"00000000",
    72 => x"0b0b0b88",
    73 => x"c4040000",
    74 => x"00000000",
    75 => x"00000000",
    76 => x"00000000",
    77 => x"00000000",
    78 => x"00000000",
    79 => x"00000000",
    80 => x"720a722b",
    81 => x"0a535104",
    82 => x"00000000",
    83 => x"00000000",
    84 => x"00000000",
    85 => x"00000000",
    86 => x"00000000",
    87 => x"00000000",
    88 => x"72729f06",
    89 => x"0981050b",
    90 => x"0b0b88a7",
    91 => x"05040000",
    92 => x"00000000",
    93 => x"00000000",
    94 => x"00000000",
    95 => x"00000000",
    96 => x"72722aff",
    97 => x"739f062a",
    98 => x"0974090a",
    99 => x"8106ff05",
   100 => x"06075351",
   101 => x"04000000",
   102 => x"00000000",
   103 => x"00000000",
   104 => x"71715351",
   105 => x"020d0406",
   106 => x"73830609",
   107 => x"81058205",
   108 => x"832b0b2b",
   109 => x"0772fc06",
   110 => x"0c515104",
   111 => x"00000000",
   112 => x"72098105",
   113 => x"72050970",
   114 => x"81050906",
   115 => x"0a810653",
   116 => x"51040000",
   117 => x"00000000",
   118 => x"00000000",
   119 => x"00000000",
   120 => x"72098105",
   121 => x"72050970",
   122 => x"81050906",
   123 => x"0a098106",
   124 => x"53510400",
   125 => x"00000000",
   126 => x"00000000",
   127 => x"00000000",
   128 => x"71098105",
   129 => x"52040000",
   130 => x"00000000",
   131 => x"00000000",
   132 => x"00000000",
   133 => x"00000000",
   134 => x"00000000",
   135 => x"00000000",
   136 => x"72720981",
   137 => x"05055351",
   138 => x"04000000",
   139 => x"00000000",
   140 => x"00000000",
   141 => x"00000000",
   142 => x"00000000",
   143 => x"00000000",
   144 => x"72097206",
   145 => x"73730906",
   146 => x"07535104",
   147 => x"00000000",
   148 => x"00000000",
   149 => x"00000000",
   150 => x"00000000",
   151 => x"00000000",
   152 => x"71fc0608",
   153 => x"72830609",
   154 => x"81058305",
   155 => x"1010102a",
   156 => x"81ff0652",
   157 => x"04000000",
   158 => x"00000000",
   159 => x"00000000",
   160 => x"71fc0608",
   161 => x"0b0b80f0",
   162 => x"c4738306",
   163 => x"10100508",
   164 => x"060b0b0b",
   165 => x"88aa0400",
   166 => x"00000000",
   167 => x"00000000",
   168 => x"80088408",
   169 => x"88087575",
   170 => x"0b0b80db",
   171 => x"f62d5050",
   172 => x"80085688",
   173 => x"0c840c80",
   174 => x"0c510400",
   175 => x"00000000",
   176 => x"80088408",
   177 => x"88087575",
   178 => x"0b0b80dd",
   179 => x"a82d5050",
   180 => x"80085688",
   181 => x"0c840c80",
   182 => x"0c510400",
   183 => x"00000000",
   184 => x"72097081",
   185 => x"0509060a",
   186 => x"8106ff05",
   187 => x"70547106",
   188 => x"73097274",
   189 => x"05ff0506",
   190 => x"07515151",
   191 => x"04000000",
   192 => x"72097081",
   193 => x"0509060a",
   194 => x"098106ff",
   195 => x"05705471",
   196 => x"06730972",
   197 => x"7405ff05",
   198 => x"06075151",
   199 => x"51040000",
   200 => x"05ff0504",
   201 => x"00000000",
   202 => x"00000000",
   203 => x"00000000",
   204 => x"00000000",
   205 => x"00000000",
   206 => x"00000000",
   207 => x"00000000",
   208 => x"810b0b0b",
   209 => x"80f0d40c",
   210 => x"51040000",
   211 => x"00000000",
   212 => x"00000000",
   213 => x"00000000",
   214 => x"00000000",
   215 => x"00000000",
   216 => x"71810552",
   217 => x"04000000",
   218 => x"00000000",
   219 => x"00000000",
   220 => x"00000000",
   221 => x"00000000",
   222 => x"00000000",
   223 => x"00000000",
   224 => x"00000000",
   225 => x"00000000",
   226 => x"00000000",
   227 => x"00000000",
   228 => x"00000000",
   229 => x"00000000",
   230 => x"00000000",
   231 => x"00000000",
   232 => x"02840572",
   233 => x"10100552",
   234 => x"04000000",
   235 => x"00000000",
   236 => x"00000000",
   237 => x"00000000",
   238 => x"00000000",
   239 => x"00000000",
   240 => x"00000000",
   241 => x"00000000",
   242 => x"00000000",
   243 => x"00000000",
   244 => x"00000000",
   245 => x"00000000",
   246 => x"00000000",
   247 => x"00000000",
   248 => x"717105ff",
   249 => x"05715351",
   250 => x"020d0400",
   251 => x"00000000",
   252 => x"00000000",
   253 => x"00000000",
   254 => x"00000000",
   255 => x"00000000",
   256 => x"82813f80",
   257 => x"daf53f04",
   258 => x"10101010",
   259 => x"10101010",
   260 => x"10101010",
   261 => x"10101010",
   262 => x"10101010",
   263 => x"10101010",
   264 => x"10101010",
   265 => x"10101053",
   266 => x"51047381",
   267 => x"ff067383",
   268 => x"06098105",
   269 => x"83051010",
   270 => x"102b0772",
   271 => x"fc060c51",
   272 => x"51043c04",
   273 => x"72728072",
   274 => x"8106ff05",
   275 => x"09720605",
   276 => x"71105272",
   277 => x"0a100a53",
   278 => x"72ed3851",
   279 => x"51535104",
   280 => x"80f0d408",
   281 => x"802ea438",
   282 => x"80f0d808",
   283 => x"822ebd38",
   284 => x"8380800b",
   285 => x"0b0b80f8",
   286 => x"980c82a0",
   287 => x"800b80f8",
   288 => x"9c0c8290",
   289 => x"800b80f8",
   290 => x"a00c04f8",
   291 => x"808080a4",
   292 => x"0b0b0b80",
   293 => x"f8980cf8",
   294 => x"80808280",
   295 => x"0b80f89c",
   296 => x"0cf88080",
   297 => x"84800b80",
   298 => x"f8a00c04",
   299 => x"80c0a880",
   300 => x"8c0b0b0b",
   301 => x"80f8980c",
   302 => x"80c0a880",
   303 => x"940b80f8",
   304 => x"9c0c0b0b",
   305 => x"80e3a80b",
   306 => x"80f8a00c",
   307 => x"04ff3d0d",
   308 => x"80f8a433",
   309 => x"5170a738",
   310 => x"80f0e008",
   311 => x"70085252",
   312 => x"70802e94",
   313 => x"38841280",
   314 => x"f0e00c70",
   315 => x"2d80f0e0",
   316 => x"08700852",
   317 => x"5270ee38",
   318 => x"810b80f8",
   319 => x"a434833d",
   320 => x"0d040480",
   321 => x"3d0d0b0b",
   322 => x"80f89408",
   323 => x"802e8e38",
   324 => x"0b0b0b0b",
   325 => x"800b802e",
   326 => x"09810685",
   327 => x"38823d0d",
   328 => x"040b0b80",
   329 => x"f894510b",
   330 => x"0b0bf5d4",
   331 => x"3f823d0d",
   332 => x"0404f83d",
   333 => x"0d7a7c59",
   334 => x"53807356",
   335 => x"57767324",
   336 => x"80de3877",
   337 => x"17548a52",
   338 => x"745180d1",
   339 => x"843f8008",
   340 => x"b0055372",
   341 => x"74348117",
   342 => x"578a5274",
   343 => x"5180d0cc",
   344 => x"3f800855",
   345 => x"8008dc38",
   346 => x"8008779f",
   347 => x"2a187081",
   348 => x"2c5b5656",
   349 => x"8079259e",
   350 => x"387717ff",
   351 => x"05557518",
   352 => x"70335553",
   353 => x"74337334",
   354 => x"73753481",
   355 => x"16ff1656",
   356 => x"56787624",
   357 => x"e9387618",
   358 => x"56807634",
   359 => x"8a3d0d04",
   360 => x"ad787081",
   361 => x"055a3472",
   362 => x"30781855",
   363 => x"558a5274",
   364 => x"5180d09d",
   365 => x"3f8008b0",
   366 => x"05537274",
   367 => x"34811757",
   368 => x"8a527451",
   369 => x"80cfe53f",
   370 => x"80085580",
   371 => x"08fef438",
   372 => x"ff9639f9",
   373 => x"3d0d7970",
   374 => x"71337081",
   375 => x"ff065455",
   376 => x"55557080",
   377 => x"2eb13880",
   378 => x"f0fc0852",
   379 => x"7281ff06",
   380 => x"81155553",
   381 => x"728a2e80",
   382 => x"f5388412",
   383 => x"0870822a",
   384 => x"81065257",
   385 => x"70802ef2",
   386 => x"3872720c",
   387 => x"73337081",
   388 => x"ff065953",
   389 => x"77d63874",
   390 => x"75335256",
   391 => x"70802e80",
   392 => x"c9387080",
   393 => x"f0f40859",
   394 => x"53811680",
   395 => x"f8ac3370",
   396 => x"81ff0670",
   397 => x"10101180",
   398 => x"f8b03370",
   399 => x"81ff0672",
   400 => x"90291170",
   401 => x"882b7a07",
   402 => x"7f0c5359",
   403 => x"59545458",
   404 => x"56728a2e",
   405 => x"be387380",
   406 => x"cf2eb838",
   407 => x"81155372",
   408 => x"80f8b034",
   409 => x"75335372",
   410 => x"c038893d",
   411 => x"0d048412",
   412 => x"0870822a",
   413 => x"81065758",
   414 => x"75802ef2",
   415 => x"388d720c",
   416 => x"84120870",
   417 => x"822a8106",
   418 => x"52577080",
   419 => x"2efeeb38",
   420 => x"fef73971",
   421 => x"a3269938",
   422 => x"81175271",
   423 => x"80f8ac34",
   424 => x"800b80f8",
   425 => x"b0347533",
   426 => x"5372fefd",
   427 => x"38ffbb39",
   428 => x"800b80f8",
   429 => x"ac34800b",
   430 => x"80f8b034",
   431 => x"e939fd3d",
   432 => x"0d80f0f0",
   433 => x"085480d5",
   434 => x"0b84150c",
   435 => x"80f0fc08",
   436 => x"52841208",
   437 => x"81065170",
   438 => x"802ef638",
   439 => x"71087081",
   440 => x"ff06f611",
   441 => x"52545170",
   442 => x"ae268c38",
   443 => x"70101080",
   444 => x"eec40551",
   445 => x"70080484",
   446 => x"12087082",
   447 => x"2a708106",
   448 => x"51515170",
   449 => x"802ef038",
   450 => x"ab720c72",
   451 => x"8a2eaa38",
   452 => x"84120870",
   453 => x"822a7081",
   454 => x"06515151",
   455 => x"70802ef0",
   456 => x"3872720c",
   457 => x"84120870",
   458 => x"822a8106",
   459 => x"51537280",
   460 => x"2ef238ad",
   461 => x"720cff99",
   462 => x"39841208",
   463 => x"70822a70",
   464 => x"81065151",
   465 => x"5170802e",
   466 => x"f0388d72",
   467 => x"0c841208",
   468 => x"70822a70",
   469 => x"81065151",
   470 => x"5170802e",
   471 => x"ffb238c1",
   472 => x"3981ff0b",
   473 => x"84150cfe",
   474 => x"e83980ff",
   475 => x"0b84150c",
   476 => x"fedf39bf",
   477 => x"0b84150c",
   478 => x"fed7399f",
   479 => x"0b84150c",
   480 => x"fecf398f",
   481 => x"0b84150c",
   482 => x"fec73987",
   483 => x"0b84150c",
   484 => x"febf3983",
   485 => x"0b84150c",
   486 => x"feb73981",
   487 => x"0b84150c",
   488 => x"feaf3980",
   489 => x"0b84150c",
   490 => x"fea739d7",
   491 => x"3d0d80f0",
   492 => x"f4085580",
   493 => x"0b84160c",
   494 => x"fe800a0b",
   495 => x"88160c80",
   496 => x"0b80f8ac",
   497 => x"34800b80",
   498 => x"f8b034a6",
   499 => x"3d705380",
   500 => x"f0e8088c",
   501 => x"11085355",
   502 => x"5bfad73f",
   503 => x"80e6d40b",
   504 => x"80e6d433",
   505 => x"555a7380",
   506 => x"2e80cc38",
   507 => x"80f0f408",
   508 => x"74575c81",
   509 => x"1a80f8ac",
   510 => x"337081ff",
   511 => x"06701010",
   512 => x"1180f8b0",
   513 => x"337081ff",
   514 => x"06729029",
   515 => x"1170882b",
   516 => x"7d07630c",
   517 => x"445c5c42",
   518 => x"575a5a75",
   519 => x"8a2e87be",
   520 => x"387680cf",
   521 => x"2e87b738",
   522 => x"81185776",
   523 => x"80f8b034",
   524 => x"79335675",
   525 => x"ffbd387a",
   526 => x"7b33555a",
   527 => x"73802e80",
   528 => x"cc3880f0",
   529 => x"f4087457",
   530 => x"5b811a80",
   531 => x"f8ac3370",
   532 => x"81ff0670",
   533 => x"10101180",
   534 => x"f8b03370",
   535 => x"81ff0672",
   536 => x"90291170",
   537 => x"882b7d07",
   538 => x"620c465c",
   539 => x"5c44575a",
   540 => x"5a758a2e",
   541 => x"87863876",
   542 => x"80cf2e86",
   543 => x"ff388118",
   544 => x"597880f8",
   545 => x"b0347933",
   546 => x"5675ffbd",
   547 => x"3880e6ec",
   548 => x"0b80e6ec",
   549 => x"33555a73",
   550 => x"802e80cc",
   551 => x"3880f0f4",
   552 => x"0874575b",
   553 => x"811a80f8",
   554 => x"ac337081",
   555 => x"ff067010",
   556 => x"101180f8",
   557 => x"b0337081",
   558 => x"ff067290",
   559 => x"29117088",
   560 => x"2b7d0762",
   561 => x"0c495c5c",
   562 => x"57575a5a",
   563 => x"758a2e85",
   564 => x"ef387680",
   565 => x"cf2e85e8",
   566 => x"3881185d",
   567 => x"7c80f8b0",
   568 => x"34793356",
   569 => x"75ffbd38",
   570 => x"80f0e808",
   571 => x"7008a53d",
   572 => x"5b575a8b",
   573 => x"5380e3ac",
   574 => x"52785180",
   575 => x"cdf43f82",
   576 => x"02840581",
   577 => x"89055957",
   578 => x"758f0654",
   579 => x"73892685",
   580 => x"93387618",
   581 => x"b0155555",
   582 => x"73753475",
   583 => x"842aff18",
   584 => x"7081ff06",
   585 => x"595c5676",
   586 => x"df387879",
   587 => x"33555a73",
   588 => x"802e80cc",
   589 => x"3880f0f4",
   590 => x"0874575b",
   591 => x"811a80f8",
   592 => x"ac337081",
   593 => x"ff067010",
   594 => x"101180f8",
   595 => x"b0337081",
   596 => x"ff067290",
   597 => x"29117088",
   598 => x"2b7d0762",
   599 => x"0c455c5c",
   600 => x"5f575a5a",
   601 => x"758a2e87",
   602 => x"f4387680",
   603 => x"cf2e87ed",
   604 => x"38811857",
   605 => x"7680f8b0",
   606 => x"34793356",
   607 => x"75ffbd38",
   608 => x"80e6f80b",
   609 => x"80e6f833",
   610 => x"555a7380",
   611 => x"2e80cc38",
   612 => x"80f0f408",
   613 => x"74575b81",
   614 => x"1a80f8ac",
   615 => x"337081ff",
   616 => x"06701010",
   617 => x"1180f8b0",
   618 => x"337081ff",
   619 => x"06729029",
   620 => x"1170882b",
   621 => x"7d07620c",
   622 => x"475c5c45",
   623 => x"575a5a75",
   624 => x"8a2e87b7",
   625 => x"387680cf",
   626 => x"2e87b038",
   627 => x"81185978",
   628 => x"80f8b034",
   629 => x"79335675",
   630 => x"ffbd3880",
   631 => x"5f890a5c",
   632 => x"ac3d087f",
   633 => x"2e098106",
   634 => x"87cb387e",
   635 => x"a13d0288",
   636 => x"0580fd05",
   637 => x"40415d7c",
   638 => x"bf064362",
   639 => x"85d53880",
   640 => x"e6cc0b80",
   641 => x"e6cc3355",
   642 => x"5a73802e",
   643 => x"80cc3880",
   644 => x"f0f40874",
   645 => x"575b811a",
   646 => x"80f8ac33",
   647 => x"7081ff06",
   648 => x"70101011",
   649 => x"80f8b033",
   650 => x"7081ff06",
   651 => x"72902911",
   652 => x"70882b7d",
   653 => x"07620c47",
   654 => x"5c5c4557",
   655 => x"5a5a758a",
   656 => x"2e848b38",
   657 => x"7680cf2e",
   658 => x"84843881",
   659 => x"18567580",
   660 => x"f8b03479",
   661 => x"335675ff",
   662 => x"bd387b56",
   663 => x"8b5380e3",
   664 => x"ac527f51",
   665 => x"80cb8b3f",
   666 => x"8857758f",
   667 => x"06547389",
   668 => x"2683d238",
   669 => x"761eb015",
   670 => x"55557375",
   671 => x"3475842a",
   672 => x"ff187081",
   673 => x"ff06595b",
   674 => x"5676df38",
   675 => x"7f603355",
   676 => x"5a73802e",
   677 => x"85bf3880",
   678 => x"f0f40874",
   679 => x"575b811a",
   680 => x"80f8ac33",
   681 => x"7081ff06",
   682 => x"70101011",
   683 => x"80f8b033",
   684 => x"7081ff06",
   685 => x"72902911",
   686 => x"70882b7d",
   687 => x"07620c5a",
   688 => x"5c5c4457",
   689 => x"5a5a758a",
   690 => x"2e83bf38",
   691 => x"7680cf2e",
   692 => x"83b83881",
   693 => x"18597880",
   694 => x"f8b03479",
   695 => x"335675ff",
   696 => x"bd3880e6",
   697 => x"fc0b80e6",
   698 => x"fc33555a",
   699 => x"73802e80",
   700 => x"c7387356",
   701 => x"811a80f8",
   702 => x"ac337081",
   703 => x"ff067010",
   704 => x"101180f8",
   705 => x"b0337081",
   706 => x"ff067290",
   707 => x"29117088",
   708 => x"2b7d0762",
   709 => x"0c495c5c",
   710 => x"57575a5a",
   711 => x"758a2e82",
   712 => x"cb387680",
   713 => x"cf2e82c4",
   714 => x"38811855",
   715 => x"7480f8b0",
   716 => x"34793356",
   717 => x"75ffbd38",
   718 => x"7b087c32",
   719 => x"70307107",
   720 => x"709f2a70",
   721 => x"81ff06b0",
   722 => x"117081ff",
   723 => x"0680f8ac",
   724 => x"337081ff",
   725 => x"06701010",
   726 => x"1180f8b0",
   727 => x"337081ff",
   728 => x"06729029",
   729 => x"1170882b",
   730 => x"7707670c",
   731 => x"4e58595c",
   732 => x"535f465a",
   733 => x"52595b58",
   734 => x"608a2e83",
   735 => x"a4387680",
   736 => x"cf2e839d",
   737 => x"38811841",
   738 => x"6080f8b0",
   739 => x"34791f84",
   740 => x"1d811f5f",
   741 => x"5d5f8fff",
   742 => x"7d27fcdb",
   743 => x"387e800c",
   744 => x"ab3d0d04",
   745 => x"7618b715",
   746 => x"55557375",
   747 => x"3475842a",
   748 => x"ff187081",
   749 => x"ff06595c",
   750 => x"5676facc",
   751 => x"38faeb39",
   752 => x"74a32680",
   753 => x"f1388119",
   754 => x"557480f8",
   755 => x"ac34800b",
   756 => x"80f8b034",
   757 => x"79335675",
   758 => x"f9ca38fa",
   759 => x"8b3974a3",
   760 => x"2680c438",
   761 => x"81195675",
   762 => x"80f8ac34",
   763 => x"800b80f8",
   764 => x"b0347933",
   765 => x"5675f7fb",
   766 => x"38f8bc39",
   767 => x"74a32699",
   768 => x"38811958",
   769 => x"7780f8ac",
   770 => x"34800b80",
   771 => x"f8b03479",
   772 => x"335675f8",
   773 => x"b438f8f5",
   774 => x"39800b80",
   775 => x"f8ac3480",
   776 => x"0b80f8b0",
   777 => x"34e93980",
   778 => x"0b80f8ac",
   779 => x"34800b80",
   780 => x"f8b034ff",
   781 => x"bd39800b",
   782 => x"80f8ac34",
   783 => x"800b80f8",
   784 => x"b034ff90",
   785 => x"39761eb7",
   786 => x"155555fc",
   787 => x"ad3974a3",
   788 => x"2680f138",
   789 => x"81195574",
   790 => x"80f8ac34",
   791 => x"800b80f8",
   792 => x"b0347933",
   793 => x"5675fbae",
   794 => x"38fbef39",
   795 => x"74a32680",
   796 => x"c4388119",
   797 => x"587780f8",
   798 => x"ac34800b",
   799 => x"80f8b034",
   800 => x"79335675",
   801 => x"fcee38fd",
   802 => x"af3974a3",
   803 => x"26993881",
   804 => x"19577680",
   805 => x"f8ac3480",
   806 => x"0b80f8b0",
   807 => x"34793356",
   808 => x"75fbfb38",
   809 => x"fcbc3980",
   810 => x"0b80f8ac",
   811 => x"34800b80",
   812 => x"f8b034e9",
   813 => x"39800b80",
   814 => x"f8ac3480",
   815 => x"0b80f8b0",
   816 => x"34ffbd39",
   817 => x"800b80f8",
   818 => x"ac34800b",
   819 => x"80f8b034",
   820 => x"ff903980",
   821 => x"f0f4087c",
   822 => x"087d3270",
   823 => x"30710770",
   824 => x"9f2a7081",
   825 => x"ff06b011",
   826 => x"7081ff06",
   827 => x"80f8ac33",
   828 => x"7081ff06",
   829 => x"70101011",
   830 => x"80f8b033",
   831 => x"7081ff06",
   832 => x"72902911",
   833 => x"70882b77",
   834 => x"077d0c4f",
   835 => x"58595d53",
   836 => x"40475b52",
   837 => x"5a5c595b",
   838 => x"608a2e09",
   839 => x"8106fcde",
   840 => x"3875a326",
   841 => x"a2388119",
   842 => x"5b7a80f8",
   843 => x"ac34800b",
   844 => x"80f8b034",
   845 => x"791f841d",
   846 => x"811f5f5d",
   847 => x"5f8fff7d",
   848 => x"27f9b438",
   849 => x"fcd73980",
   850 => x"0b80f8ac",
   851 => x"34800b80",
   852 => x"f8b034e0",
   853 => x"3980f0f4",
   854 => x"085bfb86",
   855 => x"3974a326",
   856 => x"80c43881",
   857 => x"19567580",
   858 => x"f8ac3480",
   859 => x"0b80f8b0",
   860 => x"34793356",
   861 => x"75f7c538",
   862 => x"f8863974",
   863 => x"a3269938",
   864 => x"81195877",
   865 => x"80f8ac34",
   866 => x"800b80f8",
   867 => x"b0347933",
   868 => x"5675f883",
   869 => x"38f8c439",
   870 => x"800b80f8",
   871 => x"ac34800b",
   872 => x"80f8b034",
   873 => x"e939800b",
   874 => x"80f8ac34",
   875 => x"800b80f8",
   876 => x"b034ffbd",
   877 => x"397b7f9f",
   878 => x"3d028c05",
   879 => x"80f10598",
   880 => x"3d029405",
   881 => x"80cd0545",
   882 => x"42454344",
   883 => x"5d80e6cc",
   884 => x"0b80e6cc",
   885 => x"33555a73",
   886 => x"802e80cc",
   887 => x"3880f0f4",
   888 => x"0874575b",
   889 => x"811a80f8",
   890 => x"ac337081",
   891 => x"ff067010",
   892 => x"101180f8",
   893 => x"b0337081",
   894 => x"ff067290",
   895 => x"29117088",
   896 => x"2b7d0762",
   897 => x"0c5a5c5c",
   898 => x"5f575a5a",
   899 => x"758a2e84",
   900 => x"85387680",
   901 => x"cf2e83fe",
   902 => x"38811857",
   903 => x"7680f8b0",
   904 => x"34793356",
   905 => x"75ffbd38",
   906 => x"7c568b53",
   907 => x"80e3ac52",
   908 => x"605180c3",
   909 => x"bd3f8857",
   910 => x"758f0654",
   911 => x"73892683",
   912 => x"cc386117",
   913 => x"b0155555",
   914 => x"73753475",
   915 => x"842aff18",
   916 => x"7081ff06",
   917 => x"595b5676",
   918 => x"df386061",
   919 => x"33555a73",
   920 => x"802e84e4",
   921 => x"3880f0f4",
   922 => x"0874575b",
   923 => x"811a80f8",
   924 => x"ac337081",
   925 => x"ff067010",
   926 => x"101180f8",
   927 => x"b0337081",
   928 => x"ff067290",
   929 => x"29117088",
   930 => x"2b7d0762",
   931 => x"0c425c5c",
   932 => x"57575a5a",
   933 => x"758a2e83",
   934 => x"9b387680",
   935 => x"cf2e8394",
   936 => x"38811859",
   937 => x"7880f8b0",
   938 => x"34793356",
   939 => x"75ffbd38",
   940 => x"80f8ac33",
   941 => x"7081ff06",
   942 => x"70101011",
   943 => x"80f8b033",
   944 => x"7081ff06",
   945 => x"72902911",
   946 => x"70882ba0",
   947 => x"07610c41",
   948 => x"595a5657",
   949 => x"587480cf",
   950 => x"2e84a138",
   951 => x"81175675",
   952 => x"80f8b034",
   953 => x"7c087058",
   954 => x"5ca35380",
   955 => x"e3b8527d",
   956 => x"5180c1fe",
   957 => x"3fa0567f",
   958 => x"1677b106",
   959 => x"b0075659",
   960 => x"74793476",
   961 => x"0a100aff",
   962 => x"177081ff",
   963 => x"06585957",
   964 => x"75e5387d",
   965 => x"7e33555a",
   966 => x"73802e84",
   967 => x"883880f0",
   968 => x"f4087457",
   969 => x"5b811a80",
   970 => x"f8ac3370",
   971 => x"81ff0670",
   972 => x"10101180",
   973 => x"f8b03370",
   974 => x"81ff0672",
   975 => x"90291170",
   976 => x"882b7d07",
   977 => x"620c535c",
   978 => x"5c57575a",
   979 => x"5a758a2e",
   980 => x"82803876",
   981 => x"80cf2e81",
   982 => x"f9388118",
   983 => x"567580f8",
   984 => x"b0347933",
   985 => x"5675ffbd",
   986 => x"3880f8ac",
   987 => x"337081ff",
   988 => x"06701010",
   989 => x"1180f8b0",
   990 => x"337081ff",
   991 => x"06729029",
   992 => x"1170882b",
   993 => x"a007610c",
   994 => x"5a5e5a56",
   995 => x"57587980",
   996 => x"cf2e83c5",
   997 => x"38811758",
   998 => x"7780f8b0",
   999 => x"347c7c2e",
  1000 => x"83d43880",
  1001 => x"e7800b80",
  1002 => x"e7803355",
  1003 => x"5a73802e",
  1004 => x"80c73873",
  1005 => x"56811a80",
  1006 => x"f8ac3370",
  1007 => x"81ff0670",
  1008 => x"10101180",
  1009 => x"f8b03370",
  1010 => x"81ff0672",
  1011 => x"90291170",
  1012 => x"882b7d07",
  1013 => x"620c425c",
  1014 => x"5c57575a",
  1015 => x"5a758a2e",
  1016 => x"818d3876",
  1017 => x"80cf2e81",
  1018 => x"86388118",
  1019 => x"577680f8",
  1020 => x"b0347933",
  1021 => x"5675ffbd",
  1022 => x"38841d63",
  1023 => x"8105445d",
  1024 => x"9f6327fb",
  1025 => x"c8387e80",
  1026 => x"0cab3d0d",
  1027 => x"046117b7",
  1028 => x"155555fc",
  1029 => x"b33974a3",
  1030 => x"26818038",
  1031 => x"81195675",
  1032 => x"80f8ac34",
  1033 => x"800b80f8",
  1034 => x"b0347933",
  1035 => x"5675fbb4",
  1036 => x"38fbf539",
  1037 => x"74a32680",
  1038 => x"f1388119",
  1039 => x"587780f8",
  1040 => x"ac34800b",
  1041 => x"80f8b034",
  1042 => x"79335675",
  1043 => x"fc9e38fc",
  1044 => x"df3974a3",
  1045 => x"26b73881",
  1046 => x"19577680",
  1047 => x"f8ac3480",
  1048 => x"0b80f8b0",
  1049 => x"34793356",
  1050 => x"75fdba38",
  1051 => x"fdfb3974",
  1052 => x"a32680c5",
  1053 => x"38811955",
  1054 => x"7480f8ac",
  1055 => x"34800b80",
  1056 => x"f8b03479",
  1057 => x"335675fe",
  1058 => x"ac38feed",
  1059 => x"39800b80",
  1060 => x"f8ac3480",
  1061 => x"0b80f8b0",
  1062 => x"34cb3980",
  1063 => x"0b80f8ac",
  1064 => x"34800b80",
  1065 => x"f8b034ff",
  1066 => x"8139800b",
  1067 => x"80f8ac34",
  1068 => x"800b80f8",
  1069 => x"b034ff90",
  1070 => x"39800b80",
  1071 => x"f8ac3480",
  1072 => x"0b80f8b0",
  1073 => x"34ffbc39",
  1074 => x"80f0f408",
  1075 => x"80f8ac33",
  1076 => x"7081ff06",
  1077 => x"70101011",
  1078 => x"80f8b033",
  1079 => x"7081ff06",
  1080 => x"72902911",
  1081 => x"70882ba0",
  1082 => x"07770c42",
  1083 => x"5a5b5758",
  1084 => x"595b7480",
  1085 => x"cf2e0981",
  1086 => x"06fbe138",
  1087 => x"75a32682",
  1088 => x"b8388118",
  1089 => x"5b7a80f8",
  1090 => x"ac34800b",
  1091 => x"80f8b034",
  1092 => x"7c087058",
  1093 => x"5ca35380",
  1094 => x"e3b8527d",
  1095 => x"51bdd33f",
  1096 => x"a056fbd3",
  1097 => x"3980f0f4",
  1098 => x"0880f8ac",
  1099 => x"337081ff",
  1100 => x"06701010",
  1101 => x"1180f8b0",
  1102 => x"337081ff",
  1103 => x"06729029",
  1104 => x"1170882b",
  1105 => x"a007770c",
  1106 => x"5b5f5b57",
  1107 => x"58595b79",
  1108 => x"80cf2e09",
  1109 => x"8106fcbd",
  1110 => x"3875a326",
  1111 => x"81cc3881",
  1112 => x"18577680",
  1113 => x"f8ac3480",
  1114 => x"0b80f8b0",
  1115 => x"347c7c2e",
  1116 => x"098106fc",
  1117 => x"ae3880e7",
  1118 => x"880b80e7",
  1119 => x"8833555a",
  1120 => x"73802efc",
  1121 => x"f4387381",
  1122 => x"1b80f8ac",
  1123 => x"337081ff",
  1124 => x"06701010",
  1125 => x"1180f8b0",
  1126 => x"337081ff",
  1127 => x"06729029",
  1128 => x"1170882b",
  1129 => x"7807630c",
  1130 => x"5b5d5d40",
  1131 => x"585b5b56",
  1132 => x"758a2e80",
  1133 => x"ca387680",
  1134 => x"cf2e80c3",
  1135 => x"38811859",
  1136 => x"7880f8b0",
  1137 => x"34793356",
  1138 => x"75802efc",
  1139 => x"ac38811a",
  1140 => x"80f8ac33",
  1141 => x"7081ff06",
  1142 => x"70101011",
  1143 => x"80f8b033",
  1144 => x"7081ff06",
  1145 => x"72902911",
  1146 => x"70882b7d",
  1147 => x"07620c5a",
  1148 => x"5c5c5f57",
  1149 => x"5a5a758a",
  1150 => x"2e098106",
  1151 => x"ffb83874",
  1152 => x"a3269938",
  1153 => x"81195675",
  1154 => x"80f8ac34",
  1155 => x"800b80f8",
  1156 => x"b0347933",
  1157 => x"5675ffb6",
  1158 => x"38fbde39",
  1159 => x"800b80f8",
  1160 => x"ac34800b",
  1161 => x"80f8b034",
  1162 => x"e939800b",
  1163 => x"80f8ac34",
  1164 => x"800b80f8",
  1165 => x"b034feb5",
  1166 => x"39800b80",
  1167 => x"f8ac3480",
  1168 => x"0b80f8b0",
  1169 => x"34fdc939",
  1170 => x"dd3d0d80",
  1171 => x"e79051e7",
  1172 => x"823f80f0",
  1173 => x"e4087008",
  1174 => x"80e7a053",
  1175 => x"5d55e6f3",
  1176 => x"3fa03d70",
  1177 => x"537c81ff",
  1178 => x"ff06525d",
  1179 => x"e5c43f7c",
  1180 => x"51e6e03f",
  1181 => x"80e7b451",
  1182 => x"e6d93f7b",
  1183 => x"8f2a8106",
  1184 => x"9e3d5a56",
  1185 => x"8b5380e3",
  1186 => x"ac527851",
  1187 => x"bae43f82",
  1188 => x"02840580",
  1189 => x"f1055957",
  1190 => x"758f0654",
  1191 => x"73892687",
  1192 => x"fc387618",
  1193 => x"b0155555",
  1194 => x"73753475",
  1195 => x"842aff18",
  1196 => x"7081ff06",
  1197 => x"595b5676",
  1198 => x"df387879",
  1199 => x"33555773",
  1200 => x"802ea938",
  1201 => x"7380f0fc",
  1202 => x"08565681",
  1203 => x"1757758a",
  1204 => x"2e87e638",
  1205 => x"84150870",
  1206 => x"822a8106",
  1207 => x"5b5b7980",
  1208 => x"2ef23875",
  1209 => x"750c7633",
  1210 => x"5675e038",
  1211 => x"78793355",
  1212 => x"5a73802e",
  1213 => x"80cc3873",
  1214 => x"80f0f408",
  1215 => x"5c56811a",
  1216 => x"80f8ac33",
  1217 => x"7081ff06",
  1218 => x"70101011",
  1219 => x"80f8b033",
  1220 => x"7081ff06",
  1221 => x"72902911",
  1222 => x"70882b7d",
  1223 => x"07620c53",
  1224 => x"5c5c5757",
  1225 => x"5a5a758a",
  1226 => x"2e87cf38",
  1227 => x"7680cf2e",
  1228 => x"87c83881",
  1229 => x"18577680",
  1230 => x"f8b03479",
  1231 => x"335675ff",
  1232 => x"bd3880e7",
  1233 => x"c851e58b",
  1234 => x"3f7b902a",
  1235 => x"81069b3d",
  1236 => x"5a568b53",
  1237 => x"80e3ac52",
  1238 => x"7851b996",
  1239 => x"3f820284",
  1240 => x"0580e505",
  1241 => x"5957758f",
  1242 => x"06547389",
  1243 => x"2686ef38",
  1244 => x"7618b015",
  1245 => x"55557375",
  1246 => x"3475842a",
  1247 => x"ff187081",
  1248 => x"ff065956",
  1249 => x"5676df38",
  1250 => x"78793355",
  1251 => x"5773802e",
  1252 => x"a93880f0",
  1253 => x"fc087457",
  1254 => x"55811757",
  1255 => x"758a2e87",
  1256 => x"84388415",
  1257 => x"0870822a",
  1258 => x"81065558",
  1259 => x"73802ef2",
  1260 => x"3875750c",
  1261 => x"76335675",
  1262 => x"e0387879",
  1263 => x"33555a73",
  1264 => x"802e80cc",
  1265 => x"3880f0f4",
  1266 => x"0874575b",
  1267 => x"811a80f8",
  1268 => x"ac337081",
  1269 => x"ff067010",
  1270 => x"101180f8",
  1271 => x"b0337081",
  1272 => x"ff067290",
  1273 => x"29117088",
  1274 => x"2b7d0762",
  1275 => x"0c535c5c",
  1276 => x"57575a5a",
  1277 => x"758a2e8f",
  1278 => x"d7387680",
  1279 => x"cf2e8fd0",
  1280 => x"38811857",
  1281 => x"7680f8b0",
  1282 => x"34793356",
  1283 => x"75ffbd38",
  1284 => x"80e7dc51",
  1285 => x"e3bd3f7b",
  1286 => x"952a8306",
  1287 => x"5473812e",
  1288 => x"90bd3881",
  1289 => x"7426908f",
  1290 => x"3873822e",
  1291 => x"90cf3873",
  1292 => x"832e8ce7",
  1293 => x"3880e7f0",
  1294 => x"51e3983f",
  1295 => x"7c527b97",
  1296 => x"2a870683",
  1297 => x"0581712b",
  1298 => x"525ae1e6",
  1299 => x"3f7c51e3",
  1300 => x"823f80e8",
  1301 => x"8451e2fb",
  1302 => x"3f80e88c",
  1303 => x"51e2f43f",
  1304 => x"7c527b9a",
  1305 => x"2a810681",
  1306 => x"0551e1c6",
  1307 => x"3f7c51e2",
  1308 => x"e23f80e8",
  1309 => x"a051e2db",
  1310 => x"3f7c527b",
  1311 => x"9b2a8706",
  1312 => x"830551e1",
  1313 => x"ad3f7c51",
  1314 => x"e2c93f80",
  1315 => x"e8b451e2",
  1316 => x"c23f7c52",
  1317 => x"7b9e2a82",
  1318 => x"0751e196",
  1319 => x"3f7c51e2",
  1320 => x"b23f80e8",
  1321 => x"c851e2ab",
  1322 => x"3f7b9f2a",
  1323 => x"983d5a56",
  1324 => x"8b5380e3",
  1325 => x"ac527851",
  1326 => x"b6b83f82",
  1327 => x"02840580",
  1328 => x"d9055957",
  1329 => x"758f0654",
  1330 => x"7389268c",
  1331 => x"e7387618",
  1332 => x"b0155555",
  1333 => x"73753475",
  1334 => x"842aff18",
  1335 => x"7081ff06",
  1336 => x"595d5676",
  1337 => x"df387879",
  1338 => x"33555773",
  1339 => x"802ea938",
  1340 => x"80f0fc08",
  1341 => x"74575581",
  1342 => x"1757758a",
  1343 => x"2e84cb38",
  1344 => x"84150870",
  1345 => x"822a8106",
  1346 => x"59547780",
  1347 => x"2ef23875",
  1348 => x"750c7633",
  1349 => x"5675e038",
  1350 => x"78793355",
  1351 => x"5a73802e",
  1352 => x"80cc3880",
  1353 => x"f0f40874",
  1354 => x"575b811a",
  1355 => x"80f8ac33",
  1356 => x"7081ff06",
  1357 => x"70101011",
  1358 => x"80f8b033",
  1359 => x"7081ff06",
  1360 => x"72902911",
  1361 => x"70882b7d",
  1362 => x"07620c5a",
  1363 => x"5c5c5f57",
  1364 => x"5a5a758a",
  1365 => x"2e8c9f38",
  1366 => x"7680cf2e",
  1367 => x"8c983881",
  1368 => x"18577680",
  1369 => x"f8b03479",
  1370 => x"335675ff",
  1371 => x"bd3880f0",
  1372 => x"e4088411",
  1373 => x"0880e8dc",
  1374 => x"535658e0",
  1375 => x"d63f7c52",
  1376 => x"749fff06",
  1377 => x"51dfab3f",
  1378 => x"7c51e0c7",
  1379 => x"3f80e8f0",
  1380 => x"51e0c03f",
  1381 => x"7c52748c",
  1382 => x"2a870683",
  1383 => x"0581712b",
  1384 => x"525bdf8e",
  1385 => x"3f7c51e0",
  1386 => x"aa3f80e9",
  1387 => x"8451e0a3",
  1388 => x"3f748f2a",
  1389 => x"8106953d",
  1390 => x"5a568b53",
  1391 => x"80e3ac52",
  1392 => x"7851b4ae",
  1393 => x"3f820284",
  1394 => x"0580cd05",
  1395 => x"5957758f",
  1396 => x"06547389",
  1397 => x"268af838",
  1398 => x"7618b015",
  1399 => x"55557375",
  1400 => x"3475842a",
  1401 => x"ff187081",
  1402 => x"ff065955",
  1403 => x"5676df38",
  1404 => x"78793355",
  1405 => x"5773802e",
  1406 => x"a93880f0",
  1407 => x"fc087457",
  1408 => x"55811757",
  1409 => x"758a2e82",
  1410 => x"e6388415",
  1411 => x"0870822a",
  1412 => x"8106595c",
  1413 => x"77802ef2",
  1414 => x"3875750c",
  1415 => x"76335675",
  1416 => x"e0387879",
  1417 => x"33555a73",
  1418 => x"802e80cc",
  1419 => x"3880f0f4",
  1420 => x"0874575b",
  1421 => x"811a80f8",
  1422 => x"ac337081",
  1423 => x"ff067010",
  1424 => x"101180f8",
  1425 => x"b0337081",
  1426 => x"ff067290",
  1427 => x"29117088",
  1428 => x"2b7d0762",
  1429 => x"0c425c5c",
  1430 => x"57575a5a",
  1431 => x"758a2e89",
  1432 => x"f7387680",
  1433 => x"cf2e89f0",
  1434 => x"38811857",
  1435 => x"7680f8b0",
  1436 => x"34793356",
  1437 => x"75ffbd38",
  1438 => x"80f0e408",
  1439 => x"88110880",
  1440 => x"e9985356",
  1441 => x"59decc3f",
  1442 => x"74870654",
  1443 => x"73862682",
  1444 => x"83387310",
  1445 => x"1080f080",
  1446 => x"055b7a08",
  1447 => x"047618b7",
  1448 => x"15555573",
  1449 => x"75347584",
  1450 => x"2aff1870",
  1451 => x"81ff0659",
  1452 => x"5b5676f7",
  1453 => x"e338f882",
  1454 => x"39841508",
  1455 => x"70822a81",
  1456 => x"06595477",
  1457 => x"802ef238",
  1458 => x"8d750c84",
  1459 => x"15087082",
  1460 => x"2a81065b",
  1461 => x"5b79802e",
  1462 => x"f7fa38f8",
  1463 => x"86397618",
  1464 => x"b7155555",
  1465 => x"73753475",
  1466 => x"842aff18",
  1467 => x"7081ff06",
  1468 => x"59565676",
  1469 => x"f8f038f9",
  1470 => x"8f3974a3",
  1471 => x"26993881",
  1472 => x"19567580",
  1473 => x"f8ac3480",
  1474 => x"0b80f8b0",
  1475 => x"34793356",
  1476 => x"75f7eb38",
  1477 => x"f8ac3980",
  1478 => x"0b80f8ac",
  1479 => x"34800b80",
  1480 => x"f8b034e9",
  1481 => x"39841508",
  1482 => x"70822a81",
  1483 => x"065b5b79",
  1484 => x"802ef238",
  1485 => x"8d750c84",
  1486 => x"15087082",
  1487 => x"2a810655",
  1488 => x"5873802e",
  1489 => x"f8dc38f8",
  1490 => x"e8398415",
  1491 => x"0870822a",
  1492 => x"8106555a",
  1493 => x"73802ef2",
  1494 => x"388d750c",
  1495 => x"84150870",
  1496 => x"822a8106",
  1497 => x"59547780",
  1498 => x"2efb9538",
  1499 => x"fba13984",
  1500 => x"15087082",
  1501 => x"2a81065d",
  1502 => x"5a7b802e",
  1503 => x"f2388d75",
  1504 => x"0c841508",
  1505 => x"70822a81",
  1506 => x"06595c77",
  1507 => x"802efcfa",
  1508 => x"38fd8639",
  1509 => x"80e9ac51",
  1510 => x"dcb93f80",
  1511 => x"e9b451dc",
  1512 => x"b23f80e9",
  1513 => x"bc51dcab",
  1514 => x"3f74832a",
  1515 => x"83065473",
  1516 => x"812e89a1",
  1517 => x"38817426",
  1518 => x"89913873",
  1519 => x"822e89a9",
  1520 => x"3873832e",
  1521 => x"85a73880",
  1522 => x"e9d051dc",
  1523 => x"863f80e9",
  1524 => x"d451dbff",
  1525 => x"3f74852a",
  1526 => x"87065473",
  1527 => x"812e85b1",
  1528 => x"38817426",
  1529 => x"88db3873",
  1530 => x"822e8987",
  1531 => x"3873832e",
  1532 => x"84f13880",
  1533 => x"e9e851db",
  1534 => x"da3f7490",
  1535 => x"2a870654",
  1536 => x"7385268c",
  1537 => x"38731010",
  1538 => x"80f09c05",
  1539 => x"54730804",
  1540 => x"80e9ac51",
  1541 => x"dbbd3f80",
  1542 => x"e9fc51db",
  1543 => x"b63f7c52",
  1544 => x"74932a83",
  1545 => x"06820751",
  1546 => x"da883f7c",
  1547 => x"51dba43f",
  1548 => x"80ea9051",
  1549 => x"db9d3f7c",
  1550 => x"5274942a",
  1551 => x"8f0651d9",
  1552 => x"f13f7c51",
  1553 => x"db8d3f80",
  1554 => x"eaa451db",
  1555 => x"863f7c52",
  1556 => x"74982a81",
  1557 => x"06810551",
  1558 => x"d9d83f7c",
  1559 => x"51daf43f",
  1560 => x"80eab851",
  1561 => x"daed3f7c",
  1562 => x"52749e2a",
  1563 => x"820751d9",
  1564 => x"c13f7c51",
  1565 => x"dadd3f80",
  1566 => x"eacc51da",
  1567 => x"d63f749f",
  1568 => x"2a923d5a",
  1569 => x"568b5380",
  1570 => x"e3ac5278",
  1571 => x"51aee33f",
  1572 => x"82028405",
  1573 => x"80c10559",
  1574 => x"57758f06",
  1575 => x"54738926",
  1576 => x"85a43876",
  1577 => x"18b01555",
  1578 => x"55737534",
  1579 => x"75842aff",
  1580 => x"187081ff",
  1581 => x"06595e56",
  1582 => x"76df3878",
  1583 => x"79335557",
  1584 => x"73802ea9",
  1585 => x"3880f0fc",
  1586 => x"08745755",
  1587 => x"81175775",
  1588 => x"8a2e82c5",
  1589 => x"38841508",
  1590 => x"70822a81",
  1591 => x"065d5d7b",
  1592 => x"802ef238",
  1593 => x"75750c76",
  1594 => x"335675e0",
  1595 => x"38787933",
  1596 => x"555a7380",
  1597 => x"2e80cc38",
  1598 => x"80f0f408",
  1599 => x"74575b81",
  1600 => x"1a80f8ac",
  1601 => x"337081ff",
  1602 => x"06701010",
  1603 => x"1180f8b0",
  1604 => x"337081ff",
  1605 => x"06729029",
  1606 => x"1170882b",
  1607 => x"7d07620c",
  1608 => x"5a5c5c40",
  1609 => x"575a5a75",
  1610 => x"8a2e8586",
  1611 => x"387680cf",
  1612 => x"2e84ff38",
  1613 => x"81185675",
  1614 => x"80f8b034",
  1615 => x"79335675",
  1616 => x"ffbd3880",
  1617 => x"f0e40890",
  1618 => x"110880ea",
  1619 => x"e0535859",
  1620 => x"d9813f76",
  1621 => x"8f3d5a56",
  1622 => x"8b5380e3",
  1623 => x"ac527851",
  1624 => x"ad903f88",
  1625 => x"028405b5",
  1626 => x"05595775",
  1627 => x"8f065473",
  1628 => x"892683c9",
  1629 => x"387618b0",
  1630 => x"15555573",
  1631 => x"75347584",
  1632 => x"2aff1870",
  1633 => x"81ff0659",
  1634 => x"5c5676df",
  1635 => x"38787933",
  1636 => x"55577380",
  1637 => x"2ea93880",
  1638 => x"f0fc0874",
  1639 => x"57558117",
  1640 => x"57758a2e",
  1641 => x"81983884",
  1642 => x"15087082",
  1643 => x"2a810655",
  1644 => x"5b73802e",
  1645 => x"f2387575",
  1646 => x"0c763356",
  1647 => x"75e03878",
  1648 => x"7933555a",
  1649 => x"73802e80",
  1650 => x"cc3880f0",
  1651 => x"f4087457",
  1652 => x"5b811a80",
  1653 => x"f8ac3370",
  1654 => x"81ff0670",
  1655 => x"10101180",
  1656 => x"f8b03370",
  1657 => x"81ff0672",
  1658 => x"90291170",
  1659 => x"882b7d07",
  1660 => x"620c5a5c",
  1661 => x"5c40575a",
  1662 => x"5a758a2e",
  1663 => x"83963876",
  1664 => x"80cf2e83",
  1665 => x"8f388118",
  1666 => x"567580f8",
  1667 => x"b0347933",
  1668 => x"5675ffbd",
  1669 => x"38a53d0d",
  1670 => x"04841508",
  1671 => x"70822a81",
  1672 => x"065c587a",
  1673 => x"802ef238",
  1674 => x"8d750c84",
  1675 => x"15087082",
  1676 => x"2a81065d",
  1677 => x"5d7b802e",
  1678 => x"fd9b38fd",
  1679 => x"a7398415",
  1680 => x"0870822a",
  1681 => x"81065b5c",
  1682 => x"79802ef2",
  1683 => x"388d750c",
  1684 => x"84150870",
  1685 => x"822a8106",
  1686 => x"555b7380",
  1687 => x"2efec838",
  1688 => x"fed43980",
  1689 => x"eaf451d6",
  1690 => x"ea3ffb87",
  1691 => x"3980eaf8",
  1692 => x"51d6e03f",
  1693 => x"80e9d051",
  1694 => x"d6d93f80",
  1695 => x"e9d451d6",
  1696 => x"d23f7485",
  1697 => x"2a870654",
  1698 => x"73812e09",
  1699 => x"8106fad1",
  1700 => x"3880eafc",
  1701 => x"51d6bc3f",
  1702 => x"fad93980",
  1703 => x"eb8451d6",
  1704 => x"b23f80e7",
  1705 => x"f051d6ab",
  1706 => x"3f7c527b",
  1707 => x"972a8706",
  1708 => x"83058171",
  1709 => x"2b525ad4",
  1710 => x"f93f7c51",
  1711 => x"d6953f80",
  1712 => x"e88451d6",
  1713 => x"8e3f80e8",
  1714 => x"8c51d687",
  1715 => x"3f7c527b",
  1716 => x"9a2a8106",
  1717 => x"810551d4",
  1718 => x"d93f7c51",
  1719 => x"d5f53f80",
  1720 => x"e8a051d5",
  1721 => x"ee3f7c52",
  1722 => x"7b9b2a87",
  1723 => x"06830551",
  1724 => x"d4c03f7c",
  1725 => x"51d5dc3f",
  1726 => x"80e8b451",
  1727 => x"d5d53f7c",
  1728 => x"527b9e2a",
  1729 => x"820751d4",
  1730 => x"a93f7c51",
  1731 => x"d5c53f80",
  1732 => x"e8c851d5",
  1733 => x"be3f7b9f",
  1734 => x"2a983d5a",
  1735 => x"568b5380",
  1736 => x"e3ac5278",
  1737 => x"51a9cb3f",
  1738 => x"82028405",
  1739 => x"80d90559",
  1740 => x"57f39139",
  1741 => x"7618b715",
  1742 => x"5555f398",
  1743 => x"397618b7",
  1744 => x"155555fc",
  1745 => x"b6397618",
  1746 => x"b7155555",
  1747 => x"fadb3976",
  1748 => x"18b71555",
  1749 => x"55f58739",
  1750 => x"74a32681",
  1751 => x"cb388119",
  1752 => x"567580f8",
  1753 => x"ac34800b",
  1754 => x"80f8b034",
  1755 => x"79335675",
  1756 => x"f5c238f6",
  1757 => x"833974a3",
  1758 => x"26819e38",
  1759 => x"81195675",
  1760 => x"80f8ac34",
  1761 => x"800b80f8",
  1762 => x"b0347933",
  1763 => x"5675f39a",
  1764 => x"38f3db39",
  1765 => x"74a32680",
  1766 => x"f1388119",
  1767 => x"557480f8",
  1768 => x"ac34800b",
  1769 => x"80f8b034",
  1770 => x"79335675",
  1771 => x"fca338fc",
  1772 => x"e43974a3",
  1773 => x"2680c438",
  1774 => x"81195574",
  1775 => x"80f8ac34",
  1776 => x"800b80f8",
  1777 => x"b0347933",
  1778 => x"5675fab3",
  1779 => x"38faf439",
  1780 => x"74a32699",
  1781 => x"38811956",
  1782 => x"7580f8ac",
  1783 => x"34800b80",
  1784 => x"f8b03479",
  1785 => x"335675ef",
  1786 => x"e338f0a4",
  1787 => x"39800b80",
  1788 => x"f8ac3480",
  1789 => x"0b80f8b0",
  1790 => x"34e93980",
  1791 => x"0b80f8ac",
  1792 => x"34800b80",
  1793 => x"f8b034ff",
  1794 => x"bd39800b",
  1795 => x"80f8ac34",
  1796 => x"800b80f8",
  1797 => x"b034ff90",
  1798 => x"39800b80",
  1799 => x"f8ac3480",
  1800 => x"0b80f8b0",
  1801 => x"34fee339",
  1802 => x"800b80f8",
  1803 => x"ac34800b",
  1804 => x"80f8b034",
  1805 => x"feb63980",
  1806 => x"eb8c51d3",
  1807 => x"963ffce2",
  1808 => x"3980eb94",
  1809 => x"51d38c3f",
  1810 => x"f7a93980",
  1811 => x"eb9c51d3",
  1812 => x"823ffca0",
  1813 => x"3980eba0",
  1814 => x"51d2f83f",
  1815 => x"fc963980",
  1816 => x"eba451d2",
  1817 => x"ee3ffcba",
  1818 => x"3980ebac",
  1819 => x"51d2e43f",
  1820 => x"fc823980",
  1821 => x"ebb051d2",
  1822 => x"da3ff6f7",
  1823 => x"3980ebb4",
  1824 => x"51d2d03f",
  1825 => x"fc9c3980",
  1826 => x"ebbc51f6",
  1827 => x"8b3980eb",
  1828 => x"b051f684",
  1829 => x"3980ebc0",
  1830 => x"51f5fd39",
  1831 => x"80ebc451",
  1832 => x"f5f63980",
  1833 => x"ebc851d2",
  1834 => x"aa3f80e9",
  1835 => x"fc51d2a3",
  1836 => x"3f7c5274",
  1837 => x"932a8306",
  1838 => x"820751d0",
  1839 => x"f53f7c51",
  1840 => x"d2913f80",
  1841 => x"ea9051d2",
  1842 => x"8a3f7c52",
  1843 => x"74942a8f",
  1844 => x"0651d0de",
  1845 => x"3f7c51d1",
  1846 => x"fa3f80ea",
  1847 => x"a451d1f3",
  1848 => x"3f7c5274",
  1849 => x"982a8106",
  1850 => x"810551d0",
  1851 => x"c53f7c51",
  1852 => x"d1e13f80",
  1853 => x"eab851d1",
  1854 => x"da3f7c52",
  1855 => x"749e2a82",
  1856 => x"0751d0ae",
  1857 => x"3f7c51d1",
  1858 => x"ca3f80ea",
  1859 => x"cc51d1c3",
  1860 => x"3f749f2a",
  1861 => x"923d5a56",
  1862 => x"8b5380e3",
  1863 => x"ac527851",
  1864 => x"a5d03f82",
  1865 => x"02840580",
  1866 => x"c1055957",
  1867 => x"f6eb3980",
  1868 => x"ebd851d1",
  1869 => x"9e3f80e9",
  1870 => x"fc51d197",
  1871 => x"3f7c5274",
  1872 => x"932a8306",
  1873 => x"820751cf",
  1874 => x"e93f7c51",
  1875 => x"d1853f80",
  1876 => x"ea9051d0",
  1877 => x"fe3f7c52",
  1878 => x"74942a8f",
  1879 => x"0651cfd2",
  1880 => x"3f7c51d0",
  1881 => x"ee3f80ea",
  1882 => x"a451d0e7",
  1883 => x"3f7c5274",
  1884 => x"982a8106",
  1885 => x"810551cf",
  1886 => x"b93f7c51",
  1887 => x"d0d53f80",
  1888 => x"eab851d0",
  1889 => x"ce3f7c52",
  1890 => x"749e2a82",
  1891 => x"0751cfa2",
  1892 => x"3f7c51d0",
  1893 => x"be3f80ea",
  1894 => x"cc51d0b7",
  1895 => x"3f749f2a",
  1896 => x"923d5a56",
  1897 => x"8b5380e3",
  1898 => x"ac527851",
  1899 => x"a4c43f82",
  1900 => x"02840580",
  1901 => x"c1055957",
  1902 => x"f5df3980",
  1903 => x"ebe451d0",
  1904 => x"923f80e9",
  1905 => x"fc51d08b",
  1906 => x"3f7c5274",
  1907 => x"932a8306",
  1908 => x"820751ce",
  1909 => x"dd3f7c51",
  1910 => x"cff93f80",
  1911 => x"ea9051cf",
  1912 => x"f23f7c52",
  1913 => x"74942a8f",
  1914 => x"0651cec6",
  1915 => x"3f7c51cf",
  1916 => x"e23f80ea",
  1917 => x"a451cfdb",
  1918 => x"3f7c5274",
  1919 => x"982a8106",
  1920 => x"810551ce",
  1921 => x"ad3f7c51",
  1922 => x"cfc93f80",
  1923 => x"eab851cf",
  1924 => x"c23f7c52",
  1925 => x"749e2a82",
  1926 => x"0751ce96",
  1927 => x"3f7c51cf",
  1928 => x"b23f80ea",
  1929 => x"cc51cfab",
  1930 => x"3f749f2a",
  1931 => x"923d5a56",
  1932 => x"8b5380e3",
  1933 => x"ac527851",
  1934 => x"a3b83f82",
  1935 => x"02840580",
  1936 => x"c1055957",
  1937 => x"f4d33980",
  1938 => x"ebf451cf",
  1939 => x"863f80e9",
  1940 => x"fc51ceff",
  1941 => x"3f7c5274",
  1942 => x"932a8306",
  1943 => x"820751cd",
  1944 => x"d13f7c51",
  1945 => x"ceed3f80",
  1946 => x"ea9051ce",
  1947 => x"e63f7c52",
  1948 => x"74942a8f",
  1949 => x"0651cdba",
  1950 => x"3f7c51ce",
  1951 => x"d63f80ea",
  1952 => x"a451cecf",
  1953 => x"3f7c5274",
  1954 => x"982a8106",
  1955 => x"810551cd",
  1956 => x"a13f7c51",
  1957 => x"cebd3f80",
  1958 => x"eab851ce",
  1959 => x"b63f7c52",
  1960 => x"749e2a82",
  1961 => x"0751cd8a",
  1962 => x"3f7c51ce",
  1963 => x"a63f80ea",
  1964 => x"cc51ce9f",
  1965 => x"3f749f2a",
  1966 => x"923d5a56",
  1967 => x"8b5380e3",
  1968 => x"ac527851",
  1969 => x"a2ac3f82",
  1970 => x"02840580",
  1971 => x"c1055957",
  1972 => x"f3c73980",
  1973 => x"ec8051cd",
  1974 => x"fa3f80e9",
  1975 => x"fc51cdf3",
  1976 => x"3f7c5274",
  1977 => x"932a8306",
  1978 => x"820751cc",
  1979 => x"c53f7c51",
  1980 => x"cde13f80",
  1981 => x"ea9051cd",
  1982 => x"da3f7c52",
  1983 => x"74942a8f",
  1984 => x"0651ccae",
  1985 => x"3f7c51cd",
  1986 => x"ca3f80ea",
  1987 => x"a451cdc3",
  1988 => x"3f7c5274",
  1989 => x"982a8106",
  1990 => x"810551cc",
  1991 => x"953f7c51",
  1992 => x"cdb13f80",
  1993 => x"eab851cd",
  1994 => x"aa3f7c52",
  1995 => x"749e2a82",
  1996 => x"0751cbfe",
  1997 => x"3f7c51cd",
  1998 => x"9a3f80ea",
  1999 => x"cc51cd93",
  2000 => x"3f749f2a",
  2001 => x"923d5a56",
  2002 => x"8b5380e3",
  2003 => x"ac527851",
  2004 => x"a1a03f82",
  2005 => x"02840580",
  2006 => x"c1055957",
  2007 => x"f2bb39e5",
  2008 => x"3d0d80f0",
  2009 => x"e4088411",
  2010 => x"08709fff",
  2011 => x"06515555",
  2012 => x"8a55bb74",
  2013 => x"2783388f",
  2014 => x"55735287",
  2015 => x"e8519cac",
  2016 => x"3f8008fd",
  2017 => x"05752970",
  2018 => x"83ffff06",
  2019 => x"80ec9c53",
  2020 => x"4058ccbf",
  2021 => x"3f8051d0",
  2022 => x"923f8008",
  2023 => x"83ffff06",
  2024 => x"80ecb852",
  2025 => x"57ccac3f",
  2026 => x"983d7053",
  2027 => x"80f0e808",
  2028 => x"8c110853",
  2029 => x"575dcafa",
  2030 => x"3f7c51cc",
  2031 => x"963f80e6",
  2032 => x"fc51cc8f",
  2033 => x"3f76963d",
  2034 => x"5a568b53",
  2035 => x"80e3ac52",
  2036 => x"7851a09e",
  2037 => x"3f880284",
  2038 => x"0580d105",
  2039 => x"5957758f",
  2040 => x"06547389",
  2041 => x"2687d638",
  2042 => x"7618b015",
  2043 => x"55557375",
  2044 => x"3475842a",
  2045 => x"ff187081",
  2046 => x"ff06595b",
  2047 => x"5676df38",
  2048 => x"78793355",
  2049 => x"5773802e",
  2050 => x"a9387380",
  2051 => x"f0fc0856",
  2052 => x"56811757",
  2053 => x"758a2e87",
  2054 => x"c0388415",
  2055 => x"0870822a",
  2056 => x"81064142",
  2057 => x"7f802ef2",
  2058 => x"3875750c",
  2059 => x"76335675",
  2060 => x"e0387879",
  2061 => x"33555a73",
  2062 => x"802e80cc",
  2063 => x"387380f0",
  2064 => x"f4085c56",
  2065 => x"811a80f8",
  2066 => x"ac337081",
  2067 => x"ff067010",
  2068 => x"101180f8",
  2069 => x"b0337081",
  2070 => x"ff067290",
  2071 => x"29117088",
  2072 => x"2b7d0762",
  2073 => x"0c4a5c5c",
  2074 => x"57575a5a",
  2075 => x"758a2e87",
  2076 => x"8d387680",
  2077 => x"cf2e8786",
  2078 => x"38811859",
  2079 => x"7880f8b0",
  2080 => x"34793356",
  2081 => x"75ffbd38",
  2082 => x"80f0e808",
  2083 => x"7f305755",
  2084 => x"8c150857",
  2085 => x"75772596",
  2086 => x"38800b84",
  2087 => x"160c7408",
  2088 => x"5877ed38",
  2089 => x"74085877",
  2090 => x"802ef338",
  2091 => x"e339800b",
  2092 => x"88160c74",
  2093 => x"08567580",
  2094 => x"2ef93880",
  2095 => x"750c8251",
  2096 => x"8dce3f83",
  2097 => x"ffff0b80",
  2098 => x"f0e8088c",
  2099 => x"11084356",
  2100 => x"40805ed4",
  2101 => x"cd7e4542",
  2102 => x"abb30b8c",
  2103 => x"16085b43",
  2104 => x"797f2583",
  2105 => x"c238800b",
  2106 => x"88160c74",
  2107 => x"085b7a80",
  2108 => x"2ef93880",
  2109 => x"51cdb43f",
  2110 => x"800883ff",
  2111 => x"ff0680e6",
  2112 => x"cc0b80e6",
  2113 => x"cc33565b",
  2114 => x"5c73802e",
  2115 => x"80cc3880",
  2116 => x"f0f40874",
  2117 => x"575b811a",
  2118 => x"80f8ac33",
  2119 => x"7081ff06",
  2120 => x"70101011",
  2121 => x"80f8b033",
  2122 => x"7081ff06",
  2123 => x"72902911",
  2124 => x"70882b7d",
  2125 => x"07620c53",
  2126 => x"5c5c5757",
  2127 => x"5a5a758a",
  2128 => x"2e86ce38",
  2129 => x"7680cf2e",
  2130 => x"86c73881",
  2131 => x"18597880",
  2132 => x"f8b03479",
  2133 => x"335675ff",
  2134 => x"bd387b60",
  2135 => x"278c387b",
  2136 => x"80f0e808",
  2137 => x"8c110843",
  2138 => x"58407b30",
  2139 => x"70802555",
  2140 => x"587d9738",
  2141 => x"81707506",
  2142 => x"57557580",
  2143 => x"2e8c3874",
  2144 => x"80f0e808",
  2145 => x"8c110844",
  2146 => x"5b5e7b30",
  2147 => x"70802555",
  2148 => x"5b7d802e",
  2149 => x"97388170",
  2150 => x"75065555",
  2151 => x"73802e8c",
  2152 => x"387480f0",
  2153 => x"e8088c11",
  2154 => x"08455644",
  2155 => x"80e6cc51",
  2156 => x"c8a13f82",
  2157 => x"52805193",
  2158 => x"8a3f7c52",
  2159 => x"80f0e808",
  2160 => x"8c110852",
  2161 => x"59c6eb3f",
  2162 => x"7c7d3355",
  2163 => x"5773802e",
  2164 => x"a93880f0",
  2165 => x"fc087457",
  2166 => x"55811757",
  2167 => x"758a2e84",
  2168 => x"c8388415",
  2169 => x"0870822a",
  2170 => x"81065558",
  2171 => x"73802ef2",
  2172 => x"3875750c",
  2173 => x"76335675",
  2174 => x"e03880ec",
  2175 => x"c40b80ec",
  2176 => x"c4335557",
  2177 => x"73802ea9",
  2178 => x"3880f0fc",
  2179 => x"08745755",
  2180 => x"81175775",
  2181 => x"8a2e84b6",
  2182 => x"38841508",
  2183 => x"70822a81",
  2184 => x"065a5a78",
  2185 => x"802ef238",
  2186 => x"75750c76",
  2187 => x"335675e0",
  2188 => x"387c527b",
  2189 => x"51c5fb3f",
  2190 => x"7c51c797",
  2191 => x"3f80ecc8",
  2192 => x"0b80ecc8",
  2193 => x"33555a73",
  2194 => x"802e80cc",
  2195 => x"3880f0f4",
  2196 => x"0874575b",
  2197 => x"811a80f8",
  2198 => x"ac337081",
  2199 => x"ff067010",
  2200 => x"101180f8",
  2201 => x"b0337081",
  2202 => x"ff067290",
  2203 => x"29117088",
  2204 => x"2b7d0762",
  2205 => x"0c5a5c5c",
  2206 => x"5f575a5a",
  2207 => x"758a2e83",
  2208 => x"f2387680",
  2209 => x"cf2e83eb",
  2210 => x"38811856",
  2211 => x"7580f8b0",
  2212 => x"34793356",
  2213 => x"75ffbd38",
  2214 => x"80f0e808",
  2215 => x"8c11085b",
  2216 => x"557e7a24",
  2217 => x"fcc03863",
  2218 => x"802e849f",
  2219 => x"387d802e",
  2220 => x"84993862",
  2221 => x"6231709f",
  2222 => x"2a117081",
  2223 => x"2c657131",
  2224 => x"8c190870",
  2225 => x"7231525d",
  2226 => x"59415c57",
  2227 => x"80762599",
  2228 => x"38ff1656",
  2229 => x"800b8416",
  2230 => x"0c740858",
  2231 => x"77ee3874",
  2232 => x"08587780",
  2233 => x"2ef338e4",
  2234 => x"3980e6cc",
  2235 => x"51c5e43f",
  2236 => x"7d802e85",
  2237 => x"9e3880ec",
  2238 => x"d051c5d7",
  2239 => x"3f80e6cc",
  2240 => x"51c5d03f",
  2241 => x"63802e83",
  2242 => x"d33880ec",
  2243 => x"dc51c5c3",
  2244 => x"3f80ece8",
  2245 => x"51c5bc3f",
  2246 => x"7c526151",
  2247 => x"c4943f7c",
  2248 => x"51c5b03f",
  2249 => x"80ecf851",
  2250 => x"c5a93f7c",
  2251 => x"526251c4",
  2252 => x"813f7c51",
  2253 => x"c59d3f80",
  2254 => x"e6cc51c5",
  2255 => x"963f80ed",
  2256 => x"8851c58f",
  2257 => x"3f7c5276",
  2258 => x"51c3e73f",
  2259 => x"7c51c583",
  2260 => x"3f80ed98",
  2261 => x"51c4fc3f",
  2262 => x"7c52769f",
  2263 => x"2a177081",
  2264 => x"2c5242c3",
  2265 => x"cd3f7c51",
  2266 => x"c4e93f80",
  2267 => x"e6cc51c4",
  2268 => x"e23f80ed",
  2269 => x"a851c4db",
  2270 => x"3f7c527f",
  2271 => x"51c3b33f",
  2272 => x"7c51c4cf",
  2273 => x"3f80edb8",
  2274 => x"51c4c83f",
  2275 => x"7c526051",
  2276 => x"c3a03f7c",
  2277 => x"51c4bc3f",
  2278 => x"80e6cc51",
  2279 => x"c4b53f80",
  2280 => x"edc851c4",
  2281 => x"ae3f7c52",
  2282 => x"80f0e808",
  2283 => x"8c110852",
  2284 => x"5ec2ff3f",
  2285 => x"7c51c49b",
  2286 => x"3f9d3d0d",
  2287 => x"047618b7",
  2288 => x"15555573",
  2289 => x"75347584",
  2290 => x"2aff1870",
  2291 => x"81ff0659",
  2292 => x"5b5676f8",
  2293 => x"8938f8a8",
  2294 => x"39841508",
  2295 => x"70822a81",
  2296 => x"065c5e7a",
  2297 => x"802ef238",
  2298 => x"8d750c84",
  2299 => x"15087082",
  2300 => x"2a810641",
  2301 => x"427f802e",
  2302 => x"f8a038f8",
  2303 => x"ac3974a3",
  2304 => x"26993881",
  2305 => x"19557480",
  2306 => x"f8ac3480",
  2307 => x"0b80f8b0",
  2308 => x"34793356",
  2309 => x"75f8ad38",
  2310 => x"f8ee3980",
  2311 => x"0b80f8ac",
  2312 => x"34800b80",
  2313 => x"f8b034e9",
  2314 => x"39841508",
  2315 => x"70822a81",
  2316 => x"06595b77",
  2317 => x"802ef238",
  2318 => x"8d750c84",
  2319 => x"15087082",
  2320 => x"2a810655",
  2321 => x"5873802e",
  2322 => x"fb9838fb",
  2323 => x"a4398415",
  2324 => x"0870822a",
  2325 => x"81065b54",
  2326 => x"79802ef2",
  2327 => x"388d750c",
  2328 => x"84150870",
  2329 => x"822a8106",
  2330 => x"5a5a7880",
  2331 => x"2efbaa38",
  2332 => x"fbb63974",
  2333 => x"a32680c4",
  2334 => x"38811957",
  2335 => x"7680f8ac",
  2336 => x"34800b80",
  2337 => x"f8b03479",
  2338 => x"335675fb",
  2339 => x"c738fc88",
  2340 => x"3974a326",
  2341 => x"99388119",
  2342 => x"557480f8",
  2343 => x"ac34800b",
  2344 => x"80f8b034",
  2345 => x"79335675",
  2346 => x"f8ec38f9",
  2347 => x"ad39800b",
  2348 => x"80f8ac34",
  2349 => x"800b80f8",
  2350 => x"b034e939",
  2351 => x"800b80f8",
  2352 => x"ac34800b",
  2353 => x"80f8b034",
  2354 => x"ffbd3960",
  2355 => x"6363318c",
  2356 => x"17087073",
  2357 => x"31535b58",
  2358 => x"56fbf139",
  2359 => x"80edd851",
  2360 => x"c1f13f80",
  2361 => x"ece851c1",
  2362 => x"ea3f7c52",
  2363 => x"6151c0c2",
  2364 => x"3f7c51c1",
  2365 => x"de3f80ec",
  2366 => x"f851c1d7",
  2367 => x"3f7c5262",
  2368 => x"51c0af3f",
  2369 => x"7c51c1cb",
  2370 => x"3f80e6cc",
  2371 => x"51c1c43f",
  2372 => x"80ed8851",
  2373 => x"c1bd3f7c",
  2374 => x"527651c0",
  2375 => x"953f7c51",
  2376 => x"c1b13f80",
  2377 => x"ed9851c1",
  2378 => x"aa3f7c52",
  2379 => x"769f2a17",
  2380 => x"70812c52",
  2381 => x"42ffbffa",
  2382 => x"3f7c51c1",
  2383 => x"963f80e6",
  2384 => x"cc51c18f",
  2385 => x"3f80eda8",
  2386 => x"51c1883f",
  2387 => x"7c527f51",
  2388 => x"ffbfdf3f",
  2389 => x"7c51c0fb",
  2390 => x"3f80edb8",
  2391 => x"51c0f43f",
  2392 => x"7c526051",
  2393 => x"ffbfcb3f",
  2394 => x"7c51c0e7",
  2395 => x"3f80e6cc",
  2396 => x"51c0e03f",
  2397 => x"80edc851",
  2398 => x"c0d93f7c",
  2399 => x"5280f0e8",
  2400 => x"088c1108",
  2401 => x"525effbf",
  2402 => x"a93f7c51",
  2403 => x"c0c53f9d",
  2404 => x"3d0d0480",
  2405 => x"ede851fa",
  2406 => x"e139f73d",
  2407 => x"0d800b80",
  2408 => x"f0f00870",
  2409 => x"08810a06",
  2410 => x"80f8a80c",
  2411 => x"545585ae",
  2412 => x"3f85bc3f",
  2413 => x"80f0f408",
  2414 => x"7584120c",
  2415 => x"52fe800a",
  2416 => x"0b88130c",
  2417 => x"7480f8ac",
  2418 => x"347480f8",
  2419 => x"b03480f0",
  2420 => x"fc0853b6",
  2421 => x"0b8c140c",
  2422 => x"830b8814",
  2423 => x"0c80f0f0",
  2424 => x"08881108",
  2425 => x"81ff0788",
  2426 => x"120c5380",
  2427 => x"f0ec0853",
  2428 => x"ff0b8414",
  2429 => x"0cfc9480",
  2430 => x"0b88140c",
  2431 => x"82d0affd",
  2432 => x"fb0b8c14",
  2433 => x"0c80c073",
  2434 => x"0c720870",
  2435 => x"862a8106",
  2436 => x"515271f5",
  2437 => x"38901308",
  2438 => x"70832a81",
  2439 => x"06515473",
  2440 => x"f43881fc",
  2441 => x"80810b90",
  2442 => x"140c9013",
  2443 => x"0870832a",
  2444 => x"81065152",
  2445 => x"71f43880",
  2446 => x"fdc0810b",
  2447 => x"90140c89",
  2448 => x"0a5283ff",
  2449 => x"ff537172",
  2450 => x"0c8412ff",
  2451 => x"14545272",
  2452 => x"8025f338",
  2453 => x"80e69c51",
  2454 => x"ffbef83f",
  2455 => x"800b80f0",
  2456 => x"f4085553",
  2457 => x"72882b74",
  2458 => x"0c811353",
  2459 => x"97907326",
  2460 => x"f338800b",
  2461 => x"80f8ac34",
  2462 => x"800b80f8",
  2463 => x"b03480ed",
  2464 => x"f851ffbe",
  2465 => x"ce3f80f8",
  2466 => x"a808802e",
  2467 => x"81d83880",
  2468 => x"ee8051ff",
  2469 => x"bebd3f80",
  2470 => x"ee9051ff",
  2471 => x"beb53fd7",
  2472 => x"a73f8551",
  2473 => x"81ea3ff1",
  2474 => x"b63f8a51",
  2475 => x"81e23f80",
  2476 => x"0b80f0f4",
  2477 => x"08555372",
  2478 => x"882b740c",
  2479 => x"81135397",
  2480 => x"907326f3",
  2481 => x"38800b80",
  2482 => x"f8ac3480",
  2483 => x"0b80f8b0",
  2484 => x"347451c1",
  2485 => x"d63f80f0",
  2486 => x"f0087008",
  2487 => x"70872a81",
  2488 => x"06515454",
  2489 => x"72802e8b",
  2490 => x"3880f0e8",
  2491 => x"0852800b",
  2492 => x"84130c73",
  2493 => x"0870842a",
  2494 => x"81065153",
  2495 => x"72802e8b",
  2496 => x"3880f0e8",
  2497 => x"0852800b",
  2498 => x"88130c73",
  2499 => x"0870852a",
  2500 => x"81065153",
  2501 => x"72802e96",
  2502 => x"38890a52",
  2503 => x"83ffff53",
  2504 => x"71720c84",
  2505 => x"12ff1454",
  2506 => x"52728025",
  2507 => x"f3387308",
  2508 => x"70862a81",
  2509 => x"06555373",
  2510 => x"802eff95",
  2511 => x"38800b80",
  2512 => x"f0f40855",
  2513 => x"5372882b",
  2514 => x"740c8113",
  2515 => x"53979073",
  2516 => x"26f33880",
  2517 => x"0b80f8ac",
  2518 => x"34800b80",
  2519 => x"f8b03474",
  2520 => x"813255fe",
  2521 => x"ec3980ee",
  2522 => x"b451fea7",
  2523 => x"39fd3d0d",
  2524 => x"80f0f808",
  2525 => x"76b0ea29",
  2526 => x"94120c54",
  2527 => x"850b9815",
  2528 => x"0c981408",
  2529 => x"70810651",
  2530 => x"5372f638",
  2531 => x"853d0d04",
  2532 => x"fb3d0d77",
  2533 => x"56805574",
  2534 => x"76278199",
  2535 => x"3880f0f8",
  2536 => x"0854bfa9",
  2537 => x"bc0b9415",
  2538 => x"0c850b98",
  2539 => x"150c9814",
  2540 => x"08708106",
  2541 => x"515372f6",
  2542 => x"38bfa9bc",
  2543 => x"0b94150c",
  2544 => x"850b9815",
  2545 => x"0c981408",
  2546 => x"70810651",
  2547 => x"5372f638",
  2548 => x"bfa9bc0b",
  2549 => x"94150c85",
  2550 => x"0b98150c",
  2551 => x"98140870",
  2552 => x"81065153",
  2553 => x"72f638bf",
  2554 => x"a9bc0b94",
  2555 => x"150c850b",
  2556 => x"98150c98",
  2557 => x"14087081",
  2558 => x"06515372",
  2559 => x"f638bfa9",
  2560 => x"bc0b9415",
  2561 => x"0c850b98",
  2562 => x"150c9814",
  2563 => x"08708106",
  2564 => x"515372f6",
  2565 => x"38bfa9bc",
  2566 => x"0b94150c",
  2567 => x"850b9815",
  2568 => x"0c981408",
  2569 => x"70810651",
  2570 => x"5372f638",
  2571 => x"81155575",
  2572 => x"7526feee",
  2573 => x"38873d0d",
  2574 => x"04ff3d0d",
  2575 => x"80f0f808",
  2576 => x"74101075",
  2577 => x"10059412",
  2578 => x"0c52850b",
  2579 => x"98130c98",
  2580 => x"12087081",
  2581 => x"06515170",
  2582 => x"f638833d",
  2583 => x"0d04803d",
  2584 => x"0d80f0f8",
  2585 => x"0851870b",
  2586 => x"84120c82",
  2587 => x"3d0d04fd",
  2588 => x"3d0d80f0",
  2589 => x"f0088811",
  2590 => x"0883de80",
  2591 => x"0788120c",
  2592 => x"841108fc",
  2593 => x"a1ff0684",
  2594 => x"120c538f",
  2595 => x"51fdde3f",
  2596 => x"80f0f008",
  2597 => x"841108e1",
  2598 => x"ff068412",
  2599 => x"0c841108",
  2600 => x"86800784",
  2601 => x"120c8411",
  2602 => x"0880c080",
  2603 => x"0784120c",
  2604 => x"538151ff",
  2605 => x"843f80f0",
  2606 => x"f0088411",
  2607 => x"08ffbfff",
  2608 => x"0684120c",
  2609 => x"538551fd",
  2610 => x"a43f80f0",
  2611 => x"f0088411",
  2612 => x"0880c080",
  2613 => x"0784120c",
  2614 => x"538151fe",
  2615 => x"dc3f80f0",
  2616 => x"f0088411",
  2617 => x"08ffbfff",
  2618 => x"0684120c",
  2619 => x"538151fc",
  2620 => x"fc3f80f0",
  2621 => x"f0088411",
  2622 => x"0880c080",
  2623 => x"0784120c",
  2624 => x"538151fe",
  2625 => x"b43f80f0",
  2626 => x"f0088411",
  2627 => x"08ffbfff",
  2628 => x"0684120c",
  2629 => x"538151fc",
  2630 => x"d43f80f0",
  2631 => x"f0088411",
  2632 => x"08e1ff06",
  2633 => x"84120c53",
  2634 => x"84800b84",
  2635 => x"14087072",
  2636 => x"0784160c",
  2637 => x"53841408",
  2638 => x"7080c080",
  2639 => x"0784160c",
  2640 => x"53548151",
  2641 => x"fdf33f80",
  2642 => x"f0f00884",
  2643 => x"110870ff",
  2644 => x"bfff0684",
  2645 => x"130c5353",
  2646 => x"8551fc91",
  2647 => x"3f80f0f0",
  2648 => x"08841108",
  2649 => x"70feffff",
  2650 => x"0684130c",
  2651 => x"53841108",
  2652 => x"70e1ff06",
  2653 => x"84130c53",
  2654 => x"84110870",
  2655 => x"76078413",
  2656 => x"0c538411",
  2657 => x"0880c080",
  2658 => x"0784120c",
  2659 => x"538151fd",
  2660 => x"a83f80f0",
  2661 => x"f0088411",
  2662 => x"08ffbfff",
  2663 => x"0684120c",
  2664 => x"841108e1",
  2665 => x"ff068412",
  2666 => x"0c841108",
  2667 => x"90800784",
  2668 => x"120c8411",
  2669 => x"0880c080",
  2670 => x"0784120c",
  2671 => x"548151fc",
  2672 => x"f83f80f0",
  2673 => x"f0088411",
  2674 => x"08ffbfff",
  2675 => x"0684120c",
  2676 => x"54aa51fc",
  2677 => x"e43f80f0",
  2678 => x"f0088411",
  2679 => x"08feffff",
  2680 => x"0684120c",
  2681 => x"841108e1",
  2682 => x"ff068412",
  2683 => x"0c841108",
  2684 => x"84120c84",
  2685 => x"110880c0",
  2686 => x"80078412",
  2687 => x"0c548151",
  2688 => x"fcb73f80",
  2689 => x"f0f00884",
  2690 => x"1108ffbf",
  2691 => x"ff068412",
  2692 => x"0c841108",
  2693 => x"e1ff0684",
  2694 => x"120c8411",
  2695 => x"08988007",
  2696 => x"84120c84",
  2697 => x"110880c0",
  2698 => x"80078412",
  2699 => x"0c548151",
  2700 => x"fc873f80",
  2701 => x"f0f00884",
  2702 => x"1108ffbf",
  2703 => x"ff068412",
  2704 => x"0c54aa51",
  2705 => x"fbf33f80",
  2706 => x"f0f00884",
  2707 => x"1108feff",
  2708 => x"ff068412",
  2709 => x"0c841108",
  2710 => x"e1ff0684",
  2711 => x"120c8411",
  2712 => x"0884120c",
  2713 => x"84110880",
  2714 => x"c0800784",
  2715 => x"120c5481",
  2716 => x"51fbc63f",
  2717 => x"80f0f008",
  2718 => x"841108ff",
  2719 => x"bfff0684",
  2720 => x"120c8411",
  2721 => x"08e1ff06",
  2722 => x"84120c84",
  2723 => x"11088c80",
  2724 => x"0784120c",
  2725 => x"84110880",
  2726 => x"c0800784",
  2727 => x"120c5481",
  2728 => x"51fb963f",
  2729 => x"80f0f008",
  2730 => x"841108ff",
  2731 => x"bfff0684",
  2732 => x"120c54aa",
  2733 => x"51fb823f",
  2734 => x"810b80f0",
  2735 => x"f0088411",
  2736 => x"0870feff",
  2737 => x"ff068413",
  2738 => x"0c548411",
  2739 => x"0870e1ff",
  2740 => x"0684130c",
  2741 => x"54841108",
  2742 => x"84120c84",
  2743 => x"11087080",
  2744 => x"c0800784",
  2745 => x"130c5454",
  2746 => x"705254fa",
  2747 => x"cc3f80f0",
  2748 => x"f0088411",
  2749 => x"0870ffbf",
  2750 => x"ff068413",
  2751 => x"0c538411",
  2752 => x"0870e1ff",
  2753 => x"0684130c",
  2754 => x"53841108",
  2755 => x"70828007",
  2756 => x"84130c53",
  2757 => x"84110870",
  2758 => x"80c08007",
  2759 => x"84130c53",
  2760 => x"537351fa",
  2761 => x"943f80f0",
  2762 => x"f0088411",
  2763 => x"08ffbfff",
  2764 => x"0684120c",
  2765 => x"53aa51fa",
  2766 => x"803f8251",
  2767 => x"f8af3f85",
  2768 => x"3d0d04fc",
  2769 => x"3d0d029b",
  2770 => x"05330284",
  2771 => x"059f0533",
  2772 => x"54527282",
  2773 => x"2e81ad38",
  2774 => x"82732591",
  2775 => x"3872832e",
  2776 => x"83bc3872",
  2777 => x"842e82a9",
  2778 => x"38863d0d",
  2779 => x"0472812e",
  2780 => x"098106f5",
  2781 => x"38ff8012",
  2782 => x"7081ff06",
  2783 => x"80f0f008",
  2784 => x"841108fe",
  2785 => x"ffff0684",
  2786 => x"120c8411",
  2787 => x"08e1ff06",
  2788 => x"84120c71",
  2789 => x"842b9e80",
  2790 => x"06841208",
  2791 => x"70720784",
  2792 => x"140c5484",
  2793 => x"120880c0",
  2794 => x"80078413",
  2795 => x"0c575556",
  2796 => x"528151f9",
  2797 => x"843f80f0",
  2798 => x"f0088411",
  2799 => x"08ffbfff",
  2800 => x"0684120c",
  2801 => x"841108e1",
  2802 => x"ff068412",
  2803 => x"0c75882b",
  2804 => x"9e800684",
  2805 => x"12087107",
  2806 => x"84130c84",
  2807 => x"120880c0",
  2808 => x"80078413",
  2809 => x"0c555381",
  2810 => x"51f8ce3f",
  2811 => x"80f0f008",
  2812 => x"841108ff",
  2813 => x"bfff0684",
  2814 => x"120c53aa",
  2815 => x"51f8ba3f",
  2816 => x"863d0d04",
  2817 => x"c0127081",
  2818 => x"ff0680f0",
  2819 => x"f0088411",
  2820 => x"08feffff",
  2821 => x"0684120c",
  2822 => x"841108e1",
  2823 => x"ff068412",
  2824 => x"0c71842b",
  2825 => x"9e800684",
  2826 => x"12087072",
  2827 => x"0784140c",
  2828 => x"54841208",
  2829 => x"80c08007",
  2830 => x"84130c57",
  2831 => x"55565281",
  2832 => x"51f7f63f",
  2833 => x"80f0f008",
  2834 => x"841108ff",
  2835 => x"bfff0684",
  2836 => x"120c8411",
  2837 => x"08e1ff06",
  2838 => x"84120c75",
  2839 => x"882b9e80",
  2840 => x"06841208",
  2841 => x"71078413",
  2842 => x"0c841208",
  2843 => x"80c08007",
  2844 => x"84130c55",
  2845 => x"538151f7",
  2846 => x"c03f80f0",
  2847 => x"f0088411",
  2848 => x"08ffbfff",
  2849 => x"0684120c",
  2850 => x"53aa51f7",
  2851 => x"ac3ffef0",
  2852 => x"39d01270",
  2853 => x"81ff0680",
  2854 => x"f0f00884",
  2855 => x"1108feff",
  2856 => x"ff068412",
  2857 => x"0c841108",
  2858 => x"e1ff0684",
  2859 => x"120c7184",
  2860 => x"2b9e8006",
  2861 => x"84120870",
  2862 => x"72078414",
  2863 => x"0c548412",
  2864 => x"0880c080",
  2865 => x"0784130c",
  2866 => x"57555652",
  2867 => x"8151f6e9",
  2868 => x"3f80f0f0",
  2869 => x"08841108",
  2870 => x"ffbfff06",
  2871 => x"84120c84",
  2872 => x"1108e1ff",
  2873 => x"0684120c",
  2874 => x"75882b9e",
  2875 => x"80068412",
  2876 => x"08710784",
  2877 => x"130c8412",
  2878 => x"0880c080",
  2879 => x"0784130c",
  2880 => x"55538151",
  2881 => x"f6b33f80",
  2882 => x"f0f00884",
  2883 => x"1108ffbf",
  2884 => x"ff068412",
  2885 => x"0c53aa51",
  2886 => x"f69f3ffd",
  2887 => x"e339ff90",
  2888 => x"127081ff",
  2889 => x"0680f0f0",
  2890 => x"08841108",
  2891 => x"feffff06",
  2892 => x"84120c84",
  2893 => x"1108e1ff",
  2894 => x"0684120c",
  2895 => x"71842b9e",
  2896 => x"80068412",
  2897 => x"08707207",
  2898 => x"84140c54",
  2899 => x"84120880",
  2900 => x"c0800784",
  2901 => x"130c5755",
  2902 => x"56528151",
  2903 => x"f5db3f80",
  2904 => x"f0f00884",
  2905 => x"1108ffbf",
  2906 => x"ff068412",
  2907 => x"0c841108",
  2908 => x"e1ff0684",
  2909 => x"120c7588",
  2910 => x"2b9e8006",
  2911 => x"84120871",
  2912 => x"0784130c",
  2913 => x"84120880",
  2914 => x"c0800784",
  2915 => x"130c5553",
  2916 => x"8151f5a5",
  2917 => x"3f80f0f0",
  2918 => x"08841108",
  2919 => x"ffbfff06",
  2920 => x"84120c53",
  2921 => x"aa51f591",
  2922 => x"3ffcd539",
  2923 => x"8c08028c",
  2924 => x"0cfd3d0d",
  2925 => x"80538c08",
  2926 => x"8c050852",
  2927 => x"8c088805",
  2928 => x"085182de",
  2929 => x"3f800870",
  2930 => x"800c5485",
  2931 => x"3d0d8c0c",
  2932 => x"048c0802",
  2933 => x"8c0cfd3d",
  2934 => x"0d81538c",
  2935 => x"088c0508",
  2936 => x"528c0888",
  2937 => x"05085182",
  2938 => x"b93f8008",
  2939 => x"70800c54",
  2940 => x"853d0d8c",
  2941 => x"0c048c08",
  2942 => x"028c0cf9",
  2943 => x"3d0d800b",
  2944 => x"8c08fc05",
  2945 => x"0c8c0888",
  2946 => x"05088025",
  2947 => x"ab388c08",
  2948 => x"88050830",
  2949 => x"8c088805",
  2950 => x"0c800b8c",
  2951 => x"08f4050c",
  2952 => x"8c08fc05",
  2953 => x"08883881",
  2954 => x"0b8c08f4",
  2955 => x"050c8c08",
  2956 => x"f405088c",
  2957 => x"08fc050c",
  2958 => x"8c088c05",
  2959 => x"088025ab",
  2960 => x"388c088c",
  2961 => x"0508308c",
  2962 => x"088c050c",
  2963 => x"800b8c08",
  2964 => x"f0050c8c",
  2965 => x"08fc0508",
  2966 => x"8838810b",
  2967 => x"8c08f005",
  2968 => x"0c8c08f0",
  2969 => x"05088c08",
  2970 => x"fc050c80",
  2971 => x"538c088c",
  2972 => x"0508528c",
  2973 => x"08880508",
  2974 => x"5181a73f",
  2975 => x"8008708c",
  2976 => x"08f8050c",
  2977 => x"548c08fc",
  2978 => x"0508802e",
  2979 => x"8c388c08",
  2980 => x"f8050830",
  2981 => x"8c08f805",
  2982 => x"0c8c08f8",
  2983 => x"05087080",
  2984 => x"0c54893d",
  2985 => x"0d8c0c04",
  2986 => x"8c08028c",
  2987 => x"0cfb3d0d",
  2988 => x"800b8c08",
  2989 => x"fc050c8c",
  2990 => x"08880508",
  2991 => x"80259338",
  2992 => x"8c088805",
  2993 => x"08308c08",
  2994 => x"88050c81",
  2995 => x"0b8c08fc",
  2996 => x"050c8c08",
  2997 => x"8c050880",
  2998 => x"258c388c",
  2999 => x"088c0508",
  3000 => x"308c088c",
  3001 => x"050c8153",
  3002 => x"8c088c05",
  3003 => x"08528c08",
  3004 => x"88050851",
  3005 => x"ad3f8008",
  3006 => x"708c08f8",
  3007 => x"050c548c",
  3008 => x"08fc0508",
  3009 => x"802e8c38",
  3010 => x"8c08f805",
  3011 => x"08308c08",
  3012 => x"f8050c8c",
  3013 => x"08f80508",
  3014 => x"70800c54",
  3015 => x"873d0d8c",
  3016 => x"0c048c08",
  3017 => x"028c0cfd",
  3018 => x"3d0d810b",
  3019 => x"8c08fc05",
  3020 => x"0c800b8c",
  3021 => x"08f8050c",
  3022 => x"8c088c05",
  3023 => x"088c0888",
  3024 => x"050827ac",
  3025 => x"388c08fc",
  3026 => x"0508802e",
  3027 => x"a338800b",
  3028 => x"8c088c05",
  3029 => x"08249938",
  3030 => x"8c088c05",
  3031 => x"08108c08",
  3032 => x"8c050c8c",
  3033 => x"08fc0508",
  3034 => x"108c08fc",
  3035 => x"050cc939",
  3036 => x"8c08fc05",
  3037 => x"08802e80",
  3038 => x"c9388c08",
  3039 => x"8c05088c",
  3040 => x"08880508",
  3041 => x"26a1388c",
  3042 => x"08880508",
  3043 => x"8c088c05",
  3044 => x"08318c08",
  3045 => x"88050c8c",
  3046 => x"08f80508",
  3047 => x"8c08fc05",
  3048 => x"08078c08",
  3049 => x"f8050c8c",
  3050 => x"08fc0508",
  3051 => x"812a8c08",
  3052 => x"fc050c8c",
  3053 => x"088c0508",
  3054 => x"812a8c08",
  3055 => x"8c050cff",
  3056 => x"af398c08",
  3057 => x"90050880",
  3058 => x"2e8f388c",
  3059 => x"08880508",
  3060 => x"708c08f4",
  3061 => x"050c518d",
  3062 => x"398c08f8",
  3063 => x"0508708c",
  3064 => x"08f4050c",
  3065 => x"518c08f4",
  3066 => x"0508800c",
  3067 => x"853d0d8c",
  3068 => x"0c04fc3d",
  3069 => x"0d767079",
  3070 => x"7b555555",
  3071 => x"558f7227",
  3072 => x"8c387275",
  3073 => x"07830651",
  3074 => x"70802ea7",
  3075 => x"38ff1252",
  3076 => x"71ff2e98",
  3077 => x"38727081",
  3078 => x"05543374",
  3079 => x"70810556",
  3080 => x"34ff1252",
  3081 => x"71ff2e09",
  3082 => x"8106ea38",
  3083 => x"74800c86",
  3084 => x"3d0d0474",
  3085 => x"51727084",
  3086 => x"05540871",
  3087 => x"70840553",
  3088 => x"0c727084",
  3089 => x"05540871",
  3090 => x"70840553",
  3091 => x"0c727084",
  3092 => x"05540871",
  3093 => x"70840553",
  3094 => x"0c727084",
  3095 => x"05540871",
  3096 => x"70840553",
  3097 => x"0cf01252",
  3098 => x"718f26c9",
  3099 => x"38837227",
  3100 => x"95387270",
  3101 => x"84055408",
  3102 => x"71708405",
  3103 => x"530cfc12",
  3104 => x"52718326",
  3105 => x"ed387054",
  3106 => x"ff8339fd",
  3107 => x"3d0d800b",
  3108 => x"80f0d808",
  3109 => x"54547281",
  3110 => x"2e9c3873",
  3111 => x"80f8b40c",
  3112 => x"ffa7bd3f",
  3113 => x"ffa6d93f",
  3114 => x"80f18052",
  3115 => x"8151e9ea",
  3116 => x"3f800851",
  3117 => x"a23f7280",
  3118 => x"f8b40cff",
  3119 => x"a7a23fff",
  3120 => x"a6be3f80",
  3121 => x"f1805281",
  3122 => x"51e9cf3f",
  3123 => x"80085187",
  3124 => x"3f00ff39",
  3125 => x"00ff39f7",
  3126 => x"3d0d7b80",
  3127 => x"f1840882",
  3128 => x"c811085a",
  3129 => x"545a7780",
  3130 => x"2e80da38",
  3131 => x"81881884",
  3132 => x"1908ff05",
  3133 => x"81712b59",
  3134 => x"55598074",
  3135 => x"2480ea38",
  3136 => x"807424b5",
  3137 => x"3873822b",
  3138 => x"78118805",
  3139 => x"56568180",
  3140 => x"19087706",
  3141 => x"5372802e",
  3142 => x"b6387816",
  3143 => x"70085353",
  3144 => x"79517408",
  3145 => x"53722dff",
  3146 => x"14fc17fc",
  3147 => x"1779812c",
  3148 => x"5a575754",
  3149 => x"738025d6",
  3150 => x"38770858",
  3151 => x"77ffad38",
  3152 => x"80f18408",
  3153 => x"53bc1308",
  3154 => x"a5387951",
  3155 => x"ff833f74",
  3156 => x"0853722d",
  3157 => x"ff14fc17",
  3158 => x"fc177981",
  3159 => x"2c5a5757",
  3160 => x"54738025",
  3161 => x"ffa838d1",
  3162 => x"398057ff",
  3163 => x"93397251",
  3164 => x"bc130853",
  3165 => x"722d7951",
  3166 => x"fed73fff",
  3167 => x"3d0d80f8",
  3168 => x"880bfc05",
  3169 => x"70085252",
  3170 => x"70ff2e91",
  3171 => x"38702dfc",
  3172 => x"12700852",
  3173 => x"5270ff2e",
  3174 => x"098106f1",
  3175 => x"38833d0d",
  3176 => x"0404ffa6",
  3177 => x"a83f0400",
  3178 => x"00000040",
  3179 => x"30782020",
  3180 => x"20202020",
  3181 => x"20200000",
  3182 => x"30622020",
  3183 => x"20202020",
  3184 => x"20202020",
  3185 => x"20202020",
  3186 => x"20202020",
  3187 => x"20202020",
  3188 => x"20202020",
  3189 => x"20202020",
  3190 => x"20200000",
  3191 => x"0a677265",
  3192 => x"74682072",
  3193 => x"65676973",
  3194 => x"74657273",
  3195 => x"3a000000",
  3196 => x"0a636f6e",
  3197 => x"74726f6c",
  3198 => x"3a202020",
  3199 => x"20202000",
  3200 => x"0a737461",
  3201 => x"7475733a",
  3202 => x"20202020",
  3203 => x"20202000",
  3204 => x"0a6d6163",
  3205 => x"5f6d7362",
  3206 => x"3a202020",
  3207 => x"20202000",
  3208 => x"0a6d6163",
  3209 => x"5f6c7362",
  3210 => x"3a202020",
  3211 => x"20202000",
  3212 => x"0a6d6469",
  3213 => x"6f5f636f",
  3214 => x"6e74726f",
  3215 => x"6c3a2000",
  3216 => x"0a74785f",
  3217 => x"706f696e",
  3218 => x"7465723a",
  3219 => x"20202000",
  3220 => x"0a72785f",
  3221 => x"706f696e",
  3222 => x"7465723a",
  3223 => x"20202000",
  3224 => x"0a656463",
  3225 => x"6c5f6970",
  3226 => x"3a202020",
  3227 => x"20202000",
  3228 => x"0a686173",
  3229 => x"685f6d73",
  3230 => x"623a2020",
  3231 => x"20202000",
  3232 => x"0a686173",
  3233 => x"685f6c73",
  3234 => x"623a2020",
  3235 => x"20202000",
  3236 => x"0a6d6469",
  3237 => x"6f207068",
  3238 => x"79207265",
  3239 => x"67697374",
  3240 => x"65727300",
  3241 => x"0a206d64",
  3242 => x"696f2070",
  3243 => x"68793a20",
  3244 => x"00000000",
  3245 => x"0a202072",
  3246 => x"65673a20",
  3247 => x"00000000",
  3248 => x"2d3e2000",
  3249 => x"0a677265",
  3250 => x"74682d3e",
  3251 => x"636f6e74",
  3252 => x"726f6c20",
  3253 => x"3a000000",
  3254 => x"0a677265",
  3255 => x"74682d3e",
  3256 => x"73746174",
  3257 => x"75732020",
  3258 => x"3a000000",
  3259 => x"0a646573",
  3260 => x"63722d3e",
  3261 => x"636f6e74",
  3262 => x"726f6c20",
  3263 => x"3a000000",
  3264 => x"77726974",
  3265 => x"65206164",
  3266 => x"64726573",
  3267 => x"733a2000",
  3268 => x"20206c65",
  3269 => x"6e677468",
  3270 => x"3a200000",
  3271 => x"0a0a0000",
  3272 => x"72656164",
  3273 => x"20206164",
  3274 => x"64726573",
  3275 => x"733a2000",
  3276 => x"20206578",
  3277 => x"70656374",
  3278 => x"3a200000",
  3279 => x"2020676f",
  3280 => x"743a2000",
  3281 => x"20657272",
  3282 => x"6f720000",
  3283 => x"0a000000",
  3284 => x"206f6b00",
  3285 => x"70686173",
  3286 => x"65207368",
  3287 => x"69667420",
  3288 => x"202d2020",
  3289 => x"76616c75",
  3290 => x"653a2000",
  3291 => x"20207374",
  3292 => x"61747573",
  3293 => x"3a200000",
  3294 => x"20202020",
  3295 => x"20000000",
  3296 => x"4641494c",
  3297 => x"00000000",
  3298 => x"6f6b2020",
  3299 => x"00000000",
  3300 => x"44445220",
  3301 => x"6d656d6f",
  3302 => x"72792069",
  3303 => x"6e666f00",
  3304 => x"0a617574",
  3305 => x"6f20745f",
  3306 => x"52455245",
  3307 => x"5348203a",
  3308 => x"00000000",
  3309 => x"0a636c6f",
  3310 => x"636b2065",
  3311 => x"6e61626c",
  3312 => x"6520203a",
  3313 => x"00000000",
  3314 => x"0a696e69",
  3315 => x"74616c69",
  3316 => x"7a652020",
  3317 => x"2020203a",
  3318 => x"00000000",
  3319 => x"0a636f6c",
  3320 => x"756d6e20",
  3321 => x"73697a65",
  3322 => x"2020203a",
  3323 => x"00000000",
  3324 => x"0a62616e",
  3325 => x"6b73697a",
  3326 => x"65202020",
  3327 => x"2020203a",
  3328 => x"00000000",
  3329 => x"4d627974",
  3330 => x"65000000",
  3331 => x"0a745f52",
  3332 => x"43442020",
  3333 => x"20202020",
  3334 => x"2020203a",
  3335 => x"00000000",
  3336 => x"0a745f52",
  3337 => x"46432020",
  3338 => x"20202020",
  3339 => x"2020203a",
  3340 => x"00000000",
  3341 => x"0a745f52",
  3342 => x"50202020",
  3343 => x"20202020",
  3344 => x"2020203a",
  3345 => x"00000000",
  3346 => x"0a726566",
  3347 => x"72657368",
  3348 => x"20656e2e",
  3349 => x"2020203a",
  3350 => x"00000000",
  3351 => x"0a444452",
  3352 => x"20667265",
  3353 => x"7175656e",
  3354 => x"6379203a",
  3355 => x"00000000",
  3356 => x"0a444452",
  3357 => x"20646174",
  3358 => x"61207769",
  3359 => x"6474683a",
  3360 => x"00000000",
  3361 => x"0a6d6f62",
  3362 => x"696c6520",
  3363 => x"73757070",
  3364 => x"6f72743a",
  3365 => x"00000000",
  3366 => x"0a73656c",
  3367 => x"66207265",
  3368 => x"66726573",
  3369 => x"6820203a",
  3370 => x"00000000",
  3371 => x"756e6b6e",
  3372 => x"6f776e00",
  3373 => x"20617272",
  3374 => x"61790000",
  3375 => x"0a74656d",
  3376 => x"702d636f",
  3377 => x"6d702072",
  3378 => x"6566723a",
  3379 => x"00000000",
  3380 => x"c2b04300",
  3381 => x"0a647269",
  3382 => x"76652073",
  3383 => x"7472656e",
  3384 => x"6774683a",
  3385 => x"00000000",
  3386 => x"0a706f77",
  3387 => x"65722073",
  3388 => x"6176696e",
  3389 => x"6720203a",
  3390 => x"00000000",
  3391 => x"0a745f58",
  3392 => x"50202020",
  3393 => x"20202020",
  3394 => x"2020203a",
  3395 => x"00000000",
  3396 => x"0a745f58",
  3397 => x"53522020",
  3398 => x"20202020",
  3399 => x"2020203a",
  3400 => x"00000000",
  3401 => x"0a745f43",
  3402 => x"4b452020",
  3403 => x"20202020",
  3404 => x"2020203a",
  3405 => x"00000000",
  3406 => x"0a434153",
  3407 => x"206c6174",
  3408 => x"656e6379",
  3409 => x"2020203a",
  3410 => x"00000000",
  3411 => x"0a6d6f62",
  3412 => x"696c6520",
  3413 => x"656e6162",
  3414 => x"6c65643a",
  3415 => x"00000000",
  3416 => x"0a737461",
  3417 => x"74757320",
  3418 => x"72656164",
  3419 => x"2020203a",
  3420 => x"00000000",
  3421 => x"332f3400",
  3422 => x"38350000",
  3423 => x"68616c66",
  3424 => x"00000000",
  3425 => x"34303639",
  3426 => x"00000000",
  3427 => x"20353132",
  3428 => x"00000000",
  3429 => x"66756c6c",
  3430 => x"00000000",
  3431 => x"37300000",
  3432 => x"34350000",
  3433 => x"31303234",
  3434 => x"00000000",
  3435 => x"31350000",
  3436 => x"312f3400",
  3437 => x"32303438",
  3438 => x"00000000",
  3439 => x"312f3800",
  3440 => x"312f3200",
  3441 => x"312f3100",
  3442 => x"64656570",
  3443 => x"20706f77",
  3444 => x"65722064",
  3445 => x"6f776e00",
  3446 => x"636c6f63",
  3447 => x"6b207374",
  3448 => x"6f700000",
  3449 => x"73656c66",
  3450 => x"20726566",
  3451 => x"72657368",
  3452 => x"00000000",
  3453 => x"706f7765",
  3454 => x"7220646f",
  3455 => x"776e0000",
  3456 => x"6e6f6e65",
  3457 => x"00000000",
  3458 => x"61646472",
  3459 => x"6573733a",
  3460 => x"20000000",
  3461 => x"20646174",
  3462 => x"613a2000",
  3463 => x"0a0a4443",
  3464 => x"4d207068",
  3465 => x"61736520",
  3466 => x"73686966",
  3467 => x"74207465",
  3468 => x"7374696e",
  3469 => x"67000000",
  3470 => x"0a696e69",
  3471 => x"7469616c",
  3472 => x"3a200000",
  3473 => x"09000000",
  3474 => x"20202020",
  3475 => x"00000000",
  3476 => x"6c6f7720",
  3477 => x"666f756e",
  3478 => x"64000000",
  3479 => x"68696768",
  3480 => x"20666f75",
  3481 => x"6e640000",
  3482 => x"0a6c6f77",
  3483 => x"3a202020",
  3484 => x"20202020",
  3485 => x"20200000",
  3486 => x"0a686967",
  3487 => x"683a2020",
  3488 => x"20202020",
  3489 => x"20200000",
  3490 => x"0a646966",
  3491 => x"663a2020",
  3492 => x"20202020",
  3493 => x"20200000",
  3494 => x"0a646966",
  3495 => x"662f323a",
  3496 => x"20202020",
  3497 => x"20200000",
  3498 => x"0a6d696e",
  3499 => x"5f657272",
  3500 => x"3a202020",
  3501 => x"20200000",
  3502 => x"0a6d696e",
  3503 => x"5f657272",
  3504 => x"5f706f73",
  3505 => x"3a200000",
  3506 => x"0a66696e",
  3507 => x"616c3a20",
  3508 => x"20202020",
  3509 => x"20200000",
  3510 => x"68696768",
  3511 => x"204e4f54",
  3512 => x"20666f75",
  3513 => x"6e640000",
  3514 => x"6c6f7720",
  3515 => x"4e4f5420",
  3516 => x"666f756e",
  3517 => x"64000000",
  3518 => x"74657374",
  3519 => x"2e632000",
  3520 => x"286f6e20",
  3521 => x"73696d75",
  3522 => x"6c61746f",
  3523 => x"72290a00",
  3524 => x"636f6d70",
  3525 => x"696c6564",
  3526 => x"3a204f63",
  3527 => x"74203134",
  3528 => x"20323031",
  3529 => x"30202031",
  3530 => x"323a3334",
  3531 => x"3a35350a",
  3532 => x"00000000",
  3533 => x"286f6e20",
  3534 => x"68617264",
  3535 => x"77617265",
  3536 => x"290a0000",
  3537 => x"000006d1",
  3538 => x"000006f7",
  3539 => x"000006f7",
  3540 => x"000006d1",
  3541 => x"000006f7",
  3542 => x"000006f7",
  3543 => x"000006f7",
  3544 => x"000006f7",
  3545 => x"000006f7",
  3546 => x"000006f7",
  3547 => x"000006f7",
  3548 => x"000006f7",
  3549 => x"000006f7",
  3550 => x"000006f7",
  3551 => x"000006f7",
  3552 => x"000006f7",
  3553 => x"000006f7",
  3554 => x"000006f7",
  3555 => x"000006f7",
  3556 => x"000006f7",
  3557 => x"000006f7",
  3558 => x"000006f7",
  3559 => x"000006f7",
  3560 => x"000006f7",
  3561 => x"000006f7",
  3562 => x"000006f7",
  3563 => x"000006f7",
  3564 => x"000006f7",
  3565 => x"000006f7",
  3566 => x"000006f7",
  3567 => x"000006f7",
  3568 => x"000006f7",
  3569 => x"000006f7",
  3570 => x"000006f7",
  3571 => x"000006f7",
  3572 => x"000006f7",
  3573 => x"000006f7",
  3574 => x"000006f7",
  3575 => x"000007a3",
  3576 => x"0000079b",
  3577 => x"00000793",
  3578 => x"0000078b",
  3579 => x"00000783",
  3580 => x"0000077b",
  3581 => x"00000773",
  3582 => x"0000076a",
  3583 => x"00000761",
  3584 => x"00001c9c",
  3585 => x"00001c95",
  3586 => x"00001c8e",
  3587 => x"00001794",
  3588 => x"00001794",
  3589 => x"00001c87",
  3590 => x"00001c87",
  3591 => x"00001ed3",
  3592 => x"00001e47",
  3593 => x"00001dbb",
  3594 => x"00001810",
  3595 => x"00001d2f",
  3596 => x"00001ca3",
  3597 => x"64756d6d",
  3598 => x"792e6578",
  3599 => x"65000000",
  3600 => x"43000000",
  3601 => x"00ffffff",
  3602 => x"ff00ffff",
  3603 => x"ffff00ff",
  3604 => x"ffffff00",
  3605 => x"00000000",
  3606 => x"00000000",
  3607 => x"00000000",
  3608 => x"00003c10",
  3609 => x"fff00000",
  3610 => x"80000e00",
  3611 => x"80000c00",
  3612 => x"80000800",
  3613 => x"80000600",
  3614 => x"80000200",
  3615 => x"80000100",
  3616 => x"00003834",
  3617 => x"00003888",
  3618 => x"00000000",
  3619 => x"00003af0",
  3620 => x"00003b4c",
  3621 => x"00003ba8",
  3622 => x"00000000",
  3623 => x"00000000",
  3624 => x"00000000",
  3625 => x"00000000",
  3626 => x"00000000",
  3627 => x"00000000",
  3628 => x"00000000",
  3629 => x"00000000",
  3630 => x"00000000",
  3631 => x"00003840",
  3632 => x"00000000",
  3633 => x"00000000",
  3634 => x"00000000",
  3635 => x"00000000",
  3636 => x"00000000",
  3637 => x"00000000",
  3638 => x"00000000",
  3639 => x"00000000",
  3640 => x"00000000",
  3641 => x"00000000",
  3642 => x"00000000",
  3643 => x"00000000",
  3644 => x"00000000",
  3645 => x"00000000",
  3646 => x"00000000",
  3647 => x"00000000",
  3648 => x"00000000",
  3649 => x"00000000",
  3650 => x"00000000",
  3651 => x"00000000",
  3652 => x"00000000",
  3653 => x"00000000",
  3654 => x"00000000",
  3655 => x"00000000",
  3656 => x"00000000",
  3657 => x"00000000",
  3658 => x"00000000",
  3659 => x"00000000",
  3660 => x"00000001",
  3661 => x"330eabcd",
  3662 => x"1234e66d",
  3663 => x"deec0005",
  3664 => x"000b0000",
  3665 => x"00000000",
  3666 => x"00000000",
  3667 => x"00000000",
  3668 => x"00000000",
  3669 => x"00000000",
  3670 => x"00000000",
  3671 => x"00000000",
  3672 => x"00000000",
  3673 => x"00000000",
  3674 => x"00000000",
  3675 => x"00000000",
  3676 => x"00000000",
  3677 => x"00000000",
  3678 => x"00000000",
  3679 => x"00000000",
  3680 => x"00000000",
  3681 => x"00000000",
  3682 => x"00000000",
  3683 => x"00000000",
  3684 => x"00000000",
  3685 => x"00000000",
  3686 => x"00000000",
  3687 => x"00000000",
  3688 => x"00000000",
  3689 => x"00000000",
  3690 => x"00000000",
  3691 => x"00000000",
  3692 => x"00000000",
  3693 => x"00000000",
  3694 => x"00000000",
  3695 => x"00000000",
  3696 => x"00000000",
  3697 => x"00000000",
  3698 => x"00000000",
  3699 => x"00000000",
  3700 => x"00000000",
  3701 => x"00000000",
  3702 => x"00000000",
  3703 => x"00000000",
  3704 => x"00000000",
  3705 => x"00000000",
  3706 => x"00000000",
  3707 => x"00000000",
  3708 => x"00000000",
  3709 => x"00000000",
  3710 => x"00000000",
  3711 => x"00000000",
  3712 => x"00000000",
  3713 => x"00000000",
  3714 => x"00000000",
  3715 => x"00000000",
  3716 => x"00000000",
  3717 => x"00000000",
  3718 => x"00000000",
  3719 => x"00000000",
  3720 => x"00000000",
  3721 => x"00000000",
  3722 => x"00000000",
  3723 => x"00000000",
  3724 => x"00000000",
  3725 => x"00000000",
  3726 => x"00000000",
  3727 => x"00000000",
  3728 => x"00000000",
  3729 => x"00000000",
  3730 => x"00000000",
  3731 => x"00000000",
  3732 => x"00000000",
  3733 => x"00000000",
  3734 => x"00000000",
  3735 => x"00000000",
  3736 => x"00000000",
  3737 => x"00000000",
  3738 => x"00000000",
  3739 => x"00000000",
  3740 => x"00000000",
  3741 => x"00000000",
  3742 => x"00000000",
  3743 => x"00000000",
  3744 => x"00000000",
  3745 => x"00000000",
  3746 => x"00000000",
  3747 => x"00000000",
  3748 => x"00000000",
  3749 => x"00000000",
  3750 => x"00000000",
  3751 => x"00000000",
  3752 => x"00000000",
  3753 => x"00000000",
  3754 => x"00000000",
  3755 => x"00000000",
  3756 => x"00000000",
  3757 => x"00000000",
  3758 => x"00000000",
  3759 => x"00000000",
  3760 => x"00000000",
  3761 => x"00000000",
  3762 => x"00000000",
  3763 => x"00000000",
  3764 => x"00000000",
  3765 => x"00000000",
  3766 => x"00000000",
  3767 => x"00000000",
  3768 => x"00000000",
  3769 => x"00000000",
  3770 => x"00000000",
  3771 => x"00000000",
  3772 => x"00000000",
  3773 => x"00000000",
  3774 => x"00000000",
  3775 => x"00000000",
  3776 => x"00000000",
  3777 => x"00000000",
  3778 => x"00000000",
  3779 => x"00000000",
  3780 => x"00000000",
  3781 => x"00000000",
  3782 => x"00000000",
  3783 => x"00000000",
  3784 => x"00000000",
  3785 => x"00000000",
  3786 => x"00000000",
  3787 => x"00000000",
  3788 => x"00000000",
  3789 => x"00000000",
  3790 => x"00000000",
  3791 => x"00000000",
  3792 => x"00000000",
  3793 => x"00000000",
  3794 => x"00000000",
  3795 => x"00000000",
  3796 => x"00000000",
  3797 => x"00000000",
  3798 => x"00000000",
  3799 => x"00000000",
  3800 => x"00000000",
  3801 => x"00000000",
  3802 => x"00000000",
  3803 => x"00000000",
  3804 => x"00000000",
  3805 => x"00000000",
  3806 => x"00000000",
  3807 => x"00000000",
  3808 => x"00000000",
  3809 => x"00000000",
  3810 => x"00000000",
  3811 => x"00000000",
  3812 => x"00000000",
  3813 => x"00000000",
  3814 => x"00000000",
  3815 => x"00000000",
  3816 => x"00000000",
  3817 => x"00000000",
  3818 => x"00000000",
  3819 => x"00000000",
  3820 => x"00000000",
  3821 => x"00000000",
  3822 => x"00000000",
  3823 => x"00000000",
  3824 => x"00000000",
  3825 => x"00000000",
  3826 => x"00000000",
  3827 => x"00000000",
  3828 => x"00000000",
  3829 => x"00000000",
  3830 => x"00000000",
  3831 => x"00000000",
  3832 => x"00000000",
  3833 => x"00000000",
  3834 => x"00000000",
  3835 => x"00000000",
  3836 => x"00000000",
  3837 => x"00000000",
  3838 => x"00000000",
  3839 => x"00000000",
  3840 => x"00000000",
  3841 => x"ffffffff",
  3842 => x"00000000",
  3843 => x"ffffffff",
  3844 => x"00000000",
  3845 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (memAWriteEnable = '1') then
			ram(to_integer(unsigned(memAAddr))) := memAWrite;
			memARead <= memAWrite;
		else
			memARead <= ram(to_integer(unsigned(memAAddr)));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (memBWriteEnable = '1') then
			ram(to_integer(unsigned(memBAddr))) := memBWrite;
			memBRead <= memBWrite;
		else
			memBRead <= ram(to_integer(unsigned(memBAddr)));
		end if;
	end if;
end process;




end dualport_ram_arch;
